module Regfile(
  input         clock,
  input  [5:0]  io_readPorts_0_addr,
  output [63:0] io_readPorts_0_data,
  input  [5:0]  io_readPorts_1_addr,
  output [63:0] io_readPorts_1_data,
  input  [5:0]  io_readPorts_2_addr,
  output [63:0] io_readPorts_2_data,
  input  [5:0]  io_readPorts_3_addr,
  output [63:0] io_readPorts_3_data,
  input  [5:0]  io_readPorts_4_addr,
  output [63:0] io_readPorts_4_data,
  input  [5:0]  io_readPorts_5_addr,
  output [63:0] io_readPorts_5_data,
  input  [5:0]  io_readPorts_6_addr,
  output [63:0] io_readPorts_6_data,
  input  [5:0]  io_readPorts_7_addr,
  output [63:0] io_readPorts_7_data,
  input  [5:0]  io_readPorts_8_addr,
  output [63:0] io_readPorts_8_data,
  input  [5:0]  io_readPorts_9_addr,
  output [63:0] io_readPorts_9_data,
  input         io_writePorts_0_wen,
  input  [5:0]  io_writePorts_0_addr,
  input  [63:0] io_writePorts_0_data,
  input         io_writePorts_1_wen,
  input  [5:0]  io_writePorts_1_addr,
  input  [63:0] io_writePorts_1_data,
  input         io_writePorts_2_wen,
  input  [5:0]  io_writePorts_2_addr,
  input  [63:0] io_writePorts_2_data,
  input         io_writePorts_3_wen,
  input  [5:0]  io_writePorts_3_addr,
  input  [63:0] io_writePorts_3_data,
  input         io_writePorts_4_wen,
  input  [5:0]  io_writePorts_4_addr,
  input  [63:0] io_writePorts_4_data,
  input  [5:0]  io_debug_rports_0_addr,
  output [63:0] io_debug_rports_0_data,
  input  [5:0]  io_debug_rports_1_addr,
  output [63:0] io_debug_rports_1_data,
  input  [5:0]  io_debug_rports_2_addr,
  output [63:0] io_debug_rports_2_data,
  input  [5:0]  io_debug_rports_3_addr,
  output [63:0] io_debug_rports_3_data,
  input  [5:0]  io_debug_rports_4_addr,
  output [63:0] io_debug_rports_4_data,
  input  [5:0]  io_debug_rports_5_addr,
  output [63:0] io_debug_rports_5_data,
  input  [5:0]  io_debug_rports_6_addr,
  output [63:0] io_debug_rports_6_data,
  input  [5:0]  io_debug_rports_7_addr,
  output [63:0] io_debug_rports_7_data,
  input  [5:0]  io_debug_rports_8_addr,
  output [63:0] io_debug_rports_8_data,
  input  [5:0]  io_debug_rports_9_addr,
  output [63:0] io_debug_rports_9_data,
  input  [5:0]  io_debug_rports_10_addr,
  output [63:0] io_debug_rports_10_data,
  input  [5:0]  io_debug_rports_11_addr,
  output [63:0] io_debug_rports_11_data,
  input  [5:0]  io_debug_rports_12_addr,
  output [63:0] io_debug_rports_12_data,
  input  [5:0]  io_debug_rports_13_addr,
  output [63:0] io_debug_rports_13_data,
  input  [5:0]  io_debug_rports_14_addr,
  output [63:0] io_debug_rports_14_data,
  input  [5:0]  io_debug_rports_15_addr,
  output [63:0] io_debug_rports_15_data,
  input  [5:0]  io_debug_rports_16_addr,
  output [63:0] io_debug_rports_16_data,
  input  [5:0]  io_debug_rports_17_addr,
  output [63:0] io_debug_rports_17_data,
  input  [5:0]  io_debug_rports_18_addr,
  output [63:0] io_debug_rports_18_data,
  input  [5:0]  io_debug_rports_19_addr,
  output [63:0] io_debug_rports_19_data,
  input  [5:0]  io_debug_rports_20_addr,
  output [63:0] io_debug_rports_20_data,
  input  [5:0]  io_debug_rports_21_addr,
  output [63:0] io_debug_rports_21_data,
  input  [5:0]  io_debug_rports_22_addr,
  output [63:0] io_debug_rports_22_data,
  input  [5:0]  io_debug_rports_23_addr,
  output [63:0] io_debug_rports_23_data,
  input  [5:0]  io_debug_rports_24_addr,
  output [63:0] io_debug_rports_24_data,
  input  [5:0]  io_debug_rports_25_addr,
  output [63:0] io_debug_rports_25_data,
  input  [5:0]  io_debug_rports_26_addr,
  output [63:0] io_debug_rports_26_data,
  input  [5:0]  io_debug_rports_27_addr,
  output [63:0] io_debug_rports_27_data,
  input  [5:0]  io_debug_rports_28_addr,
  output [63:0] io_debug_rports_28_data,
  input  [5:0]  io_debug_rports_29_addr,
  output [63:0] io_debug_rports_29_data,
  input  [5:0]  io_debug_rports_30_addr,
  output [63:0] io_debug_rports_30_data,
  input  [5:0]  io_debug_rports_31_addr,
  output [63:0] io_debug_rports_31_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [63:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [63:0] _RAND_39;
  reg [63:0] _RAND_40;
  reg [63:0] _RAND_41;
  reg [63:0] _RAND_42;
  reg [63:0] _RAND_43;
  reg [63:0] _RAND_44;
  reg [63:0] _RAND_45;
  reg [63:0] _RAND_46;
  reg [63:0] _RAND_47;
  reg [63:0] _RAND_48;
  reg [63:0] _RAND_49;
  reg [63:0] _RAND_50;
  reg [63:0] _RAND_51;
  reg [63:0] _RAND_52;
  reg [63:0] _RAND_53;
  reg [63:0] _RAND_54;
  reg [63:0] _RAND_55;
  reg [63:0] _RAND_56;
  reg [63:0] _RAND_57;
  reg [63:0] _RAND_58;
  reg [63:0] _RAND_59;
  reg [63:0] _RAND_60;
  reg [63:0] _RAND_61;
  reg [63:0] _RAND_62;
  reg [63:0] _RAND_63;
  reg [63:0] _RAND_64;
  reg [63:0] _RAND_65;
  reg [63:0] _RAND_66;
  reg [63:0] _RAND_67;
  reg [63:0] _RAND_68;
  reg [63:0] _RAND_69;
  reg [63:0] _RAND_70;
  reg [63:0] _RAND_71;
  reg [63:0] _RAND_72;
  reg [63:0] _RAND_73;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] mem_0; // @[Regfile.scala 51:16]
  reg [63:0] mem_1; // @[Regfile.scala 51:16]
  reg [63:0] mem_2; // @[Regfile.scala 51:16]
  reg [63:0] mem_3; // @[Regfile.scala 51:16]
  reg [63:0] mem_4; // @[Regfile.scala 51:16]
  reg [63:0] mem_5; // @[Regfile.scala 51:16]
  reg [63:0] mem_6; // @[Regfile.scala 51:16]
  reg [63:0] mem_7; // @[Regfile.scala 51:16]
  reg [63:0] mem_8; // @[Regfile.scala 51:16]
  reg [63:0] mem_9; // @[Regfile.scala 51:16]
  reg [63:0] mem_10; // @[Regfile.scala 51:16]
  reg [63:0] mem_11; // @[Regfile.scala 51:16]
  reg [63:0] mem_12; // @[Regfile.scala 51:16]
  reg [63:0] mem_13; // @[Regfile.scala 51:16]
  reg [63:0] mem_14; // @[Regfile.scala 51:16]
  reg [63:0] mem_15; // @[Regfile.scala 51:16]
  reg [63:0] mem_16; // @[Regfile.scala 51:16]
  reg [63:0] mem_17; // @[Regfile.scala 51:16]
  reg [63:0] mem_18; // @[Regfile.scala 51:16]
  reg [63:0] mem_19; // @[Regfile.scala 51:16]
  reg [63:0] mem_20; // @[Regfile.scala 51:16]
  reg [63:0] mem_21; // @[Regfile.scala 51:16]
  reg [63:0] mem_22; // @[Regfile.scala 51:16]
  reg [63:0] mem_23; // @[Regfile.scala 51:16]
  reg [63:0] mem_24; // @[Regfile.scala 51:16]
  reg [63:0] mem_25; // @[Regfile.scala 51:16]
  reg [63:0] mem_26; // @[Regfile.scala 51:16]
  reg [63:0] mem_27; // @[Regfile.scala 51:16]
  reg [63:0] mem_28; // @[Regfile.scala 51:16]
  reg [63:0] mem_29; // @[Regfile.scala 51:16]
  reg [63:0] mem_30; // @[Regfile.scala 51:16]
  reg [63:0] mem_31; // @[Regfile.scala 51:16]
  reg [63:0] mem_32; // @[Regfile.scala 51:16]
  reg [63:0] mem_33; // @[Regfile.scala 51:16]
  reg [63:0] mem_34; // @[Regfile.scala 51:16]
  reg [63:0] mem_35; // @[Regfile.scala 51:16]
  reg [63:0] mem_36; // @[Regfile.scala 51:16]
  reg [63:0] mem_37; // @[Regfile.scala 51:16]
  reg [63:0] mem_38; // @[Regfile.scala 51:16]
  reg [63:0] mem_39; // @[Regfile.scala 51:16]
  reg [63:0] mem_40; // @[Regfile.scala 51:16]
  reg [63:0] mem_41; // @[Regfile.scala 51:16]
  reg [63:0] mem_42; // @[Regfile.scala 51:16]
  reg [63:0] mem_43; // @[Regfile.scala 51:16]
  reg [63:0] mem_44; // @[Regfile.scala 51:16]
  reg [63:0] mem_45; // @[Regfile.scala 51:16]
  reg [63:0] mem_46; // @[Regfile.scala 51:16]
  reg [63:0] mem_47; // @[Regfile.scala 51:16]
  reg [63:0] mem_48; // @[Regfile.scala 51:16]
  reg [63:0] mem_49; // @[Regfile.scala 51:16]
  reg [63:0] mem_50; // @[Regfile.scala 51:16]
  reg [63:0] mem_51; // @[Regfile.scala 51:16]
  reg [63:0] mem_52; // @[Regfile.scala 51:16]
  reg [63:0] mem_53; // @[Regfile.scala 51:16]
  reg [63:0] mem_54; // @[Regfile.scala 51:16]
  reg [63:0] mem_55; // @[Regfile.scala 51:16]
  reg [63:0] mem_56; // @[Regfile.scala 51:16]
  reg [63:0] mem_57; // @[Regfile.scala 51:16]
  reg [63:0] mem_58; // @[Regfile.scala 51:16]
  reg [63:0] mem_59; // @[Regfile.scala 51:16]
  reg [63:0] mem_60; // @[Regfile.scala 51:16]
  reg [63:0] mem_61; // @[Regfile.scala 51:16]
  reg [63:0] mem_62; // @[Regfile.scala 51:16]
  reg [63:0] mem_63; // @[Regfile.scala 51:16]
  wire [63:0] _GEN_1 = 6'h1 == io_readPorts_0_addr ? mem_1 : mem_0; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_2 = 6'h2 == io_readPorts_0_addr ? mem_2 : _GEN_1; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_3 = 6'h3 == io_readPorts_0_addr ? mem_3 : _GEN_2; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_4 = 6'h4 == io_readPorts_0_addr ? mem_4 : _GEN_3; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_5 = 6'h5 == io_readPorts_0_addr ? mem_5 : _GEN_4; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_6 = 6'h6 == io_readPorts_0_addr ? mem_6 : _GEN_5; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_7 = 6'h7 == io_readPorts_0_addr ? mem_7 : _GEN_6; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_8 = 6'h8 == io_readPorts_0_addr ? mem_8 : _GEN_7; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_9 = 6'h9 == io_readPorts_0_addr ? mem_9 : _GEN_8; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_10 = 6'ha == io_readPorts_0_addr ? mem_10 : _GEN_9; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_11 = 6'hb == io_readPorts_0_addr ? mem_11 : _GEN_10; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_12 = 6'hc == io_readPorts_0_addr ? mem_12 : _GEN_11; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_13 = 6'hd == io_readPorts_0_addr ? mem_13 : _GEN_12; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_14 = 6'he == io_readPorts_0_addr ? mem_14 : _GEN_13; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_15 = 6'hf == io_readPorts_0_addr ? mem_15 : _GEN_14; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_16 = 6'h10 == io_readPorts_0_addr ? mem_16 : _GEN_15; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_17 = 6'h11 == io_readPorts_0_addr ? mem_17 : _GEN_16; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_18 = 6'h12 == io_readPorts_0_addr ? mem_18 : _GEN_17; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_19 = 6'h13 == io_readPorts_0_addr ? mem_19 : _GEN_18; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_20 = 6'h14 == io_readPorts_0_addr ? mem_20 : _GEN_19; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_21 = 6'h15 == io_readPorts_0_addr ? mem_21 : _GEN_20; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_22 = 6'h16 == io_readPorts_0_addr ? mem_22 : _GEN_21; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_23 = 6'h17 == io_readPorts_0_addr ? mem_23 : _GEN_22; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_24 = 6'h18 == io_readPorts_0_addr ? mem_24 : _GEN_23; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_25 = 6'h19 == io_readPorts_0_addr ? mem_25 : _GEN_24; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_26 = 6'h1a == io_readPorts_0_addr ? mem_26 : _GEN_25; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_27 = 6'h1b == io_readPorts_0_addr ? mem_27 : _GEN_26; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_28 = 6'h1c == io_readPorts_0_addr ? mem_28 : _GEN_27; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_29 = 6'h1d == io_readPorts_0_addr ? mem_29 : _GEN_28; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_30 = 6'h1e == io_readPorts_0_addr ? mem_30 : _GEN_29; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_31 = 6'h1f == io_readPorts_0_addr ? mem_31 : _GEN_30; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_32 = 6'h20 == io_readPorts_0_addr ? mem_32 : _GEN_31; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_33 = 6'h21 == io_readPorts_0_addr ? mem_33 : _GEN_32; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_34 = 6'h22 == io_readPorts_0_addr ? mem_34 : _GEN_33; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_35 = 6'h23 == io_readPorts_0_addr ? mem_35 : _GEN_34; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_36 = 6'h24 == io_readPorts_0_addr ? mem_36 : _GEN_35; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_37 = 6'h25 == io_readPorts_0_addr ? mem_37 : _GEN_36; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_38 = 6'h26 == io_readPorts_0_addr ? mem_38 : _GEN_37; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_39 = 6'h27 == io_readPorts_0_addr ? mem_39 : _GEN_38; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_40 = 6'h28 == io_readPorts_0_addr ? mem_40 : _GEN_39; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_41 = 6'h29 == io_readPorts_0_addr ? mem_41 : _GEN_40; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_42 = 6'h2a == io_readPorts_0_addr ? mem_42 : _GEN_41; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_43 = 6'h2b == io_readPorts_0_addr ? mem_43 : _GEN_42; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_44 = 6'h2c == io_readPorts_0_addr ? mem_44 : _GEN_43; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_45 = 6'h2d == io_readPorts_0_addr ? mem_45 : _GEN_44; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_46 = 6'h2e == io_readPorts_0_addr ? mem_46 : _GEN_45; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_47 = 6'h2f == io_readPorts_0_addr ? mem_47 : _GEN_46; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_48 = 6'h30 == io_readPorts_0_addr ? mem_48 : _GEN_47; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_49 = 6'h31 == io_readPorts_0_addr ? mem_49 : _GEN_48; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_50 = 6'h32 == io_readPorts_0_addr ? mem_50 : _GEN_49; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_51 = 6'h33 == io_readPorts_0_addr ? mem_51 : _GEN_50; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_52 = 6'h34 == io_readPorts_0_addr ? mem_52 : _GEN_51; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_53 = 6'h35 == io_readPorts_0_addr ? mem_53 : _GEN_52; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_54 = 6'h36 == io_readPorts_0_addr ? mem_54 : _GEN_53; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_55 = 6'h37 == io_readPorts_0_addr ? mem_55 : _GEN_54; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_56 = 6'h38 == io_readPorts_0_addr ? mem_56 : _GEN_55; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_57 = 6'h39 == io_readPorts_0_addr ? mem_57 : _GEN_56; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_58 = 6'h3a == io_readPorts_0_addr ? mem_58 : _GEN_57; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_59 = 6'h3b == io_readPorts_0_addr ? mem_59 : _GEN_58; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_60 = 6'h3c == io_readPorts_0_addr ? mem_60 : _GEN_59; // @[Regfile.scala 53:{33,33}]
  reg [63:0] io_readPorts_0_data_REG; // @[Regfile.scala 54:22]
  wire [63:0] _GEN_65 = 6'h1 == io_readPorts_1_addr ? mem_1 : mem_0; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_66 = 6'h2 == io_readPorts_1_addr ? mem_2 : _GEN_65; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_67 = 6'h3 == io_readPorts_1_addr ? mem_3 : _GEN_66; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_68 = 6'h4 == io_readPorts_1_addr ? mem_4 : _GEN_67; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_69 = 6'h5 == io_readPorts_1_addr ? mem_5 : _GEN_68; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_70 = 6'h6 == io_readPorts_1_addr ? mem_6 : _GEN_69; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_71 = 6'h7 == io_readPorts_1_addr ? mem_7 : _GEN_70; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_72 = 6'h8 == io_readPorts_1_addr ? mem_8 : _GEN_71; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_73 = 6'h9 == io_readPorts_1_addr ? mem_9 : _GEN_72; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_74 = 6'ha == io_readPorts_1_addr ? mem_10 : _GEN_73; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_75 = 6'hb == io_readPorts_1_addr ? mem_11 : _GEN_74; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_76 = 6'hc == io_readPorts_1_addr ? mem_12 : _GEN_75; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_77 = 6'hd == io_readPorts_1_addr ? mem_13 : _GEN_76; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_78 = 6'he == io_readPorts_1_addr ? mem_14 : _GEN_77; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_79 = 6'hf == io_readPorts_1_addr ? mem_15 : _GEN_78; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_80 = 6'h10 == io_readPorts_1_addr ? mem_16 : _GEN_79; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_81 = 6'h11 == io_readPorts_1_addr ? mem_17 : _GEN_80; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_82 = 6'h12 == io_readPorts_1_addr ? mem_18 : _GEN_81; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_83 = 6'h13 == io_readPorts_1_addr ? mem_19 : _GEN_82; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_84 = 6'h14 == io_readPorts_1_addr ? mem_20 : _GEN_83; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_85 = 6'h15 == io_readPorts_1_addr ? mem_21 : _GEN_84; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_86 = 6'h16 == io_readPorts_1_addr ? mem_22 : _GEN_85; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_87 = 6'h17 == io_readPorts_1_addr ? mem_23 : _GEN_86; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_88 = 6'h18 == io_readPorts_1_addr ? mem_24 : _GEN_87; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_89 = 6'h19 == io_readPorts_1_addr ? mem_25 : _GEN_88; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_90 = 6'h1a == io_readPorts_1_addr ? mem_26 : _GEN_89; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_91 = 6'h1b == io_readPorts_1_addr ? mem_27 : _GEN_90; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_92 = 6'h1c == io_readPorts_1_addr ? mem_28 : _GEN_91; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_93 = 6'h1d == io_readPorts_1_addr ? mem_29 : _GEN_92; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_94 = 6'h1e == io_readPorts_1_addr ? mem_30 : _GEN_93; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_95 = 6'h1f == io_readPorts_1_addr ? mem_31 : _GEN_94; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_96 = 6'h20 == io_readPorts_1_addr ? mem_32 : _GEN_95; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_97 = 6'h21 == io_readPorts_1_addr ? mem_33 : _GEN_96; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_98 = 6'h22 == io_readPorts_1_addr ? mem_34 : _GEN_97; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_99 = 6'h23 == io_readPorts_1_addr ? mem_35 : _GEN_98; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_100 = 6'h24 == io_readPorts_1_addr ? mem_36 : _GEN_99; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_101 = 6'h25 == io_readPorts_1_addr ? mem_37 : _GEN_100; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_102 = 6'h26 == io_readPorts_1_addr ? mem_38 : _GEN_101; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_103 = 6'h27 == io_readPorts_1_addr ? mem_39 : _GEN_102; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_104 = 6'h28 == io_readPorts_1_addr ? mem_40 : _GEN_103; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_105 = 6'h29 == io_readPorts_1_addr ? mem_41 : _GEN_104; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_106 = 6'h2a == io_readPorts_1_addr ? mem_42 : _GEN_105; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_107 = 6'h2b == io_readPorts_1_addr ? mem_43 : _GEN_106; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_108 = 6'h2c == io_readPorts_1_addr ? mem_44 : _GEN_107; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_109 = 6'h2d == io_readPorts_1_addr ? mem_45 : _GEN_108; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_110 = 6'h2e == io_readPorts_1_addr ? mem_46 : _GEN_109; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_111 = 6'h2f == io_readPorts_1_addr ? mem_47 : _GEN_110; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_112 = 6'h30 == io_readPorts_1_addr ? mem_48 : _GEN_111; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_113 = 6'h31 == io_readPorts_1_addr ? mem_49 : _GEN_112; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_114 = 6'h32 == io_readPorts_1_addr ? mem_50 : _GEN_113; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_115 = 6'h33 == io_readPorts_1_addr ? mem_51 : _GEN_114; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_116 = 6'h34 == io_readPorts_1_addr ? mem_52 : _GEN_115; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_117 = 6'h35 == io_readPorts_1_addr ? mem_53 : _GEN_116; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_118 = 6'h36 == io_readPorts_1_addr ? mem_54 : _GEN_117; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_119 = 6'h37 == io_readPorts_1_addr ? mem_55 : _GEN_118; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_120 = 6'h38 == io_readPorts_1_addr ? mem_56 : _GEN_119; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_121 = 6'h39 == io_readPorts_1_addr ? mem_57 : _GEN_120; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_122 = 6'h3a == io_readPorts_1_addr ? mem_58 : _GEN_121; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_123 = 6'h3b == io_readPorts_1_addr ? mem_59 : _GEN_122; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_124 = 6'h3c == io_readPorts_1_addr ? mem_60 : _GEN_123; // @[Regfile.scala 53:{33,33}]
  reg [63:0] io_readPorts_1_data_REG; // @[Regfile.scala 54:22]
  wire [63:0] _GEN_129 = 6'h1 == io_readPorts_2_addr ? mem_1 : mem_0; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_130 = 6'h2 == io_readPorts_2_addr ? mem_2 : _GEN_129; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_131 = 6'h3 == io_readPorts_2_addr ? mem_3 : _GEN_130; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_132 = 6'h4 == io_readPorts_2_addr ? mem_4 : _GEN_131; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_133 = 6'h5 == io_readPorts_2_addr ? mem_5 : _GEN_132; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_134 = 6'h6 == io_readPorts_2_addr ? mem_6 : _GEN_133; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_135 = 6'h7 == io_readPorts_2_addr ? mem_7 : _GEN_134; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_136 = 6'h8 == io_readPorts_2_addr ? mem_8 : _GEN_135; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_137 = 6'h9 == io_readPorts_2_addr ? mem_9 : _GEN_136; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_138 = 6'ha == io_readPorts_2_addr ? mem_10 : _GEN_137; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_139 = 6'hb == io_readPorts_2_addr ? mem_11 : _GEN_138; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_140 = 6'hc == io_readPorts_2_addr ? mem_12 : _GEN_139; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_141 = 6'hd == io_readPorts_2_addr ? mem_13 : _GEN_140; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_142 = 6'he == io_readPorts_2_addr ? mem_14 : _GEN_141; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_143 = 6'hf == io_readPorts_2_addr ? mem_15 : _GEN_142; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_144 = 6'h10 == io_readPorts_2_addr ? mem_16 : _GEN_143; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_145 = 6'h11 == io_readPorts_2_addr ? mem_17 : _GEN_144; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_146 = 6'h12 == io_readPorts_2_addr ? mem_18 : _GEN_145; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_147 = 6'h13 == io_readPorts_2_addr ? mem_19 : _GEN_146; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_148 = 6'h14 == io_readPorts_2_addr ? mem_20 : _GEN_147; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_149 = 6'h15 == io_readPorts_2_addr ? mem_21 : _GEN_148; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_150 = 6'h16 == io_readPorts_2_addr ? mem_22 : _GEN_149; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_151 = 6'h17 == io_readPorts_2_addr ? mem_23 : _GEN_150; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_152 = 6'h18 == io_readPorts_2_addr ? mem_24 : _GEN_151; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_153 = 6'h19 == io_readPorts_2_addr ? mem_25 : _GEN_152; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_154 = 6'h1a == io_readPorts_2_addr ? mem_26 : _GEN_153; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_155 = 6'h1b == io_readPorts_2_addr ? mem_27 : _GEN_154; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_156 = 6'h1c == io_readPorts_2_addr ? mem_28 : _GEN_155; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_157 = 6'h1d == io_readPorts_2_addr ? mem_29 : _GEN_156; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_158 = 6'h1e == io_readPorts_2_addr ? mem_30 : _GEN_157; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_159 = 6'h1f == io_readPorts_2_addr ? mem_31 : _GEN_158; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_160 = 6'h20 == io_readPorts_2_addr ? mem_32 : _GEN_159; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_161 = 6'h21 == io_readPorts_2_addr ? mem_33 : _GEN_160; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_162 = 6'h22 == io_readPorts_2_addr ? mem_34 : _GEN_161; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_163 = 6'h23 == io_readPorts_2_addr ? mem_35 : _GEN_162; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_164 = 6'h24 == io_readPorts_2_addr ? mem_36 : _GEN_163; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_165 = 6'h25 == io_readPorts_2_addr ? mem_37 : _GEN_164; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_166 = 6'h26 == io_readPorts_2_addr ? mem_38 : _GEN_165; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_167 = 6'h27 == io_readPorts_2_addr ? mem_39 : _GEN_166; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_168 = 6'h28 == io_readPorts_2_addr ? mem_40 : _GEN_167; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_169 = 6'h29 == io_readPorts_2_addr ? mem_41 : _GEN_168; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_170 = 6'h2a == io_readPorts_2_addr ? mem_42 : _GEN_169; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_171 = 6'h2b == io_readPorts_2_addr ? mem_43 : _GEN_170; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_172 = 6'h2c == io_readPorts_2_addr ? mem_44 : _GEN_171; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_173 = 6'h2d == io_readPorts_2_addr ? mem_45 : _GEN_172; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_174 = 6'h2e == io_readPorts_2_addr ? mem_46 : _GEN_173; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_175 = 6'h2f == io_readPorts_2_addr ? mem_47 : _GEN_174; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_176 = 6'h30 == io_readPorts_2_addr ? mem_48 : _GEN_175; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_177 = 6'h31 == io_readPorts_2_addr ? mem_49 : _GEN_176; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_178 = 6'h32 == io_readPorts_2_addr ? mem_50 : _GEN_177; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_179 = 6'h33 == io_readPorts_2_addr ? mem_51 : _GEN_178; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_180 = 6'h34 == io_readPorts_2_addr ? mem_52 : _GEN_179; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_181 = 6'h35 == io_readPorts_2_addr ? mem_53 : _GEN_180; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_182 = 6'h36 == io_readPorts_2_addr ? mem_54 : _GEN_181; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_183 = 6'h37 == io_readPorts_2_addr ? mem_55 : _GEN_182; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_184 = 6'h38 == io_readPorts_2_addr ? mem_56 : _GEN_183; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_185 = 6'h39 == io_readPorts_2_addr ? mem_57 : _GEN_184; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_186 = 6'h3a == io_readPorts_2_addr ? mem_58 : _GEN_185; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_187 = 6'h3b == io_readPorts_2_addr ? mem_59 : _GEN_186; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_188 = 6'h3c == io_readPorts_2_addr ? mem_60 : _GEN_187; // @[Regfile.scala 53:{33,33}]
  reg [63:0] io_readPorts_2_data_REG; // @[Regfile.scala 54:22]
  wire [63:0] _GEN_193 = 6'h1 == io_readPorts_3_addr ? mem_1 : mem_0; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_194 = 6'h2 == io_readPorts_3_addr ? mem_2 : _GEN_193; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_195 = 6'h3 == io_readPorts_3_addr ? mem_3 : _GEN_194; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_196 = 6'h4 == io_readPorts_3_addr ? mem_4 : _GEN_195; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_197 = 6'h5 == io_readPorts_3_addr ? mem_5 : _GEN_196; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_198 = 6'h6 == io_readPorts_3_addr ? mem_6 : _GEN_197; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_199 = 6'h7 == io_readPorts_3_addr ? mem_7 : _GEN_198; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_200 = 6'h8 == io_readPorts_3_addr ? mem_8 : _GEN_199; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_201 = 6'h9 == io_readPorts_3_addr ? mem_9 : _GEN_200; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_202 = 6'ha == io_readPorts_3_addr ? mem_10 : _GEN_201; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_203 = 6'hb == io_readPorts_3_addr ? mem_11 : _GEN_202; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_204 = 6'hc == io_readPorts_3_addr ? mem_12 : _GEN_203; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_205 = 6'hd == io_readPorts_3_addr ? mem_13 : _GEN_204; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_206 = 6'he == io_readPorts_3_addr ? mem_14 : _GEN_205; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_207 = 6'hf == io_readPorts_3_addr ? mem_15 : _GEN_206; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_208 = 6'h10 == io_readPorts_3_addr ? mem_16 : _GEN_207; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_209 = 6'h11 == io_readPorts_3_addr ? mem_17 : _GEN_208; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_210 = 6'h12 == io_readPorts_3_addr ? mem_18 : _GEN_209; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_211 = 6'h13 == io_readPorts_3_addr ? mem_19 : _GEN_210; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_212 = 6'h14 == io_readPorts_3_addr ? mem_20 : _GEN_211; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_213 = 6'h15 == io_readPorts_3_addr ? mem_21 : _GEN_212; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_214 = 6'h16 == io_readPorts_3_addr ? mem_22 : _GEN_213; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_215 = 6'h17 == io_readPorts_3_addr ? mem_23 : _GEN_214; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_216 = 6'h18 == io_readPorts_3_addr ? mem_24 : _GEN_215; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_217 = 6'h19 == io_readPorts_3_addr ? mem_25 : _GEN_216; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_218 = 6'h1a == io_readPorts_3_addr ? mem_26 : _GEN_217; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_219 = 6'h1b == io_readPorts_3_addr ? mem_27 : _GEN_218; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_220 = 6'h1c == io_readPorts_3_addr ? mem_28 : _GEN_219; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_221 = 6'h1d == io_readPorts_3_addr ? mem_29 : _GEN_220; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_222 = 6'h1e == io_readPorts_3_addr ? mem_30 : _GEN_221; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_223 = 6'h1f == io_readPorts_3_addr ? mem_31 : _GEN_222; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_224 = 6'h20 == io_readPorts_3_addr ? mem_32 : _GEN_223; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_225 = 6'h21 == io_readPorts_3_addr ? mem_33 : _GEN_224; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_226 = 6'h22 == io_readPorts_3_addr ? mem_34 : _GEN_225; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_227 = 6'h23 == io_readPorts_3_addr ? mem_35 : _GEN_226; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_228 = 6'h24 == io_readPorts_3_addr ? mem_36 : _GEN_227; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_229 = 6'h25 == io_readPorts_3_addr ? mem_37 : _GEN_228; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_230 = 6'h26 == io_readPorts_3_addr ? mem_38 : _GEN_229; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_231 = 6'h27 == io_readPorts_3_addr ? mem_39 : _GEN_230; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_232 = 6'h28 == io_readPorts_3_addr ? mem_40 : _GEN_231; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_233 = 6'h29 == io_readPorts_3_addr ? mem_41 : _GEN_232; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_234 = 6'h2a == io_readPorts_3_addr ? mem_42 : _GEN_233; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_235 = 6'h2b == io_readPorts_3_addr ? mem_43 : _GEN_234; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_236 = 6'h2c == io_readPorts_3_addr ? mem_44 : _GEN_235; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_237 = 6'h2d == io_readPorts_3_addr ? mem_45 : _GEN_236; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_238 = 6'h2e == io_readPorts_3_addr ? mem_46 : _GEN_237; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_239 = 6'h2f == io_readPorts_3_addr ? mem_47 : _GEN_238; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_240 = 6'h30 == io_readPorts_3_addr ? mem_48 : _GEN_239; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_241 = 6'h31 == io_readPorts_3_addr ? mem_49 : _GEN_240; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_242 = 6'h32 == io_readPorts_3_addr ? mem_50 : _GEN_241; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_243 = 6'h33 == io_readPorts_3_addr ? mem_51 : _GEN_242; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_244 = 6'h34 == io_readPorts_3_addr ? mem_52 : _GEN_243; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_245 = 6'h35 == io_readPorts_3_addr ? mem_53 : _GEN_244; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_246 = 6'h36 == io_readPorts_3_addr ? mem_54 : _GEN_245; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_247 = 6'h37 == io_readPorts_3_addr ? mem_55 : _GEN_246; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_248 = 6'h38 == io_readPorts_3_addr ? mem_56 : _GEN_247; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_249 = 6'h39 == io_readPorts_3_addr ? mem_57 : _GEN_248; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_250 = 6'h3a == io_readPorts_3_addr ? mem_58 : _GEN_249; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_251 = 6'h3b == io_readPorts_3_addr ? mem_59 : _GEN_250; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_252 = 6'h3c == io_readPorts_3_addr ? mem_60 : _GEN_251; // @[Regfile.scala 53:{33,33}]
  reg [63:0] io_readPorts_3_data_REG; // @[Regfile.scala 54:22]
  wire [63:0] _GEN_257 = 6'h1 == io_readPorts_4_addr ? mem_1 : mem_0; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_258 = 6'h2 == io_readPorts_4_addr ? mem_2 : _GEN_257; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_259 = 6'h3 == io_readPorts_4_addr ? mem_3 : _GEN_258; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_260 = 6'h4 == io_readPorts_4_addr ? mem_4 : _GEN_259; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_261 = 6'h5 == io_readPorts_4_addr ? mem_5 : _GEN_260; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_262 = 6'h6 == io_readPorts_4_addr ? mem_6 : _GEN_261; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_263 = 6'h7 == io_readPorts_4_addr ? mem_7 : _GEN_262; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_264 = 6'h8 == io_readPorts_4_addr ? mem_8 : _GEN_263; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_265 = 6'h9 == io_readPorts_4_addr ? mem_9 : _GEN_264; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_266 = 6'ha == io_readPorts_4_addr ? mem_10 : _GEN_265; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_267 = 6'hb == io_readPorts_4_addr ? mem_11 : _GEN_266; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_268 = 6'hc == io_readPorts_4_addr ? mem_12 : _GEN_267; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_269 = 6'hd == io_readPorts_4_addr ? mem_13 : _GEN_268; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_270 = 6'he == io_readPorts_4_addr ? mem_14 : _GEN_269; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_271 = 6'hf == io_readPorts_4_addr ? mem_15 : _GEN_270; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_272 = 6'h10 == io_readPorts_4_addr ? mem_16 : _GEN_271; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_273 = 6'h11 == io_readPorts_4_addr ? mem_17 : _GEN_272; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_274 = 6'h12 == io_readPorts_4_addr ? mem_18 : _GEN_273; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_275 = 6'h13 == io_readPorts_4_addr ? mem_19 : _GEN_274; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_276 = 6'h14 == io_readPorts_4_addr ? mem_20 : _GEN_275; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_277 = 6'h15 == io_readPorts_4_addr ? mem_21 : _GEN_276; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_278 = 6'h16 == io_readPorts_4_addr ? mem_22 : _GEN_277; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_279 = 6'h17 == io_readPorts_4_addr ? mem_23 : _GEN_278; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_280 = 6'h18 == io_readPorts_4_addr ? mem_24 : _GEN_279; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_281 = 6'h19 == io_readPorts_4_addr ? mem_25 : _GEN_280; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_282 = 6'h1a == io_readPorts_4_addr ? mem_26 : _GEN_281; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_283 = 6'h1b == io_readPorts_4_addr ? mem_27 : _GEN_282; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_284 = 6'h1c == io_readPorts_4_addr ? mem_28 : _GEN_283; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_285 = 6'h1d == io_readPorts_4_addr ? mem_29 : _GEN_284; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_286 = 6'h1e == io_readPorts_4_addr ? mem_30 : _GEN_285; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_287 = 6'h1f == io_readPorts_4_addr ? mem_31 : _GEN_286; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_288 = 6'h20 == io_readPorts_4_addr ? mem_32 : _GEN_287; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_289 = 6'h21 == io_readPorts_4_addr ? mem_33 : _GEN_288; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_290 = 6'h22 == io_readPorts_4_addr ? mem_34 : _GEN_289; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_291 = 6'h23 == io_readPorts_4_addr ? mem_35 : _GEN_290; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_292 = 6'h24 == io_readPorts_4_addr ? mem_36 : _GEN_291; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_293 = 6'h25 == io_readPorts_4_addr ? mem_37 : _GEN_292; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_294 = 6'h26 == io_readPorts_4_addr ? mem_38 : _GEN_293; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_295 = 6'h27 == io_readPorts_4_addr ? mem_39 : _GEN_294; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_296 = 6'h28 == io_readPorts_4_addr ? mem_40 : _GEN_295; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_297 = 6'h29 == io_readPorts_4_addr ? mem_41 : _GEN_296; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_298 = 6'h2a == io_readPorts_4_addr ? mem_42 : _GEN_297; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_299 = 6'h2b == io_readPorts_4_addr ? mem_43 : _GEN_298; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_300 = 6'h2c == io_readPorts_4_addr ? mem_44 : _GEN_299; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_301 = 6'h2d == io_readPorts_4_addr ? mem_45 : _GEN_300; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_302 = 6'h2e == io_readPorts_4_addr ? mem_46 : _GEN_301; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_303 = 6'h2f == io_readPorts_4_addr ? mem_47 : _GEN_302; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_304 = 6'h30 == io_readPorts_4_addr ? mem_48 : _GEN_303; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_305 = 6'h31 == io_readPorts_4_addr ? mem_49 : _GEN_304; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_306 = 6'h32 == io_readPorts_4_addr ? mem_50 : _GEN_305; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_307 = 6'h33 == io_readPorts_4_addr ? mem_51 : _GEN_306; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_308 = 6'h34 == io_readPorts_4_addr ? mem_52 : _GEN_307; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_309 = 6'h35 == io_readPorts_4_addr ? mem_53 : _GEN_308; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_310 = 6'h36 == io_readPorts_4_addr ? mem_54 : _GEN_309; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_311 = 6'h37 == io_readPorts_4_addr ? mem_55 : _GEN_310; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_312 = 6'h38 == io_readPorts_4_addr ? mem_56 : _GEN_311; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_313 = 6'h39 == io_readPorts_4_addr ? mem_57 : _GEN_312; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_314 = 6'h3a == io_readPorts_4_addr ? mem_58 : _GEN_313; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_315 = 6'h3b == io_readPorts_4_addr ? mem_59 : _GEN_314; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_316 = 6'h3c == io_readPorts_4_addr ? mem_60 : _GEN_315; // @[Regfile.scala 53:{33,33}]
  reg [63:0] io_readPorts_4_data_REG; // @[Regfile.scala 54:22]
  wire [63:0] _GEN_321 = 6'h1 == io_readPorts_5_addr ? mem_1 : mem_0; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_322 = 6'h2 == io_readPorts_5_addr ? mem_2 : _GEN_321; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_323 = 6'h3 == io_readPorts_5_addr ? mem_3 : _GEN_322; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_324 = 6'h4 == io_readPorts_5_addr ? mem_4 : _GEN_323; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_325 = 6'h5 == io_readPorts_5_addr ? mem_5 : _GEN_324; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_326 = 6'h6 == io_readPorts_5_addr ? mem_6 : _GEN_325; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_327 = 6'h7 == io_readPorts_5_addr ? mem_7 : _GEN_326; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_328 = 6'h8 == io_readPorts_5_addr ? mem_8 : _GEN_327; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_329 = 6'h9 == io_readPorts_5_addr ? mem_9 : _GEN_328; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_330 = 6'ha == io_readPorts_5_addr ? mem_10 : _GEN_329; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_331 = 6'hb == io_readPorts_5_addr ? mem_11 : _GEN_330; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_332 = 6'hc == io_readPorts_5_addr ? mem_12 : _GEN_331; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_333 = 6'hd == io_readPorts_5_addr ? mem_13 : _GEN_332; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_334 = 6'he == io_readPorts_5_addr ? mem_14 : _GEN_333; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_335 = 6'hf == io_readPorts_5_addr ? mem_15 : _GEN_334; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_336 = 6'h10 == io_readPorts_5_addr ? mem_16 : _GEN_335; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_337 = 6'h11 == io_readPorts_5_addr ? mem_17 : _GEN_336; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_338 = 6'h12 == io_readPorts_5_addr ? mem_18 : _GEN_337; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_339 = 6'h13 == io_readPorts_5_addr ? mem_19 : _GEN_338; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_340 = 6'h14 == io_readPorts_5_addr ? mem_20 : _GEN_339; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_341 = 6'h15 == io_readPorts_5_addr ? mem_21 : _GEN_340; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_342 = 6'h16 == io_readPorts_5_addr ? mem_22 : _GEN_341; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_343 = 6'h17 == io_readPorts_5_addr ? mem_23 : _GEN_342; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_344 = 6'h18 == io_readPorts_5_addr ? mem_24 : _GEN_343; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_345 = 6'h19 == io_readPorts_5_addr ? mem_25 : _GEN_344; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_346 = 6'h1a == io_readPorts_5_addr ? mem_26 : _GEN_345; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_347 = 6'h1b == io_readPorts_5_addr ? mem_27 : _GEN_346; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_348 = 6'h1c == io_readPorts_5_addr ? mem_28 : _GEN_347; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_349 = 6'h1d == io_readPorts_5_addr ? mem_29 : _GEN_348; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_350 = 6'h1e == io_readPorts_5_addr ? mem_30 : _GEN_349; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_351 = 6'h1f == io_readPorts_5_addr ? mem_31 : _GEN_350; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_352 = 6'h20 == io_readPorts_5_addr ? mem_32 : _GEN_351; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_353 = 6'h21 == io_readPorts_5_addr ? mem_33 : _GEN_352; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_354 = 6'h22 == io_readPorts_5_addr ? mem_34 : _GEN_353; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_355 = 6'h23 == io_readPorts_5_addr ? mem_35 : _GEN_354; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_356 = 6'h24 == io_readPorts_5_addr ? mem_36 : _GEN_355; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_357 = 6'h25 == io_readPorts_5_addr ? mem_37 : _GEN_356; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_358 = 6'h26 == io_readPorts_5_addr ? mem_38 : _GEN_357; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_359 = 6'h27 == io_readPorts_5_addr ? mem_39 : _GEN_358; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_360 = 6'h28 == io_readPorts_5_addr ? mem_40 : _GEN_359; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_361 = 6'h29 == io_readPorts_5_addr ? mem_41 : _GEN_360; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_362 = 6'h2a == io_readPorts_5_addr ? mem_42 : _GEN_361; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_363 = 6'h2b == io_readPorts_5_addr ? mem_43 : _GEN_362; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_364 = 6'h2c == io_readPorts_5_addr ? mem_44 : _GEN_363; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_365 = 6'h2d == io_readPorts_5_addr ? mem_45 : _GEN_364; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_366 = 6'h2e == io_readPorts_5_addr ? mem_46 : _GEN_365; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_367 = 6'h2f == io_readPorts_5_addr ? mem_47 : _GEN_366; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_368 = 6'h30 == io_readPorts_5_addr ? mem_48 : _GEN_367; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_369 = 6'h31 == io_readPorts_5_addr ? mem_49 : _GEN_368; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_370 = 6'h32 == io_readPorts_5_addr ? mem_50 : _GEN_369; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_371 = 6'h33 == io_readPorts_5_addr ? mem_51 : _GEN_370; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_372 = 6'h34 == io_readPorts_5_addr ? mem_52 : _GEN_371; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_373 = 6'h35 == io_readPorts_5_addr ? mem_53 : _GEN_372; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_374 = 6'h36 == io_readPorts_5_addr ? mem_54 : _GEN_373; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_375 = 6'h37 == io_readPorts_5_addr ? mem_55 : _GEN_374; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_376 = 6'h38 == io_readPorts_5_addr ? mem_56 : _GEN_375; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_377 = 6'h39 == io_readPorts_5_addr ? mem_57 : _GEN_376; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_378 = 6'h3a == io_readPorts_5_addr ? mem_58 : _GEN_377; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_379 = 6'h3b == io_readPorts_5_addr ? mem_59 : _GEN_378; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_380 = 6'h3c == io_readPorts_5_addr ? mem_60 : _GEN_379; // @[Regfile.scala 53:{33,33}]
  reg [63:0] io_readPorts_5_data_REG; // @[Regfile.scala 54:22]
  wire [63:0] _GEN_385 = 6'h1 == io_readPorts_6_addr ? mem_1 : mem_0; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_386 = 6'h2 == io_readPorts_6_addr ? mem_2 : _GEN_385; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_387 = 6'h3 == io_readPorts_6_addr ? mem_3 : _GEN_386; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_388 = 6'h4 == io_readPorts_6_addr ? mem_4 : _GEN_387; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_389 = 6'h5 == io_readPorts_6_addr ? mem_5 : _GEN_388; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_390 = 6'h6 == io_readPorts_6_addr ? mem_6 : _GEN_389; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_391 = 6'h7 == io_readPorts_6_addr ? mem_7 : _GEN_390; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_392 = 6'h8 == io_readPorts_6_addr ? mem_8 : _GEN_391; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_393 = 6'h9 == io_readPorts_6_addr ? mem_9 : _GEN_392; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_394 = 6'ha == io_readPorts_6_addr ? mem_10 : _GEN_393; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_395 = 6'hb == io_readPorts_6_addr ? mem_11 : _GEN_394; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_396 = 6'hc == io_readPorts_6_addr ? mem_12 : _GEN_395; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_397 = 6'hd == io_readPorts_6_addr ? mem_13 : _GEN_396; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_398 = 6'he == io_readPorts_6_addr ? mem_14 : _GEN_397; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_399 = 6'hf == io_readPorts_6_addr ? mem_15 : _GEN_398; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_400 = 6'h10 == io_readPorts_6_addr ? mem_16 : _GEN_399; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_401 = 6'h11 == io_readPorts_6_addr ? mem_17 : _GEN_400; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_402 = 6'h12 == io_readPorts_6_addr ? mem_18 : _GEN_401; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_403 = 6'h13 == io_readPorts_6_addr ? mem_19 : _GEN_402; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_404 = 6'h14 == io_readPorts_6_addr ? mem_20 : _GEN_403; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_405 = 6'h15 == io_readPorts_6_addr ? mem_21 : _GEN_404; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_406 = 6'h16 == io_readPorts_6_addr ? mem_22 : _GEN_405; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_407 = 6'h17 == io_readPorts_6_addr ? mem_23 : _GEN_406; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_408 = 6'h18 == io_readPorts_6_addr ? mem_24 : _GEN_407; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_409 = 6'h19 == io_readPorts_6_addr ? mem_25 : _GEN_408; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_410 = 6'h1a == io_readPorts_6_addr ? mem_26 : _GEN_409; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_411 = 6'h1b == io_readPorts_6_addr ? mem_27 : _GEN_410; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_412 = 6'h1c == io_readPorts_6_addr ? mem_28 : _GEN_411; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_413 = 6'h1d == io_readPorts_6_addr ? mem_29 : _GEN_412; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_414 = 6'h1e == io_readPorts_6_addr ? mem_30 : _GEN_413; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_415 = 6'h1f == io_readPorts_6_addr ? mem_31 : _GEN_414; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_416 = 6'h20 == io_readPorts_6_addr ? mem_32 : _GEN_415; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_417 = 6'h21 == io_readPorts_6_addr ? mem_33 : _GEN_416; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_418 = 6'h22 == io_readPorts_6_addr ? mem_34 : _GEN_417; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_419 = 6'h23 == io_readPorts_6_addr ? mem_35 : _GEN_418; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_420 = 6'h24 == io_readPorts_6_addr ? mem_36 : _GEN_419; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_421 = 6'h25 == io_readPorts_6_addr ? mem_37 : _GEN_420; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_422 = 6'h26 == io_readPorts_6_addr ? mem_38 : _GEN_421; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_423 = 6'h27 == io_readPorts_6_addr ? mem_39 : _GEN_422; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_424 = 6'h28 == io_readPorts_6_addr ? mem_40 : _GEN_423; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_425 = 6'h29 == io_readPorts_6_addr ? mem_41 : _GEN_424; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_426 = 6'h2a == io_readPorts_6_addr ? mem_42 : _GEN_425; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_427 = 6'h2b == io_readPorts_6_addr ? mem_43 : _GEN_426; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_428 = 6'h2c == io_readPorts_6_addr ? mem_44 : _GEN_427; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_429 = 6'h2d == io_readPorts_6_addr ? mem_45 : _GEN_428; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_430 = 6'h2e == io_readPorts_6_addr ? mem_46 : _GEN_429; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_431 = 6'h2f == io_readPorts_6_addr ? mem_47 : _GEN_430; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_432 = 6'h30 == io_readPorts_6_addr ? mem_48 : _GEN_431; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_433 = 6'h31 == io_readPorts_6_addr ? mem_49 : _GEN_432; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_434 = 6'h32 == io_readPorts_6_addr ? mem_50 : _GEN_433; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_435 = 6'h33 == io_readPorts_6_addr ? mem_51 : _GEN_434; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_436 = 6'h34 == io_readPorts_6_addr ? mem_52 : _GEN_435; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_437 = 6'h35 == io_readPorts_6_addr ? mem_53 : _GEN_436; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_438 = 6'h36 == io_readPorts_6_addr ? mem_54 : _GEN_437; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_439 = 6'h37 == io_readPorts_6_addr ? mem_55 : _GEN_438; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_440 = 6'h38 == io_readPorts_6_addr ? mem_56 : _GEN_439; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_441 = 6'h39 == io_readPorts_6_addr ? mem_57 : _GEN_440; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_442 = 6'h3a == io_readPorts_6_addr ? mem_58 : _GEN_441; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_443 = 6'h3b == io_readPorts_6_addr ? mem_59 : _GEN_442; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_444 = 6'h3c == io_readPorts_6_addr ? mem_60 : _GEN_443; // @[Regfile.scala 53:{33,33}]
  reg [63:0] io_readPorts_6_data_REG; // @[Regfile.scala 54:22]
  wire [63:0] _GEN_449 = 6'h1 == io_readPorts_7_addr ? mem_1 : mem_0; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_450 = 6'h2 == io_readPorts_7_addr ? mem_2 : _GEN_449; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_451 = 6'h3 == io_readPorts_7_addr ? mem_3 : _GEN_450; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_452 = 6'h4 == io_readPorts_7_addr ? mem_4 : _GEN_451; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_453 = 6'h5 == io_readPorts_7_addr ? mem_5 : _GEN_452; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_454 = 6'h6 == io_readPorts_7_addr ? mem_6 : _GEN_453; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_455 = 6'h7 == io_readPorts_7_addr ? mem_7 : _GEN_454; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_456 = 6'h8 == io_readPorts_7_addr ? mem_8 : _GEN_455; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_457 = 6'h9 == io_readPorts_7_addr ? mem_9 : _GEN_456; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_458 = 6'ha == io_readPorts_7_addr ? mem_10 : _GEN_457; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_459 = 6'hb == io_readPorts_7_addr ? mem_11 : _GEN_458; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_460 = 6'hc == io_readPorts_7_addr ? mem_12 : _GEN_459; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_461 = 6'hd == io_readPorts_7_addr ? mem_13 : _GEN_460; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_462 = 6'he == io_readPorts_7_addr ? mem_14 : _GEN_461; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_463 = 6'hf == io_readPorts_7_addr ? mem_15 : _GEN_462; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_464 = 6'h10 == io_readPorts_7_addr ? mem_16 : _GEN_463; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_465 = 6'h11 == io_readPorts_7_addr ? mem_17 : _GEN_464; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_466 = 6'h12 == io_readPorts_7_addr ? mem_18 : _GEN_465; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_467 = 6'h13 == io_readPorts_7_addr ? mem_19 : _GEN_466; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_468 = 6'h14 == io_readPorts_7_addr ? mem_20 : _GEN_467; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_469 = 6'h15 == io_readPorts_7_addr ? mem_21 : _GEN_468; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_470 = 6'h16 == io_readPorts_7_addr ? mem_22 : _GEN_469; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_471 = 6'h17 == io_readPorts_7_addr ? mem_23 : _GEN_470; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_472 = 6'h18 == io_readPorts_7_addr ? mem_24 : _GEN_471; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_473 = 6'h19 == io_readPorts_7_addr ? mem_25 : _GEN_472; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_474 = 6'h1a == io_readPorts_7_addr ? mem_26 : _GEN_473; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_475 = 6'h1b == io_readPorts_7_addr ? mem_27 : _GEN_474; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_476 = 6'h1c == io_readPorts_7_addr ? mem_28 : _GEN_475; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_477 = 6'h1d == io_readPorts_7_addr ? mem_29 : _GEN_476; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_478 = 6'h1e == io_readPorts_7_addr ? mem_30 : _GEN_477; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_479 = 6'h1f == io_readPorts_7_addr ? mem_31 : _GEN_478; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_480 = 6'h20 == io_readPorts_7_addr ? mem_32 : _GEN_479; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_481 = 6'h21 == io_readPorts_7_addr ? mem_33 : _GEN_480; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_482 = 6'h22 == io_readPorts_7_addr ? mem_34 : _GEN_481; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_483 = 6'h23 == io_readPorts_7_addr ? mem_35 : _GEN_482; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_484 = 6'h24 == io_readPorts_7_addr ? mem_36 : _GEN_483; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_485 = 6'h25 == io_readPorts_7_addr ? mem_37 : _GEN_484; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_486 = 6'h26 == io_readPorts_7_addr ? mem_38 : _GEN_485; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_487 = 6'h27 == io_readPorts_7_addr ? mem_39 : _GEN_486; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_488 = 6'h28 == io_readPorts_7_addr ? mem_40 : _GEN_487; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_489 = 6'h29 == io_readPorts_7_addr ? mem_41 : _GEN_488; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_490 = 6'h2a == io_readPorts_7_addr ? mem_42 : _GEN_489; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_491 = 6'h2b == io_readPorts_7_addr ? mem_43 : _GEN_490; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_492 = 6'h2c == io_readPorts_7_addr ? mem_44 : _GEN_491; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_493 = 6'h2d == io_readPorts_7_addr ? mem_45 : _GEN_492; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_494 = 6'h2e == io_readPorts_7_addr ? mem_46 : _GEN_493; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_495 = 6'h2f == io_readPorts_7_addr ? mem_47 : _GEN_494; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_496 = 6'h30 == io_readPorts_7_addr ? mem_48 : _GEN_495; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_497 = 6'h31 == io_readPorts_7_addr ? mem_49 : _GEN_496; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_498 = 6'h32 == io_readPorts_7_addr ? mem_50 : _GEN_497; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_499 = 6'h33 == io_readPorts_7_addr ? mem_51 : _GEN_498; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_500 = 6'h34 == io_readPorts_7_addr ? mem_52 : _GEN_499; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_501 = 6'h35 == io_readPorts_7_addr ? mem_53 : _GEN_500; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_502 = 6'h36 == io_readPorts_7_addr ? mem_54 : _GEN_501; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_503 = 6'h37 == io_readPorts_7_addr ? mem_55 : _GEN_502; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_504 = 6'h38 == io_readPorts_7_addr ? mem_56 : _GEN_503; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_505 = 6'h39 == io_readPorts_7_addr ? mem_57 : _GEN_504; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_506 = 6'h3a == io_readPorts_7_addr ? mem_58 : _GEN_505; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_507 = 6'h3b == io_readPorts_7_addr ? mem_59 : _GEN_506; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_508 = 6'h3c == io_readPorts_7_addr ? mem_60 : _GEN_507; // @[Regfile.scala 53:{33,33}]
  reg [63:0] io_readPorts_7_data_REG; // @[Regfile.scala 54:22]
  wire [63:0] _GEN_513 = 6'h1 == io_readPorts_8_addr ? mem_1 : mem_0; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_514 = 6'h2 == io_readPorts_8_addr ? mem_2 : _GEN_513; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_515 = 6'h3 == io_readPorts_8_addr ? mem_3 : _GEN_514; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_516 = 6'h4 == io_readPorts_8_addr ? mem_4 : _GEN_515; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_517 = 6'h5 == io_readPorts_8_addr ? mem_5 : _GEN_516; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_518 = 6'h6 == io_readPorts_8_addr ? mem_6 : _GEN_517; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_519 = 6'h7 == io_readPorts_8_addr ? mem_7 : _GEN_518; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_520 = 6'h8 == io_readPorts_8_addr ? mem_8 : _GEN_519; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_521 = 6'h9 == io_readPorts_8_addr ? mem_9 : _GEN_520; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_522 = 6'ha == io_readPorts_8_addr ? mem_10 : _GEN_521; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_523 = 6'hb == io_readPorts_8_addr ? mem_11 : _GEN_522; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_524 = 6'hc == io_readPorts_8_addr ? mem_12 : _GEN_523; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_525 = 6'hd == io_readPorts_8_addr ? mem_13 : _GEN_524; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_526 = 6'he == io_readPorts_8_addr ? mem_14 : _GEN_525; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_527 = 6'hf == io_readPorts_8_addr ? mem_15 : _GEN_526; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_528 = 6'h10 == io_readPorts_8_addr ? mem_16 : _GEN_527; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_529 = 6'h11 == io_readPorts_8_addr ? mem_17 : _GEN_528; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_530 = 6'h12 == io_readPorts_8_addr ? mem_18 : _GEN_529; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_531 = 6'h13 == io_readPorts_8_addr ? mem_19 : _GEN_530; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_532 = 6'h14 == io_readPorts_8_addr ? mem_20 : _GEN_531; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_533 = 6'h15 == io_readPorts_8_addr ? mem_21 : _GEN_532; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_534 = 6'h16 == io_readPorts_8_addr ? mem_22 : _GEN_533; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_535 = 6'h17 == io_readPorts_8_addr ? mem_23 : _GEN_534; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_536 = 6'h18 == io_readPorts_8_addr ? mem_24 : _GEN_535; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_537 = 6'h19 == io_readPorts_8_addr ? mem_25 : _GEN_536; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_538 = 6'h1a == io_readPorts_8_addr ? mem_26 : _GEN_537; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_539 = 6'h1b == io_readPorts_8_addr ? mem_27 : _GEN_538; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_540 = 6'h1c == io_readPorts_8_addr ? mem_28 : _GEN_539; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_541 = 6'h1d == io_readPorts_8_addr ? mem_29 : _GEN_540; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_542 = 6'h1e == io_readPorts_8_addr ? mem_30 : _GEN_541; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_543 = 6'h1f == io_readPorts_8_addr ? mem_31 : _GEN_542; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_544 = 6'h20 == io_readPorts_8_addr ? mem_32 : _GEN_543; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_545 = 6'h21 == io_readPorts_8_addr ? mem_33 : _GEN_544; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_546 = 6'h22 == io_readPorts_8_addr ? mem_34 : _GEN_545; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_547 = 6'h23 == io_readPorts_8_addr ? mem_35 : _GEN_546; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_548 = 6'h24 == io_readPorts_8_addr ? mem_36 : _GEN_547; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_549 = 6'h25 == io_readPorts_8_addr ? mem_37 : _GEN_548; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_550 = 6'h26 == io_readPorts_8_addr ? mem_38 : _GEN_549; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_551 = 6'h27 == io_readPorts_8_addr ? mem_39 : _GEN_550; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_552 = 6'h28 == io_readPorts_8_addr ? mem_40 : _GEN_551; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_553 = 6'h29 == io_readPorts_8_addr ? mem_41 : _GEN_552; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_554 = 6'h2a == io_readPorts_8_addr ? mem_42 : _GEN_553; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_555 = 6'h2b == io_readPorts_8_addr ? mem_43 : _GEN_554; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_556 = 6'h2c == io_readPorts_8_addr ? mem_44 : _GEN_555; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_557 = 6'h2d == io_readPorts_8_addr ? mem_45 : _GEN_556; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_558 = 6'h2e == io_readPorts_8_addr ? mem_46 : _GEN_557; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_559 = 6'h2f == io_readPorts_8_addr ? mem_47 : _GEN_558; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_560 = 6'h30 == io_readPorts_8_addr ? mem_48 : _GEN_559; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_561 = 6'h31 == io_readPorts_8_addr ? mem_49 : _GEN_560; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_562 = 6'h32 == io_readPorts_8_addr ? mem_50 : _GEN_561; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_563 = 6'h33 == io_readPorts_8_addr ? mem_51 : _GEN_562; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_564 = 6'h34 == io_readPorts_8_addr ? mem_52 : _GEN_563; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_565 = 6'h35 == io_readPorts_8_addr ? mem_53 : _GEN_564; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_566 = 6'h36 == io_readPorts_8_addr ? mem_54 : _GEN_565; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_567 = 6'h37 == io_readPorts_8_addr ? mem_55 : _GEN_566; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_568 = 6'h38 == io_readPorts_8_addr ? mem_56 : _GEN_567; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_569 = 6'h39 == io_readPorts_8_addr ? mem_57 : _GEN_568; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_570 = 6'h3a == io_readPorts_8_addr ? mem_58 : _GEN_569; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_571 = 6'h3b == io_readPorts_8_addr ? mem_59 : _GEN_570; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_572 = 6'h3c == io_readPorts_8_addr ? mem_60 : _GEN_571; // @[Regfile.scala 53:{33,33}]
  reg [63:0] io_readPorts_8_data_REG; // @[Regfile.scala 54:22]
  wire [63:0] _GEN_577 = 6'h1 == io_readPorts_9_addr ? mem_1 : mem_0; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_578 = 6'h2 == io_readPorts_9_addr ? mem_2 : _GEN_577; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_579 = 6'h3 == io_readPorts_9_addr ? mem_3 : _GEN_578; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_580 = 6'h4 == io_readPorts_9_addr ? mem_4 : _GEN_579; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_581 = 6'h5 == io_readPorts_9_addr ? mem_5 : _GEN_580; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_582 = 6'h6 == io_readPorts_9_addr ? mem_6 : _GEN_581; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_583 = 6'h7 == io_readPorts_9_addr ? mem_7 : _GEN_582; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_584 = 6'h8 == io_readPorts_9_addr ? mem_8 : _GEN_583; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_585 = 6'h9 == io_readPorts_9_addr ? mem_9 : _GEN_584; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_586 = 6'ha == io_readPorts_9_addr ? mem_10 : _GEN_585; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_587 = 6'hb == io_readPorts_9_addr ? mem_11 : _GEN_586; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_588 = 6'hc == io_readPorts_9_addr ? mem_12 : _GEN_587; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_589 = 6'hd == io_readPorts_9_addr ? mem_13 : _GEN_588; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_590 = 6'he == io_readPorts_9_addr ? mem_14 : _GEN_589; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_591 = 6'hf == io_readPorts_9_addr ? mem_15 : _GEN_590; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_592 = 6'h10 == io_readPorts_9_addr ? mem_16 : _GEN_591; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_593 = 6'h11 == io_readPorts_9_addr ? mem_17 : _GEN_592; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_594 = 6'h12 == io_readPorts_9_addr ? mem_18 : _GEN_593; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_595 = 6'h13 == io_readPorts_9_addr ? mem_19 : _GEN_594; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_596 = 6'h14 == io_readPorts_9_addr ? mem_20 : _GEN_595; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_597 = 6'h15 == io_readPorts_9_addr ? mem_21 : _GEN_596; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_598 = 6'h16 == io_readPorts_9_addr ? mem_22 : _GEN_597; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_599 = 6'h17 == io_readPorts_9_addr ? mem_23 : _GEN_598; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_600 = 6'h18 == io_readPorts_9_addr ? mem_24 : _GEN_599; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_601 = 6'h19 == io_readPorts_9_addr ? mem_25 : _GEN_600; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_602 = 6'h1a == io_readPorts_9_addr ? mem_26 : _GEN_601; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_603 = 6'h1b == io_readPorts_9_addr ? mem_27 : _GEN_602; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_604 = 6'h1c == io_readPorts_9_addr ? mem_28 : _GEN_603; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_605 = 6'h1d == io_readPorts_9_addr ? mem_29 : _GEN_604; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_606 = 6'h1e == io_readPorts_9_addr ? mem_30 : _GEN_605; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_607 = 6'h1f == io_readPorts_9_addr ? mem_31 : _GEN_606; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_608 = 6'h20 == io_readPorts_9_addr ? mem_32 : _GEN_607; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_609 = 6'h21 == io_readPorts_9_addr ? mem_33 : _GEN_608; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_610 = 6'h22 == io_readPorts_9_addr ? mem_34 : _GEN_609; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_611 = 6'h23 == io_readPorts_9_addr ? mem_35 : _GEN_610; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_612 = 6'h24 == io_readPorts_9_addr ? mem_36 : _GEN_611; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_613 = 6'h25 == io_readPorts_9_addr ? mem_37 : _GEN_612; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_614 = 6'h26 == io_readPorts_9_addr ? mem_38 : _GEN_613; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_615 = 6'h27 == io_readPorts_9_addr ? mem_39 : _GEN_614; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_616 = 6'h28 == io_readPorts_9_addr ? mem_40 : _GEN_615; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_617 = 6'h29 == io_readPorts_9_addr ? mem_41 : _GEN_616; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_618 = 6'h2a == io_readPorts_9_addr ? mem_42 : _GEN_617; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_619 = 6'h2b == io_readPorts_9_addr ? mem_43 : _GEN_618; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_620 = 6'h2c == io_readPorts_9_addr ? mem_44 : _GEN_619; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_621 = 6'h2d == io_readPorts_9_addr ? mem_45 : _GEN_620; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_622 = 6'h2e == io_readPorts_9_addr ? mem_46 : _GEN_621; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_623 = 6'h2f == io_readPorts_9_addr ? mem_47 : _GEN_622; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_624 = 6'h30 == io_readPorts_9_addr ? mem_48 : _GEN_623; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_625 = 6'h31 == io_readPorts_9_addr ? mem_49 : _GEN_624; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_626 = 6'h32 == io_readPorts_9_addr ? mem_50 : _GEN_625; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_627 = 6'h33 == io_readPorts_9_addr ? mem_51 : _GEN_626; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_628 = 6'h34 == io_readPorts_9_addr ? mem_52 : _GEN_627; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_629 = 6'h35 == io_readPorts_9_addr ? mem_53 : _GEN_628; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_630 = 6'h36 == io_readPorts_9_addr ? mem_54 : _GEN_629; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_631 = 6'h37 == io_readPorts_9_addr ? mem_55 : _GEN_630; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_632 = 6'h38 == io_readPorts_9_addr ? mem_56 : _GEN_631; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_633 = 6'h39 == io_readPorts_9_addr ? mem_57 : _GEN_632; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_634 = 6'h3a == io_readPorts_9_addr ? mem_58 : _GEN_633; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_635 = 6'h3b == io_readPorts_9_addr ? mem_59 : _GEN_634; // @[Regfile.scala 53:{33,33}]
  wire [63:0] _GEN_636 = 6'h3c == io_readPorts_9_addr ? mem_60 : _GEN_635; // @[Regfile.scala 53:{33,33}]
  reg [63:0] io_readPorts_9_data_REG; // @[Regfile.scala 54:22]
  wire [63:0] _GEN_640 = 6'h0 == io_writePorts_0_addr ? io_writePorts_0_data : mem_0; // @[Regfile.scala 51:16 58:{19,19}]
  wire [63:0] _GEN_641 = 6'h1 == io_writePorts_0_addr ? io_writePorts_0_data : mem_1; // @[Regfile.scala 51:16 58:{19,19}]
  wire [63:0] _GEN_642 = 6'h2 == io_writePorts_0_addr ? io_writePorts_0_data : mem_2; // @[Regfile.scala 51:16 58:{19,19}]
  wire [63:0] _GEN_643 = 6'h3 == io_writePorts_0_addr ? io_writePorts_0_data : mem_3; // @[Regfile.scala 51:16 58:{19,19}]
  wire [63:0] _GEN_644 = 6'h4 == io_writePorts_0_addr ? io_writePorts_0_data : mem_4; // @[Regfile.scala 51:16 58:{19,19}]
  wire [63:0] _GEN_645 = 6'h5 == io_writePorts_0_addr ? io_writePorts_0_data : mem_5; // @[Regfile.scala 51:16 58:{19,19}]
  wire [63:0] _GEN_646 = 6'h6 == io_writePorts_0_addr ? io_writePorts_0_data : mem_6; // @[Regfile.scala 51:16 58:{19,19}]
  wire [63:0] _GEN_647 = 6'h7 == io_writePorts_0_addr ? io_writePorts_0_data : mem_7; // @[Regfile.scala 51:16 58:{19,19}]
  wire [63:0] _GEN_648 = 6'h8 == io_writePorts_0_addr ? io_writePorts_0_data : mem_8; // @[Regfile.scala 51:16 58:{19,19}]
  wire [63:0] _GEN_649 = 6'h9 == io_writePorts_0_addr ? io_writePorts_0_data : mem_9; // @[Regfile.scala 51:16 58:{19,19}]
  wire [63:0] _GEN_650 = 6'ha == io_writePorts_0_addr ? io_writePorts_0_data : mem_10; // @[Regfile.scala 51:16 58:{19,19}]
  wire [63:0] _GEN_651 = 6'hb == io_writePorts_0_addr ? io_writePorts_0_data : mem_11; // @[Regfile.scala 51:16 58:{19,19}]
  wire [63:0] _GEN_652 = 6'hc == io_writePorts_0_addr ? io_writePorts_0_data : mem_12; // @[Regfile.scala 51:16 58:{19,19}]
  wire [63:0] _GEN_653 = 6'hd == io_writePorts_0_addr ? io_writePorts_0_data : mem_13; // @[Regfile.scala 51:16 58:{19,19}]
  wire [63:0] _GEN_654 = 6'he == io_writePorts_0_addr ? io_writePorts_0_data : mem_14; // @[Regfile.scala 51:16 58:{19,19}]
  wire [63:0] _GEN_655 = 6'hf == io_writePorts_0_addr ? io_writePorts_0_data : mem_15; // @[Regfile.scala 51:16 58:{19,19}]
  wire [63:0] _GEN_656 = 6'h10 == io_writePorts_0_addr ? io_writePorts_0_data : mem_16; // @[Regfile.scala 51:16 58:{19,19}]
  wire [63:0] _GEN_657 = 6'h11 == io_writePorts_0_addr ? io_writePorts_0_data : mem_17; // @[Regfile.scala 51:16 58:{19,19}]
  wire [63:0] _GEN_658 = 6'h12 == io_writePorts_0_addr ? io_writePorts_0_data : mem_18; // @[Regfile.scala 51:16 58:{19,19}]
  wire [63:0] _GEN_659 = 6'h13 == io_writePorts_0_addr ? io_writePorts_0_data : mem_19; // @[Regfile.scala 51:16 58:{19,19}]
  wire [63:0] _GEN_660 = 6'h14 == io_writePorts_0_addr ? io_writePorts_0_data : mem_20; // @[Regfile.scala 51:16 58:{19,19}]
  wire [63:0] _GEN_661 = 6'h15 == io_writePorts_0_addr ? io_writePorts_0_data : mem_21; // @[Regfile.scala 51:16 58:{19,19}]
  wire [63:0] _GEN_662 = 6'h16 == io_writePorts_0_addr ? io_writePorts_0_data : mem_22; // @[Regfile.scala 51:16 58:{19,19}]
  wire [63:0] _GEN_663 = 6'h17 == io_writePorts_0_addr ? io_writePorts_0_data : mem_23; // @[Regfile.scala 51:16 58:{19,19}]
  wire [63:0] _GEN_664 = 6'h18 == io_writePorts_0_addr ? io_writePorts_0_data : mem_24; // @[Regfile.scala 51:16 58:{19,19}]
  wire [63:0] _GEN_665 = 6'h19 == io_writePorts_0_addr ? io_writePorts_0_data : mem_25; // @[Regfile.scala 51:16 58:{19,19}]
  wire [63:0] _GEN_666 = 6'h1a == io_writePorts_0_addr ? io_writePorts_0_data : mem_26; // @[Regfile.scala 51:16 58:{19,19}]
  wire [63:0] _GEN_667 = 6'h1b == io_writePorts_0_addr ? io_writePorts_0_data : mem_27; // @[Regfile.scala 51:16 58:{19,19}]
  wire [63:0] _GEN_668 = 6'h1c == io_writePorts_0_addr ? io_writePorts_0_data : mem_28; // @[Regfile.scala 51:16 58:{19,19}]
  wire [63:0] _GEN_669 = 6'h1d == io_writePorts_0_addr ? io_writePorts_0_data : mem_29; // @[Regfile.scala 51:16 58:{19,19}]
  wire [63:0] _GEN_670 = 6'h1e == io_writePorts_0_addr ? io_writePorts_0_data : mem_30; // @[Regfile.scala 51:16 58:{19,19}]
  wire [63:0] _GEN_671 = 6'h1f == io_writePorts_0_addr ? io_writePorts_0_data : mem_31; // @[Regfile.scala 51:16 58:{19,19}]
  wire [63:0] _GEN_672 = 6'h20 == io_writePorts_0_addr ? io_writePorts_0_data : mem_32; // @[Regfile.scala 51:16 58:{19,19}]
  wire [63:0] _GEN_673 = 6'h21 == io_writePorts_0_addr ? io_writePorts_0_data : mem_33; // @[Regfile.scala 51:16 58:{19,19}]
  wire [63:0] _GEN_674 = 6'h22 == io_writePorts_0_addr ? io_writePorts_0_data : mem_34; // @[Regfile.scala 51:16 58:{19,19}]
  wire [63:0] _GEN_675 = 6'h23 == io_writePorts_0_addr ? io_writePorts_0_data : mem_35; // @[Regfile.scala 51:16 58:{19,19}]
  wire [63:0] _GEN_676 = 6'h24 == io_writePorts_0_addr ? io_writePorts_0_data : mem_36; // @[Regfile.scala 51:16 58:{19,19}]
  wire [63:0] _GEN_677 = 6'h25 == io_writePorts_0_addr ? io_writePorts_0_data : mem_37; // @[Regfile.scala 51:16 58:{19,19}]
  wire [63:0] _GEN_678 = 6'h26 == io_writePorts_0_addr ? io_writePorts_0_data : mem_38; // @[Regfile.scala 51:16 58:{19,19}]
  wire [63:0] _GEN_679 = 6'h27 == io_writePorts_0_addr ? io_writePorts_0_data : mem_39; // @[Regfile.scala 51:16 58:{19,19}]
  wire [63:0] _GEN_680 = 6'h28 == io_writePorts_0_addr ? io_writePorts_0_data : mem_40; // @[Regfile.scala 51:16 58:{19,19}]
  wire [63:0] _GEN_681 = 6'h29 == io_writePorts_0_addr ? io_writePorts_0_data : mem_41; // @[Regfile.scala 51:16 58:{19,19}]
  wire [63:0] _GEN_682 = 6'h2a == io_writePorts_0_addr ? io_writePorts_0_data : mem_42; // @[Regfile.scala 51:16 58:{19,19}]
  wire [63:0] _GEN_683 = 6'h2b == io_writePorts_0_addr ? io_writePorts_0_data : mem_43; // @[Regfile.scala 51:16 58:{19,19}]
  wire [63:0] _GEN_684 = 6'h2c == io_writePorts_0_addr ? io_writePorts_0_data : mem_44; // @[Regfile.scala 51:16 58:{19,19}]
  wire [63:0] _GEN_685 = 6'h2d == io_writePorts_0_addr ? io_writePorts_0_data : mem_45; // @[Regfile.scala 51:16 58:{19,19}]
  wire [63:0] _GEN_686 = 6'h2e == io_writePorts_0_addr ? io_writePorts_0_data : mem_46; // @[Regfile.scala 51:16 58:{19,19}]
  wire [63:0] _GEN_687 = 6'h2f == io_writePorts_0_addr ? io_writePorts_0_data : mem_47; // @[Regfile.scala 51:16 58:{19,19}]
  wire [63:0] _GEN_688 = 6'h30 == io_writePorts_0_addr ? io_writePorts_0_data : mem_48; // @[Regfile.scala 51:16 58:{19,19}]
  wire [63:0] _GEN_689 = 6'h31 == io_writePorts_0_addr ? io_writePorts_0_data : mem_49; // @[Regfile.scala 51:16 58:{19,19}]
  wire [63:0] _GEN_690 = 6'h32 == io_writePorts_0_addr ? io_writePorts_0_data : mem_50; // @[Regfile.scala 51:16 58:{19,19}]
  wire [63:0] _GEN_691 = 6'h33 == io_writePorts_0_addr ? io_writePorts_0_data : mem_51; // @[Regfile.scala 51:16 58:{19,19}]
  wire [63:0] _GEN_692 = 6'h34 == io_writePorts_0_addr ? io_writePorts_0_data : mem_52; // @[Regfile.scala 51:16 58:{19,19}]
  wire [63:0] _GEN_693 = 6'h35 == io_writePorts_0_addr ? io_writePorts_0_data : mem_53; // @[Regfile.scala 51:16 58:{19,19}]
  wire [63:0] _GEN_694 = 6'h36 == io_writePorts_0_addr ? io_writePorts_0_data : mem_54; // @[Regfile.scala 51:16 58:{19,19}]
  wire [63:0] _GEN_695 = 6'h37 == io_writePorts_0_addr ? io_writePorts_0_data : mem_55; // @[Regfile.scala 51:16 58:{19,19}]
  wire [63:0] _GEN_696 = 6'h38 == io_writePorts_0_addr ? io_writePorts_0_data : mem_56; // @[Regfile.scala 51:16 58:{19,19}]
  wire [63:0] _GEN_697 = 6'h39 == io_writePorts_0_addr ? io_writePorts_0_data : mem_57; // @[Regfile.scala 51:16 58:{19,19}]
  wire [63:0] _GEN_698 = 6'h3a == io_writePorts_0_addr ? io_writePorts_0_data : mem_58; // @[Regfile.scala 51:16 58:{19,19}]
  wire [63:0] _GEN_699 = 6'h3b == io_writePorts_0_addr ? io_writePorts_0_data : mem_59; // @[Regfile.scala 51:16 58:{19,19}]
  wire [63:0] _GEN_700 = 6'h3c == io_writePorts_0_addr ? io_writePorts_0_data : mem_60; // @[Regfile.scala 51:16 58:{19,19}]
  wire [63:0] _GEN_701 = 6'h3d == io_writePorts_0_addr ? io_writePorts_0_data : mem_61; // @[Regfile.scala 51:16 58:{19,19}]
  wire [63:0] _GEN_702 = 6'h3e == io_writePorts_0_addr ? io_writePorts_0_data : mem_62; // @[Regfile.scala 51:16 58:{19,19}]
  wire [63:0] _GEN_703 = 6'h3f == io_writePorts_0_addr ? io_writePorts_0_data : mem_63; // @[Regfile.scala 51:16 58:{19,19}]
  wire [63:0] _GEN_704 = io_writePorts_0_wen ? _GEN_640 : mem_0; // @[Regfile.scala 51:16 57:17]
  wire [63:0] _GEN_705 = io_writePorts_0_wen ? _GEN_641 : mem_1; // @[Regfile.scala 51:16 57:17]
  wire [63:0] _GEN_706 = io_writePorts_0_wen ? _GEN_642 : mem_2; // @[Regfile.scala 51:16 57:17]
  wire [63:0] _GEN_707 = io_writePorts_0_wen ? _GEN_643 : mem_3; // @[Regfile.scala 51:16 57:17]
  wire [63:0] _GEN_708 = io_writePorts_0_wen ? _GEN_644 : mem_4; // @[Regfile.scala 51:16 57:17]
  wire [63:0] _GEN_709 = io_writePorts_0_wen ? _GEN_645 : mem_5; // @[Regfile.scala 51:16 57:17]
  wire [63:0] _GEN_710 = io_writePorts_0_wen ? _GEN_646 : mem_6; // @[Regfile.scala 51:16 57:17]
  wire [63:0] _GEN_711 = io_writePorts_0_wen ? _GEN_647 : mem_7; // @[Regfile.scala 51:16 57:17]
  wire [63:0] _GEN_712 = io_writePorts_0_wen ? _GEN_648 : mem_8; // @[Regfile.scala 51:16 57:17]
  wire [63:0] _GEN_713 = io_writePorts_0_wen ? _GEN_649 : mem_9; // @[Regfile.scala 51:16 57:17]
  wire [63:0] _GEN_714 = io_writePorts_0_wen ? _GEN_650 : mem_10; // @[Regfile.scala 51:16 57:17]
  wire [63:0] _GEN_715 = io_writePorts_0_wen ? _GEN_651 : mem_11; // @[Regfile.scala 51:16 57:17]
  wire [63:0] _GEN_716 = io_writePorts_0_wen ? _GEN_652 : mem_12; // @[Regfile.scala 51:16 57:17]
  wire [63:0] _GEN_717 = io_writePorts_0_wen ? _GEN_653 : mem_13; // @[Regfile.scala 51:16 57:17]
  wire [63:0] _GEN_718 = io_writePorts_0_wen ? _GEN_654 : mem_14; // @[Regfile.scala 51:16 57:17]
  wire [63:0] _GEN_719 = io_writePorts_0_wen ? _GEN_655 : mem_15; // @[Regfile.scala 51:16 57:17]
  wire [63:0] _GEN_720 = io_writePorts_0_wen ? _GEN_656 : mem_16; // @[Regfile.scala 51:16 57:17]
  wire [63:0] _GEN_721 = io_writePorts_0_wen ? _GEN_657 : mem_17; // @[Regfile.scala 51:16 57:17]
  wire [63:0] _GEN_722 = io_writePorts_0_wen ? _GEN_658 : mem_18; // @[Regfile.scala 51:16 57:17]
  wire [63:0] _GEN_723 = io_writePorts_0_wen ? _GEN_659 : mem_19; // @[Regfile.scala 51:16 57:17]
  wire [63:0] _GEN_724 = io_writePorts_0_wen ? _GEN_660 : mem_20; // @[Regfile.scala 51:16 57:17]
  wire [63:0] _GEN_725 = io_writePorts_0_wen ? _GEN_661 : mem_21; // @[Regfile.scala 51:16 57:17]
  wire [63:0] _GEN_726 = io_writePorts_0_wen ? _GEN_662 : mem_22; // @[Regfile.scala 51:16 57:17]
  wire [63:0] _GEN_727 = io_writePorts_0_wen ? _GEN_663 : mem_23; // @[Regfile.scala 51:16 57:17]
  wire [63:0] _GEN_728 = io_writePorts_0_wen ? _GEN_664 : mem_24; // @[Regfile.scala 51:16 57:17]
  wire [63:0] _GEN_729 = io_writePorts_0_wen ? _GEN_665 : mem_25; // @[Regfile.scala 51:16 57:17]
  wire [63:0] _GEN_730 = io_writePorts_0_wen ? _GEN_666 : mem_26; // @[Regfile.scala 51:16 57:17]
  wire [63:0] _GEN_731 = io_writePorts_0_wen ? _GEN_667 : mem_27; // @[Regfile.scala 51:16 57:17]
  wire [63:0] _GEN_732 = io_writePorts_0_wen ? _GEN_668 : mem_28; // @[Regfile.scala 51:16 57:17]
  wire [63:0] _GEN_733 = io_writePorts_0_wen ? _GEN_669 : mem_29; // @[Regfile.scala 51:16 57:17]
  wire [63:0] _GEN_734 = io_writePorts_0_wen ? _GEN_670 : mem_30; // @[Regfile.scala 51:16 57:17]
  wire [63:0] _GEN_735 = io_writePorts_0_wen ? _GEN_671 : mem_31; // @[Regfile.scala 51:16 57:17]
  wire [63:0] _GEN_736 = io_writePorts_0_wen ? _GEN_672 : mem_32; // @[Regfile.scala 51:16 57:17]
  wire [63:0] _GEN_737 = io_writePorts_0_wen ? _GEN_673 : mem_33; // @[Regfile.scala 51:16 57:17]
  wire [63:0] _GEN_738 = io_writePorts_0_wen ? _GEN_674 : mem_34; // @[Regfile.scala 51:16 57:17]
  wire [63:0] _GEN_739 = io_writePorts_0_wen ? _GEN_675 : mem_35; // @[Regfile.scala 51:16 57:17]
  wire [63:0] _GEN_740 = io_writePorts_0_wen ? _GEN_676 : mem_36; // @[Regfile.scala 51:16 57:17]
  wire [63:0] _GEN_741 = io_writePorts_0_wen ? _GEN_677 : mem_37; // @[Regfile.scala 51:16 57:17]
  wire [63:0] _GEN_742 = io_writePorts_0_wen ? _GEN_678 : mem_38; // @[Regfile.scala 51:16 57:17]
  wire [63:0] _GEN_743 = io_writePorts_0_wen ? _GEN_679 : mem_39; // @[Regfile.scala 51:16 57:17]
  wire [63:0] _GEN_744 = io_writePorts_0_wen ? _GEN_680 : mem_40; // @[Regfile.scala 51:16 57:17]
  wire [63:0] _GEN_745 = io_writePorts_0_wen ? _GEN_681 : mem_41; // @[Regfile.scala 51:16 57:17]
  wire [63:0] _GEN_746 = io_writePorts_0_wen ? _GEN_682 : mem_42; // @[Regfile.scala 51:16 57:17]
  wire [63:0] _GEN_747 = io_writePorts_0_wen ? _GEN_683 : mem_43; // @[Regfile.scala 51:16 57:17]
  wire [63:0] _GEN_748 = io_writePorts_0_wen ? _GEN_684 : mem_44; // @[Regfile.scala 51:16 57:17]
  wire [63:0] _GEN_749 = io_writePorts_0_wen ? _GEN_685 : mem_45; // @[Regfile.scala 51:16 57:17]
  wire [63:0] _GEN_750 = io_writePorts_0_wen ? _GEN_686 : mem_46; // @[Regfile.scala 51:16 57:17]
  wire [63:0] _GEN_751 = io_writePorts_0_wen ? _GEN_687 : mem_47; // @[Regfile.scala 51:16 57:17]
  wire [63:0] _GEN_752 = io_writePorts_0_wen ? _GEN_688 : mem_48; // @[Regfile.scala 51:16 57:17]
  wire [63:0] _GEN_753 = io_writePorts_0_wen ? _GEN_689 : mem_49; // @[Regfile.scala 51:16 57:17]
  wire [63:0] _GEN_754 = io_writePorts_0_wen ? _GEN_690 : mem_50; // @[Regfile.scala 51:16 57:17]
  wire [63:0] _GEN_755 = io_writePorts_0_wen ? _GEN_691 : mem_51; // @[Regfile.scala 51:16 57:17]
  wire [63:0] _GEN_756 = io_writePorts_0_wen ? _GEN_692 : mem_52; // @[Regfile.scala 51:16 57:17]
  wire [63:0] _GEN_757 = io_writePorts_0_wen ? _GEN_693 : mem_53; // @[Regfile.scala 51:16 57:17]
  wire [63:0] _GEN_758 = io_writePorts_0_wen ? _GEN_694 : mem_54; // @[Regfile.scala 51:16 57:17]
  wire [63:0] _GEN_759 = io_writePorts_0_wen ? _GEN_695 : mem_55; // @[Regfile.scala 51:16 57:17]
  wire [63:0] _GEN_760 = io_writePorts_0_wen ? _GEN_696 : mem_56; // @[Regfile.scala 51:16 57:17]
  wire [63:0] _GEN_761 = io_writePorts_0_wen ? _GEN_697 : mem_57; // @[Regfile.scala 51:16 57:17]
  wire [63:0] _GEN_762 = io_writePorts_0_wen ? _GEN_698 : mem_58; // @[Regfile.scala 51:16 57:17]
  wire [63:0] _GEN_763 = io_writePorts_0_wen ? _GEN_699 : mem_59; // @[Regfile.scala 51:16 57:17]
  wire [63:0] _GEN_764 = io_writePorts_0_wen ? _GEN_700 : mem_60; // @[Regfile.scala 51:16 57:17]
  wire [63:0] _GEN_765 = io_writePorts_0_wen ? _GEN_701 : mem_61; // @[Regfile.scala 51:16 57:17]
  wire [63:0] _GEN_766 = io_writePorts_0_wen ? _GEN_702 : mem_62; // @[Regfile.scala 51:16 57:17]
  wire [63:0] _GEN_767 = io_writePorts_0_wen ? _GEN_703 : mem_63; // @[Regfile.scala 51:16 57:17]
  wire [63:0] _GEN_768 = 6'h0 == io_writePorts_1_addr ? io_writePorts_1_data : _GEN_704; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_769 = 6'h1 == io_writePorts_1_addr ? io_writePorts_1_data : _GEN_705; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_770 = 6'h2 == io_writePorts_1_addr ? io_writePorts_1_data : _GEN_706; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_771 = 6'h3 == io_writePorts_1_addr ? io_writePorts_1_data : _GEN_707; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_772 = 6'h4 == io_writePorts_1_addr ? io_writePorts_1_data : _GEN_708; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_773 = 6'h5 == io_writePorts_1_addr ? io_writePorts_1_data : _GEN_709; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_774 = 6'h6 == io_writePorts_1_addr ? io_writePorts_1_data : _GEN_710; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_775 = 6'h7 == io_writePorts_1_addr ? io_writePorts_1_data : _GEN_711; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_776 = 6'h8 == io_writePorts_1_addr ? io_writePorts_1_data : _GEN_712; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_777 = 6'h9 == io_writePorts_1_addr ? io_writePorts_1_data : _GEN_713; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_778 = 6'ha == io_writePorts_1_addr ? io_writePorts_1_data : _GEN_714; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_779 = 6'hb == io_writePorts_1_addr ? io_writePorts_1_data : _GEN_715; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_780 = 6'hc == io_writePorts_1_addr ? io_writePorts_1_data : _GEN_716; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_781 = 6'hd == io_writePorts_1_addr ? io_writePorts_1_data : _GEN_717; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_782 = 6'he == io_writePorts_1_addr ? io_writePorts_1_data : _GEN_718; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_783 = 6'hf == io_writePorts_1_addr ? io_writePorts_1_data : _GEN_719; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_784 = 6'h10 == io_writePorts_1_addr ? io_writePorts_1_data : _GEN_720; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_785 = 6'h11 == io_writePorts_1_addr ? io_writePorts_1_data : _GEN_721; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_786 = 6'h12 == io_writePorts_1_addr ? io_writePorts_1_data : _GEN_722; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_787 = 6'h13 == io_writePorts_1_addr ? io_writePorts_1_data : _GEN_723; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_788 = 6'h14 == io_writePorts_1_addr ? io_writePorts_1_data : _GEN_724; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_789 = 6'h15 == io_writePorts_1_addr ? io_writePorts_1_data : _GEN_725; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_790 = 6'h16 == io_writePorts_1_addr ? io_writePorts_1_data : _GEN_726; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_791 = 6'h17 == io_writePorts_1_addr ? io_writePorts_1_data : _GEN_727; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_792 = 6'h18 == io_writePorts_1_addr ? io_writePorts_1_data : _GEN_728; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_793 = 6'h19 == io_writePorts_1_addr ? io_writePorts_1_data : _GEN_729; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_794 = 6'h1a == io_writePorts_1_addr ? io_writePorts_1_data : _GEN_730; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_795 = 6'h1b == io_writePorts_1_addr ? io_writePorts_1_data : _GEN_731; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_796 = 6'h1c == io_writePorts_1_addr ? io_writePorts_1_data : _GEN_732; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_797 = 6'h1d == io_writePorts_1_addr ? io_writePorts_1_data : _GEN_733; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_798 = 6'h1e == io_writePorts_1_addr ? io_writePorts_1_data : _GEN_734; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_799 = 6'h1f == io_writePorts_1_addr ? io_writePorts_1_data : _GEN_735; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_800 = 6'h20 == io_writePorts_1_addr ? io_writePorts_1_data : _GEN_736; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_801 = 6'h21 == io_writePorts_1_addr ? io_writePorts_1_data : _GEN_737; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_802 = 6'h22 == io_writePorts_1_addr ? io_writePorts_1_data : _GEN_738; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_803 = 6'h23 == io_writePorts_1_addr ? io_writePorts_1_data : _GEN_739; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_804 = 6'h24 == io_writePorts_1_addr ? io_writePorts_1_data : _GEN_740; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_805 = 6'h25 == io_writePorts_1_addr ? io_writePorts_1_data : _GEN_741; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_806 = 6'h26 == io_writePorts_1_addr ? io_writePorts_1_data : _GEN_742; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_807 = 6'h27 == io_writePorts_1_addr ? io_writePorts_1_data : _GEN_743; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_808 = 6'h28 == io_writePorts_1_addr ? io_writePorts_1_data : _GEN_744; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_809 = 6'h29 == io_writePorts_1_addr ? io_writePorts_1_data : _GEN_745; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_810 = 6'h2a == io_writePorts_1_addr ? io_writePorts_1_data : _GEN_746; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_811 = 6'h2b == io_writePorts_1_addr ? io_writePorts_1_data : _GEN_747; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_812 = 6'h2c == io_writePorts_1_addr ? io_writePorts_1_data : _GEN_748; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_813 = 6'h2d == io_writePorts_1_addr ? io_writePorts_1_data : _GEN_749; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_814 = 6'h2e == io_writePorts_1_addr ? io_writePorts_1_data : _GEN_750; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_815 = 6'h2f == io_writePorts_1_addr ? io_writePorts_1_data : _GEN_751; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_816 = 6'h30 == io_writePorts_1_addr ? io_writePorts_1_data : _GEN_752; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_817 = 6'h31 == io_writePorts_1_addr ? io_writePorts_1_data : _GEN_753; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_818 = 6'h32 == io_writePorts_1_addr ? io_writePorts_1_data : _GEN_754; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_819 = 6'h33 == io_writePorts_1_addr ? io_writePorts_1_data : _GEN_755; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_820 = 6'h34 == io_writePorts_1_addr ? io_writePorts_1_data : _GEN_756; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_821 = 6'h35 == io_writePorts_1_addr ? io_writePorts_1_data : _GEN_757; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_822 = 6'h36 == io_writePorts_1_addr ? io_writePorts_1_data : _GEN_758; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_823 = 6'h37 == io_writePorts_1_addr ? io_writePorts_1_data : _GEN_759; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_824 = 6'h38 == io_writePorts_1_addr ? io_writePorts_1_data : _GEN_760; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_825 = 6'h39 == io_writePorts_1_addr ? io_writePorts_1_data : _GEN_761; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_826 = 6'h3a == io_writePorts_1_addr ? io_writePorts_1_data : _GEN_762; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_827 = 6'h3b == io_writePorts_1_addr ? io_writePorts_1_data : _GEN_763; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_828 = 6'h3c == io_writePorts_1_addr ? io_writePorts_1_data : _GEN_764; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_829 = 6'h3d == io_writePorts_1_addr ? io_writePorts_1_data : _GEN_765; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_830 = 6'h3e == io_writePorts_1_addr ? io_writePorts_1_data : _GEN_766; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_831 = 6'h3f == io_writePorts_1_addr ? io_writePorts_1_data : _GEN_767; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_832 = io_writePorts_1_wen ? _GEN_768 : _GEN_704; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_833 = io_writePorts_1_wen ? _GEN_769 : _GEN_705; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_834 = io_writePorts_1_wen ? _GEN_770 : _GEN_706; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_835 = io_writePorts_1_wen ? _GEN_771 : _GEN_707; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_836 = io_writePorts_1_wen ? _GEN_772 : _GEN_708; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_837 = io_writePorts_1_wen ? _GEN_773 : _GEN_709; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_838 = io_writePorts_1_wen ? _GEN_774 : _GEN_710; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_839 = io_writePorts_1_wen ? _GEN_775 : _GEN_711; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_840 = io_writePorts_1_wen ? _GEN_776 : _GEN_712; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_841 = io_writePorts_1_wen ? _GEN_777 : _GEN_713; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_842 = io_writePorts_1_wen ? _GEN_778 : _GEN_714; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_843 = io_writePorts_1_wen ? _GEN_779 : _GEN_715; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_844 = io_writePorts_1_wen ? _GEN_780 : _GEN_716; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_845 = io_writePorts_1_wen ? _GEN_781 : _GEN_717; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_846 = io_writePorts_1_wen ? _GEN_782 : _GEN_718; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_847 = io_writePorts_1_wen ? _GEN_783 : _GEN_719; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_848 = io_writePorts_1_wen ? _GEN_784 : _GEN_720; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_849 = io_writePorts_1_wen ? _GEN_785 : _GEN_721; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_850 = io_writePorts_1_wen ? _GEN_786 : _GEN_722; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_851 = io_writePorts_1_wen ? _GEN_787 : _GEN_723; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_852 = io_writePorts_1_wen ? _GEN_788 : _GEN_724; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_853 = io_writePorts_1_wen ? _GEN_789 : _GEN_725; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_854 = io_writePorts_1_wen ? _GEN_790 : _GEN_726; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_855 = io_writePorts_1_wen ? _GEN_791 : _GEN_727; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_856 = io_writePorts_1_wen ? _GEN_792 : _GEN_728; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_857 = io_writePorts_1_wen ? _GEN_793 : _GEN_729; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_858 = io_writePorts_1_wen ? _GEN_794 : _GEN_730; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_859 = io_writePorts_1_wen ? _GEN_795 : _GEN_731; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_860 = io_writePorts_1_wen ? _GEN_796 : _GEN_732; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_861 = io_writePorts_1_wen ? _GEN_797 : _GEN_733; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_862 = io_writePorts_1_wen ? _GEN_798 : _GEN_734; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_863 = io_writePorts_1_wen ? _GEN_799 : _GEN_735; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_864 = io_writePorts_1_wen ? _GEN_800 : _GEN_736; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_865 = io_writePorts_1_wen ? _GEN_801 : _GEN_737; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_866 = io_writePorts_1_wen ? _GEN_802 : _GEN_738; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_867 = io_writePorts_1_wen ? _GEN_803 : _GEN_739; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_868 = io_writePorts_1_wen ? _GEN_804 : _GEN_740; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_869 = io_writePorts_1_wen ? _GEN_805 : _GEN_741; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_870 = io_writePorts_1_wen ? _GEN_806 : _GEN_742; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_871 = io_writePorts_1_wen ? _GEN_807 : _GEN_743; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_872 = io_writePorts_1_wen ? _GEN_808 : _GEN_744; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_873 = io_writePorts_1_wen ? _GEN_809 : _GEN_745; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_874 = io_writePorts_1_wen ? _GEN_810 : _GEN_746; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_875 = io_writePorts_1_wen ? _GEN_811 : _GEN_747; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_876 = io_writePorts_1_wen ? _GEN_812 : _GEN_748; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_877 = io_writePorts_1_wen ? _GEN_813 : _GEN_749; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_878 = io_writePorts_1_wen ? _GEN_814 : _GEN_750; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_879 = io_writePorts_1_wen ? _GEN_815 : _GEN_751; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_880 = io_writePorts_1_wen ? _GEN_816 : _GEN_752; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_881 = io_writePorts_1_wen ? _GEN_817 : _GEN_753; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_882 = io_writePorts_1_wen ? _GEN_818 : _GEN_754; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_883 = io_writePorts_1_wen ? _GEN_819 : _GEN_755; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_884 = io_writePorts_1_wen ? _GEN_820 : _GEN_756; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_885 = io_writePorts_1_wen ? _GEN_821 : _GEN_757; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_886 = io_writePorts_1_wen ? _GEN_822 : _GEN_758; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_887 = io_writePorts_1_wen ? _GEN_823 : _GEN_759; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_888 = io_writePorts_1_wen ? _GEN_824 : _GEN_760; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_889 = io_writePorts_1_wen ? _GEN_825 : _GEN_761; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_890 = io_writePorts_1_wen ? _GEN_826 : _GEN_762; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_891 = io_writePorts_1_wen ? _GEN_827 : _GEN_763; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_892 = io_writePorts_1_wen ? _GEN_828 : _GEN_764; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_893 = io_writePorts_1_wen ? _GEN_829 : _GEN_765; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_894 = io_writePorts_1_wen ? _GEN_830 : _GEN_766; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_895 = io_writePorts_1_wen ? _GEN_831 : _GEN_767; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_896 = 6'h0 == io_writePorts_2_addr ? io_writePorts_2_data : _GEN_832; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_897 = 6'h1 == io_writePorts_2_addr ? io_writePorts_2_data : _GEN_833; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_898 = 6'h2 == io_writePorts_2_addr ? io_writePorts_2_data : _GEN_834; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_899 = 6'h3 == io_writePorts_2_addr ? io_writePorts_2_data : _GEN_835; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_900 = 6'h4 == io_writePorts_2_addr ? io_writePorts_2_data : _GEN_836; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_901 = 6'h5 == io_writePorts_2_addr ? io_writePorts_2_data : _GEN_837; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_902 = 6'h6 == io_writePorts_2_addr ? io_writePorts_2_data : _GEN_838; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_903 = 6'h7 == io_writePorts_2_addr ? io_writePorts_2_data : _GEN_839; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_904 = 6'h8 == io_writePorts_2_addr ? io_writePorts_2_data : _GEN_840; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_905 = 6'h9 == io_writePorts_2_addr ? io_writePorts_2_data : _GEN_841; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_906 = 6'ha == io_writePorts_2_addr ? io_writePorts_2_data : _GEN_842; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_907 = 6'hb == io_writePorts_2_addr ? io_writePorts_2_data : _GEN_843; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_908 = 6'hc == io_writePorts_2_addr ? io_writePorts_2_data : _GEN_844; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_909 = 6'hd == io_writePorts_2_addr ? io_writePorts_2_data : _GEN_845; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_910 = 6'he == io_writePorts_2_addr ? io_writePorts_2_data : _GEN_846; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_911 = 6'hf == io_writePorts_2_addr ? io_writePorts_2_data : _GEN_847; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_912 = 6'h10 == io_writePorts_2_addr ? io_writePorts_2_data : _GEN_848; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_913 = 6'h11 == io_writePorts_2_addr ? io_writePorts_2_data : _GEN_849; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_914 = 6'h12 == io_writePorts_2_addr ? io_writePorts_2_data : _GEN_850; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_915 = 6'h13 == io_writePorts_2_addr ? io_writePorts_2_data : _GEN_851; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_916 = 6'h14 == io_writePorts_2_addr ? io_writePorts_2_data : _GEN_852; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_917 = 6'h15 == io_writePorts_2_addr ? io_writePorts_2_data : _GEN_853; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_918 = 6'h16 == io_writePorts_2_addr ? io_writePorts_2_data : _GEN_854; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_919 = 6'h17 == io_writePorts_2_addr ? io_writePorts_2_data : _GEN_855; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_920 = 6'h18 == io_writePorts_2_addr ? io_writePorts_2_data : _GEN_856; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_921 = 6'h19 == io_writePorts_2_addr ? io_writePorts_2_data : _GEN_857; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_922 = 6'h1a == io_writePorts_2_addr ? io_writePorts_2_data : _GEN_858; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_923 = 6'h1b == io_writePorts_2_addr ? io_writePorts_2_data : _GEN_859; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_924 = 6'h1c == io_writePorts_2_addr ? io_writePorts_2_data : _GEN_860; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_925 = 6'h1d == io_writePorts_2_addr ? io_writePorts_2_data : _GEN_861; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_926 = 6'h1e == io_writePorts_2_addr ? io_writePorts_2_data : _GEN_862; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_927 = 6'h1f == io_writePorts_2_addr ? io_writePorts_2_data : _GEN_863; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_928 = 6'h20 == io_writePorts_2_addr ? io_writePorts_2_data : _GEN_864; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_929 = 6'h21 == io_writePorts_2_addr ? io_writePorts_2_data : _GEN_865; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_930 = 6'h22 == io_writePorts_2_addr ? io_writePorts_2_data : _GEN_866; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_931 = 6'h23 == io_writePorts_2_addr ? io_writePorts_2_data : _GEN_867; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_932 = 6'h24 == io_writePorts_2_addr ? io_writePorts_2_data : _GEN_868; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_933 = 6'h25 == io_writePorts_2_addr ? io_writePorts_2_data : _GEN_869; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_934 = 6'h26 == io_writePorts_2_addr ? io_writePorts_2_data : _GEN_870; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_935 = 6'h27 == io_writePorts_2_addr ? io_writePorts_2_data : _GEN_871; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_936 = 6'h28 == io_writePorts_2_addr ? io_writePorts_2_data : _GEN_872; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_937 = 6'h29 == io_writePorts_2_addr ? io_writePorts_2_data : _GEN_873; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_938 = 6'h2a == io_writePorts_2_addr ? io_writePorts_2_data : _GEN_874; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_939 = 6'h2b == io_writePorts_2_addr ? io_writePorts_2_data : _GEN_875; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_940 = 6'h2c == io_writePorts_2_addr ? io_writePorts_2_data : _GEN_876; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_941 = 6'h2d == io_writePorts_2_addr ? io_writePorts_2_data : _GEN_877; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_942 = 6'h2e == io_writePorts_2_addr ? io_writePorts_2_data : _GEN_878; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_943 = 6'h2f == io_writePorts_2_addr ? io_writePorts_2_data : _GEN_879; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_944 = 6'h30 == io_writePorts_2_addr ? io_writePorts_2_data : _GEN_880; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_945 = 6'h31 == io_writePorts_2_addr ? io_writePorts_2_data : _GEN_881; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_946 = 6'h32 == io_writePorts_2_addr ? io_writePorts_2_data : _GEN_882; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_947 = 6'h33 == io_writePorts_2_addr ? io_writePorts_2_data : _GEN_883; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_948 = 6'h34 == io_writePorts_2_addr ? io_writePorts_2_data : _GEN_884; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_949 = 6'h35 == io_writePorts_2_addr ? io_writePorts_2_data : _GEN_885; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_950 = 6'h36 == io_writePorts_2_addr ? io_writePorts_2_data : _GEN_886; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_951 = 6'h37 == io_writePorts_2_addr ? io_writePorts_2_data : _GEN_887; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_952 = 6'h38 == io_writePorts_2_addr ? io_writePorts_2_data : _GEN_888; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_953 = 6'h39 == io_writePorts_2_addr ? io_writePorts_2_data : _GEN_889; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_954 = 6'h3a == io_writePorts_2_addr ? io_writePorts_2_data : _GEN_890; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_955 = 6'h3b == io_writePorts_2_addr ? io_writePorts_2_data : _GEN_891; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_956 = 6'h3c == io_writePorts_2_addr ? io_writePorts_2_data : _GEN_892; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_957 = 6'h3d == io_writePorts_2_addr ? io_writePorts_2_data : _GEN_893; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_958 = 6'h3e == io_writePorts_2_addr ? io_writePorts_2_data : _GEN_894; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_959 = 6'h3f == io_writePorts_2_addr ? io_writePorts_2_data : _GEN_895; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_960 = io_writePorts_2_wen ? _GEN_896 : _GEN_832; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_961 = io_writePorts_2_wen ? _GEN_897 : _GEN_833; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_962 = io_writePorts_2_wen ? _GEN_898 : _GEN_834; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_963 = io_writePorts_2_wen ? _GEN_899 : _GEN_835; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_964 = io_writePorts_2_wen ? _GEN_900 : _GEN_836; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_965 = io_writePorts_2_wen ? _GEN_901 : _GEN_837; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_966 = io_writePorts_2_wen ? _GEN_902 : _GEN_838; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_967 = io_writePorts_2_wen ? _GEN_903 : _GEN_839; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_968 = io_writePorts_2_wen ? _GEN_904 : _GEN_840; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_969 = io_writePorts_2_wen ? _GEN_905 : _GEN_841; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_970 = io_writePorts_2_wen ? _GEN_906 : _GEN_842; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_971 = io_writePorts_2_wen ? _GEN_907 : _GEN_843; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_972 = io_writePorts_2_wen ? _GEN_908 : _GEN_844; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_973 = io_writePorts_2_wen ? _GEN_909 : _GEN_845; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_974 = io_writePorts_2_wen ? _GEN_910 : _GEN_846; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_975 = io_writePorts_2_wen ? _GEN_911 : _GEN_847; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_976 = io_writePorts_2_wen ? _GEN_912 : _GEN_848; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_977 = io_writePorts_2_wen ? _GEN_913 : _GEN_849; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_978 = io_writePorts_2_wen ? _GEN_914 : _GEN_850; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_979 = io_writePorts_2_wen ? _GEN_915 : _GEN_851; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_980 = io_writePorts_2_wen ? _GEN_916 : _GEN_852; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_981 = io_writePorts_2_wen ? _GEN_917 : _GEN_853; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_982 = io_writePorts_2_wen ? _GEN_918 : _GEN_854; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_983 = io_writePorts_2_wen ? _GEN_919 : _GEN_855; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_984 = io_writePorts_2_wen ? _GEN_920 : _GEN_856; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_985 = io_writePorts_2_wen ? _GEN_921 : _GEN_857; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_986 = io_writePorts_2_wen ? _GEN_922 : _GEN_858; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_987 = io_writePorts_2_wen ? _GEN_923 : _GEN_859; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_988 = io_writePorts_2_wen ? _GEN_924 : _GEN_860; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_989 = io_writePorts_2_wen ? _GEN_925 : _GEN_861; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_990 = io_writePorts_2_wen ? _GEN_926 : _GEN_862; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_991 = io_writePorts_2_wen ? _GEN_927 : _GEN_863; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_992 = io_writePorts_2_wen ? _GEN_928 : _GEN_864; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_993 = io_writePorts_2_wen ? _GEN_929 : _GEN_865; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_994 = io_writePorts_2_wen ? _GEN_930 : _GEN_866; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_995 = io_writePorts_2_wen ? _GEN_931 : _GEN_867; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_996 = io_writePorts_2_wen ? _GEN_932 : _GEN_868; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_997 = io_writePorts_2_wen ? _GEN_933 : _GEN_869; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_998 = io_writePorts_2_wen ? _GEN_934 : _GEN_870; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_999 = io_writePorts_2_wen ? _GEN_935 : _GEN_871; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1000 = io_writePorts_2_wen ? _GEN_936 : _GEN_872; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1001 = io_writePorts_2_wen ? _GEN_937 : _GEN_873; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1002 = io_writePorts_2_wen ? _GEN_938 : _GEN_874; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1003 = io_writePorts_2_wen ? _GEN_939 : _GEN_875; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1004 = io_writePorts_2_wen ? _GEN_940 : _GEN_876; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1005 = io_writePorts_2_wen ? _GEN_941 : _GEN_877; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1006 = io_writePorts_2_wen ? _GEN_942 : _GEN_878; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1007 = io_writePorts_2_wen ? _GEN_943 : _GEN_879; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1008 = io_writePorts_2_wen ? _GEN_944 : _GEN_880; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1009 = io_writePorts_2_wen ? _GEN_945 : _GEN_881; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1010 = io_writePorts_2_wen ? _GEN_946 : _GEN_882; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1011 = io_writePorts_2_wen ? _GEN_947 : _GEN_883; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1012 = io_writePorts_2_wen ? _GEN_948 : _GEN_884; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1013 = io_writePorts_2_wen ? _GEN_949 : _GEN_885; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1014 = io_writePorts_2_wen ? _GEN_950 : _GEN_886; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1015 = io_writePorts_2_wen ? _GEN_951 : _GEN_887; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1016 = io_writePorts_2_wen ? _GEN_952 : _GEN_888; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1017 = io_writePorts_2_wen ? _GEN_953 : _GEN_889; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1018 = io_writePorts_2_wen ? _GEN_954 : _GEN_890; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1019 = io_writePorts_2_wen ? _GEN_955 : _GEN_891; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1020 = io_writePorts_2_wen ? _GEN_956 : _GEN_892; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1021 = io_writePorts_2_wen ? _GEN_957 : _GEN_893; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1022 = io_writePorts_2_wen ? _GEN_958 : _GEN_894; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1023 = io_writePorts_2_wen ? _GEN_959 : _GEN_895; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1024 = 6'h0 == io_writePorts_3_addr ? io_writePorts_3_data : _GEN_960; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_1025 = 6'h1 == io_writePorts_3_addr ? io_writePorts_3_data : _GEN_961; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_1026 = 6'h2 == io_writePorts_3_addr ? io_writePorts_3_data : _GEN_962; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_1027 = 6'h3 == io_writePorts_3_addr ? io_writePorts_3_data : _GEN_963; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_1028 = 6'h4 == io_writePorts_3_addr ? io_writePorts_3_data : _GEN_964; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_1029 = 6'h5 == io_writePorts_3_addr ? io_writePorts_3_data : _GEN_965; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_1030 = 6'h6 == io_writePorts_3_addr ? io_writePorts_3_data : _GEN_966; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_1031 = 6'h7 == io_writePorts_3_addr ? io_writePorts_3_data : _GEN_967; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_1032 = 6'h8 == io_writePorts_3_addr ? io_writePorts_3_data : _GEN_968; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_1033 = 6'h9 == io_writePorts_3_addr ? io_writePorts_3_data : _GEN_969; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_1034 = 6'ha == io_writePorts_3_addr ? io_writePorts_3_data : _GEN_970; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_1035 = 6'hb == io_writePorts_3_addr ? io_writePorts_3_data : _GEN_971; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_1036 = 6'hc == io_writePorts_3_addr ? io_writePorts_3_data : _GEN_972; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_1037 = 6'hd == io_writePorts_3_addr ? io_writePorts_3_data : _GEN_973; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_1038 = 6'he == io_writePorts_3_addr ? io_writePorts_3_data : _GEN_974; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_1039 = 6'hf == io_writePorts_3_addr ? io_writePorts_3_data : _GEN_975; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_1040 = 6'h10 == io_writePorts_3_addr ? io_writePorts_3_data : _GEN_976; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_1041 = 6'h11 == io_writePorts_3_addr ? io_writePorts_3_data : _GEN_977; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_1042 = 6'h12 == io_writePorts_3_addr ? io_writePorts_3_data : _GEN_978; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_1043 = 6'h13 == io_writePorts_3_addr ? io_writePorts_3_data : _GEN_979; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_1044 = 6'h14 == io_writePorts_3_addr ? io_writePorts_3_data : _GEN_980; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_1045 = 6'h15 == io_writePorts_3_addr ? io_writePorts_3_data : _GEN_981; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_1046 = 6'h16 == io_writePorts_3_addr ? io_writePorts_3_data : _GEN_982; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_1047 = 6'h17 == io_writePorts_3_addr ? io_writePorts_3_data : _GEN_983; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_1048 = 6'h18 == io_writePorts_3_addr ? io_writePorts_3_data : _GEN_984; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_1049 = 6'h19 == io_writePorts_3_addr ? io_writePorts_3_data : _GEN_985; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_1050 = 6'h1a == io_writePorts_3_addr ? io_writePorts_3_data : _GEN_986; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_1051 = 6'h1b == io_writePorts_3_addr ? io_writePorts_3_data : _GEN_987; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_1052 = 6'h1c == io_writePorts_3_addr ? io_writePorts_3_data : _GEN_988; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_1053 = 6'h1d == io_writePorts_3_addr ? io_writePorts_3_data : _GEN_989; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_1054 = 6'h1e == io_writePorts_3_addr ? io_writePorts_3_data : _GEN_990; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_1055 = 6'h1f == io_writePorts_3_addr ? io_writePorts_3_data : _GEN_991; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_1056 = 6'h20 == io_writePorts_3_addr ? io_writePorts_3_data : _GEN_992; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_1057 = 6'h21 == io_writePorts_3_addr ? io_writePorts_3_data : _GEN_993; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_1058 = 6'h22 == io_writePorts_3_addr ? io_writePorts_3_data : _GEN_994; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_1059 = 6'h23 == io_writePorts_3_addr ? io_writePorts_3_data : _GEN_995; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_1060 = 6'h24 == io_writePorts_3_addr ? io_writePorts_3_data : _GEN_996; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_1061 = 6'h25 == io_writePorts_3_addr ? io_writePorts_3_data : _GEN_997; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_1062 = 6'h26 == io_writePorts_3_addr ? io_writePorts_3_data : _GEN_998; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_1063 = 6'h27 == io_writePorts_3_addr ? io_writePorts_3_data : _GEN_999; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_1064 = 6'h28 == io_writePorts_3_addr ? io_writePorts_3_data : _GEN_1000; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_1065 = 6'h29 == io_writePorts_3_addr ? io_writePorts_3_data : _GEN_1001; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_1066 = 6'h2a == io_writePorts_3_addr ? io_writePorts_3_data : _GEN_1002; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_1067 = 6'h2b == io_writePorts_3_addr ? io_writePorts_3_data : _GEN_1003; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_1068 = 6'h2c == io_writePorts_3_addr ? io_writePorts_3_data : _GEN_1004; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_1069 = 6'h2d == io_writePorts_3_addr ? io_writePorts_3_data : _GEN_1005; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_1070 = 6'h2e == io_writePorts_3_addr ? io_writePorts_3_data : _GEN_1006; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_1071 = 6'h2f == io_writePorts_3_addr ? io_writePorts_3_data : _GEN_1007; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_1072 = 6'h30 == io_writePorts_3_addr ? io_writePorts_3_data : _GEN_1008; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_1073 = 6'h31 == io_writePorts_3_addr ? io_writePorts_3_data : _GEN_1009; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_1074 = 6'h32 == io_writePorts_3_addr ? io_writePorts_3_data : _GEN_1010; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_1075 = 6'h33 == io_writePorts_3_addr ? io_writePorts_3_data : _GEN_1011; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_1076 = 6'h34 == io_writePorts_3_addr ? io_writePorts_3_data : _GEN_1012; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_1077 = 6'h35 == io_writePorts_3_addr ? io_writePorts_3_data : _GEN_1013; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_1078 = 6'h36 == io_writePorts_3_addr ? io_writePorts_3_data : _GEN_1014; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_1079 = 6'h37 == io_writePorts_3_addr ? io_writePorts_3_data : _GEN_1015; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_1080 = 6'h38 == io_writePorts_3_addr ? io_writePorts_3_data : _GEN_1016; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_1081 = 6'h39 == io_writePorts_3_addr ? io_writePorts_3_data : _GEN_1017; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_1082 = 6'h3a == io_writePorts_3_addr ? io_writePorts_3_data : _GEN_1018; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_1083 = 6'h3b == io_writePorts_3_addr ? io_writePorts_3_data : _GEN_1019; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_1084 = 6'h3c == io_writePorts_3_addr ? io_writePorts_3_data : _GEN_1020; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_1085 = 6'h3d == io_writePorts_3_addr ? io_writePorts_3_data : _GEN_1021; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_1086 = 6'h3e == io_writePorts_3_addr ? io_writePorts_3_data : _GEN_1022; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_1087 = 6'h3f == io_writePorts_3_addr ? io_writePorts_3_data : _GEN_1023; // @[Regfile.scala 58:{19,19}]
  wire [63:0] _GEN_1088 = io_writePorts_3_wen ? _GEN_1024 : _GEN_960; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1089 = io_writePorts_3_wen ? _GEN_1025 : _GEN_961; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1090 = io_writePorts_3_wen ? _GEN_1026 : _GEN_962; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1091 = io_writePorts_3_wen ? _GEN_1027 : _GEN_963; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1092 = io_writePorts_3_wen ? _GEN_1028 : _GEN_964; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1093 = io_writePorts_3_wen ? _GEN_1029 : _GEN_965; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1094 = io_writePorts_3_wen ? _GEN_1030 : _GEN_966; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1095 = io_writePorts_3_wen ? _GEN_1031 : _GEN_967; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1096 = io_writePorts_3_wen ? _GEN_1032 : _GEN_968; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1097 = io_writePorts_3_wen ? _GEN_1033 : _GEN_969; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1098 = io_writePorts_3_wen ? _GEN_1034 : _GEN_970; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1099 = io_writePorts_3_wen ? _GEN_1035 : _GEN_971; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1100 = io_writePorts_3_wen ? _GEN_1036 : _GEN_972; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1101 = io_writePorts_3_wen ? _GEN_1037 : _GEN_973; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1102 = io_writePorts_3_wen ? _GEN_1038 : _GEN_974; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1103 = io_writePorts_3_wen ? _GEN_1039 : _GEN_975; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1104 = io_writePorts_3_wen ? _GEN_1040 : _GEN_976; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1105 = io_writePorts_3_wen ? _GEN_1041 : _GEN_977; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1106 = io_writePorts_3_wen ? _GEN_1042 : _GEN_978; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1107 = io_writePorts_3_wen ? _GEN_1043 : _GEN_979; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1108 = io_writePorts_3_wen ? _GEN_1044 : _GEN_980; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1109 = io_writePorts_3_wen ? _GEN_1045 : _GEN_981; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1110 = io_writePorts_3_wen ? _GEN_1046 : _GEN_982; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1111 = io_writePorts_3_wen ? _GEN_1047 : _GEN_983; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1112 = io_writePorts_3_wen ? _GEN_1048 : _GEN_984; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1113 = io_writePorts_3_wen ? _GEN_1049 : _GEN_985; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1114 = io_writePorts_3_wen ? _GEN_1050 : _GEN_986; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1115 = io_writePorts_3_wen ? _GEN_1051 : _GEN_987; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1116 = io_writePorts_3_wen ? _GEN_1052 : _GEN_988; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1117 = io_writePorts_3_wen ? _GEN_1053 : _GEN_989; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1118 = io_writePorts_3_wen ? _GEN_1054 : _GEN_990; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1119 = io_writePorts_3_wen ? _GEN_1055 : _GEN_991; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1120 = io_writePorts_3_wen ? _GEN_1056 : _GEN_992; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1121 = io_writePorts_3_wen ? _GEN_1057 : _GEN_993; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1122 = io_writePorts_3_wen ? _GEN_1058 : _GEN_994; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1123 = io_writePorts_3_wen ? _GEN_1059 : _GEN_995; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1124 = io_writePorts_3_wen ? _GEN_1060 : _GEN_996; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1125 = io_writePorts_3_wen ? _GEN_1061 : _GEN_997; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1126 = io_writePorts_3_wen ? _GEN_1062 : _GEN_998; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1127 = io_writePorts_3_wen ? _GEN_1063 : _GEN_999; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1128 = io_writePorts_3_wen ? _GEN_1064 : _GEN_1000; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1129 = io_writePorts_3_wen ? _GEN_1065 : _GEN_1001; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1130 = io_writePorts_3_wen ? _GEN_1066 : _GEN_1002; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1131 = io_writePorts_3_wen ? _GEN_1067 : _GEN_1003; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1132 = io_writePorts_3_wen ? _GEN_1068 : _GEN_1004; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1133 = io_writePorts_3_wen ? _GEN_1069 : _GEN_1005; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1134 = io_writePorts_3_wen ? _GEN_1070 : _GEN_1006; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1135 = io_writePorts_3_wen ? _GEN_1071 : _GEN_1007; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1136 = io_writePorts_3_wen ? _GEN_1072 : _GEN_1008; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1137 = io_writePorts_3_wen ? _GEN_1073 : _GEN_1009; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1138 = io_writePorts_3_wen ? _GEN_1074 : _GEN_1010; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1139 = io_writePorts_3_wen ? _GEN_1075 : _GEN_1011; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1140 = io_writePorts_3_wen ? _GEN_1076 : _GEN_1012; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1141 = io_writePorts_3_wen ? _GEN_1077 : _GEN_1013; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1142 = io_writePorts_3_wen ? _GEN_1078 : _GEN_1014; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1143 = io_writePorts_3_wen ? _GEN_1079 : _GEN_1015; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1144 = io_writePorts_3_wen ? _GEN_1080 : _GEN_1016; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1145 = io_writePorts_3_wen ? _GEN_1081 : _GEN_1017; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1146 = io_writePorts_3_wen ? _GEN_1082 : _GEN_1018; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1147 = io_writePorts_3_wen ? _GEN_1083 : _GEN_1019; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1148 = io_writePorts_3_wen ? _GEN_1084 : _GEN_1020; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1149 = io_writePorts_3_wen ? _GEN_1085 : _GEN_1021; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1150 = io_writePorts_3_wen ? _GEN_1086 : _GEN_1022; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1151 = io_writePorts_3_wen ? _GEN_1087 : _GEN_1023; // @[Regfile.scala 57:17]
  wire [63:0] _GEN_1281 = 6'h1 == io_debug_rports_0_addr ? mem_1 : mem_0; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1282 = 6'h2 == io_debug_rports_0_addr ? mem_2 : _GEN_1281; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1283 = 6'h3 == io_debug_rports_0_addr ? mem_3 : _GEN_1282; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1284 = 6'h4 == io_debug_rports_0_addr ? mem_4 : _GEN_1283; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1285 = 6'h5 == io_debug_rports_0_addr ? mem_5 : _GEN_1284; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1286 = 6'h6 == io_debug_rports_0_addr ? mem_6 : _GEN_1285; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1287 = 6'h7 == io_debug_rports_0_addr ? mem_7 : _GEN_1286; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1288 = 6'h8 == io_debug_rports_0_addr ? mem_8 : _GEN_1287; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1289 = 6'h9 == io_debug_rports_0_addr ? mem_9 : _GEN_1288; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1290 = 6'ha == io_debug_rports_0_addr ? mem_10 : _GEN_1289; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1291 = 6'hb == io_debug_rports_0_addr ? mem_11 : _GEN_1290; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1292 = 6'hc == io_debug_rports_0_addr ? mem_12 : _GEN_1291; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1293 = 6'hd == io_debug_rports_0_addr ? mem_13 : _GEN_1292; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1294 = 6'he == io_debug_rports_0_addr ? mem_14 : _GEN_1293; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1295 = 6'hf == io_debug_rports_0_addr ? mem_15 : _GEN_1294; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1296 = 6'h10 == io_debug_rports_0_addr ? mem_16 : _GEN_1295; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1297 = 6'h11 == io_debug_rports_0_addr ? mem_17 : _GEN_1296; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1298 = 6'h12 == io_debug_rports_0_addr ? mem_18 : _GEN_1297; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1299 = 6'h13 == io_debug_rports_0_addr ? mem_19 : _GEN_1298; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1300 = 6'h14 == io_debug_rports_0_addr ? mem_20 : _GEN_1299; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1301 = 6'h15 == io_debug_rports_0_addr ? mem_21 : _GEN_1300; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1302 = 6'h16 == io_debug_rports_0_addr ? mem_22 : _GEN_1301; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1303 = 6'h17 == io_debug_rports_0_addr ? mem_23 : _GEN_1302; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1304 = 6'h18 == io_debug_rports_0_addr ? mem_24 : _GEN_1303; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1305 = 6'h19 == io_debug_rports_0_addr ? mem_25 : _GEN_1304; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1306 = 6'h1a == io_debug_rports_0_addr ? mem_26 : _GEN_1305; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1307 = 6'h1b == io_debug_rports_0_addr ? mem_27 : _GEN_1306; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1308 = 6'h1c == io_debug_rports_0_addr ? mem_28 : _GEN_1307; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1309 = 6'h1d == io_debug_rports_0_addr ? mem_29 : _GEN_1308; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1310 = 6'h1e == io_debug_rports_0_addr ? mem_30 : _GEN_1309; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1311 = 6'h1f == io_debug_rports_0_addr ? mem_31 : _GEN_1310; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1312 = 6'h20 == io_debug_rports_0_addr ? mem_32 : _GEN_1311; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1313 = 6'h21 == io_debug_rports_0_addr ? mem_33 : _GEN_1312; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1314 = 6'h22 == io_debug_rports_0_addr ? mem_34 : _GEN_1313; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1315 = 6'h23 == io_debug_rports_0_addr ? mem_35 : _GEN_1314; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1316 = 6'h24 == io_debug_rports_0_addr ? mem_36 : _GEN_1315; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1317 = 6'h25 == io_debug_rports_0_addr ? mem_37 : _GEN_1316; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1318 = 6'h26 == io_debug_rports_0_addr ? mem_38 : _GEN_1317; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1319 = 6'h27 == io_debug_rports_0_addr ? mem_39 : _GEN_1318; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1320 = 6'h28 == io_debug_rports_0_addr ? mem_40 : _GEN_1319; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1321 = 6'h29 == io_debug_rports_0_addr ? mem_41 : _GEN_1320; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1322 = 6'h2a == io_debug_rports_0_addr ? mem_42 : _GEN_1321; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1323 = 6'h2b == io_debug_rports_0_addr ? mem_43 : _GEN_1322; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1324 = 6'h2c == io_debug_rports_0_addr ? mem_44 : _GEN_1323; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1325 = 6'h2d == io_debug_rports_0_addr ? mem_45 : _GEN_1324; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1326 = 6'h2e == io_debug_rports_0_addr ? mem_46 : _GEN_1325; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1327 = 6'h2f == io_debug_rports_0_addr ? mem_47 : _GEN_1326; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1328 = 6'h30 == io_debug_rports_0_addr ? mem_48 : _GEN_1327; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1329 = 6'h31 == io_debug_rports_0_addr ? mem_49 : _GEN_1328; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1330 = 6'h32 == io_debug_rports_0_addr ? mem_50 : _GEN_1329; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1331 = 6'h33 == io_debug_rports_0_addr ? mem_51 : _GEN_1330; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1332 = 6'h34 == io_debug_rports_0_addr ? mem_52 : _GEN_1331; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1333 = 6'h35 == io_debug_rports_0_addr ? mem_53 : _GEN_1332; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1334 = 6'h36 == io_debug_rports_0_addr ? mem_54 : _GEN_1333; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1335 = 6'h37 == io_debug_rports_0_addr ? mem_55 : _GEN_1334; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1336 = 6'h38 == io_debug_rports_0_addr ? mem_56 : _GEN_1335; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1337 = 6'h39 == io_debug_rports_0_addr ? mem_57 : _GEN_1336; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1338 = 6'h3a == io_debug_rports_0_addr ? mem_58 : _GEN_1337; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1339 = 6'h3b == io_debug_rports_0_addr ? mem_59 : _GEN_1338; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1340 = 6'h3c == io_debug_rports_0_addr ? mem_60 : _GEN_1339; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1341 = 6'h3d == io_debug_rports_0_addr ? mem_61 : _GEN_1340; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1342 = 6'h3e == io_debug_rports_0_addr ? mem_62 : _GEN_1341; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1343 = 6'h3f == io_debug_rports_0_addr ? mem_63 : _GEN_1342; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1345 = 6'h1 == io_debug_rports_1_addr ? mem_1 : mem_0; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1346 = 6'h2 == io_debug_rports_1_addr ? mem_2 : _GEN_1345; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1347 = 6'h3 == io_debug_rports_1_addr ? mem_3 : _GEN_1346; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1348 = 6'h4 == io_debug_rports_1_addr ? mem_4 : _GEN_1347; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1349 = 6'h5 == io_debug_rports_1_addr ? mem_5 : _GEN_1348; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1350 = 6'h6 == io_debug_rports_1_addr ? mem_6 : _GEN_1349; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1351 = 6'h7 == io_debug_rports_1_addr ? mem_7 : _GEN_1350; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1352 = 6'h8 == io_debug_rports_1_addr ? mem_8 : _GEN_1351; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1353 = 6'h9 == io_debug_rports_1_addr ? mem_9 : _GEN_1352; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1354 = 6'ha == io_debug_rports_1_addr ? mem_10 : _GEN_1353; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1355 = 6'hb == io_debug_rports_1_addr ? mem_11 : _GEN_1354; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1356 = 6'hc == io_debug_rports_1_addr ? mem_12 : _GEN_1355; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1357 = 6'hd == io_debug_rports_1_addr ? mem_13 : _GEN_1356; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1358 = 6'he == io_debug_rports_1_addr ? mem_14 : _GEN_1357; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1359 = 6'hf == io_debug_rports_1_addr ? mem_15 : _GEN_1358; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1360 = 6'h10 == io_debug_rports_1_addr ? mem_16 : _GEN_1359; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1361 = 6'h11 == io_debug_rports_1_addr ? mem_17 : _GEN_1360; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1362 = 6'h12 == io_debug_rports_1_addr ? mem_18 : _GEN_1361; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1363 = 6'h13 == io_debug_rports_1_addr ? mem_19 : _GEN_1362; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1364 = 6'h14 == io_debug_rports_1_addr ? mem_20 : _GEN_1363; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1365 = 6'h15 == io_debug_rports_1_addr ? mem_21 : _GEN_1364; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1366 = 6'h16 == io_debug_rports_1_addr ? mem_22 : _GEN_1365; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1367 = 6'h17 == io_debug_rports_1_addr ? mem_23 : _GEN_1366; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1368 = 6'h18 == io_debug_rports_1_addr ? mem_24 : _GEN_1367; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1369 = 6'h19 == io_debug_rports_1_addr ? mem_25 : _GEN_1368; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1370 = 6'h1a == io_debug_rports_1_addr ? mem_26 : _GEN_1369; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1371 = 6'h1b == io_debug_rports_1_addr ? mem_27 : _GEN_1370; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1372 = 6'h1c == io_debug_rports_1_addr ? mem_28 : _GEN_1371; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1373 = 6'h1d == io_debug_rports_1_addr ? mem_29 : _GEN_1372; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1374 = 6'h1e == io_debug_rports_1_addr ? mem_30 : _GEN_1373; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1375 = 6'h1f == io_debug_rports_1_addr ? mem_31 : _GEN_1374; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1376 = 6'h20 == io_debug_rports_1_addr ? mem_32 : _GEN_1375; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1377 = 6'h21 == io_debug_rports_1_addr ? mem_33 : _GEN_1376; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1378 = 6'h22 == io_debug_rports_1_addr ? mem_34 : _GEN_1377; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1379 = 6'h23 == io_debug_rports_1_addr ? mem_35 : _GEN_1378; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1380 = 6'h24 == io_debug_rports_1_addr ? mem_36 : _GEN_1379; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1381 = 6'h25 == io_debug_rports_1_addr ? mem_37 : _GEN_1380; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1382 = 6'h26 == io_debug_rports_1_addr ? mem_38 : _GEN_1381; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1383 = 6'h27 == io_debug_rports_1_addr ? mem_39 : _GEN_1382; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1384 = 6'h28 == io_debug_rports_1_addr ? mem_40 : _GEN_1383; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1385 = 6'h29 == io_debug_rports_1_addr ? mem_41 : _GEN_1384; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1386 = 6'h2a == io_debug_rports_1_addr ? mem_42 : _GEN_1385; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1387 = 6'h2b == io_debug_rports_1_addr ? mem_43 : _GEN_1386; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1388 = 6'h2c == io_debug_rports_1_addr ? mem_44 : _GEN_1387; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1389 = 6'h2d == io_debug_rports_1_addr ? mem_45 : _GEN_1388; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1390 = 6'h2e == io_debug_rports_1_addr ? mem_46 : _GEN_1389; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1391 = 6'h2f == io_debug_rports_1_addr ? mem_47 : _GEN_1390; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1392 = 6'h30 == io_debug_rports_1_addr ? mem_48 : _GEN_1391; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1393 = 6'h31 == io_debug_rports_1_addr ? mem_49 : _GEN_1392; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1394 = 6'h32 == io_debug_rports_1_addr ? mem_50 : _GEN_1393; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1395 = 6'h33 == io_debug_rports_1_addr ? mem_51 : _GEN_1394; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1396 = 6'h34 == io_debug_rports_1_addr ? mem_52 : _GEN_1395; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1397 = 6'h35 == io_debug_rports_1_addr ? mem_53 : _GEN_1396; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1398 = 6'h36 == io_debug_rports_1_addr ? mem_54 : _GEN_1397; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1399 = 6'h37 == io_debug_rports_1_addr ? mem_55 : _GEN_1398; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1400 = 6'h38 == io_debug_rports_1_addr ? mem_56 : _GEN_1399; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1401 = 6'h39 == io_debug_rports_1_addr ? mem_57 : _GEN_1400; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1402 = 6'h3a == io_debug_rports_1_addr ? mem_58 : _GEN_1401; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1403 = 6'h3b == io_debug_rports_1_addr ? mem_59 : _GEN_1402; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1404 = 6'h3c == io_debug_rports_1_addr ? mem_60 : _GEN_1403; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1405 = 6'h3d == io_debug_rports_1_addr ? mem_61 : _GEN_1404; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1406 = 6'h3e == io_debug_rports_1_addr ? mem_62 : _GEN_1405; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1407 = 6'h3f == io_debug_rports_1_addr ? mem_63 : _GEN_1406; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1409 = 6'h1 == io_debug_rports_2_addr ? mem_1 : mem_0; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1410 = 6'h2 == io_debug_rports_2_addr ? mem_2 : _GEN_1409; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1411 = 6'h3 == io_debug_rports_2_addr ? mem_3 : _GEN_1410; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1412 = 6'h4 == io_debug_rports_2_addr ? mem_4 : _GEN_1411; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1413 = 6'h5 == io_debug_rports_2_addr ? mem_5 : _GEN_1412; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1414 = 6'h6 == io_debug_rports_2_addr ? mem_6 : _GEN_1413; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1415 = 6'h7 == io_debug_rports_2_addr ? mem_7 : _GEN_1414; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1416 = 6'h8 == io_debug_rports_2_addr ? mem_8 : _GEN_1415; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1417 = 6'h9 == io_debug_rports_2_addr ? mem_9 : _GEN_1416; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1418 = 6'ha == io_debug_rports_2_addr ? mem_10 : _GEN_1417; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1419 = 6'hb == io_debug_rports_2_addr ? mem_11 : _GEN_1418; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1420 = 6'hc == io_debug_rports_2_addr ? mem_12 : _GEN_1419; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1421 = 6'hd == io_debug_rports_2_addr ? mem_13 : _GEN_1420; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1422 = 6'he == io_debug_rports_2_addr ? mem_14 : _GEN_1421; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1423 = 6'hf == io_debug_rports_2_addr ? mem_15 : _GEN_1422; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1424 = 6'h10 == io_debug_rports_2_addr ? mem_16 : _GEN_1423; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1425 = 6'h11 == io_debug_rports_2_addr ? mem_17 : _GEN_1424; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1426 = 6'h12 == io_debug_rports_2_addr ? mem_18 : _GEN_1425; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1427 = 6'h13 == io_debug_rports_2_addr ? mem_19 : _GEN_1426; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1428 = 6'h14 == io_debug_rports_2_addr ? mem_20 : _GEN_1427; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1429 = 6'h15 == io_debug_rports_2_addr ? mem_21 : _GEN_1428; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1430 = 6'h16 == io_debug_rports_2_addr ? mem_22 : _GEN_1429; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1431 = 6'h17 == io_debug_rports_2_addr ? mem_23 : _GEN_1430; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1432 = 6'h18 == io_debug_rports_2_addr ? mem_24 : _GEN_1431; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1433 = 6'h19 == io_debug_rports_2_addr ? mem_25 : _GEN_1432; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1434 = 6'h1a == io_debug_rports_2_addr ? mem_26 : _GEN_1433; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1435 = 6'h1b == io_debug_rports_2_addr ? mem_27 : _GEN_1434; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1436 = 6'h1c == io_debug_rports_2_addr ? mem_28 : _GEN_1435; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1437 = 6'h1d == io_debug_rports_2_addr ? mem_29 : _GEN_1436; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1438 = 6'h1e == io_debug_rports_2_addr ? mem_30 : _GEN_1437; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1439 = 6'h1f == io_debug_rports_2_addr ? mem_31 : _GEN_1438; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1440 = 6'h20 == io_debug_rports_2_addr ? mem_32 : _GEN_1439; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1441 = 6'h21 == io_debug_rports_2_addr ? mem_33 : _GEN_1440; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1442 = 6'h22 == io_debug_rports_2_addr ? mem_34 : _GEN_1441; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1443 = 6'h23 == io_debug_rports_2_addr ? mem_35 : _GEN_1442; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1444 = 6'h24 == io_debug_rports_2_addr ? mem_36 : _GEN_1443; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1445 = 6'h25 == io_debug_rports_2_addr ? mem_37 : _GEN_1444; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1446 = 6'h26 == io_debug_rports_2_addr ? mem_38 : _GEN_1445; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1447 = 6'h27 == io_debug_rports_2_addr ? mem_39 : _GEN_1446; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1448 = 6'h28 == io_debug_rports_2_addr ? mem_40 : _GEN_1447; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1449 = 6'h29 == io_debug_rports_2_addr ? mem_41 : _GEN_1448; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1450 = 6'h2a == io_debug_rports_2_addr ? mem_42 : _GEN_1449; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1451 = 6'h2b == io_debug_rports_2_addr ? mem_43 : _GEN_1450; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1452 = 6'h2c == io_debug_rports_2_addr ? mem_44 : _GEN_1451; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1453 = 6'h2d == io_debug_rports_2_addr ? mem_45 : _GEN_1452; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1454 = 6'h2e == io_debug_rports_2_addr ? mem_46 : _GEN_1453; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1455 = 6'h2f == io_debug_rports_2_addr ? mem_47 : _GEN_1454; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1456 = 6'h30 == io_debug_rports_2_addr ? mem_48 : _GEN_1455; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1457 = 6'h31 == io_debug_rports_2_addr ? mem_49 : _GEN_1456; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1458 = 6'h32 == io_debug_rports_2_addr ? mem_50 : _GEN_1457; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1459 = 6'h33 == io_debug_rports_2_addr ? mem_51 : _GEN_1458; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1460 = 6'h34 == io_debug_rports_2_addr ? mem_52 : _GEN_1459; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1461 = 6'h35 == io_debug_rports_2_addr ? mem_53 : _GEN_1460; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1462 = 6'h36 == io_debug_rports_2_addr ? mem_54 : _GEN_1461; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1463 = 6'h37 == io_debug_rports_2_addr ? mem_55 : _GEN_1462; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1464 = 6'h38 == io_debug_rports_2_addr ? mem_56 : _GEN_1463; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1465 = 6'h39 == io_debug_rports_2_addr ? mem_57 : _GEN_1464; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1466 = 6'h3a == io_debug_rports_2_addr ? mem_58 : _GEN_1465; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1467 = 6'h3b == io_debug_rports_2_addr ? mem_59 : _GEN_1466; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1468 = 6'h3c == io_debug_rports_2_addr ? mem_60 : _GEN_1467; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1469 = 6'h3d == io_debug_rports_2_addr ? mem_61 : _GEN_1468; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1470 = 6'h3e == io_debug_rports_2_addr ? mem_62 : _GEN_1469; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1471 = 6'h3f == io_debug_rports_2_addr ? mem_63 : _GEN_1470; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1473 = 6'h1 == io_debug_rports_3_addr ? mem_1 : mem_0; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1474 = 6'h2 == io_debug_rports_3_addr ? mem_2 : _GEN_1473; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1475 = 6'h3 == io_debug_rports_3_addr ? mem_3 : _GEN_1474; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1476 = 6'h4 == io_debug_rports_3_addr ? mem_4 : _GEN_1475; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1477 = 6'h5 == io_debug_rports_3_addr ? mem_5 : _GEN_1476; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1478 = 6'h6 == io_debug_rports_3_addr ? mem_6 : _GEN_1477; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1479 = 6'h7 == io_debug_rports_3_addr ? mem_7 : _GEN_1478; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1480 = 6'h8 == io_debug_rports_3_addr ? mem_8 : _GEN_1479; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1481 = 6'h9 == io_debug_rports_3_addr ? mem_9 : _GEN_1480; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1482 = 6'ha == io_debug_rports_3_addr ? mem_10 : _GEN_1481; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1483 = 6'hb == io_debug_rports_3_addr ? mem_11 : _GEN_1482; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1484 = 6'hc == io_debug_rports_3_addr ? mem_12 : _GEN_1483; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1485 = 6'hd == io_debug_rports_3_addr ? mem_13 : _GEN_1484; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1486 = 6'he == io_debug_rports_3_addr ? mem_14 : _GEN_1485; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1487 = 6'hf == io_debug_rports_3_addr ? mem_15 : _GEN_1486; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1488 = 6'h10 == io_debug_rports_3_addr ? mem_16 : _GEN_1487; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1489 = 6'h11 == io_debug_rports_3_addr ? mem_17 : _GEN_1488; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1490 = 6'h12 == io_debug_rports_3_addr ? mem_18 : _GEN_1489; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1491 = 6'h13 == io_debug_rports_3_addr ? mem_19 : _GEN_1490; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1492 = 6'h14 == io_debug_rports_3_addr ? mem_20 : _GEN_1491; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1493 = 6'h15 == io_debug_rports_3_addr ? mem_21 : _GEN_1492; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1494 = 6'h16 == io_debug_rports_3_addr ? mem_22 : _GEN_1493; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1495 = 6'h17 == io_debug_rports_3_addr ? mem_23 : _GEN_1494; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1496 = 6'h18 == io_debug_rports_3_addr ? mem_24 : _GEN_1495; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1497 = 6'h19 == io_debug_rports_3_addr ? mem_25 : _GEN_1496; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1498 = 6'h1a == io_debug_rports_3_addr ? mem_26 : _GEN_1497; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1499 = 6'h1b == io_debug_rports_3_addr ? mem_27 : _GEN_1498; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1500 = 6'h1c == io_debug_rports_3_addr ? mem_28 : _GEN_1499; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1501 = 6'h1d == io_debug_rports_3_addr ? mem_29 : _GEN_1500; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1502 = 6'h1e == io_debug_rports_3_addr ? mem_30 : _GEN_1501; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1503 = 6'h1f == io_debug_rports_3_addr ? mem_31 : _GEN_1502; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1504 = 6'h20 == io_debug_rports_3_addr ? mem_32 : _GEN_1503; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1505 = 6'h21 == io_debug_rports_3_addr ? mem_33 : _GEN_1504; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1506 = 6'h22 == io_debug_rports_3_addr ? mem_34 : _GEN_1505; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1507 = 6'h23 == io_debug_rports_3_addr ? mem_35 : _GEN_1506; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1508 = 6'h24 == io_debug_rports_3_addr ? mem_36 : _GEN_1507; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1509 = 6'h25 == io_debug_rports_3_addr ? mem_37 : _GEN_1508; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1510 = 6'h26 == io_debug_rports_3_addr ? mem_38 : _GEN_1509; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1511 = 6'h27 == io_debug_rports_3_addr ? mem_39 : _GEN_1510; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1512 = 6'h28 == io_debug_rports_3_addr ? mem_40 : _GEN_1511; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1513 = 6'h29 == io_debug_rports_3_addr ? mem_41 : _GEN_1512; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1514 = 6'h2a == io_debug_rports_3_addr ? mem_42 : _GEN_1513; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1515 = 6'h2b == io_debug_rports_3_addr ? mem_43 : _GEN_1514; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1516 = 6'h2c == io_debug_rports_3_addr ? mem_44 : _GEN_1515; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1517 = 6'h2d == io_debug_rports_3_addr ? mem_45 : _GEN_1516; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1518 = 6'h2e == io_debug_rports_3_addr ? mem_46 : _GEN_1517; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1519 = 6'h2f == io_debug_rports_3_addr ? mem_47 : _GEN_1518; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1520 = 6'h30 == io_debug_rports_3_addr ? mem_48 : _GEN_1519; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1521 = 6'h31 == io_debug_rports_3_addr ? mem_49 : _GEN_1520; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1522 = 6'h32 == io_debug_rports_3_addr ? mem_50 : _GEN_1521; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1523 = 6'h33 == io_debug_rports_3_addr ? mem_51 : _GEN_1522; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1524 = 6'h34 == io_debug_rports_3_addr ? mem_52 : _GEN_1523; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1525 = 6'h35 == io_debug_rports_3_addr ? mem_53 : _GEN_1524; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1526 = 6'h36 == io_debug_rports_3_addr ? mem_54 : _GEN_1525; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1527 = 6'h37 == io_debug_rports_3_addr ? mem_55 : _GEN_1526; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1528 = 6'h38 == io_debug_rports_3_addr ? mem_56 : _GEN_1527; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1529 = 6'h39 == io_debug_rports_3_addr ? mem_57 : _GEN_1528; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1530 = 6'h3a == io_debug_rports_3_addr ? mem_58 : _GEN_1529; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1531 = 6'h3b == io_debug_rports_3_addr ? mem_59 : _GEN_1530; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1532 = 6'h3c == io_debug_rports_3_addr ? mem_60 : _GEN_1531; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1533 = 6'h3d == io_debug_rports_3_addr ? mem_61 : _GEN_1532; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1534 = 6'h3e == io_debug_rports_3_addr ? mem_62 : _GEN_1533; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1535 = 6'h3f == io_debug_rports_3_addr ? mem_63 : _GEN_1534; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1537 = 6'h1 == io_debug_rports_4_addr ? mem_1 : mem_0; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1538 = 6'h2 == io_debug_rports_4_addr ? mem_2 : _GEN_1537; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1539 = 6'h3 == io_debug_rports_4_addr ? mem_3 : _GEN_1538; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1540 = 6'h4 == io_debug_rports_4_addr ? mem_4 : _GEN_1539; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1541 = 6'h5 == io_debug_rports_4_addr ? mem_5 : _GEN_1540; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1542 = 6'h6 == io_debug_rports_4_addr ? mem_6 : _GEN_1541; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1543 = 6'h7 == io_debug_rports_4_addr ? mem_7 : _GEN_1542; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1544 = 6'h8 == io_debug_rports_4_addr ? mem_8 : _GEN_1543; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1545 = 6'h9 == io_debug_rports_4_addr ? mem_9 : _GEN_1544; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1546 = 6'ha == io_debug_rports_4_addr ? mem_10 : _GEN_1545; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1547 = 6'hb == io_debug_rports_4_addr ? mem_11 : _GEN_1546; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1548 = 6'hc == io_debug_rports_4_addr ? mem_12 : _GEN_1547; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1549 = 6'hd == io_debug_rports_4_addr ? mem_13 : _GEN_1548; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1550 = 6'he == io_debug_rports_4_addr ? mem_14 : _GEN_1549; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1551 = 6'hf == io_debug_rports_4_addr ? mem_15 : _GEN_1550; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1552 = 6'h10 == io_debug_rports_4_addr ? mem_16 : _GEN_1551; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1553 = 6'h11 == io_debug_rports_4_addr ? mem_17 : _GEN_1552; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1554 = 6'h12 == io_debug_rports_4_addr ? mem_18 : _GEN_1553; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1555 = 6'h13 == io_debug_rports_4_addr ? mem_19 : _GEN_1554; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1556 = 6'h14 == io_debug_rports_4_addr ? mem_20 : _GEN_1555; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1557 = 6'h15 == io_debug_rports_4_addr ? mem_21 : _GEN_1556; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1558 = 6'h16 == io_debug_rports_4_addr ? mem_22 : _GEN_1557; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1559 = 6'h17 == io_debug_rports_4_addr ? mem_23 : _GEN_1558; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1560 = 6'h18 == io_debug_rports_4_addr ? mem_24 : _GEN_1559; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1561 = 6'h19 == io_debug_rports_4_addr ? mem_25 : _GEN_1560; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1562 = 6'h1a == io_debug_rports_4_addr ? mem_26 : _GEN_1561; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1563 = 6'h1b == io_debug_rports_4_addr ? mem_27 : _GEN_1562; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1564 = 6'h1c == io_debug_rports_4_addr ? mem_28 : _GEN_1563; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1565 = 6'h1d == io_debug_rports_4_addr ? mem_29 : _GEN_1564; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1566 = 6'h1e == io_debug_rports_4_addr ? mem_30 : _GEN_1565; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1567 = 6'h1f == io_debug_rports_4_addr ? mem_31 : _GEN_1566; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1568 = 6'h20 == io_debug_rports_4_addr ? mem_32 : _GEN_1567; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1569 = 6'h21 == io_debug_rports_4_addr ? mem_33 : _GEN_1568; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1570 = 6'h22 == io_debug_rports_4_addr ? mem_34 : _GEN_1569; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1571 = 6'h23 == io_debug_rports_4_addr ? mem_35 : _GEN_1570; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1572 = 6'h24 == io_debug_rports_4_addr ? mem_36 : _GEN_1571; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1573 = 6'h25 == io_debug_rports_4_addr ? mem_37 : _GEN_1572; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1574 = 6'h26 == io_debug_rports_4_addr ? mem_38 : _GEN_1573; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1575 = 6'h27 == io_debug_rports_4_addr ? mem_39 : _GEN_1574; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1576 = 6'h28 == io_debug_rports_4_addr ? mem_40 : _GEN_1575; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1577 = 6'h29 == io_debug_rports_4_addr ? mem_41 : _GEN_1576; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1578 = 6'h2a == io_debug_rports_4_addr ? mem_42 : _GEN_1577; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1579 = 6'h2b == io_debug_rports_4_addr ? mem_43 : _GEN_1578; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1580 = 6'h2c == io_debug_rports_4_addr ? mem_44 : _GEN_1579; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1581 = 6'h2d == io_debug_rports_4_addr ? mem_45 : _GEN_1580; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1582 = 6'h2e == io_debug_rports_4_addr ? mem_46 : _GEN_1581; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1583 = 6'h2f == io_debug_rports_4_addr ? mem_47 : _GEN_1582; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1584 = 6'h30 == io_debug_rports_4_addr ? mem_48 : _GEN_1583; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1585 = 6'h31 == io_debug_rports_4_addr ? mem_49 : _GEN_1584; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1586 = 6'h32 == io_debug_rports_4_addr ? mem_50 : _GEN_1585; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1587 = 6'h33 == io_debug_rports_4_addr ? mem_51 : _GEN_1586; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1588 = 6'h34 == io_debug_rports_4_addr ? mem_52 : _GEN_1587; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1589 = 6'h35 == io_debug_rports_4_addr ? mem_53 : _GEN_1588; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1590 = 6'h36 == io_debug_rports_4_addr ? mem_54 : _GEN_1589; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1591 = 6'h37 == io_debug_rports_4_addr ? mem_55 : _GEN_1590; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1592 = 6'h38 == io_debug_rports_4_addr ? mem_56 : _GEN_1591; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1593 = 6'h39 == io_debug_rports_4_addr ? mem_57 : _GEN_1592; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1594 = 6'h3a == io_debug_rports_4_addr ? mem_58 : _GEN_1593; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1595 = 6'h3b == io_debug_rports_4_addr ? mem_59 : _GEN_1594; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1596 = 6'h3c == io_debug_rports_4_addr ? mem_60 : _GEN_1595; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1597 = 6'h3d == io_debug_rports_4_addr ? mem_61 : _GEN_1596; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1598 = 6'h3e == io_debug_rports_4_addr ? mem_62 : _GEN_1597; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1599 = 6'h3f == io_debug_rports_4_addr ? mem_63 : _GEN_1598; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1601 = 6'h1 == io_debug_rports_5_addr ? mem_1 : mem_0; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1602 = 6'h2 == io_debug_rports_5_addr ? mem_2 : _GEN_1601; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1603 = 6'h3 == io_debug_rports_5_addr ? mem_3 : _GEN_1602; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1604 = 6'h4 == io_debug_rports_5_addr ? mem_4 : _GEN_1603; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1605 = 6'h5 == io_debug_rports_5_addr ? mem_5 : _GEN_1604; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1606 = 6'h6 == io_debug_rports_5_addr ? mem_6 : _GEN_1605; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1607 = 6'h7 == io_debug_rports_5_addr ? mem_7 : _GEN_1606; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1608 = 6'h8 == io_debug_rports_5_addr ? mem_8 : _GEN_1607; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1609 = 6'h9 == io_debug_rports_5_addr ? mem_9 : _GEN_1608; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1610 = 6'ha == io_debug_rports_5_addr ? mem_10 : _GEN_1609; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1611 = 6'hb == io_debug_rports_5_addr ? mem_11 : _GEN_1610; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1612 = 6'hc == io_debug_rports_5_addr ? mem_12 : _GEN_1611; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1613 = 6'hd == io_debug_rports_5_addr ? mem_13 : _GEN_1612; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1614 = 6'he == io_debug_rports_5_addr ? mem_14 : _GEN_1613; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1615 = 6'hf == io_debug_rports_5_addr ? mem_15 : _GEN_1614; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1616 = 6'h10 == io_debug_rports_5_addr ? mem_16 : _GEN_1615; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1617 = 6'h11 == io_debug_rports_5_addr ? mem_17 : _GEN_1616; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1618 = 6'h12 == io_debug_rports_5_addr ? mem_18 : _GEN_1617; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1619 = 6'h13 == io_debug_rports_5_addr ? mem_19 : _GEN_1618; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1620 = 6'h14 == io_debug_rports_5_addr ? mem_20 : _GEN_1619; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1621 = 6'h15 == io_debug_rports_5_addr ? mem_21 : _GEN_1620; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1622 = 6'h16 == io_debug_rports_5_addr ? mem_22 : _GEN_1621; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1623 = 6'h17 == io_debug_rports_5_addr ? mem_23 : _GEN_1622; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1624 = 6'h18 == io_debug_rports_5_addr ? mem_24 : _GEN_1623; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1625 = 6'h19 == io_debug_rports_5_addr ? mem_25 : _GEN_1624; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1626 = 6'h1a == io_debug_rports_5_addr ? mem_26 : _GEN_1625; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1627 = 6'h1b == io_debug_rports_5_addr ? mem_27 : _GEN_1626; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1628 = 6'h1c == io_debug_rports_5_addr ? mem_28 : _GEN_1627; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1629 = 6'h1d == io_debug_rports_5_addr ? mem_29 : _GEN_1628; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1630 = 6'h1e == io_debug_rports_5_addr ? mem_30 : _GEN_1629; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1631 = 6'h1f == io_debug_rports_5_addr ? mem_31 : _GEN_1630; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1632 = 6'h20 == io_debug_rports_5_addr ? mem_32 : _GEN_1631; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1633 = 6'h21 == io_debug_rports_5_addr ? mem_33 : _GEN_1632; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1634 = 6'h22 == io_debug_rports_5_addr ? mem_34 : _GEN_1633; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1635 = 6'h23 == io_debug_rports_5_addr ? mem_35 : _GEN_1634; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1636 = 6'h24 == io_debug_rports_5_addr ? mem_36 : _GEN_1635; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1637 = 6'h25 == io_debug_rports_5_addr ? mem_37 : _GEN_1636; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1638 = 6'h26 == io_debug_rports_5_addr ? mem_38 : _GEN_1637; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1639 = 6'h27 == io_debug_rports_5_addr ? mem_39 : _GEN_1638; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1640 = 6'h28 == io_debug_rports_5_addr ? mem_40 : _GEN_1639; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1641 = 6'h29 == io_debug_rports_5_addr ? mem_41 : _GEN_1640; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1642 = 6'h2a == io_debug_rports_5_addr ? mem_42 : _GEN_1641; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1643 = 6'h2b == io_debug_rports_5_addr ? mem_43 : _GEN_1642; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1644 = 6'h2c == io_debug_rports_5_addr ? mem_44 : _GEN_1643; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1645 = 6'h2d == io_debug_rports_5_addr ? mem_45 : _GEN_1644; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1646 = 6'h2e == io_debug_rports_5_addr ? mem_46 : _GEN_1645; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1647 = 6'h2f == io_debug_rports_5_addr ? mem_47 : _GEN_1646; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1648 = 6'h30 == io_debug_rports_5_addr ? mem_48 : _GEN_1647; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1649 = 6'h31 == io_debug_rports_5_addr ? mem_49 : _GEN_1648; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1650 = 6'h32 == io_debug_rports_5_addr ? mem_50 : _GEN_1649; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1651 = 6'h33 == io_debug_rports_5_addr ? mem_51 : _GEN_1650; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1652 = 6'h34 == io_debug_rports_5_addr ? mem_52 : _GEN_1651; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1653 = 6'h35 == io_debug_rports_5_addr ? mem_53 : _GEN_1652; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1654 = 6'h36 == io_debug_rports_5_addr ? mem_54 : _GEN_1653; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1655 = 6'h37 == io_debug_rports_5_addr ? mem_55 : _GEN_1654; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1656 = 6'h38 == io_debug_rports_5_addr ? mem_56 : _GEN_1655; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1657 = 6'h39 == io_debug_rports_5_addr ? mem_57 : _GEN_1656; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1658 = 6'h3a == io_debug_rports_5_addr ? mem_58 : _GEN_1657; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1659 = 6'h3b == io_debug_rports_5_addr ? mem_59 : _GEN_1658; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1660 = 6'h3c == io_debug_rports_5_addr ? mem_60 : _GEN_1659; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1661 = 6'h3d == io_debug_rports_5_addr ? mem_61 : _GEN_1660; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1662 = 6'h3e == io_debug_rports_5_addr ? mem_62 : _GEN_1661; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1663 = 6'h3f == io_debug_rports_5_addr ? mem_63 : _GEN_1662; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1665 = 6'h1 == io_debug_rports_6_addr ? mem_1 : mem_0; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1666 = 6'h2 == io_debug_rports_6_addr ? mem_2 : _GEN_1665; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1667 = 6'h3 == io_debug_rports_6_addr ? mem_3 : _GEN_1666; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1668 = 6'h4 == io_debug_rports_6_addr ? mem_4 : _GEN_1667; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1669 = 6'h5 == io_debug_rports_6_addr ? mem_5 : _GEN_1668; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1670 = 6'h6 == io_debug_rports_6_addr ? mem_6 : _GEN_1669; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1671 = 6'h7 == io_debug_rports_6_addr ? mem_7 : _GEN_1670; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1672 = 6'h8 == io_debug_rports_6_addr ? mem_8 : _GEN_1671; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1673 = 6'h9 == io_debug_rports_6_addr ? mem_9 : _GEN_1672; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1674 = 6'ha == io_debug_rports_6_addr ? mem_10 : _GEN_1673; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1675 = 6'hb == io_debug_rports_6_addr ? mem_11 : _GEN_1674; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1676 = 6'hc == io_debug_rports_6_addr ? mem_12 : _GEN_1675; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1677 = 6'hd == io_debug_rports_6_addr ? mem_13 : _GEN_1676; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1678 = 6'he == io_debug_rports_6_addr ? mem_14 : _GEN_1677; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1679 = 6'hf == io_debug_rports_6_addr ? mem_15 : _GEN_1678; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1680 = 6'h10 == io_debug_rports_6_addr ? mem_16 : _GEN_1679; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1681 = 6'h11 == io_debug_rports_6_addr ? mem_17 : _GEN_1680; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1682 = 6'h12 == io_debug_rports_6_addr ? mem_18 : _GEN_1681; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1683 = 6'h13 == io_debug_rports_6_addr ? mem_19 : _GEN_1682; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1684 = 6'h14 == io_debug_rports_6_addr ? mem_20 : _GEN_1683; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1685 = 6'h15 == io_debug_rports_6_addr ? mem_21 : _GEN_1684; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1686 = 6'h16 == io_debug_rports_6_addr ? mem_22 : _GEN_1685; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1687 = 6'h17 == io_debug_rports_6_addr ? mem_23 : _GEN_1686; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1688 = 6'h18 == io_debug_rports_6_addr ? mem_24 : _GEN_1687; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1689 = 6'h19 == io_debug_rports_6_addr ? mem_25 : _GEN_1688; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1690 = 6'h1a == io_debug_rports_6_addr ? mem_26 : _GEN_1689; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1691 = 6'h1b == io_debug_rports_6_addr ? mem_27 : _GEN_1690; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1692 = 6'h1c == io_debug_rports_6_addr ? mem_28 : _GEN_1691; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1693 = 6'h1d == io_debug_rports_6_addr ? mem_29 : _GEN_1692; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1694 = 6'h1e == io_debug_rports_6_addr ? mem_30 : _GEN_1693; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1695 = 6'h1f == io_debug_rports_6_addr ? mem_31 : _GEN_1694; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1696 = 6'h20 == io_debug_rports_6_addr ? mem_32 : _GEN_1695; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1697 = 6'h21 == io_debug_rports_6_addr ? mem_33 : _GEN_1696; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1698 = 6'h22 == io_debug_rports_6_addr ? mem_34 : _GEN_1697; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1699 = 6'h23 == io_debug_rports_6_addr ? mem_35 : _GEN_1698; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1700 = 6'h24 == io_debug_rports_6_addr ? mem_36 : _GEN_1699; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1701 = 6'h25 == io_debug_rports_6_addr ? mem_37 : _GEN_1700; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1702 = 6'h26 == io_debug_rports_6_addr ? mem_38 : _GEN_1701; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1703 = 6'h27 == io_debug_rports_6_addr ? mem_39 : _GEN_1702; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1704 = 6'h28 == io_debug_rports_6_addr ? mem_40 : _GEN_1703; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1705 = 6'h29 == io_debug_rports_6_addr ? mem_41 : _GEN_1704; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1706 = 6'h2a == io_debug_rports_6_addr ? mem_42 : _GEN_1705; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1707 = 6'h2b == io_debug_rports_6_addr ? mem_43 : _GEN_1706; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1708 = 6'h2c == io_debug_rports_6_addr ? mem_44 : _GEN_1707; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1709 = 6'h2d == io_debug_rports_6_addr ? mem_45 : _GEN_1708; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1710 = 6'h2e == io_debug_rports_6_addr ? mem_46 : _GEN_1709; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1711 = 6'h2f == io_debug_rports_6_addr ? mem_47 : _GEN_1710; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1712 = 6'h30 == io_debug_rports_6_addr ? mem_48 : _GEN_1711; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1713 = 6'h31 == io_debug_rports_6_addr ? mem_49 : _GEN_1712; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1714 = 6'h32 == io_debug_rports_6_addr ? mem_50 : _GEN_1713; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1715 = 6'h33 == io_debug_rports_6_addr ? mem_51 : _GEN_1714; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1716 = 6'h34 == io_debug_rports_6_addr ? mem_52 : _GEN_1715; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1717 = 6'h35 == io_debug_rports_6_addr ? mem_53 : _GEN_1716; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1718 = 6'h36 == io_debug_rports_6_addr ? mem_54 : _GEN_1717; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1719 = 6'h37 == io_debug_rports_6_addr ? mem_55 : _GEN_1718; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1720 = 6'h38 == io_debug_rports_6_addr ? mem_56 : _GEN_1719; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1721 = 6'h39 == io_debug_rports_6_addr ? mem_57 : _GEN_1720; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1722 = 6'h3a == io_debug_rports_6_addr ? mem_58 : _GEN_1721; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1723 = 6'h3b == io_debug_rports_6_addr ? mem_59 : _GEN_1722; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1724 = 6'h3c == io_debug_rports_6_addr ? mem_60 : _GEN_1723; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1725 = 6'h3d == io_debug_rports_6_addr ? mem_61 : _GEN_1724; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1726 = 6'h3e == io_debug_rports_6_addr ? mem_62 : _GEN_1725; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1727 = 6'h3f == io_debug_rports_6_addr ? mem_63 : _GEN_1726; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1729 = 6'h1 == io_debug_rports_7_addr ? mem_1 : mem_0; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1730 = 6'h2 == io_debug_rports_7_addr ? mem_2 : _GEN_1729; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1731 = 6'h3 == io_debug_rports_7_addr ? mem_3 : _GEN_1730; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1732 = 6'h4 == io_debug_rports_7_addr ? mem_4 : _GEN_1731; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1733 = 6'h5 == io_debug_rports_7_addr ? mem_5 : _GEN_1732; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1734 = 6'h6 == io_debug_rports_7_addr ? mem_6 : _GEN_1733; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1735 = 6'h7 == io_debug_rports_7_addr ? mem_7 : _GEN_1734; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1736 = 6'h8 == io_debug_rports_7_addr ? mem_8 : _GEN_1735; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1737 = 6'h9 == io_debug_rports_7_addr ? mem_9 : _GEN_1736; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1738 = 6'ha == io_debug_rports_7_addr ? mem_10 : _GEN_1737; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1739 = 6'hb == io_debug_rports_7_addr ? mem_11 : _GEN_1738; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1740 = 6'hc == io_debug_rports_7_addr ? mem_12 : _GEN_1739; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1741 = 6'hd == io_debug_rports_7_addr ? mem_13 : _GEN_1740; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1742 = 6'he == io_debug_rports_7_addr ? mem_14 : _GEN_1741; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1743 = 6'hf == io_debug_rports_7_addr ? mem_15 : _GEN_1742; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1744 = 6'h10 == io_debug_rports_7_addr ? mem_16 : _GEN_1743; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1745 = 6'h11 == io_debug_rports_7_addr ? mem_17 : _GEN_1744; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1746 = 6'h12 == io_debug_rports_7_addr ? mem_18 : _GEN_1745; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1747 = 6'h13 == io_debug_rports_7_addr ? mem_19 : _GEN_1746; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1748 = 6'h14 == io_debug_rports_7_addr ? mem_20 : _GEN_1747; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1749 = 6'h15 == io_debug_rports_7_addr ? mem_21 : _GEN_1748; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1750 = 6'h16 == io_debug_rports_7_addr ? mem_22 : _GEN_1749; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1751 = 6'h17 == io_debug_rports_7_addr ? mem_23 : _GEN_1750; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1752 = 6'h18 == io_debug_rports_7_addr ? mem_24 : _GEN_1751; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1753 = 6'h19 == io_debug_rports_7_addr ? mem_25 : _GEN_1752; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1754 = 6'h1a == io_debug_rports_7_addr ? mem_26 : _GEN_1753; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1755 = 6'h1b == io_debug_rports_7_addr ? mem_27 : _GEN_1754; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1756 = 6'h1c == io_debug_rports_7_addr ? mem_28 : _GEN_1755; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1757 = 6'h1d == io_debug_rports_7_addr ? mem_29 : _GEN_1756; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1758 = 6'h1e == io_debug_rports_7_addr ? mem_30 : _GEN_1757; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1759 = 6'h1f == io_debug_rports_7_addr ? mem_31 : _GEN_1758; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1760 = 6'h20 == io_debug_rports_7_addr ? mem_32 : _GEN_1759; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1761 = 6'h21 == io_debug_rports_7_addr ? mem_33 : _GEN_1760; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1762 = 6'h22 == io_debug_rports_7_addr ? mem_34 : _GEN_1761; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1763 = 6'h23 == io_debug_rports_7_addr ? mem_35 : _GEN_1762; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1764 = 6'h24 == io_debug_rports_7_addr ? mem_36 : _GEN_1763; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1765 = 6'h25 == io_debug_rports_7_addr ? mem_37 : _GEN_1764; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1766 = 6'h26 == io_debug_rports_7_addr ? mem_38 : _GEN_1765; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1767 = 6'h27 == io_debug_rports_7_addr ? mem_39 : _GEN_1766; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1768 = 6'h28 == io_debug_rports_7_addr ? mem_40 : _GEN_1767; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1769 = 6'h29 == io_debug_rports_7_addr ? mem_41 : _GEN_1768; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1770 = 6'h2a == io_debug_rports_7_addr ? mem_42 : _GEN_1769; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1771 = 6'h2b == io_debug_rports_7_addr ? mem_43 : _GEN_1770; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1772 = 6'h2c == io_debug_rports_7_addr ? mem_44 : _GEN_1771; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1773 = 6'h2d == io_debug_rports_7_addr ? mem_45 : _GEN_1772; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1774 = 6'h2e == io_debug_rports_7_addr ? mem_46 : _GEN_1773; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1775 = 6'h2f == io_debug_rports_7_addr ? mem_47 : _GEN_1774; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1776 = 6'h30 == io_debug_rports_7_addr ? mem_48 : _GEN_1775; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1777 = 6'h31 == io_debug_rports_7_addr ? mem_49 : _GEN_1776; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1778 = 6'h32 == io_debug_rports_7_addr ? mem_50 : _GEN_1777; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1779 = 6'h33 == io_debug_rports_7_addr ? mem_51 : _GEN_1778; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1780 = 6'h34 == io_debug_rports_7_addr ? mem_52 : _GEN_1779; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1781 = 6'h35 == io_debug_rports_7_addr ? mem_53 : _GEN_1780; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1782 = 6'h36 == io_debug_rports_7_addr ? mem_54 : _GEN_1781; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1783 = 6'h37 == io_debug_rports_7_addr ? mem_55 : _GEN_1782; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1784 = 6'h38 == io_debug_rports_7_addr ? mem_56 : _GEN_1783; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1785 = 6'h39 == io_debug_rports_7_addr ? mem_57 : _GEN_1784; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1786 = 6'h3a == io_debug_rports_7_addr ? mem_58 : _GEN_1785; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1787 = 6'h3b == io_debug_rports_7_addr ? mem_59 : _GEN_1786; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1788 = 6'h3c == io_debug_rports_7_addr ? mem_60 : _GEN_1787; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1789 = 6'h3d == io_debug_rports_7_addr ? mem_61 : _GEN_1788; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1790 = 6'h3e == io_debug_rports_7_addr ? mem_62 : _GEN_1789; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1791 = 6'h3f == io_debug_rports_7_addr ? mem_63 : _GEN_1790; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1793 = 6'h1 == io_debug_rports_8_addr ? mem_1 : mem_0; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1794 = 6'h2 == io_debug_rports_8_addr ? mem_2 : _GEN_1793; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1795 = 6'h3 == io_debug_rports_8_addr ? mem_3 : _GEN_1794; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1796 = 6'h4 == io_debug_rports_8_addr ? mem_4 : _GEN_1795; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1797 = 6'h5 == io_debug_rports_8_addr ? mem_5 : _GEN_1796; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1798 = 6'h6 == io_debug_rports_8_addr ? mem_6 : _GEN_1797; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1799 = 6'h7 == io_debug_rports_8_addr ? mem_7 : _GEN_1798; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1800 = 6'h8 == io_debug_rports_8_addr ? mem_8 : _GEN_1799; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1801 = 6'h9 == io_debug_rports_8_addr ? mem_9 : _GEN_1800; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1802 = 6'ha == io_debug_rports_8_addr ? mem_10 : _GEN_1801; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1803 = 6'hb == io_debug_rports_8_addr ? mem_11 : _GEN_1802; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1804 = 6'hc == io_debug_rports_8_addr ? mem_12 : _GEN_1803; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1805 = 6'hd == io_debug_rports_8_addr ? mem_13 : _GEN_1804; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1806 = 6'he == io_debug_rports_8_addr ? mem_14 : _GEN_1805; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1807 = 6'hf == io_debug_rports_8_addr ? mem_15 : _GEN_1806; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1808 = 6'h10 == io_debug_rports_8_addr ? mem_16 : _GEN_1807; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1809 = 6'h11 == io_debug_rports_8_addr ? mem_17 : _GEN_1808; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1810 = 6'h12 == io_debug_rports_8_addr ? mem_18 : _GEN_1809; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1811 = 6'h13 == io_debug_rports_8_addr ? mem_19 : _GEN_1810; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1812 = 6'h14 == io_debug_rports_8_addr ? mem_20 : _GEN_1811; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1813 = 6'h15 == io_debug_rports_8_addr ? mem_21 : _GEN_1812; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1814 = 6'h16 == io_debug_rports_8_addr ? mem_22 : _GEN_1813; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1815 = 6'h17 == io_debug_rports_8_addr ? mem_23 : _GEN_1814; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1816 = 6'h18 == io_debug_rports_8_addr ? mem_24 : _GEN_1815; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1817 = 6'h19 == io_debug_rports_8_addr ? mem_25 : _GEN_1816; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1818 = 6'h1a == io_debug_rports_8_addr ? mem_26 : _GEN_1817; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1819 = 6'h1b == io_debug_rports_8_addr ? mem_27 : _GEN_1818; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1820 = 6'h1c == io_debug_rports_8_addr ? mem_28 : _GEN_1819; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1821 = 6'h1d == io_debug_rports_8_addr ? mem_29 : _GEN_1820; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1822 = 6'h1e == io_debug_rports_8_addr ? mem_30 : _GEN_1821; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1823 = 6'h1f == io_debug_rports_8_addr ? mem_31 : _GEN_1822; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1824 = 6'h20 == io_debug_rports_8_addr ? mem_32 : _GEN_1823; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1825 = 6'h21 == io_debug_rports_8_addr ? mem_33 : _GEN_1824; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1826 = 6'h22 == io_debug_rports_8_addr ? mem_34 : _GEN_1825; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1827 = 6'h23 == io_debug_rports_8_addr ? mem_35 : _GEN_1826; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1828 = 6'h24 == io_debug_rports_8_addr ? mem_36 : _GEN_1827; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1829 = 6'h25 == io_debug_rports_8_addr ? mem_37 : _GEN_1828; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1830 = 6'h26 == io_debug_rports_8_addr ? mem_38 : _GEN_1829; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1831 = 6'h27 == io_debug_rports_8_addr ? mem_39 : _GEN_1830; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1832 = 6'h28 == io_debug_rports_8_addr ? mem_40 : _GEN_1831; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1833 = 6'h29 == io_debug_rports_8_addr ? mem_41 : _GEN_1832; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1834 = 6'h2a == io_debug_rports_8_addr ? mem_42 : _GEN_1833; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1835 = 6'h2b == io_debug_rports_8_addr ? mem_43 : _GEN_1834; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1836 = 6'h2c == io_debug_rports_8_addr ? mem_44 : _GEN_1835; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1837 = 6'h2d == io_debug_rports_8_addr ? mem_45 : _GEN_1836; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1838 = 6'h2e == io_debug_rports_8_addr ? mem_46 : _GEN_1837; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1839 = 6'h2f == io_debug_rports_8_addr ? mem_47 : _GEN_1838; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1840 = 6'h30 == io_debug_rports_8_addr ? mem_48 : _GEN_1839; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1841 = 6'h31 == io_debug_rports_8_addr ? mem_49 : _GEN_1840; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1842 = 6'h32 == io_debug_rports_8_addr ? mem_50 : _GEN_1841; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1843 = 6'h33 == io_debug_rports_8_addr ? mem_51 : _GEN_1842; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1844 = 6'h34 == io_debug_rports_8_addr ? mem_52 : _GEN_1843; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1845 = 6'h35 == io_debug_rports_8_addr ? mem_53 : _GEN_1844; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1846 = 6'h36 == io_debug_rports_8_addr ? mem_54 : _GEN_1845; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1847 = 6'h37 == io_debug_rports_8_addr ? mem_55 : _GEN_1846; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1848 = 6'h38 == io_debug_rports_8_addr ? mem_56 : _GEN_1847; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1849 = 6'h39 == io_debug_rports_8_addr ? mem_57 : _GEN_1848; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1850 = 6'h3a == io_debug_rports_8_addr ? mem_58 : _GEN_1849; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1851 = 6'h3b == io_debug_rports_8_addr ? mem_59 : _GEN_1850; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1852 = 6'h3c == io_debug_rports_8_addr ? mem_60 : _GEN_1851; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1853 = 6'h3d == io_debug_rports_8_addr ? mem_61 : _GEN_1852; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1854 = 6'h3e == io_debug_rports_8_addr ? mem_62 : _GEN_1853; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1855 = 6'h3f == io_debug_rports_8_addr ? mem_63 : _GEN_1854; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1857 = 6'h1 == io_debug_rports_9_addr ? mem_1 : mem_0; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1858 = 6'h2 == io_debug_rports_9_addr ? mem_2 : _GEN_1857; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1859 = 6'h3 == io_debug_rports_9_addr ? mem_3 : _GEN_1858; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1860 = 6'h4 == io_debug_rports_9_addr ? mem_4 : _GEN_1859; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1861 = 6'h5 == io_debug_rports_9_addr ? mem_5 : _GEN_1860; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1862 = 6'h6 == io_debug_rports_9_addr ? mem_6 : _GEN_1861; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1863 = 6'h7 == io_debug_rports_9_addr ? mem_7 : _GEN_1862; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1864 = 6'h8 == io_debug_rports_9_addr ? mem_8 : _GEN_1863; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1865 = 6'h9 == io_debug_rports_9_addr ? mem_9 : _GEN_1864; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1866 = 6'ha == io_debug_rports_9_addr ? mem_10 : _GEN_1865; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1867 = 6'hb == io_debug_rports_9_addr ? mem_11 : _GEN_1866; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1868 = 6'hc == io_debug_rports_9_addr ? mem_12 : _GEN_1867; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1869 = 6'hd == io_debug_rports_9_addr ? mem_13 : _GEN_1868; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1870 = 6'he == io_debug_rports_9_addr ? mem_14 : _GEN_1869; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1871 = 6'hf == io_debug_rports_9_addr ? mem_15 : _GEN_1870; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1872 = 6'h10 == io_debug_rports_9_addr ? mem_16 : _GEN_1871; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1873 = 6'h11 == io_debug_rports_9_addr ? mem_17 : _GEN_1872; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1874 = 6'h12 == io_debug_rports_9_addr ? mem_18 : _GEN_1873; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1875 = 6'h13 == io_debug_rports_9_addr ? mem_19 : _GEN_1874; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1876 = 6'h14 == io_debug_rports_9_addr ? mem_20 : _GEN_1875; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1877 = 6'h15 == io_debug_rports_9_addr ? mem_21 : _GEN_1876; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1878 = 6'h16 == io_debug_rports_9_addr ? mem_22 : _GEN_1877; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1879 = 6'h17 == io_debug_rports_9_addr ? mem_23 : _GEN_1878; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1880 = 6'h18 == io_debug_rports_9_addr ? mem_24 : _GEN_1879; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1881 = 6'h19 == io_debug_rports_9_addr ? mem_25 : _GEN_1880; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1882 = 6'h1a == io_debug_rports_9_addr ? mem_26 : _GEN_1881; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1883 = 6'h1b == io_debug_rports_9_addr ? mem_27 : _GEN_1882; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1884 = 6'h1c == io_debug_rports_9_addr ? mem_28 : _GEN_1883; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1885 = 6'h1d == io_debug_rports_9_addr ? mem_29 : _GEN_1884; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1886 = 6'h1e == io_debug_rports_9_addr ? mem_30 : _GEN_1885; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1887 = 6'h1f == io_debug_rports_9_addr ? mem_31 : _GEN_1886; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1888 = 6'h20 == io_debug_rports_9_addr ? mem_32 : _GEN_1887; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1889 = 6'h21 == io_debug_rports_9_addr ? mem_33 : _GEN_1888; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1890 = 6'h22 == io_debug_rports_9_addr ? mem_34 : _GEN_1889; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1891 = 6'h23 == io_debug_rports_9_addr ? mem_35 : _GEN_1890; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1892 = 6'h24 == io_debug_rports_9_addr ? mem_36 : _GEN_1891; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1893 = 6'h25 == io_debug_rports_9_addr ? mem_37 : _GEN_1892; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1894 = 6'h26 == io_debug_rports_9_addr ? mem_38 : _GEN_1893; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1895 = 6'h27 == io_debug_rports_9_addr ? mem_39 : _GEN_1894; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1896 = 6'h28 == io_debug_rports_9_addr ? mem_40 : _GEN_1895; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1897 = 6'h29 == io_debug_rports_9_addr ? mem_41 : _GEN_1896; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1898 = 6'h2a == io_debug_rports_9_addr ? mem_42 : _GEN_1897; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1899 = 6'h2b == io_debug_rports_9_addr ? mem_43 : _GEN_1898; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1900 = 6'h2c == io_debug_rports_9_addr ? mem_44 : _GEN_1899; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1901 = 6'h2d == io_debug_rports_9_addr ? mem_45 : _GEN_1900; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1902 = 6'h2e == io_debug_rports_9_addr ? mem_46 : _GEN_1901; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1903 = 6'h2f == io_debug_rports_9_addr ? mem_47 : _GEN_1902; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1904 = 6'h30 == io_debug_rports_9_addr ? mem_48 : _GEN_1903; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1905 = 6'h31 == io_debug_rports_9_addr ? mem_49 : _GEN_1904; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1906 = 6'h32 == io_debug_rports_9_addr ? mem_50 : _GEN_1905; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1907 = 6'h33 == io_debug_rports_9_addr ? mem_51 : _GEN_1906; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1908 = 6'h34 == io_debug_rports_9_addr ? mem_52 : _GEN_1907; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1909 = 6'h35 == io_debug_rports_9_addr ? mem_53 : _GEN_1908; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1910 = 6'h36 == io_debug_rports_9_addr ? mem_54 : _GEN_1909; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1911 = 6'h37 == io_debug_rports_9_addr ? mem_55 : _GEN_1910; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1912 = 6'h38 == io_debug_rports_9_addr ? mem_56 : _GEN_1911; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1913 = 6'h39 == io_debug_rports_9_addr ? mem_57 : _GEN_1912; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1914 = 6'h3a == io_debug_rports_9_addr ? mem_58 : _GEN_1913; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1915 = 6'h3b == io_debug_rports_9_addr ? mem_59 : _GEN_1914; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1916 = 6'h3c == io_debug_rports_9_addr ? mem_60 : _GEN_1915; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1917 = 6'h3d == io_debug_rports_9_addr ? mem_61 : _GEN_1916; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1918 = 6'h3e == io_debug_rports_9_addr ? mem_62 : _GEN_1917; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1919 = 6'h3f == io_debug_rports_9_addr ? mem_63 : _GEN_1918; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1921 = 6'h1 == io_debug_rports_10_addr ? mem_1 : mem_0; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1922 = 6'h2 == io_debug_rports_10_addr ? mem_2 : _GEN_1921; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1923 = 6'h3 == io_debug_rports_10_addr ? mem_3 : _GEN_1922; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1924 = 6'h4 == io_debug_rports_10_addr ? mem_4 : _GEN_1923; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1925 = 6'h5 == io_debug_rports_10_addr ? mem_5 : _GEN_1924; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1926 = 6'h6 == io_debug_rports_10_addr ? mem_6 : _GEN_1925; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1927 = 6'h7 == io_debug_rports_10_addr ? mem_7 : _GEN_1926; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1928 = 6'h8 == io_debug_rports_10_addr ? mem_8 : _GEN_1927; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1929 = 6'h9 == io_debug_rports_10_addr ? mem_9 : _GEN_1928; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1930 = 6'ha == io_debug_rports_10_addr ? mem_10 : _GEN_1929; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1931 = 6'hb == io_debug_rports_10_addr ? mem_11 : _GEN_1930; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1932 = 6'hc == io_debug_rports_10_addr ? mem_12 : _GEN_1931; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1933 = 6'hd == io_debug_rports_10_addr ? mem_13 : _GEN_1932; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1934 = 6'he == io_debug_rports_10_addr ? mem_14 : _GEN_1933; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1935 = 6'hf == io_debug_rports_10_addr ? mem_15 : _GEN_1934; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1936 = 6'h10 == io_debug_rports_10_addr ? mem_16 : _GEN_1935; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1937 = 6'h11 == io_debug_rports_10_addr ? mem_17 : _GEN_1936; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1938 = 6'h12 == io_debug_rports_10_addr ? mem_18 : _GEN_1937; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1939 = 6'h13 == io_debug_rports_10_addr ? mem_19 : _GEN_1938; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1940 = 6'h14 == io_debug_rports_10_addr ? mem_20 : _GEN_1939; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1941 = 6'h15 == io_debug_rports_10_addr ? mem_21 : _GEN_1940; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1942 = 6'h16 == io_debug_rports_10_addr ? mem_22 : _GEN_1941; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1943 = 6'h17 == io_debug_rports_10_addr ? mem_23 : _GEN_1942; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1944 = 6'h18 == io_debug_rports_10_addr ? mem_24 : _GEN_1943; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1945 = 6'h19 == io_debug_rports_10_addr ? mem_25 : _GEN_1944; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1946 = 6'h1a == io_debug_rports_10_addr ? mem_26 : _GEN_1945; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1947 = 6'h1b == io_debug_rports_10_addr ? mem_27 : _GEN_1946; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1948 = 6'h1c == io_debug_rports_10_addr ? mem_28 : _GEN_1947; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1949 = 6'h1d == io_debug_rports_10_addr ? mem_29 : _GEN_1948; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1950 = 6'h1e == io_debug_rports_10_addr ? mem_30 : _GEN_1949; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1951 = 6'h1f == io_debug_rports_10_addr ? mem_31 : _GEN_1950; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1952 = 6'h20 == io_debug_rports_10_addr ? mem_32 : _GEN_1951; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1953 = 6'h21 == io_debug_rports_10_addr ? mem_33 : _GEN_1952; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1954 = 6'h22 == io_debug_rports_10_addr ? mem_34 : _GEN_1953; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1955 = 6'h23 == io_debug_rports_10_addr ? mem_35 : _GEN_1954; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1956 = 6'h24 == io_debug_rports_10_addr ? mem_36 : _GEN_1955; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1957 = 6'h25 == io_debug_rports_10_addr ? mem_37 : _GEN_1956; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1958 = 6'h26 == io_debug_rports_10_addr ? mem_38 : _GEN_1957; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1959 = 6'h27 == io_debug_rports_10_addr ? mem_39 : _GEN_1958; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1960 = 6'h28 == io_debug_rports_10_addr ? mem_40 : _GEN_1959; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1961 = 6'h29 == io_debug_rports_10_addr ? mem_41 : _GEN_1960; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1962 = 6'h2a == io_debug_rports_10_addr ? mem_42 : _GEN_1961; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1963 = 6'h2b == io_debug_rports_10_addr ? mem_43 : _GEN_1962; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1964 = 6'h2c == io_debug_rports_10_addr ? mem_44 : _GEN_1963; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1965 = 6'h2d == io_debug_rports_10_addr ? mem_45 : _GEN_1964; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1966 = 6'h2e == io_debug_rports_10_addr ? mem_46 : _GEN_1965; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1967 = 6'h2f == io_debug_rports_10_addr ? mem_47 : _GEN_1966; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1968 = 6'h30 == io_debug_rports_10_addr ? mem_48 : _GEN_1967; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1969 = 6'h31 == io_debug_rports_10_addr ? mem_49 : _GEN_1968; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1970 = 6'h32 == io_debug_rports_10_addr ? mem_50 : _GEN_1969; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1971 = 6'h33 == io_debug_rports_10_addr ? mem_51 : _GEN_1970; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1972 = 6'h34 == io_debug_rports_10_addr ? mem_52 : _GEN_1971; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1973 = 6'h35 == io_debug_rports_10_addr ? mem_53 : _GEN_1972; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1974 = 6'h36 == io_debug_rports_10_addr ? mem_54 : _GEN_1973; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1975 = 6'h37 == io_debug_rports_10_addr ? mem_55 : _GEN_1974; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1976 = 6'h38 == io_debug_rports_10_addr ? mem_56 : _GEN_1975; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1977 = 6'h39 == io_debug_rports_10_addr ? mem_57 : _GEN_1976; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1978 = 6'h3a == io_debug_rports_10_addr ? mem_58 : _GEN_1977; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1979 = 6'h3b == io_debug_rports_10_addr ? mem_59 : _GEN_1978; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1980 = 6'h3c == io_debug_rports_10_addr ? mem_60 : _GEN_1979; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1981 = 6'h3d == io_debug_rports_10_addr ? mem_61 : _GEN_1980; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1982 = 6'h3e == io_debug_rports_10_addr ? mem_62 : _GEN_1981; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1983 = 6'h3f == io_debug_rports_10_addr ? mem_63 : _GEN_1982; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1985 = 6'h1 == io_debug_rports_11_addr ? mem_1 : mem_0; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1986 = 6'h2 == io_debug_rports_11_addr ? mem_2 : _GEN_1985; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1987 = 6'h3 == io_debug_rports_11_addr ? mem_3 : _GEN_1986; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1988 = 6'h4 == io_debug_rports_11_addr ? mem_4 : _GEN_1987; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1989 = 6'h5 == io_debug_rports_11_addr ? mem_5 : _GEN_1988; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1990 = 6'h6 == io_debug_rports_11_addr ? mem_6 : _GEN_1989; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1991 = 6'h7 == io_debug_rports_11_addr ? mem_7 : _GEN_1990; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1992 = 6'h8 == io_debug_rports_11_addr ? mem_8 : _GEN_1991; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1993 = 6'h9 == io_debug_rports_11_addr ? mem_9 : _GEN_1992; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1994 = 6'ha == io_debug_rports_11_addr ? mem_10 : _GEN_1993; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1995 = 6'hb == io_debug_rports_11_addr ? mem_11 : _GEN_1994; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1996 = 6'hc == io_debug_rports_11_addr ? mem_12 : _GEN_1995; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1997 = 6'hd == io_debug_rports_11_addr ? mem_13 : _GEN_1996; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1998 = 6'he == io_debug_rports_11_addr ? mem_14 : _GEN_1997; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_1999 = 6'hf == io_debug_rports_11_addr ? mem_15 : _GEN_1998; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2000 = 6'h10 == io_debug_rports_11_addr ? mem_16 : _GEN_1999; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2001 = 6'h11 == io_debug_rports_11_addr ? mem_17 : _GEN_2000; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2002 = 6'h12 == io_debug_rports_11_addr ? mem_18 : _GEN_2001; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2003 = 6'h13 == io_debug_rports_11_addr ? mem_19 : _GEN_2002; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2004 = 6'h14 == io_debug_rports_11_addr ? mem_20 : _GEN_2003; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2005 = 6'h15 == io_debug_rports_11_addr ? mem_21 : _GEN_2004; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2006 = 6'h16 == io_debug_rports_11_addr ? mem_22 : _GEN_2005; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2007 = 6'h17 == io_debug_rports_11_addr ? mem_23 : _GEN_2006; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2008 = 6'h18 == io_debug_rports_11_addr ? mem_24 : _GEN_2007; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2009 = 6'h19 == io_debug_rports_11_addr ? mem_25 : _GEN_2008; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2010 = 6'h1a == io_debug_rports_11_addr ? mem_26 : _GEN_2009; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2011 = 6'h1b == io_debug_rports_11_addr ? mem_27 : _GEN_2010; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2012 = 6'h1c == io_debug_rports_11_addr ? mem_28 : _GEN_2011; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2013 = 6'h1d == io_debug_rports_11_addr ? mem_29 : _GEN_2012; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2014 = 6'h1e == io_debug_rports_11_addr ? mem_30 : _GEN_2013; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2015 = 6'h1f == io_debug_rports_11_addr ? mem_31 : _GEN_2014; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2016 = 6'h20 == io_debug_rports_11_addr ? mem_32 : _GEN_2015; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2017 = 6'h21 == io_debug_rports_11_addr ? mem_33 : _GEN_2016; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2018 = 6'h22 == io_debug_rports_11_addr ? mem_34 : _GEN_2017; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2019 = 6'h23 == io_debug_rports_11_addr ? mem_35 : _GEN_2018; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2020 = 6'h24 == io_debug_rports_11_addr ? mem_36 : _GEN_2019; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2021 = 6'h25 == io_debug_rports_11_addr ? mem_37 : _GEN_2020; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2022 = 6'h26 == io_debug_rports_11_addr ? mem_38 : _GEN_2021; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2023 = 6'h27 == io_debug_rports_11_addr ? mem_39 : _GEN_2022; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2024 = 6'h28 == io_debug_rports_11_addr ? mem_40 : _GEN_2023; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2025 = 6'h29 == io_debug_rports_11_addr ? mem_41 : _GEN_2024; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2026 = 6'h2a == io_debug_rports_11_addr ? mem_42 : _GEN_2025; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2027 = 6'h2b == io_debug_rports_11_addr ? mem_43 : _GEN_2026; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2028 = 6'h2c == io_debug_rports_11_addr ? mem_44 : _GEN_2027; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2029 = 6'h2d == io_debug_rports_11_addr ? mem_45 : _GEN_2028; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2030 = 6'h2e == io_debug_rports_11_addr ? mem_46 : _GEN_2029; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2031 = 6'h2f == io_debug_rports_11_addr ? mem_47 : _GEN_2030; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2032 = 6'h30 == io_debug_rports_11_addr ? mem_48 : _GEN_2031; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2033 = 6'h31 == io_debug_rports_11_addr ? mem_49 : _GEN_2032; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2034 = 6'h32 == io_debug_rports_11_addr ? mem_50 : _GEN_2033; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2035 = 6'h33 == io_debug_rports_11_addr ? mem_51 : _GEN_2034; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2036 = 6'h34 == io_debug_rports_11_addr ? mem_52 : _GEN_2035; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2037 = 6'h35 == io_debug_rports_11_addr ? mem_53 : _GEN_2036; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2038 = 6'h36 == io_debug_rports_11_addr ? mem_54 : _GEN_2037; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2039 = 6'h37 == io_debug_rports_11_addr ? mem_55 : _GEN_2038; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2040 = 6'h38 == io_debug_rports_11_addr ? mem_56 : _GEN_2039; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2041 = 6'h39 == io_debug_rports_11_addr ? mem_57 : _GEN_2040; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2042 = 6'h3a == io_debug_rports_11_addr ? mem_58 : _GEN_2041; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2043 = 6'h3b == io_debug_rports_11_addr ? mem_59 : _GEN_2042; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2044 = 6'h3c == io_debug_rports_11_addr ? mem_60 : _GEN_2043; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2045 = 6'h3d == io_debug_rports_11_addr ? mem_61 : _GEN_2044; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2046 = 6'h3e == io_debug_rports_11_addr ? mem_62 : _GEN_2045; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2047 = 6'h3f == io_debug_rports_11_addr ? mem_63 : _GEN_2046; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2049 = 6'h1 == io_debug_rports_12_addr ? mem_1 : mem_0; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2050 = 6'h2 == io_debug_rports_12_addr ? mem_2 : _GEN_2049; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2051 = 6'h3 == io_debug_rports_12_addr ? mem_3 : _GEN_2050; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2052 = 6'h4 == io_debug_rports_12_addr ? mem_4 : _GEN_2051; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2053 = 6'h5 == io_debug_rports_12_addr ? mem_5 : _GEN_2052; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2054 = 6'h6 == io_debug_rports_12_addr ? mem_6 : _GEN_2053; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2055 = 6'h7 == io_debug_rports_12_addr ? mem_7 : _GEN_2054; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2056 = 6'h8 == io_debug_rports_12_addr ? mem_8 : _GEN_2055; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2057 = 6'h9 == io_debug_rports_12_addr ? mem_9 : _GEN_2056; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2058 = 6'ha == io_debug_rports_12_addr ? mem_10 : _GEN_2057; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2059 = 6'hb == io_debug_rports_12_addr ? mem_11 : _GEN_2058; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2060 = 6'hc == io_debug_rports_12_addr ? mem_12 : _GEN_2059; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2061 = 6'hd == io_debug_rports_12_addr ? mem_13 : _GEN_2060; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2062 = 6'he == io_debug_rports_12_addr ? mem_14 : _GEN_2061; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2063 = 6'hf == io_debug_rports_12_addr ? mem_15 : _GEN_2062; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2064 = 6'h10 == io_debug_rports_12_addr ? mem_16 : _GEN_2063; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2065 = 6'h11 == io_debug_rports_12_addr ? mem_17 : _GEN_2064; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2066 = 6'h12 == io_debug_rports_12_addr ? mem_18 : _GEN_2065; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2067 = 6'h13 == io_debug_rports_12_addr ? mem_19 : _GEN_2066; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2068 = 6'h14 == io_debug_rports_12_addr ? mem_20 : _GEN_2067; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2069 = 6'h15 == io_debug_rports_12_addr ? mem_21 : _GEN_2068; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2070 = 6'h16 == io_debug_rports_12_addr ? mem_22 : _GEN_2069; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2071 = 6'h17 == io_debug_rports_12_addr ? mem_23 : _GEN_2070; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2072 = 6'h18 == io_debug_rports_12_addr ? mem_24 : _GEN_2071; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2073 = 6'h19 == io_debug_rports_12_addr ? mem_25 : _GEN_2072; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2074 = 6'h1a == io_debug_rports_12_addr ? mem_26 : _GEN_2073; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2075 = 6'h1b == io_debug_rports_12_addr ? mem_27 : _GEN_2074; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2076 = 6'h1c == io_debug_rports_12_addr ? mem_28 : _GEN_2075; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2077 = 6'h1d == io_debug_rports_12_addr ? mem_29 : _GEN_2076; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2078 = 6'h1e == io_debug_rports_12_addr ? mem_30 : _GEN_2077; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2079 = 6'h1f == io_debug_rports_12_addr ? mem_31 : _GEN_2078; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2080 = 6'h20 == io_debug_rports_12_addr ? mem_32 : _GEN_2079; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2081 = 6'h21 == io_debug_rports_12_addr ? mem_33 : _GEN_2080; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2082 = 6'h22 == io_debug_rports_12_addr ? mem_34 : _GEN_2081; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2083 = 6'h23 == io_debug_rports_12_addr ? mem_35 : _GEN_2082; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2084 = 6'h24 == io_debug_rports_12_addr ? mem_36 : _GEN_2083; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2085 = 6'h25 == io_debug_rports_12_addr ? mem_37 : _GEN_2084; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2086 = 6'h26 == io_debug_rports_12_addr ? mem_38 : _GEN_2085; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2087 = 6'h27 == io_debug_rports_12_addr ? mem_39 : _GEN_2086; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2088 = 6'h28 == io_debug_rports_12_addr ? mem_40 : _GEN_2087; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2089 = 6'h29 == io_debug_rports_12_addr ? mem_41 : _GEN_2088; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2090 = 6'h2a == io_debug_rports_12_addr ? mem_42 : _GEN_2089; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2091 = 6'h2b == io_debug_rports_12_addr ? mem_43 : _GEN_2090; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2092 = 6'h2c == io_debug_rports_12_addr ? mem_44 : _GEN_2091; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2093 = 6'h2d == io_debug_rports_12_addr ? mem_45 : _GEN_2092; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2094 = 6'h2e == io_debug_rports_12_addr ? mem_46 : _GEN_2093; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2095 = 6'h2f == io_debug_rports_12_addr ? mem_47 : _GEN_2094; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2096 = 6'h30 == io_debug_rports_12_addr ? mem_48 : _GEN_2095; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2097 = 6'h31 == io_debug_rports_12_addr ? mem_49 : _GEN_2096; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2098 = 6'h32 == io_debug_rports_12_addr ? mem_50 : _GEN_2097; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2099 = 6'h33 == io_debug_rports_12_addr ? mem_51 : _GEN_2098; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2100 = 6'h34 == io_debug_rports_12_addr ? mem_52 : _GEN_2099; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2101 = 6'h35 == io_debug_rports_12_addr ? mem_53 : _GEN_2100; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2102 = 6'h36 == io_debug_rports_12_addr ? mem_54 : _GEN_2101; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2103 = 6'h37 == io_debug_rports_12_addr ? mem_55 : _GEN_2102; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2104 = 6'h38 == io_debug_rports_12_addr ? mem_56 : _GEN_2103; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2105 = 6'h39 == io_debug_rports_12_addr ? mem_57 : _GEN_2104; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2106 = 6'h3a == io_debug_rports_12_addr ? mem_58 : _GEN_2105; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2107 = 6'h3b == io_debug_rports_12_addr ? mem_59 : _GEN_2106; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2108 = 6'h3c == io_debug_rports_12_addr ? mem_60 : _GEN_2107; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2109 = 6'h3d == io_debug_rports_12_addr ? mem_61 : _GEN_2108; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2110 = 6'h3e == io_debug_rports_12_addr ? mem_62 : _GEN_2109; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2111 = 6'h3f == io_debug_rports_12_addr ? mem_63 : _GEN_2110; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2113 = 6'h1 == io_debug_rports_13_addr ? mem_1 : mem_0; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2114 = 6'h2 == io_debug_rports_13_addr ? mem_2 : _GEN_2113; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2115 = 6'h3 == io_debug_rports_13_addr ? mem_3 : _GEN_2114; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2116 = 6'h4 == io_debug_rports_13_addr ? mem_4 : _GEN_2115; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2117 = 6'h5 == io_debug_rports_13_addr ? mem_5 : _GEN_2116; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2118 = 6'h6 == io_debug_rports_13_addr ? mem_6 : _GEN_2117; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2119 = 6'h7 == io_debug_rports_13_addr ? mem_7 : _GEN_2118; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2120 = 6'h8 == io_debug_rports_13_addr ? mem_8 : _GEN_2119; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2121 = 6'h9 == io_debug_rports_13_addr ? mem_9 : _GEN_2120; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2122 = 6'ha == io_debug_rports_13_addr ? mem_10 : _GEN_2121; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2123 = 6'hb == io_debug_rports_13_addr ? mem_11 : _GEN_2122; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2124 = 6'hc == io_debug_rports_13_addr ? mem_12 : _GEN_2123; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2125 = 6'hd == io_debug_rports_13_addr ? mem_13 : _GEN_2124; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2126 = 6'he == io_debug_rports_13_addr ? mem_14 : _GEN_2125; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2127 = 6'hf == io_debug_rports_13_addr ? mem_15 : _GEN_2126; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2128 = 6'h10 == io_debug_rports_13_addr ? mem_16 : _GEN_2127; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2129 = 6'h11 == io_debug_rports_13_addr ? mem_17 : _GEN_2128; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2130 = 6'h12 == io_debug_rports_13_addr ? mem_18 : _GEN_2129; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2131 = 6'h13 == io_debug_rports_13_addr ? mem_19 : _GEN_2130; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2132 = 6'h14 == io_debug_rports_13_addr ? mem_20 : _GEN_2131; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2133 = 6'h15 == io_debug_rports_13_addr ? mem_21 : _GEN_2132; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2134 = 6'h16 == io_debug_rports_13_addr ? mem_22 : _GEN_2133; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2135 = 6'h17 == io_debug_rports_13_addr ? mem_23 : _GEN_2134; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2136 = 6'h18 == io_debug_rports_13_addr ? mem_24 : _GEN_2135; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2137 = 6'h19 == io_debug_rports_13_addr ? mem_25 : _GEN_2136; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2138 = 6'h1a == io_debug_rports_13_addr ? mem_26 : _GEN_2137; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2139 = 6'h1b == io_debug_rports_13_addr ? mem_27 : _GEN_2138; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2140 = 6'h1c == io_debug_rports_13_addr ? mem_28 : _GEN_2139; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2141 = 6'h1d == io_debug_rports_13_addr ? mem_29 : _GEN_2140; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2142 = 6'h1e == io_debug_rports_13_addr ? mem_30 : _GEN_2141; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2143 = 6'h1f == io_debug_rports_13_addr ? mem_31 : _GEN_2142; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2144 = 6'h20 == io_debug_rports_13_addr ? mem_32 : _GEN_2143; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2145 = 6'h21 == io_debug_rports_13_addr ? mem_33 : _GEN_2144; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2146 = 6'h22 == io_debug_rports_13_addr ? mem_34 : _GEN_2145; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2147 = 6'h23 == io_debug_rports_13_addr ? mem_35 : _GEN_2146; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2148 = 6'h24 == io_debug_rports_13_addr ? mem_36 : _GEN_2147; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2149 = 6'h25 == io_debug_rports_13_addr ? mem_37 : _GEN_2148; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2150 = 6'h26 == io_debug_rports_13_addr ? mem_38 : _GEN_2149; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2151 = 6'h27 == io_debug_rports_13_addr ? mem_39 : _GEN_2150; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2152 = 6'h28 == io_debug_rports_13_addr ? mem_40 : _GEN_2151; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2153 = 6'h29 == io_debug_rports_13_addr ? mem_41 : _GEN_2152; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2154 = 6'h2a == io_debug_rports_13_addr ? mem_42 : _GEN_2153; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2155 = 6'h2b == io_debug_rports_13_addr ? mem_43 : _GEN_2154; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2156 = 6'h2c == io_debug_rports_13_addr ? mem_44 : _GEN_2155; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2157 = 6'h2d == io_debug_rports_13_addr ? mem_45 : _GEN_2156; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2158 = 6'h2e == io_debug_rports_13_addr ? mem_46 : _GEN_2157; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2159 = 6'h2f == io_debug_rports_13_addr ? mem_47 : _GEN_2158; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2160 = 6'h30 == io_debug_rports_13_addr ? mem_48 : _GEN_2159; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2161 = 6'h31 == io_debug_rports_13_addr ? mem_49 : _GEN_2160; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2162 = 6'h32 == io_debug_rports_13_addr ? mem_50 : _GEN_2161; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2163 = 6'h33 == io_debug_rports_13_addr ? mem_51 : _GEN_2162; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2164 = 6'h34 == io_debug_rports_13_addr ? mem_52 : _GEN_2163; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2165 = 6'h35 == io_debug_rports_13_addr ? mem_53 : _GEN_2164; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2166 = 6'h36 == io_debug_rports_13_addr ? mem_54 : _GEN_2165; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2167 = 6'h37 == io_debug_rports_13_addr ? mem_55 : _GEN_2166; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2168 = 6'h38 == io_debug_rports_13_addr ? mem_56 : _GEN_2167; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2169 = 6'h39 == io_debug_rports_13_addr ? mem_57 : _GEN_2168; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2170 = 6'h3a == io_debug_rports_13_addr ? mem_58 : _GEN_2169; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2171 = 6'h3b == io_debug_rports_13_addr ? mem_59 : _GEN_2170; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2172 = 6'h3c == io_debug_rports_13_addr ? mem_60 : _GEN_2171; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2173 = 6'h3d == io_debug_rports_13_addr ? mem_61 : _GEN_2172; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2174 = 6'h3e == io_debug_rports_13_addr ? mem_62 : _GEN_2173; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2175 = 6'h3f == io_debug_rports_13_addr ? mem_63 : _GEN_2174; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2177 = 6'h1 == io_debug_rports_14_addr ? mem_1 : mem_0; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2178 = 6'h2 == io_debug_rports_14_addr ? mem_2 : _GEN_2177; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2179 = 6'h3 == io_debug_rports_14_addr ? mem_3 : _GEN_2178; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2180 = 6'h4 == io_debug_rports_14_addr ? mem_4 : _GEN_2179; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2181 = 6'h5 == io_debug_rports_14_addr ? mem_5 : _GEN_2180; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2182 = 6'h6 == io_debug_rports_14_addr ? mem_6 : _GEN_2181; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2183 = 6'h7 == io_debug_rports_14_addr ? mem_7 : _GEN_2182; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2184 = 6'h8 == io_debug_rports_14_addr ? mem_8 : _GEN_2183; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2185 = 6'h9 == io_debug_rports_14_addr ? mem_9 : _GEN_2184; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2186 = 6'ha == io_debug_rports_14_addr ? mem_10 : _GEN_2185; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2187 = 6'hb == io_debug_rports_14_addr ? mem_11 : _GEN_2186; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2188 = 6'hc == io_debug_rports_14_addr ? mem_12 : _GEN_2187; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2189 = 6'hd == io_debug_rports_14_addr ? mem_13 : _GEN_2188; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2190 = 6'he == io_debug_rports_14_addr ? mem_14 : _GEN_2189; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2191 = 6'hf == io_debug_rports_14_addr ? mem_15 : _GEN_2190; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2192 = 6'h10 == io_debug_rports_14_addr ? mem_16 : _GEN_2191; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2193 = 6'h11 == io_debug_rports_14_addr ? mem_17 : _GEN_2192; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2194 = 6'h12 == io_debug_rports_14_addr ? mem_18 : _GEN_2193; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2195 = 6'h13 == io_debug_rports_14_addr ? mem_19 : _GEN_2194; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2196 = 6'h14 == io_debug_rports_14_addr ? mem_20 : _GEN_2195; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2197 = 6'h15 == io_debug_rports_14_addr ? mem_21 : _GEN_2196; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2198 = 6'h16 == io_debug_rports_14_addr ? mem_22 : _GEN_2197; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2199 = 6'h17 == io_debug_rports_14_addr ? mem_23 : _GEN_2198; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2200 = 6'h18 == io_debug_rports_14_addr ? mem_24 : _GEN_2199; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2201 = 6'h19 == io_debug_rports_14_addr ? mem_25 : _GEN_2200; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2202 = 6'h1a == io_debug_rports_14_addr ? mem_26 : _GEN_2201; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2203 = 6'h1b == io_debug_rports_14_addr ? mem_27 : _GEN_2202; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2204 = 6'h1c == io_debug_rports_14_addr ? mem_28 : _GEN_2203; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2205 = 6'h1d == io_debug_rports_14_addr ? mem_29 : _GEN_2204; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2206 = 6'h1e == io_debug_rports_14_addr ? mem_30 : _GEN_2205; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2207 = 6'h1f == io_debug_rports_14_addr ? mem_31 : _GEN_2206; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2208 = 6'h20 == io_debug_rports_14_addr ? mem_32 : _GEN_2207; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2209 = 6'h21 == io_debug_rports_14_addr ? mem_33 : _GEN_2208; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2210 = 6'h22 == io_debug_rports_14_addr ? mem_34 : _GEN_2209; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2211 = 6'h23 == io_debug_rports_14_addr ? mem_35 : _GEN_2210; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2212 = 6'h24 == io_debug_rports_14_addr ? mem_36 : _GEN_2211; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2213 = 6'h25 == io_debug_rports_14_addr ? mem_37 : _GEN_2212; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2214 = 6'h26 == io_debug_rports_14_addr ? mem_38 : _GEN_2213; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2215 = 6'h27 == io_debug_rports_14_addr ? mem_39 : _GEN_2214; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2216 = 6'h28 == io_debug_rports_14_addr ? mem_40 : _GEN_2215; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2217 = 6'h29 == io_debug_rports_14_addr ? mem_41 : _GEN_2216; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2218 = 6'h2a == io_debug_rports_14_addr ? mem_42 : _GEN_2217; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2219 = 6'h2b == io_debug_rports_14_addr ? mem_43 : _GEN_2218; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2220 = 6'h2c == io_debug_rports_14_addr ? mem_44 : _GEN_2219; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2221 = 6'h2d == io_debug_rports_14_addr ? mem_45 : _GEN_2220; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2222 = 6'h2e == io_debug_rports_14_addr ? mem_46 : _GEN_2221; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2223 = 6'h2f == io_debug_rports_14_addr ? mem_47 : _GEN_2222; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2224 = 6'h30 == io_debug_rports_14_addr ? mem_48 : _GEN_2223; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2225 = 6'h31 == io_debug_rports_14_addr ? mem_49 : _GEN_2224; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2226 = 6'h32 == io_debug_rports_14_addr ? mem_50 : _GEN_2225; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2227 = 6'h33 == io_debug_rports_14_addr ? mem_51 : _GEN_2226; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2228 = 6'h34 == io_debug_rports_14_addr ? mem_52 : _GEN_2227; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2229 = 6'h35 == io_debug_rports_14_addr ? mem_53 : _GEN_2228; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2230 = 6'h36 == io_debug_rports_14_addr ? mem_54 : _GEN_2229; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2231 = 6'h37 == io_debug_rports_14_addr ? mem_55 : _GEN_2230; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2232 = 6'h38 == io_debug_rports_14_addr ? mem_56 : _GEN_2231; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2233 = 6'h39 == io_debug_rports_14_addr ? mem_57 : _GEN_2232; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2234 = 6'h3a == io_debug_rports_14_addr ? mem_58 : _GEN_2233; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2235 = 6'h3b == io_debug_rports_14_addr ? mem_59 : _GEN_2234; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2236 = 6'h3c == io_debug_rports_14_addr ? mem_60 : _GEN_2235; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2237 = 6'h3d == io_debug_rports_14_addr ? mem_61 : _GEN_2236; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2238 = 6'h3e == io_debug_rports_14_addr ? mem_62 : _GEN_2237; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2239 = 6'h3f == io_debug_rports_14_addr ? mem_63 : _GEN_2238; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2241 = 6'h1 == io_debug_rports_15_addr ? mem_1 : mem_0; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2242 = 6'h2 == io_debug_rports_15_addr ? mem_2 : _GEN_2241; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2243 = 6'h3 == io_debug_rports_15_addr ? mem_3 : _GEN_2242; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2244 = 6'h4 == io_debug_rports_15_addr ? mem_4 : _GEN_2243; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2245 = 6'h5 == io_debug_rports_15_addr ? mem_5 : _GEN_2244; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2246 = 6'h6 == io_debug_rports_15_addr ? mem_6 : _GEN_2245; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2247 = 6'h7 == io_debug_rports_15_addr ? mem_7 : _GEN_2246; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2248 = 6'h8 == io_debug_rports_15_addr ? mem_8 : _GEN_2247; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2249 = 6'h9 == io_debug_rports_15_addr ? mem_9 : _GEN_2248; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2250 = 6'ha == io_debug_rports_15_addr ? mem_10 : _GEN_2249; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2251 = 6'hb == io_debug_rports_15_addr ? mem_11 : _GEN_2250; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2252 = 6'hc == io_debug_rports_15_addr ? mem_12 : _GEN_2251; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2253 = 6'hd == io_debug_rports_15_addr ? mem_13 : _GEN_2252; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2254 = 6'he == io_debug_rports_15_addr ? mem_14 : _GEN_2253; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2255 = 6'hf == io_debug_rports_15_addr ? mem_15 : _GEN_2254; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2256 = 6'h10 == io_debug_rports_15_addr ? mem_16 : _GEN_2255; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2257 = 6'h11 == io_debug_rports_15_addr ? mem_17 : _GEN_2256; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2258 = 6'h12 == io_debug_rports_15_addr ? mem_18 : _GEN_2257; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2259 = 6'h13 == io_debug_rports_15_addr ? mem_19 : _GEN_2258; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2260 = 6'h14 == io_debug_rports_15_addr ? mem_20 : _GEN_2259; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2261 = 6'h15 == io_debug_rports_15_addr ? mem_21 : _GEN_2260; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2262 = 6'h16 == io_debug_rports_15_addr ? mem_22 : _GEN_2261; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2263 = 6'h17 == io_debug_rports_15_addr ? mem_23 : _GEN_2262; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2264 = 6'h18 == io_debug_rports_15_addr ? mem_24 : _GEN_2263; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2265 = 6'h19 == io_debug_rports_15_addr ? mem_25 : _GEN_2264; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2266 = 6'h1a == io_debug_rports_15_addr ? mem_26 : _GEN_2265; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2267 = 6'h1b == io_debug_rports_15_addr ? mem_27 : _GEN_2266; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2268 = 6'h1c == io_debug_rports_15_addr ? mem_28 : _GEN_2267; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2269 = 6'h1d == io_debug_rports_15_addr ? mem_29 : _GEN_2268; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2270 = 6'h1e == io_debug_rports_15_addr ? mem_30 : _GEN_2269; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2271 = 6'h1f == io_debug_rports_15_addr ? mem_31 : _GEN_2270; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2272 = 6'h20 == io_debug_rports_15_addr ? mem_32 : _GEN_2271; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2273 = 6'h21 == io_debug_rports_15_addr ? mem_33 : _GEN_2272; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2274 = 6'h22 == io_debug_rports_15_addr ? mem_34 : _GEN_2273; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2275 = 6'h23 == io_debug_rports_15_addr ? mem_35 : _GEN_2274; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2276 = 6'h24 == io_debug_rports_15_addr ? mem_36 : _GEN_2275; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2277 = 6'h25 == io_debug_rports_15_addr ? mem_37 : _GEN_2276; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2278 = 6'h26 == io_debug_rports_15_addr ? mem_38 : _GEN_2277; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2279 = 6'h27 == io_debug_rports_15_addr ? mem_39 : _GEN_2278; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2280 = 6'h28 == io_debug_rports_15_addr ? mem_40 : _GEN_2279; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2281 = 6'h29 == io_debug_rports_15_addr ? mem_41 : _GEN_2280; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2282 = 6'h2a == io_debug_rports_15_addr ? mem_42 : _GEN_2281; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2283 = 6'h2b == io_debug_rports_15_addr ? mem_43 : _GEN_2282; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2284 = 6'h2c == io_debug_rports_15_addr ? mem_44 : _GEN_2283; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2285 = 6'h2d == io_debug_rports_15_addr ? mem_45 : _GEN_2284; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2286 = 6'h2e == io_debug_rports_15_addr ? mem_46 : _GEN_2285; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2287 = 6'h2f == io_debug_rports_15_addr ? mem_47 : _GEN_2286; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2288 = 6'h30 == io_debug_rports_15_addr ? mem_48 : _GEN_2287; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2289 = 6'h31 == io_debug_rports_15_addr ? mem_49 : _GEN_2288; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2290 = 6'h32 == io_debug_rports_15_addr ? mem_50 : _GEN_2289; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2291 = 6'h33 == io_debug_rports_15_addr ? mem_51 : _GEN_2290; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2292 = 6'h34 == io_debug_rports_15_addr ? mem_52 : _GEN_2291; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2293 = 6'h35 == io_debug_rports_15_addr ? mem_53 : _GEN_2292; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2294 = 6'h36 == io_debug_rports_15_addr ? mem_54 : _GEN_2293; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2295 = 6'h37 == io_debug_rports_15_addr ? mem_55 : _GEN_2294; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2296 = 6'h38 == io_debug_rports_15_addr ? mem_56 : _GEN_2295; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2297 = 6'h39 == io_debug_rports_15_addr ? mem_57 : _GEN_2296; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2298 = 6'h3a == io_debug_rports_15_addr ? mem_58 : _GEN_2297; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2299 = 6'h3b == io_debug_rports_15_addr ? mem_59 : _GEN_2298; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2300 = 6'h3c == io_debug_rports_15_addr ? mem_60 : _GEN_2299; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2301 = 6'h3d == io_debug_rports_15_addr ? mem_61 : _GEN_2300; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2302 = 6'h3e == io_debug_rports_15_addr ? mem_62 : _GEN_2301; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2303 = 6'h3f == io_debug_rports_15_addr ? mem_63 : _GEN_2302; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2305 = 6'h1 == io_debug_rports_16_addr ? mem_1 : mem_0; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2306 = 6'h2 == io_debug_rports_16_addr ? mem_2 : _GEN_2305; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2307 = 6'h3 == io_debug_rports_16_addr ? mem_3 : _GEN_2306; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2308 = 6'h4 == io_debug_rports_16_addr ? mem_4 : _GEN_2307; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2309 = 6'h5 == io_debug_rports_16_addr ? mem_5 : _GEN_2308; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2310 = 6'h6 == io_debug_rports_16_addr ? mem_6 : _GEN_2309; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2311 = 6'h7 == io_debug_rports_16_addr ? mem_7 : _GEN_2310; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2312 = 6'h8 == io_debug_rports_16_addr ? mem_8 : _GEN_2311; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2313 = 6'h9 == io_debug_rports_16_addr ? mem_9 : _GEN_2312; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2314 = 6'ha == io_debug_rports_16_addr ? mem_10 : _GEN_2313; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2315 = 6'hb == io_debug_rports_16_addr ? mem_11 : _GEN_2314; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2316 = 6'hc == io_debug_rports_16_addr ? mem_12 : _GEN_2315; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2317 = 6'hd == io_debug_rports_16_addr ? mem_13 : _GEN_2316; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2318 = 6'he == io_debug_rports_16_addr ? mem_14 : _GEN_2317; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2319 = 6'hf == io_debug_rports_16_addr ? mem_15 : _GEN_2318; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2320 = 6'h10 == io_debug_rports_16_addr ? mem_16 : _GEN_2319; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2321 = 6'h11 == io_debug_rports_16_addr ? mem_17 : _GEN_2320; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2322 = 6'h12 == io_debug_rports_16_addr ? mem_18 : _GEN_2321; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2323 = 6'h13 == io_debug_rports_16_addr ? mem_19 : _GEN_2322; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2324 = 6'h14 == io_debug_rports_16_addr ? mem_20 : _GEN_2323; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2325 = 6'h15 == io_debug_rports_16_addr ? mem_21 : _GEN_2324; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2326 = 6'h16 == io_debug_rports_16_addr ? mem_22 : _GEN_2325; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2327 = 6'h17 == io_debug_rports_16_addr ? mem_23 : _GEN_2326; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2328 = 6'h18 == io_debug_rports_16_addr ? mem_24 : _GEN_2327; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2329 = 6'h19 == io_debug_rports_16_addr ? mem_25 : _GEN_2328; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2330 = 6'h1a == io_debug_rports_16_addr ? mem_26 : _GEN_2329; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2331 = 6'h1b == io_debug_rports_16_addr ? mem_27 : _GEN_2330; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2332 = 6'h1c == io_debug_rports_16_addr ? mem_28 : _GEN_2331; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2333 = 6'h1d == io_debug_rports_16_addr ? mem_29 : _GEN_2332; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2334 = 6'h1e == io_debug_rports_16_addr ? mem_30 : _GEN_2333; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2335 = 6'h1f == io_debug_rports_16_addr ? mem_31 : _GEN_2334; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2336 = 6'h20 == io_debug_rports_16_addr ? mem_32 : _GEN_2335; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2337 = 6'h21 == io_debug_rports_16_addr ? mem_33 : _GEN_2336; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2338 = 6'h22 == io_debug_rports_16_addr ? mem_34 : _GEN_2337; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2339 = 6'h23 == io_debug_rports_16_addr ? mem_35 : _GEN_2338; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2340 = 6'h24 == io_debug_rports_16_addr ? mem_36 : _GEN_2339; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2341 = 6'h25 == io_debug_rports_16_addr ? mem_37 : _GEN_2340; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2342 = 6'h26 == io_debug_rports_16_addr ? mem_38 : _GEN_2341; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2343 = 6'h27 == io_debug_rports_16_addr ? mem_39 : _GEN_2342; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2344 = 6'h28 == io_debug_rports_16_addr ? mem_40 : _GEN_2343; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2345 = 6'h29 == io_debug_rports_16_addr ? mem_41 : _GEN_2344; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2346 = 6'h2a == io_debug_rports_16_addr ? mem_42 : _GEN_2345; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2347 = 6'h2b == io_debug_rports_16_addr ? mem_43 : _GEN_2346; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2348 = 6'h2c == io_debug_rports_16_addr ? mem_44 : _GEN_2347; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2349 = 6'h2d == io_debug_rports_16_addr ? mem_45 : _GEN_2348; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2350 = 6'h2e == io_debug_rports_16_addr ? mem_46 : _GEN_2349; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2351 = 6'h2f == io_debug_rports_16_addr ? mem_47 : _GEN_2350; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2352 = 6'h30 == io_debug_rports_16_addr ? mem_48 : _GEN_2351; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2353 = 6'h31 == io_debug_rports_16_addr ? mem_49 : _GEN_2352; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2354 = 6'h32 == io_debug_rports_16_addr ? mem_50 : _GEN_2353; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2355 = 6'h33 == io_debug_rports_16_addr ? mem_51 : _GEN_2354; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2356 = 6'h34 == io_debug_rports_16_addr ? mem_52 : _GEN_2355; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2357 = 6'h35 == io_debug_rports_16_addr ? mem_53 : _GEN_2356; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2358 = 6'h36 == io_debug_rports_16_addr ? mem_54 : _GEN_2357; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2359 = 6'h37 == io_debug_rports_16_addr ? mem_55 : _GEN_2358; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2360 = 6'h38 == io_debug_rports_16_addr ? mem_56 : _GEN_2359; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2361 = 6'h39 == io_debug_rports_16_addr ? mem_57 : _GEN_2360; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2362 = 6'h3a == io_debug_rports_16_addr ? mem_58 : _GEN_2361; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2363 = 6'h3b == io_debug_rports_16_addr ? mem_59 : _GEN_2362; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2364 = 6'h3c == io_debug_rports_16_addr ? mem_60 : _GEN_2363; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2365 = 6'h3d == io_debug_rports_16_addr ? mem_61 : _GEN_2364; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2366 = 6'h3e == io_debug_rports_16_addr ? mem_62 : _GEN_2365; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2367 = 6'h3f == io_debug_rports_16_addr ? mem_63 : _GEN_2366; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2369 = 6'h1 == io_debug_rports_17_addr ? mem_1 : mem_0; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2370 = 6'h2 == io_debug_rports_17_addr ? mem_2 : _GEN_2369; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2371 = 6'h3 == io_debug_rports_17_addr ? mem_3 : _GEN_2370; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2372 = 6'h4 == io_debug_rports_17_addr ? mem_4 : _GEN_2371; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2373 = 6'h5 == io_debug_rports_17_addr ? mem_5 : _GEN_2372; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2374 = 6'h6 == io_debug_rports_17_addr ? mem_6 : _GEN_2373; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2375 = 6'h7 == io_debug_rports_17_addr ? mem_7 : _GEN_2374; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2376 = 6'h8 == io_debug_rports_17_addr ? mem_8 : _GEN_2375; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2377 = 6'h9 == io_debug_rports_17_addr ? mem_9 : _GEN_2376; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2378 = 6'ha == io_debug_rports_17_addr ? mem_10 : _GEN_2377; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2379 = 6'hb == io_debug_rports_17_addr ? mem_11 : _GEN_2378; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2380 = 6'hc == io_debug_rports_17_addr ? mem_12 : _GEN_2379; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2381 = 6'hd == io_debug_rports_17_addr ? mem_13 : _GEN_2380; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2382 = 6'he == io_debug_rports_17_addr ? mem_14 : _GEN_2381; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2383 = 6'hf == io_debug_rports_17_addr ? mem_15 : _GEN_2382; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2384 = 6'h10 == io_debug_rports_17_addr ? mem_16 : _GEN_2383; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2385 = 6'h11 == io_debug_rports_17_addr ? mem_17 : _GEN_2384; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2386 = 6'h12 == io_debug_rports_17_addr ? mem_18 : _GEN_2385; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2387 = 6'h13 == io_debug_rports_17_addr ? mem_19 : _GEN_2386; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2388 = 6'h14 == io_debug_rports_17_addr ? mem_20 : _GEN_2387; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2389 = 6'h15 == io_debug_rports_17_addr ? mem_21 : _GEN_2388; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2390 = 6'h16 == io_debug_rports_17_addr ? mem_22 : _GEN_2389; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2391 = 6'h17 == io_debug_rports_17_addr ? mem_23 : _GEN_2390; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2392 = 6'h18 == io_debug_rports_17_addr ? mem_24 : _GEN_2391; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2393 = 6'h19 == io_debug_rports_17_addr ? mem_25 : _GEN_2392; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2394 = 6'h1a == io_debug_rports_17_addr ? mem_26 : _GEN_2393; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2395 = 6'h1b == io_debug_rports_17_addr ? mem_27 : _GEN_2394; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2396 = 6'h1c == io_debug_rports_17_addr ? mem_28 : _GEN_2395; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2397 = 6'h1d == io_debug_rports_17_addr ? mem_29 : _GEN_2396; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2398 = 6'h1e == io_debug_rports_17_addr ? mem_30 : _GEN_2397; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2399 = 6'h1f == io_debug_rports_17_addr ? mem_31 : _GEN_2398; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2400 = 6'h20 == io_debug_rports_17_addr ? mem_32 : _GEN_2399; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2401 = 6'h21 == io_debug_rports_17_addr ? mem_33 : _GEN_2400; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2402 = 6'h22 == io_debug_rports_17_addr ? mem_34 : _GEN_2401; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2403 = 6'h23 == io_debug_rports_17_addr ? mem_35 : _GEN_2402; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2404 = 6'h24 == io_debug_rports_17_addr ? mem_36 : _GEN_2403; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2405 = 6'h25 == io_debug_rports_17_addr ? mem_37 : _GEN_2404; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2406 = 6'h26 == io_debug_rports_17_addr ? mem_38 : _GEN_2405; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2407 = 6'h27 == io_debug_rports_17_addr ? mem_39 : _GEN_2406; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2408 = 6'h28 == io_debug_rports_17_addr ? mem_40 : _GEN_2407; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2409 = 6'h29 == io_debug_rports_17_addr ? mem_41 : _GEN_2408; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2410 = 6'h2a == io_debug_rports_17_addr ? mem_42 : _GEN_2409; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2411 = 6'h2b == io_debug_rports_17_addr ? mem_43 : _GEN_2410; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2412 = 6'h2c == io_debug_rports_17_addr ? mem_44 : _GEN_2411; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2413 = 6'h2d == io_debug_rports_17_addr ? mem_45 : _GEN_2412; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2414 = 6'h2e == io_debug_rports_17_addr ? mem_46 : _GEN_2413; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2415 = 6'h2f == io_debug_rports_17_addr ? mem_47 : _GEN_2414; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2416 = 6'h30 == io_debug_rports_17_addr ? mem_48 : _GEN_2415; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2417 = 6'h31 == io_debug_rports_17_addr ? mem_49 : _GEN_2416; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2418 = 6'h32 == io_debug_rports_17_addr ? mem_50 : _GEN_2417; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2419 = 6'h33 == io_debug_rports_17_addr ? mem_51 : _GEN_2418; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2420 = 6'h34 == io_debug_rports_17_addr ? mem_52 : _GEN_2419; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2421 = 6'h35 == io_debug_rports_17_addr ? mem_53 : _GEN_2420; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2422 = 6'h36 == io_debug_rports_17_addr ? mem_54 : _GEN_2421; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2423 = 6'h37 == io_debug_rports_17_addr ? mem_55 : _GEN_2422; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2424 = 6'h38 == io_debug_rports_17_addr ? mem_56 : _GEN_2423; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2425 = 6'h39 == io_debug_rports_17_addr ? mem_57 : _GEN_2424; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2426 = 6'h3a == io_debug_rports_17_addr ? mem_58 : _GEN_2425; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2427 = 6'h3b == io_debug_rports_17_addr ? mem_59 : _GEN_2426; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2428 = 6'h3c == io_debug_rports_17_addr ? mem_60 : _GEN_2427; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2429 = 6'h3d == io_debug_rports_17_addr ? mem_61 : _GEN_2428; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2430 = 6'h3e == io_debug_rports_17_addr ? mem_62 : _GEN_2429; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2431 = 6'h3f == io_debug_rports_17_addr ? mem_63 : _GEN_2430; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2433 = 6'h1 == io_debug_rports_18_addr ? mem_1 : mem_0; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2434 = 6'h2 == io_debug_rports_18_addr ? mem_2 : _GEN_2433; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2435 = 6'h3 == io_debug_rports_18_addr ? mem_3 : _GEN_2434; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2436 = 6'h4 == io_debug_rports_18_addr ? mem_4 : _GEN_2435; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2437 = 6'h5 == io_debug_rports_18_addr ? mem_5 : _GEN_2436; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2438 = 6'h6 == io_debug_rports_18_addr ? mem_6 : _GEN_2437; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2439 = 6'h7 == io_debug_rports_18_addr ? mem_7 : _GEN_2438; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2440 = 6'h8 == io_debug_rports_18_addr ? mem_8 : _GEN_2439; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2441 = 6'h9 == io_debug_rports_18_addr ? mem_9 : _GEN_2440; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2442 = 6'ha == io_debug_rports_18_addr ? mem_10 : _GEN_2441; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2443 = 6'hb == io_debug_rports_18_addr ? mem_11 : _GEN_2442; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2444 = 6'hc == io_debug_rports_18_addr ? mem_12 : _GEN_2443; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2445 = 6'hd == io_debug_rports_18_addr ? mem_13 : _GEN_2444; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2446 = 6'he == io_debug_rports_18_addr ? mem_14 : _GEN_2445; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2447 = 6'hf == io_debug_rports_18_addr ? mem_15 : _GEN_2446; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2448 = 6'h10 == io_debug_rports_18_addr ? mem_16 : _GEN_2447; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2449 = 6'h11 == io_debug_rports_18_addr ? mem_17 : _GEN_2448; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2450 = 6'h12 == io_debug_rports_18_addr ? mem_18 : _GEN_2449; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2451 = 6'h13 == io_debug_rports_18_addr ? mem_19 : _GEN_2450; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2452 = 6'h14 == io_debug_rports_18_addr ? mem_20 : _GEN_2451; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2453 = 6'h15 == io_debug_rports_18_addr ? mem_21 : _GEN_2452; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2454 = 6'h16 == io_debug_rports_18_addr ? mem_22 : _GEN_2453; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2455 = 6'h17 == io_debug_rports_18_addr ? mem_23 : _GEN_2454; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2456 = 6'h18 == io_debug_rports_18_addr ? mem_24 : _GEN_2455; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2457 = 6'h19 == io_debug_rports_18_addr ? mem_25 : _GEN_2456; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2458 = 6'h1a == io_debug_rports_18_addr ? mem_26 : _GEN_2457; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2459 = 6'h1b == io_debug_rports_18_addr ? mem_27 : _GEN_2458; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2460 = 6'h1c == io_debug_rports_18_addr ? mem_28 : _GEN_2459; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2461 = 6'h1d == io_debug_rports_18_addr ? mem_29 : _GEN_2460; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2462 = 6'h1e == io_debug_rports_18_addr ? mem_30 : _GEN_2461; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2463 = 6'h1f == io_debug_rports_18_addr ? mem_31 : _GEN_2462; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2464 = 6'h20 == io_debug_rports_18_addr ? mem_32 : _GEN_2463; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2465 = 6'h21 == io_debug_rports_18_addr ? mem_33 : _GEN_2464; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2466 = 6'h22 == io_debug_rports_18_addr ? mem_34 : _GEN_2465; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2467 = 6'h23 == io_debug_rports_18_addr ? mem_35 : _GEN_2466; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2468 = 6'h24 == io_debug_rports_18_addr ? mem_36 : _GEN_2467; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2469 = 6'h25 == io_debug_rports_18_addr ? mem_37 : _GEN_2468; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2470 = 6'h26 == io_debug_rports_18_addr ? mem_38 : _GEN_2469; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2471 = 6'h27 == io_debug_rports_18_addr ? mem_39 : _GEN_2470; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2472 = 6'h28 == io_debug_rports_18_addr ? mem_40 : _GEN_2471; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2473 = 6'h29 == io_debug_rports_18_addr ? mem_41 : _GEN_2472; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2474 = 6'h2a == io_debug_rports_18_addr ? mem_42 : _GEN_2473; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2475 = 6'h2b == io_debug_rports_18_addr ? mem_43 : _GEN_2474; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2476 = 6'h2c == io_debug_rports_18_addr ? mem_44 : _GEN_2475; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2477 = 6'h2d == io_debug_rports_18_addr ? mem_45 : _GEN_2476; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2478 = 6'h2e == io_debug_rports_18_addr ? mem_46 : _GEN_2477; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2479 = 6'h2f == io_debug_rports_18_addr ? mem_47 : _GEN_2478; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2480 = 6'h30 == io_debug_rports_18_addr ? mem_48 : _GEN_2479; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2481 = 6'h31 == io_debug_rports_18_addr ? mem_49 : _GEN_2480; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2482 = 6'h32 == io_debug_rports_18_addr ? mem_50 : _GEN_2481; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2483 = 6'h33 == io_debug_rports_18_addr ? mem_51 : _GEN_2482; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2484 = 6'h34 == io_debug_rports_18_addr ? mem_52 : _GEN_2483; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2485 = 6'h35 == io_debug_rports_18_addr ? mem_53 : _GEN_2484; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2486 = 6'h36 == io_debug_rports_18_addr ? mem_54 : _GEN_2485; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2487 = 6'h37 == io_debug_rports_18_addr ? mem_55 : _GEN_2486; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2488 = 6'h38 == io_debug_rports_18_addr ? mem_56 : _GEN_2487; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2489 = 6'h39 == io_debug_rports_18_addr ? mem_57 : _GEN_2488; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2490 = 6'h3a == io_debug_rports_18_addr ? mem_58 : _GEN_2489; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2491 = 6'h3b == io_debug_rports_18_addr ? mem_59 : _GEN_2490; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2492 = 6'h3c == io_debug_rports_18_addr ? mem_60 : _GEN_2491; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2493 = 6'h3d == io_debug_rports_18_addr ? mem_61 : _GEN_2492; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2494 = 6'h3e == io_debug_rports_18_addr ? mem_62 : _GEN_2493; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2495 = 6'h3f == io_debug_rports_18_addr ? mem_63 : _GEN_2494; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2497 = 6'h1 == io_debug_rports_19_addr ? mem_1 : mem_0; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2498 = 6'h2 == io_debug_rports_19_addr ? mem_2 : _GEN_2497; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2499 = 6'h3 == io_debug_rports_19_addr ? mem_3 : _GEN_2498; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2500 = 6'h4 == io_debug_rports_19_addr ? mem_4 : _GEN_2499; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2501 = 6'h5 == io_debug_rports_19_addr ? mem_5 : _GEN_2500; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2502 = 6'h6 == io_debug_rports_19_addr ? mem_6 : _GEN_2501; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2503 = 6'h7 == io_debug_rports_19_addr ? mem_7 : _GEN_2502; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2504 = 6'h8 == io_debug_rports_19_addr ? mem_8 : _GEN_2503; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2505 = 6'h9 == io_debug_rports_19_addr ? mem_9 : _GEN_2504; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2506 = 6'ha == io_debug_rports_19_addr ? mem_10 : _GEN_2505; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2507 = 6'hb == io_debug_rports_19_addr ? mem_11 : _GEN_2506; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2508 = 6'hc == io_debug_rports_19_addr ? mem_12 : _GEN_2507; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2509 = 6'hd == io_debug_rports_19_addr ? mem_13 : _GEN_2508; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2510 = 6'he == io_debug_rports_19_addr ? mem_14 : _GEN_2509; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2511 = 6'hf == io_debug_rports_19_addr ? mem_15 : _GEN_2510; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2512 = 6'h10 == io_debug_rports_19_addr ? mem_16 : _GEN_2511; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2513 = 6'h11 == io_debug_rports_19_addr ? mem_17 : _GEN_2512; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2514 = 6'h12 == io_debug_rports_19_addr ? mem_18 : _GEN_2513; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2515 = 6'h13 == io_debug_rports_19_addr ? mem_19 : _GEN_2514; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2516 = 6'h14 == io_debug_rports_19_addr ? mem_20 : _GEN_2515; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2517 = 6'h15 == io_debug_rports_19_addr ? mem_21 : _GEN_2516; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2518 = 6'h16 == io_debug_rports_19_addr ? mem_22 : _GEN_2517; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2519 = 6'h17 == io_debug_rports_19_addr ? mem_23 : _GEN_2518; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2520 = 6'h18 == io_debug_rports_19_addr ? mem_24 : _GEN_2519; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2521 = 6'h19 == io_debug_rports_19_addr ? mem_25 : _GEN_2520; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2522 = 6'h1a == io_debug_rports_19_addr ? mem_26 : _GEN_2521; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2523 = 6'h1b == io_debug_rports_19_addr ? mem_27 : _GEN_2522; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2524 = 6'h1c == io_debug_rports_19_addr ? mem_28 : _GEN_2523; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2525 = 6'h1d == io_debug_rports_19_addr ? mem_29 : _GEN_2524; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2526 = 6'h1e == io_debug_rports_19_addr ? mem_30 : _GEN_2525; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2527 = 6'h1f == io_debug_rports_19_addr ? mem_31 : _GEN_2526; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2528 = 6'h20 == io_debug_rports_19_addr ? mem_32 : _GEN_2527; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2529 = 6'h21 == io_debug_rports_19_addr ? mem_33 : _GEN_2528; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2530 = 6'h22 == io_debug_rports_19_addr ? mem_34 : _GEN_2529; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2531 = 6'h23 == io_debug_rports_19_addr ? mem_35 : _GEN_2530; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2532 = 6'h24 == io_debug_rports_19_addr ? mem_36 : _GEN_2531; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2533 = 6'h25 == io_debug_rports_19_addr ? mem_37 : _GEN_2532; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2534 = 6'h26 == io_debug_rports_19_addr ? mem_38 : _GEN_2533; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2535 = 6'h27 == io_debug_rports_19_addr ? mem_39 : _GEN_2534; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2536 = 6'h28 == io_debug_rports_19_addr ? mem_40 : _GEN_2535; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2537 = 6'h29 == io_debug_rports_19_addr ? mem_41 : _GEN_2536; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2538 = 6'h2a == io_debug_rports_19_addr ? mem_42 : _GEN_2537; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2539 = 6'h2b == io_debug_rports_19_addr ? mem_43 : _GEN_2538; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2540 = 6'h2c == io_debug_rports_19_addr ? mem_44 : _GEN_2539; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2541 = 6'h2d == io_debug_rports_19_addr ? mem_45 : _GEN_2540; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2542 = 6'h2e == io_debug_rports_19_addr ? mem_46 : _GEN_2541; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2543 = 6'h2f == io_debug_rports_19_addr ? mem_47 : _GEN_2542; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2544 = 6'h30 == io_debug_rports_19_addr ? mem_48 : _GEN_2543; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2545 = 6'h31 == io_debug_rports_19_addr ? mem_49 : _GEN_2544; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2546 = 6'h32 == io_debug_rports_19_addr ? mem_50 : _GEN_2545; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2547 = 6'h33 == io_debug_rports_19_addr ? mem_51 : _GEN_2546; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2548 = 6'h34 == io_debug_rports_19_addr ? mem_52 : _GEN_2547; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2549 = 6'h35 == io_debug_rports_19_addr ? mem_53 : _GEN_2548; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2550 = 6'h36 == io_debug_rports_19_addr ? mem_54 : _GEN_2549; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2551 = 6'h37 == io_debug_rports_19_addr ? mem_55 : _GEN_2550; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2552 = 6'h38 == io_debug_rports_19_addr ? mem_56 : _GEN_2551; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2553 = 6'h39 == io_debug_rports_19_addr ? mem_57 : _GEN_2552; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2554 = 6'h3a == io_debug_rports_19_addr ? mem_58 : _GEN_2553; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2555 = 6'h3b == io_debug_rports_19_addr ? mem_59 : _GEN_2554; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2556 = 6'h3c == io_debug_rports_19_addr ? mem_60 : _GEN_2555; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2557 = 6'h3d == io_debug_rports_19_addr ? mem_61 : _GEN_2556; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2558 = 6'h3e == io_debug_rports_19_addr ? mem_62 : _GEN_2557; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2559 = 6'h3f == io_debug_rports_19_addr ? mem_63 : _GEN_2558; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2561 = 6'h1 == io_debug_rports_20_addr ? mem_1 : mem_0; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2562 = 6'h2 == io_debug_rports_20_addr ? mem_2 : _GEN_2561; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2563 = 6'h3 == io_debug_rports_20_addr ? mem_3 : _GEN_2562; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2564 = 6'h4 == io_debug_rports_20_addr ? mem_4 : _GEN_2563; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2565 = 6'h5 == io_debug_rports_20_addr ? mem_5 : _GEN_2564; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2566 = 6'h6 == io_debug_rports_20_addr ? mem_6 : _GEN_2565; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2567 = 6'h7 == io_debug_rports_20_addr ? mem_7 : _GEN_2566; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2568 = 6'h8 == io_debug_rports_20_addr ? mem_8 : _GEN_2567; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2569 = 6'h9 == io_debug_rports_20_addr ? mem_9 : _GEN_2568; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2570 = 6'ha == io_debug_rports_20_addr ? mem_10 : _GEN_2569; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2571 = 6'hb == io_debug_rports_20_addr ? mem_11 : _GEN_2570; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2572 = 6'hc == io_debug_rports_20_addr ? mem_12 : _GEN_2571; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2573 = 6'hd == io_debug_rports_20_addr ? mem_13 : _GEN_2572; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2574 = 6'he == io_debug_rports_20_addr ? mem_14 : _GEN_2573; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2575 = 6'hf == io_debug_rports_20_addr ? mem_15 : _GEN_2574; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2576 = 6'h10 == io_debug_rports_20_addr ? mem_16 : _GEN_2575; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2577 = 6'h11 == io_debug_rports_20_addr ? mem_17 : _GEN_2576; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2578 = 6'h12 == io_debug_rports_20_addr ? mem_18 : _GEN_2577; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2579 = 6'h13 == io_debug_rports_20_addr ? mem_19 : _GEN_2578; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2580 = 6'h14 == io_debug_rports_20_addr ? mem_20 : _GEN_2579; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2581 = 6'h15 == io_debug_rports_20_addr ? mem_21 : _GEN_2580; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2582 = 6'h16 == io_debug_rports_20_addr ? mem_22 : _GEN_2581; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2583 = 6'h17 == io_debug_rports_20_addr ? mem_23 : _GEN_2582; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2584 = 6'h18 == io_debug_rports_20_addr ? mem_24 : _GEN_2583; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2585 = 6'h19 == io_debug_rports_20_addr ? mem_25 : _GEN_2584; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2586 = 6'h1a == io_debug_rports_20_addr ? mem_26 : _GEN_2585; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2587 = 6'h1b == io_debug_rports_20_addr ? mem_27 : _GEN_2586; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2588 = 6'h1c == io_debug_rports_20_addr ? mem_28 : _GEN_2587; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2589 = 6'h1d == io_debug_rports_20_addr ? mem_29 : _GEN_2588; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2590 = 6'h1e == io_debug_rports_20_addr ? mem_30 : _GEN_2589; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2591 = 6'h1f == io_debug_rports_20_addr ? mem_31 : _GEN_2590; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2592 = 6'h20 == io_debug_rports_20_addr ? mem_32 : _GEN_2591; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2593 = 6'h21 == io_debug_rports_20_addr ? mem_33 : _GEN_2592; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2594 = 6'h22 == io_debug_rports_20_addr ? mem_34 : _GEN_2593; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2595 = 6'h23 == io_debug_rports_20_addr ? mem_35 : _GEN_2594; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2596 = 6'h24 == io_debug_rports_20_addr ? mem_36 : _GEN_2595; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2597 = 6'h25 == io_debug_rports_20_addr ? mem_37 : _GEN_2596; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2598 = 6'h26 == io_debug_rports_20_addr ? mem_38 : _GEN_2597; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2599 = 6'h27 == io_debug_rports_20_addr ? mem_39 : _GEN_2598; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2600 = 6'h28 == io_debug_rports_20_addr ? mem_40 : _GEN_2599; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2601 = 6'h29 == io_debug_rports_20_addr ? mem_41 : _GEN_2600; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2602 = 6'h2a == io_debug_rports_20_addr ? mem_42 : _GEN_2601; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2603 = 6'h2b == io_debug_rports_20_addr ? mem_43 : _GEN_2602; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2604 = 6'h2c == io_debug_rports_20_addr ? mem_44 : _GEN_2603; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2605 = 6'h2d == io_debug_rports_20_addr ? mem_45 : _GEN_2604; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2606 = 6'h2e == io_debug_rports_20_addr ? mem_46 : _GEN_2605; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2607 = 6'h2f == io_debug_rports_20_addr ? mem_47 : _GEN_2606; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2608 = 6'h30 == io_debug_rports_20_addr ? mem_48 : _GEN_2607; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2609 = 6'h31 == io_debug_rports_20_addr ? mem_49 : _GEN_2608; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2610 = 6'h32 == io_debug_rports_20_addr ? mem_50 : _GEN_2609; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2611 = 6'h33 == io_debug_rports_20_addr ? mem_51 : _GEN_2610; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2612 = 6'h34 == io_debug_rports_20_addr ? mem_52 : _GEN_2611; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2613 = 6'h35 == io_debug_rports_20_addr ? mem_53 : _GEN_2612; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2614 = 6'h36 == io_debug_rports_20_addr ? mem_54 : _GEN_2613; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2615 = 6'h37 == io_debug_rports_20_addr ? mem_55 : _GEN_2614; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2616 = 6'h38 == io_debug_rports_20_addr ? mem_56 : _GEN_2615; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2617 = 6'h39 == io_debug_rports_20_addr ? mem_57 : _GEN_2616; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2618 = 6'h3a == io_debug_rports_20_addr ? mem_58 : _GEN_2617; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2619 = 6'h3b == io_debug_rports_20_addr ? mem_59 : _GEN_2618; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2620 = 6'h3c == io_debug_rports_20_addr ? mem_60 : _GEN_2619; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2621 = 6'h3d == io_debug_rports_20_addr ? mem_61 : _GEN_2620; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2622 = 6'h3e == io_debug_rports_20_addr ? mem_62 : _GEN_2621; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2623 = 6'h3f == io_debug_rports_20_addr ? mem_63 : _GEN_2622; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2625 = 6'h1 == io_debug_rports_21_addr ? mem_1 : mem_0; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2626 = 6'h2 == io_debug_rports_21_addr ? mem_2 : _GEN_2625; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2627 = 6'h3 == io_debug_rports_21_addr ? mem_3 : _GEN_2626; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2628 = 6'h4 == io_debug_rports_21_addr ? mem_4 : _GEN_2627; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2629 = 6'h5 == io_debug_rports_21_addr ? mem_5 : _GEN_2628; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2630 = 6'h6 == io_debug_rports_21_addr ? mem_6 : _GEN_2629; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2631 = 6'h7 == io_debug_rports_21_addr ? mem_7 : _GEN_2630; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2632 = 6'h8 == io_debug_rports_21_addr ? mem_8 : _GEN_2631; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2633 = 6'h9 == io_debug_rports_21_addr ? mem_9 : _GEN_2632; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2634 = 6'ha == io_debug_rports_21_addr ? mem_10 : _GEN_2633; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2635 = 6'hb == io_debug_rports_21_addr ? mem_11 : _GEN_2634; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2636 = 6'hc == io_debug_rports_21_addr ? mem_12 : _GEN_2635; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2637 = 6'hd == io_debug_rports_21_addr ? mem_13 : _GEN_2636; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2638 = 6'he == io_debug_rports_21_addr ? mem_14 : _GEN_2637; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2639 = 6'hf == io_debug_rports_21_addr ? mem_15 : _GEN_2638; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2640 = 6'h10 == io_debug_rports_21_addr ? mem_16 : _GEN_2639; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2641 = 6'h11 == io_debug_rports_21_addr ? mem_17 : _GEN_2640; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2642 = 6'h12 == io_debug_rports_21_addr ? mem_18 : _GEN_2641; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2643 = 6'h13 == io_debug_rports_21_addr ? mem_19 : _GEN_2642; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2644 = 6'h14 == io_debug_rports_21_addr ? mem_20 : _GEN_2643; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2645 = 6'h15 == io_debug_rports_21_addr ? mem_21 : _GEN_2644; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2646 = 6'h16 == io_debug_rports_21_addr ? mem_22 : _GEN_2645; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2647 = 6'h17 == io_debug_rports_21_addr ? mem_23 : _GEN_2646; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2648 = 6'h18 == io_debug_rports_21_addr ? mem_24 : _GEN_2647; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2649 = 6'h19 == io_debug_rports_21_addr ? mem_25 : _GEN_2648; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2650 = 6'h1a == io_debug_rports_21_addr ? mem_26 : _GEN_2649; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2651 = 6'h1b == io_debug_rports_21_addr ? mem_27 : _GEN_2650; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2652 = 6'h1c == io_debug_rports_21_addr ? mem_28 : _GEN_2651; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2653 = 6'h1d == io_debug_rports_21_addr ? mem_29 : _GEN_2652; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2654 = 6'h1e == io_debug_rports_21_addr ? mem_30 : _GEN_2653; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2655 = 6'h1f == io_debug_rports_21_addr ? mem_31 : _GEN_2654; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2656 = 6'h20 == io_debug_rports_21_addr ? mem_32 : _GEN_2655; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2657 = 6'h21 == io_debug_rports_21_addr ? mem_33 : _GEN_2656; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2658 = 6'h22 == io_debug_rports_21_addr ? mem_34 : _GEN_2657; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2659 = 6'h23 == io_debug_rports_21_addr ? mem_35 : _GEN_2658; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2660 = 6'h24 == io_debug_rports_21_addr ? mem_36 : _GEN_2659; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2661 = 6'h25 == io_debug_rports_21_addr ? mem_37 : _GEN_2660; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2662 = 6'h26 == io_debug_rports_21_addr ? mem_38 : _GEN_2661; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2663 = 6'h27 == io_debug_rports_21_addr ? mem_39 : _GEN_2662; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2664 = 6'h28 == io_debug_rports_21_addr ? mem_40 : _GEN_2663; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2665 = 6'h29 == io_debug_rports_21_addr ? mem_41 : _GEN_2664; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2666 = 6'h2a == io_debug_rports_21_addr ? mem_42 : _GEN_2665; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2667 = 6'h2b == io_debug_rports_21_addr ? mem_43 : _GEN_2666; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2668 = 6'h2c == io_debug_rports_21_addr ? mem_44 : _GEN_2667; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2669 = 6'h2d == io_debug_rports_21_addr ? mem_45 : _GEN_2668; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2670 = 6'h2e == io_debug_rports_21_addr ? mem_46 : _GEN_2669; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2671 = 6'h2f == io_debug_rports_21_addr ? mem_47 : _GEN_2670; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2672 = 6'h30 == io_debug_rports_21_addr ? mem_48 : _GEN_2671; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2673 = 6'h31 == io_debug_rports_21_addr ? mem_49 : _GEN_2672; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2674 = 6'h32 == io_debug_rports_21_addr ? mem_50 : _GEN_2673; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2675 = 6'h33 == io_debug_rports_21_addr ? mem_51 : _GEN_2674; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2676 = 6'h34 == io_debug_rports_21_addr ? mem_52 : _GEN_2675; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2677 = 6'h35 == io_debug_rports_21_addr ? mem_53 : _GEN_2676; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2678 = 6'h36 == io_debug_rports_21_addr ? mem_54 : _GEN_2677; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2679 = 6'h37 == io_debug_rports_21_addr ? mem_55 : _GEN_2678; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2680 = 6'h38 == io_debug_rports_21_addr ? mem_56 : _GEN_2679; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2681 = 6'h39 == io_debug_rports_21_addr ? mem_57 : _GEN_2680; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2682 = 6'h3a == io_debug_rports_21_addr ? mem_58 : _GEN_2681; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2683 = 6'h3b == io_debug_rports_21_addr ? mem_59 : _GEN_2682; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2684 = 6'h3c == io_debug_rports_21_addr ? mem_60 : _GEN_2683; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2685 = 6'h3d == io_debug_rports_21_addr ? mem_61 : _GEN_2684; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2686 = 6'h3e == io_debug_rports_21_addr ? mem_62 : _GEN_2685; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2687 = 6'h3f == io_debug_rports_21_addr ? mem_63 : _GEN_2686; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2689 = 6'h1 == io_debug_rports_22_addr ? mem_1 : mem_0; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2690 = 6'h2 == io_debug_rports_22_addr ? mem_2 : _GEN_2689; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2691 = 6'h3 == io_debug_rports_22_addr ? mem_3 : _GEN_2690; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2692 = 6'h4 == io_debug_rports_22_addr ? mem_4 : _GEN_2691; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2693 = 6'h5 == io_debug_rports_22_addr ? mem_5 : _GEN_2692; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2694 = 6'h6 == io_debug_rports_22_addr ? mem_6 : _GEN_2693; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2695 = 6'h7 == io_debug_rports_22_addr ? mem_7 : _GEN_2694; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2696 = 6'h8 == io_debug_rports_22_addr ? mem_8 : _GEN_2695; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2697 = 6'h9 == io_debug_rports_22_addr ? mem_9 : _GEN_2696; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2698 = 6'ha == io_debug_rports_22_addr ? mem_10 : _GEN_2697; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2699 = 6'hb == io_debug_rports_22_addr ? mem_11 : _GEN_2698; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2700 = 6'hc == io_debug_rports_22_addr ? mem_12 : _GEN_2699; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2701 = 6'hd == io_debug_rports_22_addr ? mem_13 : _GEN_2700; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2702 = 6'he == io_debug_rports_22_addr ? mem_14 : _GEN_2701; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2703 = 6'hf == io_debug_rports_22_addr ? mem_15 : _GEN_2702; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2704 = 6'h10 == io_debug_rports_22_addr ? mem_16 : _GEN_2703; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2705 = 6'h11 == io_debug_rports_22_addr ? mem_17 : _GEN_2704; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2706 = 6'h12 == io_debug_rports_22_addr ? mem_18 : _GEN_2705; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2707 = 6'h13 == io_debug_rports_22_addr ? mem_19 : _GEN_2706; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2708 = 6'h14 == io_debug_rports_22_addr ? mem_20 : _GEN_2707; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2709 = 6'h15 == io_debug_rports_22_addr ? mem_21 : _GEN_2708; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2710 = 6'h16 == io_debug_rports_22_addr ? mem_22 : _GEN_2709; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2711 = 6'h17 == io_debug_rports_22_addr ? mem_23 : _GEN_2710; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2712 = 6'h18 == io_debug_rports_22_addr ? mem_24 : _GEN_2711; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2713 = 6'h19 == io_debug_rports_22_addr ? mem_25 : _GEN_2712; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2714 = 6'h1a == io_debug_rports_22_addr ? mem_26 : _GEN_2713; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2715 = 6'h1b == io_debug_rports_22_addr ? mem_27 : _GEN_2714; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2716 = 6'h1c == io_debug_rports_22_addr ? mem_28 : _GEN_2715; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2717 = 6'h1d == io_debug_rports_22_addr ? mem_29 : _GEN_2716; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2718 = 6'h1e == io_debug_rports_22_addr ? mem_30 : _GEN_2717; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2719 = 6'h1f == io_debug_rports_22_addr ? mem_31 : _GEN_2718; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2720 = 6'h20 == io_debug_rports_22_addr ? mem_32 : _GEN_2719; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2721 = 6'h21 == io_debug_rports_22_addr ? mem_33 : _GEN_2720; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2722 = 6'h22 == io_debug_rports_22_addr ? mem_34 : _GEN_2721; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2723 = 6'h23 == io_debug_rports_22_addr ? mem_35 : _GEN_2722; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2724 = 6'h24 == io_debug_rports_22_addr ? mem_36 : _GEN_2723; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2725 = 6'h25 == io_debug_rports_22_addr ? mem_37 : _GEN_2724; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2726 = 6'h26 == io_debug_rports_22_addr ? mem_38 : _GEN_2725; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2727 = 6'h27 == io_debug_rports_22_addr ? mem_39 : _GEN_2726; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2728 = 6'h28 == io_debug_rports_22_addr ? mem_40 : _GEN_2727; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2729 = 6'h29 == io_debug_rports_22_addr ? mem_41 : _GEN_2728; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2730 = 6'h2a == io_debug_rports_22_addr ? mem_42 : _GEN_2729; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2731 = 6'h2b == io_debug_rports_22_addr ? mem_43 : _GEN_2730; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2732 = 6'h2c == io_debug_rports_22_addr ? mem_44 : _GEN_2731; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2733 = 6'h2d == io_debug_rports_22_addr ? mem_45 : _GEN_2732; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2734 = 6'h2e == io_debug_rports_22_addr ? mem_46 : _GEN_2733; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2735 = 6'h2f == io_debug_rports_22_addr ? mem_47 : _GEN_2734; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2736 = 6'h30 == io_debug_rports_22_addr ? mem_48 : _GEN_2735; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2737 = 6'h31 == io_debug_rports_22_addr ? mem_49 : _GEN_2736; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2738 = 6'h32 == io_debug_rports_22_addr ? mem_50 : _GEN_2737; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2739 = 6'h33 == io_debug_rports_22_addr ? mem_51 : _GEN_2738; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2740 = 6'h34 == io_debug_rports_22_addr ? mem_52 : _GEN_2739; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2741 = 6'h35 == io_debug_rports_22_addr ? mem_53 : _GEN_2740; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2742 = 6'h36 == io_debug_rports_22_addr ? mem_54 : _GEN_2741; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2743 = 6'h37 == io_debug_rports_22_addr ? mem_55 : _GEN_2742; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2744 = 6'h38 == io_debug_rports_22_addr ? mem_56 : _GEN_2743; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2745 = 6'h39 == io_debug_rports_22_addr ? mem_57 : _GEN_2744; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2746 = 6'h3a == io_debug_rports_22_addr ? mem_58 : _GEN_2745; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2747 = 6'h3b == io_debug_rports_22_addr ? mem_59 : _GEN_2746; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2748 = 6'h3c == io_debug_rports_22_addr ? mem_60 : _GEN_2747; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2749 = 6'h3d == io_debug_rports_22_addr ? mem_61 : _GEN_2748; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2750 = 6'h3e == io_debug_rports_22_addr ? mem_62 : _GEN_2749; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2751 = 6'h3f == io_debug_rports_22_addr ? mem_63 : _GEN_2750; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2753 = 6'h1 == io_debug_rports_23_addr ? mem_1 : mem_0; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2754 = 6'h2 == io_debug_rports_23_addr ? mem_2 : _GEN_2753; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2755 = 6'h3 == io_debug_rports_23_addr ? mem_3 : _GEN_2754; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2756 = 6'h4 == io_debug_rports_23_addr ? mem_4 : _GEN_2755; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2757 = 6'h5 == io_debug_rports_23_addr ? mem_5 : _GEN_2756; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2758 = 6'h6 == io_debug_rports_23_addr ? mem_6 : _GEN_2757; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2759 = 6'h7 == io_debug_rports_23_addr ? mem_7 : _GEN_2758; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2760 = 6'h8 == io_debug_rports_23_addr ? mem_8 : _GEN_2759; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2761 = 6'h9 == io_debug_rports_23_addr ? mem_9 : _GEN_2760; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2762 = 6'ha == io_debug_rports_23_addr ? mem_10 : _GEN_2761; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2763 = 6'hb == io_debug_rports_23_addr ? mem_11 : _GEN_2762; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2764 = 6'hc == io_debug_rports_23_addr ? mem_12 : _GEN_2763; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2765 = 6'hd == io_debug_rports_23_addr ? mem_13 : _GEN_2764; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2766 = 6'he == io_debug_rports_23_addr ? mem_14 : _GEN_2765; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2767 = 6'hf == io_debug_rports_23_addr ? mem_15 : _GEN_2766; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2768 = 6'h10 == io_debug_rports_23_addr ? mem_16 : _GEN_2767; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2769 = 6'h11 == io_debug_rports_23_addr ? mem_17 : _GEN_2768; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2770 = 6'h12 == io_debug_rports_23_addr ? mem_18 : _GEN_2769; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2771 = 6'h13 == io_debug_rports_23_addr ? mem_19 : _GEN_2770; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2772 = 6'h14 == io_debug_rports_23_addr ? mem_20 : _GEN_2771; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2773 = 6'h15 == io_debug_rports_23_addr ? mem_21 : _GEN_2772; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2774 = 6'h16 == io_debug_rports_23_addr ? mem_22 : _GEN_2773; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2775 = 6'h17 == io_debug_rports_23_addr ? mem_23 : _GEN_2774; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2776 = 6'h18 == io_debug_rports_23_addr ? mem_24 : _GEN_2775; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2777 = 6'h19 == io_debug_rports_23_addr ? mem_25 : _GEN_2776; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2778 = 6'h1a == io_debug_rports_23_addr ? mem_26 : _GEN_2777; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2779 = 6'h1b == io_debug_rports_23_addr ? mem_27 : _GEN_2778; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2780 = 6'h1c == io_debug_rports_23_addr ? mem_28 : _GEN_2779; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2781 = 6'h1d == io_debug_rports_23_addr ? mem_29 : _GEN_2780; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2782 = 6'h1e == io_debug_rports_23_addr ? mem_30 : _GEN_2781; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2783 = 6'h1f == io_debug_rports_23_addr ? mem_31 : _GEN_2782; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2784 = 6'h20 == io_debug_rports_23_addr ? mem_32 : _GEN_2783; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2785 = 6'h21 == io_debug_rports_23_addr ? mem_33 : _GEN_2784; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2786 = 6'h22 == io_debug_rports_23_addr ? mem_34 : _GEN_2785; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2787 = 6'h23 == io_debug_rports_23_addr ? mem_35 : _GEN_2786; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2788 = 6'h24 == io_debug_rports_23_addr ? mem_36 : _GEN_2787; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2789 = 6'h25 == io_debug_rports_23_addr ? mem_37 : _GEN_2788; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2790 = 6'h26 == io_debug_rports_23_addr ? mem_38 : _GEN_2789; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2791 = 6'h27 == io_debug_rports_23_addr ? mem_39 : _GEN_2790; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2792 = 6'h28 == io_debug_rports_23_addr ? mem_40 : _GEN_2791; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2793 = 6'h29 == io_debug_rports_23_addr ? mem_41 : _GEN_2792; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2794 = 6'h2a == io_debug_rports_23_addr ? mem_42 : _GEN_2793; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2795 = 6'h2b == io_debug_rports_23_addr ? mem_43 : _GEN_2794; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2796 = 6'h2c == io_debug_rports_23_addr ? mem_44 : _GEN_2795; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2797 = 6'h2d == io_debug_rports_23_addr ? mem_45 : _GEN_2796; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2798 = 6'h2e == io_debug_rports_23_addr ? mem_46 : _GEN_2797; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2799 = 6'h2f == io_debug_rports_23_addr ? mem_47 : _GEN_2798; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2800 = 6'h30 == io_debug_rports_23_addr ? mem_48 : _GEN_2799; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2801 = 6'h31 == io_debug_rports_23_addr ? mem_49 : _GEN_2800; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2802 = 6'h32 == io_debug_rports_23_addr ? mem_50 : _GEN_2801; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2803 = 6'h33 == io_debug_rports_23_addr ? mem_51 : _GEN_2802; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2804 = 6'h34 == io_debug_rports_23_addr ? mem_52 : _GEN_2803; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2805 = 6'h35 == io_debug_rports_23_addr ? mem_53 : _GEN_2804; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2806 = 6'h36 == io_debug_rports_23_addr ? mem_54 : _GEN_2805; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2807 = 6'h37 == io_debug_rports_23_addr ? mem_55 : _GEN_2806; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2808 = 6'h38 == io_debug_rports_23_addr ? mem_56 : _GEN_2807; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2809 = 6'h39 == io_debug_rports_23_addr ? mem_57 : _GEN_2808; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2810 = 6'h3a == io_debug_rports_23_addr ? mem_58 : _GEN_2809; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2811 = 6'h3b == io_debug_rports_23_addr ? mem_59 : _GEN_2810; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2812 = 6'h3c == io_debug_rports_23_addr ? mem_60 : _GEN_2811; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2813 = 6'h3d == io_debug_rports_23_addr ? mem_61 : _GEN_2812; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2814 = 6'h3e == io_debug_rports_23_addr ? mem_62 : _GEN_2813; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2815 = 6'h3f == io_debug_rports_23_addr ? mem_63 : _GEN_2814; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2817 = 6'h1 == io_debug_rports_24_addr ? mem_1 : mem_0; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2818 = 6'h2 == io_debug_rports_24_addr ? mem_2 : _GEN_2817; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2819 = 6'h3 == io_debug_rports_24_addr ? mem_3 : _GEN_2818; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2820 = 6'h4 == io_debug_rports_24_addr ? mem_4 : _GEN_2819; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2821 = 6'h5 == io_debug_rports_24_addr ? mem_5 : _GEN_2820; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2822 = 6'h6 == io_debug_rports_24_addr ? mem_6 : _GEN_2821; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2823 = 6'h7 == io_debug_rports_24_addr ? mem_7 : _GEN_2822; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2824 = 6'h8 == io_debug_rports_24_addr ? mem_8 : _GEN_2823; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2825 = 6'h9 == io_debug_rports_24_addr ? mem_9 : _GEN_2824; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2826 = 6'ha == io_debug_rports_24_addr ? mem_10 : _GEN_2825; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2827 = 6'hb == io_debug_rports_24_addr ? mem_11 : _GEN_2826; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2828 = 6'hc == io_debug_rports_24_addr ? mem_12 : _GEN_2827; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2829 = 6'hd == io_debug_rports_24_addr ? mem_13 : _GEN_2828; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2830 = 6'he == io_debug_rports_24_addr ? mem_14 : _GEN_2829; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2831 = 6'hf == io_debug_rports_24_addr ? mem_15 : _GEN_2830; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2832 = 6'h10 == io_debug_rports_24_addr ? mem_16 : _GEN_2831; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2833 = 6'h11 == io_debug_rports_24_addr ? mem_17 : _GEN_2832; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2834 = 6'h12 == io_debug_rports_24_addr ? mem_18 : _GEN_2833; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2835 = 6'h13 == io_debug_rports_24_addr ? mem_19 : _GEN_2834; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2836 = 6'h14 == io_debug_rports_24_addr ? mem_20 : _GEN_2835; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2837 = 6'h15 == io_debug_rports_24_addr ? mem_21 : _GEN_2836; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2838 = 6'h16 == io_debug_rports_24_addr ? mem_22 : _GEN_2837; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2839 = 6'h17 == io_debug_rports_24_addr ? mem_23 : _GEN_2838; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2840 = 6'h18 == io_debug_rports_24_addr ? mem_24 : _GEN_2839; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2841 = 6'h19 == io_debug_rports_24_addr ? mem_25 : _GEN_2840; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2842 = 6'h1a == io_debug_rports_24_addr ? mem_26 : _GEN_2841; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2843 = 6'h1b == io_debug_rports_24_addr ? mem_27 : _GEN_2842; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2844 = 6'h1c == io_debug_rports_24_addr ? mem_28 : _GEN_2843; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2845 = 6'h1d == io_debug_rports_24_addr ? mem_29 : _GEN_2844; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2846 = 6'h1e == io_debug_rports_24_addr ? mem_30 : _GEN_2845; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2847 = 6'h1f == io_debug_rports_24_addr ? mem_31 : _GEN_2846; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2848 = 6'h20 == io_debug_rports_24_addr ? mem_32 : _GEN_2847; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2849 = 6'h21 == io_debug_rports_24_addr ? mem_33 : _GEN_2848; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2850 = 6'h22 == io_debug_rports_24_addr ? mem_34 : _GEN_2849; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2851 = 6'h23 == io_debug_rports_24_addr ? mem_35 : _GEN_2850; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2852 = 6'h24 == io_debug_rports_24_addr ? mem_36 : _GEN_2851; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2853 = 6'h25 == io_debug_rports_24_addr ? mem_37 : _GEN_2852; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2854 = 6'h26 == io_debug_rports_24_addr ? mem_38 : _GEN_2853; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2855 = 6'h27 == io_debug_rports_24_addr ? mem_39 : _GEN_2854; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2856 = 6'h28 == io_debug_rports_24_addr ? mem_40 : _GEN_2855; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2857 = 6'h29 == io_debug_rports_24_addr ? mem_41 : _GEN_2856; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2858 = 6'h2a == io_debug_rports_24_addr ? mem_42 : _GEN_2857; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2859 = 6'h2b == io_debug_rports_24_addr ? mem_43 : _GEN_2858; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2860 = 6'h2c == io_debug_rports_24_addr ? mem_44 : _GEN_2859; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2861 = 6'h2d == io_debug_rports_24_addr ? mem_45 : _GEN_2860; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2862 = 6'h2e == io_debug_rports_24_addr ? mem_46 : _GEN_2861; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2863 = 6'h2f == io_debug_rports_24_addr ? mem_47 : _GEN_2862; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2864 = 6'h30 == io_debug_rports_24_addr ? mem_48 : _GEN_2863; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2865 = 6'h31 == io_debug_rports_24_addr ? mem_49 : _GEN_2864; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2866 = 6'h32 == io_debug_rports_24_addr ? mem_50 : _GEN_2865; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2867 = 6'h33 == io_debug_rports_24_addr ? mem_51 : _GEN_2866; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2868 = 6'h34 == io_debug_rports_24_addr ? mem_52 : _GEN_2867; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2869 = 6'h35 == io_debug_rports_24_addr ? mem_53 : _GEN_2868; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2870 = 6'h36 == io_debug_rports_24_addr ? mem_54 : _GEN_2869; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2871 = 6'h37 == io_debug_rports_24_addr ? mem_55 : _GEN_2870; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2872 = 6'h38 == io_debug_rports_24_addr ? mem_56 : _GEN_2871; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2873 = 6'h39 == io_debug_rports_24_addr ? mem_57 : _GEN_2872; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2874 = 6'h3a == io_debug_rports_24_addr ? mem_58 : _GEN_2873; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2875 = 6'h3b == io_debug_rports_24_addr ? mem_59 : _GEN_2874; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2876 = 6'h3c == io_debug_rports_24_addr ? mem_60 : _GEN_2875; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2877 = 6'h3d == io_debug_rports_24_addr ? mem_61 : _GEN_2876; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2878 = 6'h3e == io_debug_rports_24_addr ? mem_62 : _GEN_2877; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2879 = 6'h3f == io_debug_rports_24_addr ? mem_63 : _GEN_2878; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2881 = 6'h1 == io_debug_rports_25_addr ? mem_1 : mem_0; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2882 = 6'h2 == io_debug_rports_25_addr ? mem_2 : _GEN_2881; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2883 = 6'h3 == io_debug_rports_25_addr ? mem_3 : _GEN_2882; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2884 = 6'h4 == io_debug_rports_25_addr ? mem_4 : _GEN_2883; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2885 = 6'h5 == io_debug_rports_25_addr ? mem_5 : _GEN_2884; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2886 = 6'h6 == io_debug_rports_25_addr ? mem_6 : _GEN_2885; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2887 = 6'h7 == io_debug_rports_25_addr ? mem_7 : _GEN_2886; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2888 = 6'h8 == io_debug_rports_25_addr ? mem_8 : _GEN_2887; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2889 = 6'h9 == io_debug_rports_25_addr ? mem_9 : _GEN_2888; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2890 = 6'ha == io_debug_rports_25_addr ? mem_10 : _GEN_2889; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2891 = 6'hb == io_debug_rports_25_addr ? mem_11 : _GEN_2890; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2892 = 6'hc == io_debug_rports_25_addr ? mem_12 : _GEN_2891; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2893 = 6'hd == io_debug_rports_25_addr ? mem_13 : _GEN_2892; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2894 = 6'he == io_debug_rports_25_addr ? mem_14 : _GEN_2893; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2895 = 6'hf == io_debug_rports_25_addr ? mem_15 : _GEN_2894; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2896 = 6'h10 == io_debug_rports_25_addr ? mem_16 : _GEN_2895; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2897 = 6'h11 == io_debug_rports_25_addr ? mem_17 : _GEN_2896; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2898 = 6'h12 == io_debug_rports_25_addr ? mem_18 : _GEN_2897; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2899 = 6'h13 == io_debug_rports_25_addr ? mem_19 : _GEN_2898; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2900 = 6'h14 == io_debug_rports_25_addr ? mem_20 : _GEN_2899; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2901 = 6'h15 == io_debug_rports_25_addr ? mem_21 : _GEN_2900; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2902 = 6'h16 == io_debug_rports_25_addr ? mem_22 : _GEN_2901; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2903 = 6'h17 == io_debug_rports_25_addr ? mem_23 : _GEN_2902; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2904 = 6'h18 == io_debug_rports_25_addr ? mem_24 : _GEN_2903; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2905 = 6'h19 == io_debug_rports_25_addr ? mem_25 : _GEN_2904; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2906 = 6'h1a == io_debug_rports_25_addr ? mem_26 : _GEN_2905; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2907 = 6'h1b == io_debug_rports_25_addr ? mem_27 : _GEN_2906; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2908 = 6'h1c == io_debug_rports_25_addr ? mem_28 : _GEN_2907; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2909 = 6'h1d == io_debug_rports_25_addr ? mem_29 : _GEN_2908; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2910 = 6'h1e == io_debug_rports_25_addr ? mem_30 : _GEN_2909; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2911 = 6'h1f == io_debug_rports_25_addr ? mem_31 : _GEN_2910; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2912 = 6'h20 == io_debug_rports_25_addr ? mem_32 : _GEN_2911; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2913 = 6'h21 == io_debug_rports_25_addr ? mem_33 : _GEN_2912; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2914 = 6'h22 == io_debug_rports_25_addr ? mem_34 : _GEN_2913; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2915 = 6'h23 == io_debug_rports_25_addr ? mem_35 : _GEN_2914; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2916 = 6'h24 == io_debug_rports_25_addr ? mem_36 : _GEN_2915; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2917 = 6'h25 == io_debug_rports_25_addr ? mem_37 : _GEN_2916; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2918 = 6'h26 == io_debug_rports_25_addr ? mem_38 : _GEN_2917; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2919 = 6'h27 == io_debug_rports_25_addr ? mem_39 : _GEN_2918; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2920 = 6'h28 == io_debug_rports_25_addr ? mem_40 : _GEN_2919; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2921 = 6'h29 == io_debug_rports_25_addr ? mem_41 : _GEN_2920; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2922 = 6'h2a == io_debug_rports_25_addr ? mem_42 : _GEN_2921; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2923 = 6'h2b == io_debug_rports_25_addr ? mem_43 : _GEN_2922; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2924 = 6'h2c == io_debug_rports_25_addr ? mem_44 : _GEN_2923; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2925 = 6'h2d == io_debug_rports_25_addr ? mem_45 : _GEN_2924; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2926 = 6'h2e == io_debug_rports_25_addr ? mem_46 : _GEN_2925; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2927 = 6'h2f == io_debug_rports_25_addr ? mem_47 : _GEN_2926; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2928 = 6'h30 == io_debug_rports_25_addr ? mem_48 : _GEN_2927; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2929 = 6'h31 == io_debug_rports_25_addr ? mem_49 : _GEN_2928; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2930 = 6'h32 == io_debug_rports_25_addr ? mem_50 : _GEN_2929; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2931 = 6'h33 == io_debug_rports_25_addr ? mem_51 : _GEN_2930; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2932 = 6'h34 == io_debug_rports_25_addr ? mem_52 : _GEN_2931; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2933 = 6'h35 == io_debug_rports_25_addr ? mem_53 : _GEN_2932; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2934 = 6'h36 == io_debug_rports_25_addr ? mem_54 : _GEN_2933; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2935 = 6'h37 == io_debug_rports_25_addr ? mem_55 : _GEN_2934; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2936 = 6'h38 == io_debug_rports_25_addr ? mem_56 : _GEN_2935; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2937 = 6'h39 == io_debug_rports_25_addr ? mem_57 : _GEN_2936; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2938 = 6'h3a == io_debug_rports_25_addr ? mem_58 : _GEN_2937; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2939 = 6'h3b == io_debug_rports_25_addr ? mem_59 : _GEN_2938; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2940 = 6'h3c == io_debug_rports_25_addr ? mem_60 : _GEN_2939; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2941 = 6'h3d == io_debug_rports_25_addr ? mem_61 : _GEN_2940; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2942 = 6'h3e == io_debug_rports_25_addr ? mem_62 : _GEN_2941; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2943 = 6'h3f == io_debug_rports_25_addr ? mem_63 : _GEN_2942; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2945 = 6'h1 == io_debug_rports_26_addr ? mem_1 : mem_0; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2946 = 6'h2 == io_debug_rports_26_addr ? mem_2 : _GEN_2945; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2947 = 6'h3 == io_debug_rports_26_addr ? mem_3 : _GEN_2946; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2948 = 6'h4 == io_debug_rports_26_addr ? mem_4 : _GEN_2947; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2949 = 6'h5 == io_debug_rports_26_addr ? mem_5 : _GEN_2948; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2950 = 6'h6 == io_debug_rports_26_addr ? mem_6 : _GEN_2949; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2951 = 6'h7 == io_debug_rports_26_addr ? mem_7 : _GEN_2950; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2952 = 6'h8 == io_debug_rports_26_addr ? mem_8 : _GEN_2951; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2953 = 6'h9 == io_debug_rports_26_addr ? mem_9 : _GEN_2952; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2954 = 6'ha == io_debug_rports_26_addr ? mem_10 : _GEN_2953; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2955 = 6'hb == io_debug_rports_26_addr ? mem_11 : _GEN_2954; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2956 = 6'hc == io_debug_rports_26_addr ? mem_12 : _GEN_2955; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2957 = 6'hd == io_debug_rports_26_addr ? mem_13 : _GEN_2956; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2958 = 6'he == io_debug_rports_26_addr ? mem_14 : _GEN_2957; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2959 = 6'hf == io_debug_rports_26_addr ? mem_15 : _GEN_2958; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2960 = 6'h10 == io_debug_rports_26_addr ? mem_16 : _GEN_2959; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2961 = 6'h11 == io_debug_rports_26_addr ? mem_17 : _GEN_2960; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2962 = 6'h12 == io_debug_rports_26_addr ? mem_18 : _GEN_2961; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2963 = 6'h13 == io_debug_rports_26_addr ? mem_19 : _GEN_2962; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2964 = 6'h14 == io_debug_rports_26_addr ? mem_20 : _GEN_2963; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2965 = 6'h15 == io_debug_rports_26_addr ? mem_21 : _GEN_2964; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2966 = 6'h16 == io_debug_rports_26_addr ? mem_22 : _GEN_2965; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2967 = 6'h17 == io_debug_rports_26_addr ? mem_23 : _GEN_2966; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2968 = 6'h18 == io_debug_rports_26_addr ? mem_24 : _GEN_2967; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2969 = 6'h19 == io_debug_rports_26_addr ? mem_25 : _GEN_2968; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2970 = 6'h1a == io_debug_rports_26_addr ? mem_26 : _GEN_2969; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2971 = 6'h1b == io_debug_rports_26_addr ? mem_27 : _GEN_2970; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2972 = 6'h1c == io_debug_rports_26_addr ? mem_28 : _GEN_2971; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2973 = 6'h1d == io_debug_rports_26_addr ? mem_29 : _GEN_2972; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2974 = 6'h1e == io_debug_rports_26_addr ? mem_30 : _GEN_2973; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2975 = 6'h1f == io_debug_rports_26_addr ? mem_31 : _GEN_2974; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2976 = 6'h20 == io_debug_rports_26_addr ? mem_32 : _GEN_2975; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2977 = 6'h21 == io_debug_rports_26_addr ? mem_33 : _GEN_2976; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2978 = 6'h22 == io_debug_rports_26_addr ? mem_34 : _GEN_2977; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2979 = 6'h23 == io_debug_rports_26_addr ? mem_35 : _GEN_2978; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2980 = 6'h24 == io_debug_rports_26_addr ? mem_36 : _GEN_2979; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2981 = 6'h25 == io_debug_rports_26_addr ? mem_37 : _GEN_2980; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2982 = 6'h26 == io_debug_rports_26_addr ? mem_38 : _GEN_2981; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2983 = 6'h27 == io_debug_rports_26_addr ? mem_39 : _GEN_2982; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2984 = 6'h28 == io_debug_rports_26_addr ? mem_40 : _GEN_2983; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2985 = 6'h29 == io_debug_rports_26_addr ? mem_41 : _GEN_2984; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2986 = 6'h2a == io_debug_rports_26_addr ? mem_42 : _GEN_2985; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2987 = 6'h2b == io_debug_rports_26_addr ? mem_43 : _GEN_2986; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2988 = 6'h2c == io_debug_rports_26_addr ? mem_44 : _GEN_2987; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2989 = 6'h2d == io_debug_rports_26_addr ? mem_45 : _GEN_2988; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2990 = 6'h2e == io_debug_rports_26_addr ? mem_46 : _GEN_2989; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2991 = 6'h2f == io_debug_rports_26_addr ? mem_47 : _GEN_2990; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2992 = 6'h30 == io_debug_rports_26_addr ? mem_48 : _GEN_2991; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2993 = 6'h31 == io_debug_rports_26_addr ? mem_49 : _GEN_2992; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2994 = 6'h32 == io_debug_rports_26_addr ? mem_50 : _GEN_2993; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2995 = 6'h33 == io_debug_rports_26_addr ? mem_51 : _GEN_2994; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2996 = 6'h34 == io_debug_rports_26_addr ? mem_52 : _GEN_2995; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2997 = 6'h35 == io_debug_rports_26_addr ? mem_53 : _GEN_2996; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2998 = 6'h36 == io_debug_rports_26_addr ? mem_54 : _GEN_2997; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_2999 = 6'h37 == io_debug_rports_26_addr ? mem_55 : _GEN_2998; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3000 = 6'h38 == io_debug_rports_26_addr ? mem_56 : _GEN_2999; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3001 = 6'h39 == io_debug_rports_26_addr ? mem_57 : _GEN_3000; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3002 = 6'h3a == io_debug_rports_26_addr ? mem_58 : _GEN_3001; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3003 = 6'h3b == io_debug_rports_26_addr ? mem_59 : _GEN_3002; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3004 = 6'h3c == io_debug_rports_26_addr ? mem_60 : _GEN_3003; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3005 = 6'h3d == io_debug_rports_26_addr ? mem_61 : _GEN_3004; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3006 = 6'h3e == io_debug_rports_26_addr ? mem_62 : _GEN_3005; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3007 = 6'h3f == io_debug_rports_26_addr ? mem_63 : _GEN_3006; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3009 = 6'h1 == io_debug_rports_27_addr ? mem_1 : mem_0; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3010 = 6'h2 == io_debug_rports_27_addr ? mem_2 : _GEN_3009; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3011 = 6'h3 == io_debug_rports_27_addr ? mem_3 : _GEN_3010; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3012 = 6'h4 == io_debug_rports_27_addr ? mem_4 : _GEN_3011; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3013 = 6'h5 == io_debug_rports_27_addr ? mem_5 : _GEN_3012; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3014 = 6'h6 == io_debug_rports_27_addr ? mem_6 : _GEN_3013; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3015 = 6'h7 == io_debug_rports_27_addr ? mem_7 : _GEN_3014; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3016 = 6'h8 == io_debug_rports_27_addr ? mem_8 : _GEN_3015; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3017 = 6'h9 == io_debug_rports_27_addr ? mem_9 : _GEN_3016; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3018 = 6'ha == io_debug_rports_27_addr ? mem_10 : _GEN_3017; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3019 = 6'hb == io_debug_rports_27_addr ? mem_11 : _GEN_3018; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3020 = 6'hc == io_debug_rports_27_addr ? mem_12 : _GEN_3019; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3021 = 6'hd == io_debug_rports_27_addr ? mem_13 : _GEN_3020; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3022 = 6'he == io_debug_rports_27_addr ? mem_14 : _GEN_3021; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3023 = 6'hf == io_debug_rports_27_addr ? mem_15 : _GEN_3022; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3024 = 6'h10 == io_debug_rports_27_addr ? mem_16 : _GEN_3023; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3025 = 6'h11 == io_debug_rports_27_addr ? mem_17 : _GEN_3024; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3026 = 6'h12 == io_debug_rports_27_addr ? mem_18 : _GEN_3025; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3027 = 6'h13 == io_debug_rports_27_addr ? mem_19 : _GEN_3026; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3028 = 6'h14 == io_debug_rports_27_addr ? mem_20 : _GEN_3027; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3029 = 6'h15 == io_debug_rports_27_addr ? mem_21 : _GEN_3028; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3030 = 6'h16 == io_debug_rports_27_addr ? mem_22 : _GEN_3029; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3031 = 6'h17 == io_debug_rports_27_addr ? mem_23 : _GEN_3030; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3032 = 6'h18 == io_debug_rports_27_addr ? mem_24 : _GEN_3031; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3033 = 6'h19 == io_debug_rports_27_addr ? mem_25 : _GEN_3032; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3034 = 6'h1a == io_debug_rports_27_addr ? mem_26 : _GEN_3033; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3035 = 6'h1b == io_debug_rports_27_addr ? mem_27 : _GEN_3034; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3036 = 6'h1c == io_debug_rports_27_addr ? mem_28 : _GEN_3035; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3037 = 6'h1d == io_debug_rports_27_addr ? mem_29 : _GEN_3036; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3038 = 6'h1e == io_debug_rports_27_addr ? mem_30 : _GEN_3037; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3039 = 6'h1f == io_debug_rports_27_addr ? mem_31 : _GEN_3038; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3040 = 6'h20 == io_debug_rports_27_addr ? mem_32 : _GEN_3039; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3041 = 6'h21 == io_debug_rports_27_addr ? mem_33 : _GEN_3040; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3042 = 6'h22 == io_debug_rports_27_addr ? mem_34 : _GEN_3041; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3043 = 6'h23 == io_debug_rports_27_addr ? mem_35 : _GEN_3042; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3044 = 6'h24 == io_debug_rports_27_addr ? mem_36 : _GEN_3043; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3045 = 6'h25 == io_debug_rports_27_addr ? mem_37 : _GEN_3044; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3046 = 6'h26 == io_debug_rports_27_addr ? mem_38 : _GEN_3045; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3047 = 6'h27 == io_debug_rports_27_addr ? mem_39 : _GEN_3046; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3048 = 6'h28 == io_debug_rports_27_addr ? mem_40 : _GEN_3047; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3049 = 6'h29 == io_debug_rports_27_addr ? mem_41 : _GEN_3048; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3050 = 6'h2a == io_debug_rports_27_addr ? mem_42 : _GEN_3049; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3051 = 6'h2b == io_debug_rports_27_addr ? mem_43 : _GEN_3050; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3052 = 6'h2c == io_debug_rports_27_addr ? mem_44 : _GEN_3051; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3053 = 6'h2d == io_debug_rports_27_addr ? mem_45 : _GEN_3052; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3054 = 6'h2e == io_debug_rports_27_addr ? mem_46 : _GEN_3053; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3055 = 6'h2f == io_debug_rports_27_addr ? mem_47 : _GEN_3054; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3056 = 6'h30 == io_debug_rports_27_addr ? mem_48 : _GEN_3055; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3057 = 6'h31 == io_debug_rports_27_addr ? mem_49 : _GEN_3056; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3058 = 6'h32 == io_debug_rports_27_addr ? mem_50 : _GEN_3057; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3059 = 6'h33 == io_debug_rports_27_addr ? mem_51 : _GEN_3058; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3060 = 6'h34 == io_debug_rports_27_addr ? mem_52 : _GEN_3059; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3061 = 6'h35 == io_debug_rports_27_addr ? mem_53 : _GEN_3060; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3062 = 6'h36 == io_debug_rports_27_addr ? mem_54 : _GEN_3061; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3063 = 6'h37 == io_debug_rports_27_addr ? mem_55 : _GEN_3062; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3064 = 6'h38 == io_debug_rports_27_addr ? mem_56 : _GEN_3063; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3065 = 6'h39 == io_debug_rports_27_addr ? mem_57 : _GEN_3064; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3066 = 6'h3a == io_debug_rports_27_addr ? mem_58 : _GEN_3065; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3067 = 6'h3b == io_debug_rports_27_addr ? mem_59 : _GEN_3066; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3068 = 6'h3c == io_debug_rports_27_addr ? mem_60 : _GEN_3067; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3069 = 6'h3d == io_debug_rports_27_addr ? mem_61 : _GEN_3068; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3070 = 6'h3e == io_debug_rports_27_addr ? mem_62 : _GEN_3069; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3071 = 6'h3f == io_debug_rports_27_addr ? mem_63 : _GEN_3070; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3073 = 6'h1 == io_debug_rports_28_addr ? mem_1 : mem_0; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3074 = 6'h2 == io_debug_rports_28_addr ? mem_2 : _GEN_3073; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3075 = 6'h3 == io_debug_rports_28_addr ? mem_3 : _GEN_3074; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3076 = 6'h4 == io_debug_rports_28_addr ? mem_4 : _GEN_3075; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3077 = 6'h5 == io_debug_rports_28_addr ? mem_5 : _GEN_3076; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3078 = 6'h6 == io_debug_rports_28_addr ? mem_6 : _GEN_3077; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3079 = 6'h7 == io_debug_rports_28_addr ? mem_7 : _GEN_3078; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3080 = 6'h8 == io_debug_rports_28_addr ? mem_8 : _GEN_3079; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3081 = 6'h9 == io_debug_rports_28_addr ? mem_9 : _GEN_3080; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3082 = 6'ha == io_debug_rports_28_addr ? mem_10 : _GEN_3081; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3083 = 6'hb == io_debug_rports_28_addr ? mem_11 : _GEN_3082; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3084 = 6'hc == io_debug_rports_28_addr ? mem_12 : _GEN_3083; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3085 = 6'hd == io_debug_rports_28_addr ? mem_13 : _GEN_3084; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3086 = 6'he == io_debug_rports_28_addr ? mem_14 : _GEN_3085; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3087 = 6'hf == io_debug_rports_28_addr ? mem_15 : _GEN_3086; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3088 = 6'h10 == io_debug_rports_28_addr ? mem_16 : _GEN_3087; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3089 = 6'h11 == io_debug_rports_28_addr ? mem_17 : _GEN_3088; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3090 = 6'h12 == io_debug_rports_28_addr ? mem_18 : _GEN_3089; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3091 = 6'h13 == io_debug_rports_28_addr ? mem_19 : _GEN_3090; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3092 = 6'h14 == io_debug_rports_28_addr ? mem_20 : _GEN_3091; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3093 = 6'h15 == io_debug_rports_28_addr ? mem_21 : _GEN_3092; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3094 = 6'h16 == io_debug_rports_28_addr ? mem_22 : _GEN_3093; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3095 = 6'h17 == io_debug_rports_28_addr ? mem_23 : _GEN_3094; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3096 = 6'h18 == io_debug_rports_28_addr ? mem_24 : _GEN_3095; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3097 = 6'h19 == io_debug_rports_28_addr ? mem_25 : _GEN_3096; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3098 = 6'h1a == io_debug_rports_28_addr ? mem_26 : _GEN_3097; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3099 = 6'h1b == io_debug_rports_28_addr ? mem_27 : _GEN_3098; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3100 = 6'h1c == io_debug_rports_28_addr ? mem_28 : _GEN_3099; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3101 = 6'h1d == io_debug_rports_28_addr ? mem_29 : _GEN_3100; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3102 = 6'h1e == io_debug_rports_28_addr ? mem_30 : _GEN_3101; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3103 = 6'h1f == io_debug_rports_28_addr ? mem_31 : _GEN_3102; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3104 = 6'h20 == io_debug_rports_28_addr ? mem_32 : _GEN_3103; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3105 = 6'h21 == io_debug_rports_28_addr ? mem_33 : _GEN_3104; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3106 = 6'h22 == io_debug_rports_28_addr ? mem_34 : _GEN_3105; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3107 = 6'h23 == io_debug_rports_28_addr ? mem_35 : _GEN_3106; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3108 = 6'h24 == io_debug_rports_28_addr ? mem_36 : _GEN_3107; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3109 = 6'h25 == io_debug_rports_28_addr ? mem_37 : _GEN_3108; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3110 = 6'h26 == io_debug_rports_28_addr ? mem_38 : _GEN_3109; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3111 = 6'h27 == io_debug_rports_28_addr ? mem_39 : _GEN_3110; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3112 = 6'h28 == io_debug_rports_28_addr ? mem_40 : _GEN_3111; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3113 = 6'h29 == io_debug_rports_28_addr ? mem_41 : _GEN_3112; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3114 = 6'h2a == io_debug_rports_28_addr ? mem_42 : _GEN_3113; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3115 = 6'h2b == io_debug_rports_28_addr ? mem_43 : _GEN_3114; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3116 = 6'h2c == io_debug_rports_28_addr ? mem_44 : _GEN_3115; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3117 = 6'h2d == io_debug_rports_28_addr ? mem_45 : _GEN_3116; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3118 = 6'h2e == io_debug_rports_28_addr ? mem_46 : _GEN_3117; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3119 = 6'h2f == io_debug_rports_28_addr ? mem_47 : _GEN_3118; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3120 = 6'h30 == io_debug_rports_28_addr ? mem_48 : _GEN_3119; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3121 = 6'h31 == io_debug_rports_28_addr ? mem_49 : _GEN_3120; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3122 = 6'h32 == io_debug_rports_28_addr ? mem_50 : _GEN_3121; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3123 = 6'h33 == io_debug_rports_28_addr ? mem_51 : _GEN_3122; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3124 = 6'h34 == io_debug_rports_28_addr ? mem_52 : _GEN_3123; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3125 = 6'h35 == io_debug_rports_28_addr ? mem_53 : _GEN_3124; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3126 = 6'h36 == io_debug_rports_28_addr ? mem_54 : _GEN_3125; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3127 = 6'h37 == io_debug_rports_28_addr ? mem_55 : _GEN_3126; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3128 = 6'h38 == io_debug_rports_28_addr ? mem_56 : _GEN_3127; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3129 = 6'h39 == io_debug_rports_28_addr ? mem_57 : _GEN_3128; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3130 = 6'h3a == io_debug_rports_28_addr ? mem_58 : _GEN_3129; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3131 = 6'h3b == io_debug_rports_28_addr ? mem_59 : _GEN_3130; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3132 = 6'h3c == io_debug_rports_28_addr ? mem_60 : _GEN_3131; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3133 = 6'h3d == io_debug_rports_28_addr ? mem_61 : _GEN_3132; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3134 = 6'h3e == io_debug_rports_28_addr ? mem_62 : _GEN_3133; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3135 = 6'h3f == io_debug_rports_28_addr ? mem_63 : _GEN_3134; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3137 = 6'h1 == io_debug_rports_29_addr ? mem_1 : mem_0; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3138 = 6'h2 == io_debug_rports_29_addr ? mem_2 : _GEN_3137; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3139 = 6'h3 == io_debug_rports_29_addr ? mem_3 : _GEN_3138; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3140 = 6'h4 == io_debug_rports_29_addr ? mem_4 : _GEN_3139; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3141 = 6'h5 == io_debug_rports_29_addr ? mem_5 : _GEN_3140; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3142 = 6'h6 == io_debug_rports_29_addr ? mem_6 : _GEN_3141; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3143 = 6'h7 == io_debug_rports_29_addr ? mem_7 : _GEN_3142; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3144 = 6'h8 == io_debug_rports_29_addr ? mem_8 : _GEN_3143; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3145 = 6'h9 == io_debug_rports_29_addr ? mem_9 : _GEN_3144; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3146 = 6'ha == io_debug_rports_29_addr ? mem_10 : _GEN_3145; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3147 = 6'hb == io_debug_rports_29_addr ? mem_11 : _GEN_3146; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3148 = 6'hc == io_debug_rports_29_addr ? mem_12 : _GEN_3147; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3149 = 6'hd == io_debug_rports_29_addr ? mem_13 : _GEN_3148; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3150 = 6'he == io_debug_rports_29_addr ? mem_14 : _GEN_3149; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3151 = 6'hf == io_debug_rports_29_addr ? mem_15 : _GEN_3150; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3152 = 6'h10 == io_debug_rports_29_addr ? mem_16 : _GEN_3151; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3153 = 6'h11 == io_debug_rports_29_addr ? mem_17 : _GEN_3152; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3154 = 6'h12 == io_debug_rports_29_addr ? mem_18 : _GEN_3153; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3155 = 6'h13 == io_debug_rports_29_addr ? mem_19 : _GEN_3154; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3156 = 6'h14 == io_debug_rports_29_addr ? mem_20 : _GEN_3155; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3157 = 6'h15 == io_debug_rports_29_addr ? mem_21 : _GEN_3156; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3158 = 6'h16 == io_debug_rports_29_addr ? mem_22 : _GEN_3157; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3159 = 6'h17 == io_debug_rports_29_addr ? mem_23 : _GEN_3158; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3160 = 6'h18 == io_debug_rports_29_addr ? mem_24 : _GEN_3159; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3161 = 6'h19 == io_debug_rports_29_addr ? mem_25 : _GEN_3160; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3162 = 6'h1a == io_debug_rports_29_addr ? mem_26 : _GEN_3161; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3163 = 6'h1b == io_debug_rports_29_addr ? mem_27 : _GEN_3162; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3164 = 6'h1c == io_debug_rports_29_addr ? mem_28 : _GEN_3163; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3165 = 6'h1d == io_debug_rports_29_addr ? mem_29 : _GEN_3164; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3166 = 6'h1e == io_debug_rports_29_addr ? mem_30 : _GEN_3165; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3167 = 6'h1f == io_debug_rports_29_addr ? mem_31 : _GEN_3166; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3168 = 6'h20 == io_debug_rports_29_addr ? mem_32 : _GEN_3167; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3169 = 6'h21 == io_debug_rports_29_addr ? mem_33 : _GEN_3168; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3170 = 6'h22 == io_debug_rports_29_addr ? mem_34 : _GEN_3169; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3171 = 6'h23 == io_debug_rports_29_addr ? mem_35 : _GEN_3170; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3172 = 6'h24 == io_debug_rports_29_addr ? mem_36 : _GEN_3171; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3173 = 6'h25 == io_debug_rports_29_addr ? mem_37 : _GEN_3172; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3174 = 6'h26 == io_debug_rports_29_addr ? mem_38 : _GEN_3173; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3175 = 6'h27 == io_debug_rports_29_addr ? mem_39 : _GEN_3174; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3176 = 6'h28 == io_debug_rports_29_addr ? mem_40 : _GEN_3175; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3177 = 6'h29 == io_debug_rports_29_addr ? mem_41 : _GEN_3176; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3178 = 6'h2a == io_debug_rports_29_addr ? mem_42 : _GEN_3177; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3179 = 6'h2b == io_debug_rports_29_addr ? mem_43 : _GEN_3178; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3180 = 6'h2c == io_debug_rports_29_addr ? mem_44 : _GEN_3179; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3181 = 6'h2d == io_debug_rports_29_addr ? mem_45 : _GEN_3180; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3182 = 6'h2e == io_debug_rports_29_addr ? mem_46 : _GEN_3181; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3183 = 6'h2f == io_debug_rports_29_addr ? mem_47 : _GEN_3182; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3184 = 6'h30 == io_debug_rports_29_addr ? mem_48 : _GEN_3183; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3185 = 6'h31 == io_debug_rports_29_addr ? mem_49 : _GEN_3184; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3186 = 6'h32 == io_debug_rports_29_addr ? mem_50 : _GEN_3185; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3187 = 6'h33 == io_debug_rports_29_addr ? mem_51 : _GEN_3186; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3188 = 6'h34 == io_debug_rports_29_addr ? mem_52 : _GEN_3187; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3189 = 6'h35 == io_debug_rports_29_addr ? mem_53 : _GEN_3188; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3190 = 6'h36 == io_debug_rports_29_addr ? mem_54 : _GEN_3189; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3191 = 6'h37 == io_debug_rports_29_addr ? mem_55 : _GEN_3190; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3192 = 6'h38 == io_debug_rports_29_addr ? mem_56 : _GEN_3191; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3193 = 6'h39 == io_debug_rports_29_addr ? mem_57 : _GEN_3192; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3194 = 6'h3a == io_debug_rports_29_addr ? mem_58 : _GEN_3193; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3195 = 6'h3b == io_debug_rports_29_addr ? mem_59 : _GEN_3194; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3196 = 6'h3c == io_debug_rports_29_addr ? mem_60 : _GEN_3195; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3197 = 6'h3d == io_debug_rports_29_addr ? mem_61 : _GEN_3196; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3198 = 6'h3e == io_debug_rports_29_addr ? mem_62 : _GEN_3197; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3199 = 6'h3f == io_debug_rports_29_addr ? mem_63 : _GEN_3198; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3201 = 6'h1 == io_debug_rports_30_addr ? mem_1 : mem_0; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3202 = 6'h2 == io_debug_rports_30_addr ? mem_2 : _GEN_3201; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3203 = 6'h3 == io_debug_rports_30_addr ? mem_3 : _GEN_3202; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3204 = 6'h4 == io_debug_rports_30_addr ? mem_4 : _GEN_3203; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3205 = 6'h5 == io_debug_rports_30_addr ? mem_5 : _GEN_3204; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3206 = 6'h6 == io_debug_rports_30_addr ? mem_6 : _GEN_3205; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3207 = 6'h7 == io_debug_rports_30_addr ? mem_7 : _GEN_3206; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3208 = 6'h8 == io_debug_rports_30_addr ? mem_8 : _GEN_3207; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3209 = 6'h9 == io_debug_rports_30_addr ? mem_9 : _GEN_3208; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3210 = 6'ha == io_debug_rports_30_addr ? mem_10 : _GEN_3209; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3211 = 6'hb == io_debug_rports_30_addr ? mem_11 : _GEN_3210; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3212 = 6'hc == io_debug_rports_30_addr ? mem_12 : _GEN_3211; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3213 = 6'hd == io_debug_rports_30_addr ? mem_13 : _GEN_3212; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3214 = 6'he == io_debug_rports_30_addr ? mem_14 : _GEN_3213; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3215 = 6'hf == io_debug_rports_30_addr ? mem_15 : _GEN_3214; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3216 = 6'h10 == io_debug_rports_30_addr ? mem_16 : _GEN_3215; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3217 = 6'h11 == io_debug_rports_30_addr ? mem_17 : _GEN_3216; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3218 = 6'h12 == io_debug_rports_30_addr ? mem_18 : _GEN_3217; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3219 = 6'h13 == io_debug_rports_30_addr ? mem_19 : _GEN_3218; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3220 = 6'h14 == io_debug_rports_30_addr ? mem_20 : _GEN_3219; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3221 = 6'h15 == io_debug_rports_30_addr ? mem_21 : _GEN_3220; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3222 = 6'h16 == io_debug_rports_30_addr ? mem_22 : _GEN_3221; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3223 = 6'h17 == io_debug_rports_30_addr ? mem_23 : _GEN_3222; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3224 = 6'h18 == io_debug_rports_30_addr ? mem_24 : _GEN_3223; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3225 = 6'h19 == io_debug_rports_30_addr ? mem_25 : _GEN_3224; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3226 = 6'h1a == io_debug_rports_30_addr ? mem_26 : _GEN_3225; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3227 = 6'h1b == io_debug_rports_30_addr ? mem_27 : _GEN_3226; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3228 = 6'h1c == io_debug_rports_30_addr ? mem_28 : _GEN_3227; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3229 = 6'h1d == io_debug_rports_30_addr ? mem_29 : _GEN_3228; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3230 = 6'h1e == io_debug_rports_30_addr ? mem_30 : _GEN_3229; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3231 = 6'h1f == io_debug_rports_30_addr ? mem_31 : _GEN_3230; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3232 = 6'h20 == io_debug_rports_30_addr ? mem_32 : _GEN_3231; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3233 = 6'h21 == io_debug_rports_30_addr ? mem_33 : _GEN_3232; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3234 = 6'h22 == io_debug_rports_30_addr ? mem_34 : _GEN_3233; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3235 = 6'h23 == io_debug_rports_30_addr ? mem_35 : _GEN_3234; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3236 = 6'h24 == io_debug_rports_30_addr ? mem_36 : _GEN_3235; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3237 = 6'h25 == io_debug_rports_30_addr ? mem_37 : _GEN_3236; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3238 = 6'h26 == io_debug_rports_30_addr ? mem_38 : _GEN_3237; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3239 = 6'h27 == io_debug_rports_30_addr ? mem_39 : _GEN_3238; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3240 = 6'h28 == io_debug_rports_30_addr ? mem_40 : _GEN_3239; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3241 = 6'h29 == io_debug_rports_30_addr ? mem_41 : _GEN_3240; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3242 = 6'h2a == io_debug_rports_30_addr ? mem_42 : _GEN_3241; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3243 = 6'h2b == io_debug_rports_30_addr ? mem_43 : _GEN_3242; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3244 = 6'h2c == io_debug_rports_30_addr ? mem_44 : _GEN_3243; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3245 = 6'h2d == io_debug_rports_30_addr ? mem_45 : _GEN_3244; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3246 = 6'h2e == io_debug_rports_30_addr ? mem_46 : _GEN_3245; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3247 = 6'h2f == io_debug_rports_30_addr ? mem_47 : _GEN_3246; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3248 = 6'h30 == io_debug_rports_30_addr ? mem_48 : _GEN_3247; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3249 = 6'h31 == io_debug_rports_30_addr ? mem_49 : _GEN_3248; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3250 = 6'h32 == io_debug_rports_30_addr ? mem_50 : _GEN_3249; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3251 = 6'h33 == io_debug_rports_30_addr ? mem_51 : _GEN_3250; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3252 = 6'h34 == io_debug_rports_30_addr ? mem_52 : _GEN_3251; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3253 = 6'h35 == io_debug_rports_30_addr ? mem_53 : _GEN_3252; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3254 = 6'h36 == io_debug_rports_30_addr ? mem_54 : _GEN_3253; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3255 = 6'h37 == io_debug_rports_30_addr ? mem_55 : _GEN_3254; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3256 = 6'h38 == io_debug_rports_30_addr ? mem_56 : _GEN_3255; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3257 = 6'h39 == io_debug_rports_30_addr ? mem_57 : _GEN_3256; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3258 = 6'h3a == io_debug_rports_30_addr ? mem_58 : _GEN_3257; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3259 = 6'h3b == io_debug_rports_30_addr ? mem_59 : _GEN_3258; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3260 = 6'h3c == io_debug_rports_30_addr ? mem_60 : _GEN_3259; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3261 = 6'h3d == io_debug_rports_30_addr ? mem_61 : _GEN_3260; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3262 = 6'h3e == io_debug_rports_30_addr ? mem_62 : _GEN_3261; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3263 = 6'h3f == io_debug_rports_30_addr ? mem_63 : _GEN_3262; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3265 = 6'h1 == io_debug_rports_31_addr ? mem_1 : mem_0; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3266 = 6'h2 == io_debug_rports_31_addr ? mem_2 : _GEN_3265; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3267 = 6'h3 == io_debug_rports_31_addr ? mem_3 : _GEN_3266; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3268 = 6'h4 == io_debug_rports_31_addr ? mem_4 : _GEN_3267; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3269 = 6'h5 == io_debug_rports_31_addr ? mem_5 : _GEN_3268; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3270 = 6'h6 == io_debug_rports_31_addr ? mem_6 : _GEN_3269; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3271 = 6'h7 == io_debug_rports_31_addr ? mem_7 : _GEN_3270; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3272 = 6'h8 == io_debug_rports_31_addr ? mem_8 : _GEN_3271; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3273 = 6'h9 == io_debug_rports_31_addr ? mem_9 : _GEN_3272; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3274 = 6'ha == io_debug_rports_31_addr ? mem_10 : _GEN_3273; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3275 = 6'hb == io_debug_rports_31_addr ? mem_11 : _GEN_3274; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3276 = 6'hc == io_debug_rports_31_addr ? mem_12 : _GEN_3275; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3277 = 6'hd == io_debug_rports_31_addr ? mem_13 : _GEN_3276; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3278 = 6'he == io_debug_rports_31_addr ? mem_14 : _GEN_3277; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3279 = 6'hf == io_debug_rports_31_addr ? mem_15 : _GEN_3278; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3280 = 6'h10 == io_debug_rports_31_addr ? mem_16 : _GEN_3279; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3281 = 6'h11 == io_debug_rports_31_addr ? mem_17 : _GEN_3280; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3282 = 6'h12 == io_debug_rports_31_addr ? mem_18 : _GEN_3281; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3283 = 6'h13 == io_debug_rports_31_addr ? mem_19 : _GEN_3282; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3284 = 6'h14 == io_debug_rports_31_addr ? mem_20 : _GEN_3283; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3285 = 6'h15 == io_debug_rports_31_addr ? mem_21 : _GEN_3284; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3286 = 6'h16 == io_debug_rports_31_addr ? mem_22 : _GEN_3285; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3287 = 6'h17 == io_debug_rports_31_addr ? mem_23 : _GEN_3286; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3288 = 6'h18 == io_debug_rports_31_addr ? mem_24 : _GEN_3287; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3289 = 6'h19 == io_debug_rports_31_addr ? mem_25 : _GEN_3288; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3290 = 6'h1a == io_debug_rports_31_addr ? mem_26 : _GEN_3289; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3291 = 6'h1b == io_debug_rports_31_addr ? mem_27 : _GEN_3290; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3292 = 6'h1c == io_debug_rports_31_addr ? mem_28 : _GEN_3291; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3293 = 6'h1d == io_debug_rports_31_addr ? mem_29 : _GEN_3292; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3294 = 6'h1e == io_debug_rports_31_addr ? mem_30 : _GEN_3293; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3295 = 6'h1f == io_debug_rports_31_addr ? mem_31 : _GEN_3294; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3296 = 6'h20 == io_debug_rports_31_addr ? mem_32 : _GEN_3295; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3297 = 6'h21 == io_debug_rports_31_addr ? mem_33 : _GEN_3296; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3298 = 6'h22 == io_debug_rports_31_addr ? mem_34 : _GEN_3297; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3299 = 6'h23 == io_debug_rports_31_addr ? mem_35 : _GEN_3298; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3300 = 6'h24 == io_debug_rports_31_addr ? mem_36 : _GEN_3299; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3301 = 6'h25 == io_debug_rports_31_addr ? mem_37 : _GEN_3300; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3302 = 6'h26 == io_debug_rports_31_addr ? mem_38 : _GEN_3301; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3303 = 6'h27 == io_debug_rports_31_addr ? mem_39 : _GEN_3302; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3304 = 6'h28 == io_debug_rports_31_addr ? mem_40 : _GEN_3303; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3305 = 6'h29 == io_debug_rports_31_addr ? mem_41 : _GEN_3304; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3306 = 6'h2a == io_debug_rports_31_addr ? mem_42 : _GEN_3305; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3307 = 6'h2b == io_debug_rports_31_addr ? mem_43 : _GEN_3306; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3308 = 6'h2c == io_debug_rports_31_addr ? mem_44 : _GEN_3307; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3309 = 6'h2d == io_debug_rports_31_addr ? mem_45 : _GEN_3308; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3310 = 6'h2e == io_debug_rports_31_addr ? mem_46 : _GEN_3309; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3311 = 6'h2f == io_debug_rports_31_addr ? mem_47 : _GEN_3310; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3312 = 6'h30 == io_debug_rports_31_addr ? mem_48 : _GEN_3311; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3313 = 6'h31 == io_debug_rports_31_addr ? mem_49 : _GEN_3312; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3314 = 6'h32 == io_debug_rports_31_addr ? mem_50 : _GEN_3313; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3315 = 6'h33 == io_debug_rports_31_addr ? mem_51 : _GEN_3314; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3316 = 6'h34 == io_debug_rports_31_addr ? mem_52 : _GEN_3315; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3317 = 6'h35 == io_debug_rports_31_addr ? mem_53 : _GEN_3316; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3318 = 6'h36 == io_debug_rports_31_addr ? mem_54 : _GEN_3317; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3319 = 6'h37 == io_debug_rports_31_addr ? mem_55 : _GEN_3318; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3320 = 6'h38 == io_debug_rports_31_addr ? mem_56 : _GEN_3319; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3321 = 6'h39 == io_debug_rports_31_addr ? mem_57 : _GEN_3320; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3322 = 6'h3a == io_debug_rports_31_addr ? mem_58 : _GEN_3321; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3323 = 6'h3b == io_debug_rports_31_addr ? mem_59 : _GEN_3322; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3324 = 6'h3c == io_debug_rports_31_addr ? mem_60 : _GEN_3323; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3325 = 6'h3d == io_debug_rports_31_addr ? mem_61 : _GEN_3324; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3326 = 6'h3e == io_debug_rports_31_addr ? mem_62 : _GEN_3325; // @[Regfile.scala 63:{25,25}]
  wire [63:0] _GEN_3327 = 6'h3f == io_debug_rports_31_addr ? mem_63 : _GEN_3326; // @[Regfile.scala 63:{25,25}]
  assign io_readPorts_0_data = io_readPorts_0_data_REG; // @[Regfile.scala 54:12]
  assign io_readPorts_1_data = io_readPorts_1_data_REG; // @[Regfile.scala 54:12]
  assign io_readPorts_2_data = io_readPorts_2_data_REG; // @[Regfile.scala 54:12]
  assign io_readPorts_3_data = io_readPorts_3_data_REG; // @[Regfile.scala 54:12]
  assign io_readPorts_4_data = io_readPorts_4_data_REG; // @[Regfile.scala 54:12]
  assign io_readPorts_5_data = io_readPorts_5_data_REG; // @[Regfile.scala 54:12]
  assign io_readPorts_6_data = io_readPorts_6_data_REG; // @[Regfile.scala 54:12]
  assign io_readPorts_7_data = io_readPorts_7_data_REG; // @[Regfile.scala 54:12]
  assign io_readPorts_8_data = io_readPorts_8_data_REG; // @[Regfile.scala 54:12]
  assign io_readPorts_9_data = io_readPorts_9_data_REG; // @[Regfile.scala 54:12]
  assign io_debug_rports_0_data = io_debug_rports_0_addr == 6'h0 ? 64'h0 : _GEN_1343; // @[Regfile.scala 63:25]
  assign io_debug_rports_1_data = io_debug_rports_1_addr == 6'h0 ? 64'h0 : _GEN_1407; // @[Regfile.scala 63:25]
  assign io_debug_rports_2_data = io_debug_rports_2_addr == 6'h0 ? 64'h0 : _GEN_1471; // @[Regfile.scala 63:25]
  assign io_debug_rports_3_data = io_debug_rports_3_addr == 6'h0 ? 64'h0 : _GEN_1535; // @[Regfile.scala 63:25]
  assign io_debug_rports_4_data = io_debug_rports_4_addr == 6'h0 ? 64'h0 : _GEN_1599; // @[Regfile.scala 63:25]
  assign io_debug_rports_5_data = io_debug_rports_5_addr == 6'h0 ? 64'h0 : _GEN_1663; // @[Regfile.scala 63:25]
  assign io_debug_rports_6_data = io_debug_rports_6_addr == 6'h0 ? 64'h0 : _GEN_1727; // @[Regfile.scala 63:25]
  assign io_debug_rports_7_data = io_debug_rports_7_addr == 6'h0 ? 64'h0 : _GEN_1791; // @[Regfile.scala 63:25]
  assign io_debug_rports_8_data = io_debug_rports_8_addr == 6'h0 ? 64'h0 : _GEN_1855; // @[Regfile.scala 63:25]
  assign io_debug_rports_9_data = io_debug_rports_9_addr == 6'h0 ? 64'h0 : _GEN_1919; // @[Regfile.scala 63:25]
  assign io_debug_rports_10_data = io_debug_rports_10_addr == 6'h0 ? 64'h0 : _GEN_1983; // @[Regfile.scala 63:25]
  assign io_debug_rports_11_data = io_debug_rports_11_addr == 6'h0 ? 64'h0 : _GEN_2047; // @[Regfile.scala 63:25]
  assign io_debug_rports_12_data = io_debug_rports_12_addr == 6'h0 ? 64'h0 : _GEN_2111; // @[Regfile.scala 63:25]
  assign io_debug_rports_13_data = io_debug_rports_13_addr == 6'h0 ? 64'h0 : _GEN_2175; // @[Regfile.scala 63:25]
  assign io_debug_rports_14_data = io_debug_rports_14_addr == 6'h0 ? 64'h0 : _GEN_2239; // @[Regfile.scala 63:25]
  assign io_debug_rports_15_data = io_debug_rports_15_addr == 6'h0 ? 64'h0 : _GEN_2303; // @[Regfile.scala 63:25]
  assign io_debug_rports_16_data = io_debug_rports_16_addr == 6'h0 ? 64'h0 : _GEN_2367; // @[Regfile.scala 63:25]
  assign io_debug_rports_17_data = io_debug_rports_17_addr == 6'h0 ? 64'h0 : _GEN_2431; // @[Regfile.scala 63:25]
  assign io_debug_rports_18_data = io_debug_rports_18_addr == 6'h0 ? 64'h0 : _GEN_2495; // @[Regfile.scala 63:25]
  assign io_debug_rports_19_data = io_debug_rports_19_addr == 6'h0 ? 64'h0 : _GEN_2559; // @[Regfile.scala 63:25]
  assign io_debug_rports_20_data = io_debug_rports_20_addr == 6'h0 ? 64'h0 : _GEN_2623; // @[Regfile.scala 63:25]
  assign io_debug_rports_21_data = io_debug_rports_21_addr == 6'h0 ? 64'h0 : _GEN_2687; // @[Regfile.scala 63:25]
  assign io_debug_rports_22_data = io_debug_rports_22_addr == 6'h0 ? 64'h0 : _GEN_2751; // @[Regfile.scala 63:25]
  assign io_debug_rports_23_data = io_debug_rports_23_addr == 6'h0 ? 64'h0 : _GEN_2815; // @[Regfile.scala 63:25]
  assign io_debug_rports_24_data = io_debug_rports_24_addr == 6'h0 ? 64'h0 : _GEN_2879; // @[Regfile.scala 63:25]
  assign io_debug_rports_25_data = io_debug_rports_25_addr == 6'h0 ? 64'h0 : _GEN_2943; // @[Regfile.scala 63:25]
  assign io_debug_rports_26_data = io_debug_rports_26_addr == 6'h0 ? 64'h0 : _GEN_3007; // @[Regfile.scala 63:25]
  assign io_debug_rports_27_data = io_debug_rports_27_addr == 6'h0 ? 64'h0 : _GEN_3071; // @[Regfile.scala 63:25]
  assign io_debug_rports_28_data = io_debug_rports_28_addr == 6'h0 ? 64'h0 : _GEN_3135; // @[Regfile.scala 63:25]
  assign io_debug_rports_29_data = io_debug_rports_29_addr == 6'h0 ? 64'h0 : _GEN_3199; // @[Regfile.scala 63:25]
  assign io_debug_rports_30_data = io_debug_rports_30_addr == 6'h0 ? 64'h0 : _GEN_3263; // @[Regfile.scala 63:25]
  assign io_debug_rports_31_data = io_debug_rports_31_addr == 6'h0 ? 64'h0 : _GEN_3327; // @[Regfile.scala 63:25]
  always @(posedge clock) begin
    if (io_writePorts_4_wen) begin // @[Regfile.scala 57:17]
      if (6'h0 == io_writePorts_4_addr) begin // @[Regfile.scala 58:19]
        mem_0 <= io_writePorts_4_data; // @[Regfile.scala 58:19]
      end else begin
        mem_0 <= _GEN_1088;
      end
    end else begin
      mem_0 <= _GEN_1088;
    end
    if (io_writePorts_4_wen) begin // @[Regfile.scala 57:17]
      if (6'h1 == io_writePorts_4_addr) begin // @[Regfile.scala 58:19]
        mem_1 <= io_writePorts_4_data; // @[Regfile.scala 58:19]
      end else begin
        mem_1 <= _GEN_1089;
      end
    end else begin
      mem_1 <= _GEN_1089;
    end
    if (io_writePorts_4_wen) begin // @[Regfile.scala 57:17]
      if (6'h2 == io_writePorts_4_addr) begin // @[Regfile.scala 58:19]
        mem_2 <= io_writePorts_4_data; // @[Regfile.scala 58:19]
      end else begin
        mem_2 <= _GEN_1090;
      end
    end else begin
      mem_2 <= _GEN_1090;
    end
    if (io_writePorts_4_wen) begin // @[Regfile.scala 57:17]
      if (6'h3 == io_writePorts_4_addr) begin // @[Regfile.scala 58:19]
        mem_3 <= io_writePorts_4_data; // @[Regfile.scala 58:19]
      end else begin
        mem_3 <= _GEN_1091;
      end
    end else begin
      mem_3 <= _GEN_1091;
    end
    if (io_writePorts_4_wen) begin // @[Regfile.scala 57:17]
      if (6'h4 == io_writePorts_4_addr) begin // @[Regfile.scala 58:19]
        mem_4 <= io_writePorts_4_data; // @[Regfile.scala 58:19]
      end else begin
        mem_4 <= _GEN_1092;
      end
    end else begin
      mem_4 <= _GEN_1092;
    end
    if (io_writePorts_4_wen) begin // @[Regfile.scala 57:17]
      if (6'h5 == io_writePorts_4_addr) begin // @[Regfile.scala 58:19]
        mem_5 <= io_writePorts_4_data; // @[Regfile.scala 58:19]
      end else begin
        mem_5 <= _GEN_1093;
      end
    end else begin
      mem_5 <= _GEN_1093;
    end
    if (io_writePorts_4_wen) begin // @[Regfile.scala 57:17]
      if (6'h6 == io_writePorts_4_addr) begin // @[Regfile.scala 58:19]
        mem_6 <= io_writePorts_4_data; // @[Regfile.scala 58:19]
      end else begin
        mem_6 <= _GEN_1094;
      end
    end else begin
      mem_6 <= _GEN_1094;
    end
    if (io_writePorts_4_wen) begin // @[Regfile.scala 57:17]
      if (6'h7 == io_writePorts_4_addr) begin // @[Regfile.scala 58:19]
        mem_7 <= io_writePorts_4_data; // @[Regfile.scala 58:19]
      end else begin
        mem_7 <= _GEN_1095;
      end
    end else begin
      mem_7 <= _GEN_1095;
    end
    if (io_writePorts_4_wen) begin // @[Regfile.scala 57:17]
      if (6'h8 == io_writePorts_4_addr) begin // @[Regfile.scala 58:19]
        mem_8 <= io_writePorts_4_data; // @[Regfile.scala 58:19]
      end else begin
        mem_8 <= _GEN_1096;
      end
    end else begin
      mem_8 <= _GEN_1096;
    end
    if (io_writePorts_4_wen) begin // @[Regfile.scala 57:17]
      if (6'h9 == io_writePorts_4_addr) begin // @[Regfile.scala 58:19]
        mem_9 <= io_writePorts_4_data; // @[Regfile.scala 58:19]
      end else begin
        mem_9 <= _GEN_1097;
      end
    end else begin
      mem_9 <= _GEN_1097;
    end
    if (io_writePorts_4_wen) begin // @[Regfile.scala 57:17]
      if (6'ha == io_writePorts_4_addr) begin // @[Regfile.scala 58:19]
        mem_10 <= io_writePorts_4_data; // @[Regfile.scala 58:19]
      end else begin
        mem_10 <= _GEN_1098;
      end
    end else begin
      mem_10 <= _GEN_1098;
    end
    if (io_writePorts_4_wen) begin // @[Regfile.scala 57:17]
      if (6'hb == io_writePorts_4_addr) begin // @[Regfile.scala 58:19]
        mem_11 <= io_writePorts_4_data; // @[Regfile.scala 58:19]
      end else begin
        mem_11 <= _GEN_1099;
      end
    end else begin
      mem_11 <= _GEN_1099;
    end
    if (io_writePorts_4_wen) begin // @[Regfile.scala 57:17]
      if (6'hc == io_writePorts_4_addr) begin // @[Regfile.scala 58:19]
        mem_12 <= io_writePorts_4_data; // @[Regfile.scala 58:19]
      end else begin
        mem_12 <= _GEN_1100;
      end
    end else begin
      mem_12 <= _GEN_1100;
    end
    if (io_writePorts_4_wen) begin // @[Regfile.scala 57:17]
      if (6'hd == io_writePorts_4_addr) begin // @[Regfile.scala 58:19]
        mem_13 <= io_writePorts_4_data; // @[Regfile.scala 58:19]
      end else begin
        mem_13 <= _GEN_1101;
      end
    end else begin
      mem_13 <= _GEN_1101;
    end
    if (io_writePorts_4_wen) begin // @[Regfile.scala 57:17]
      if (6'he == io_writePorts_4_addr) begin // @[Regfile.scala 58:19]
        mem_14 <= io_writePorts_4_data; // @[Regfile.scala 58:19]
      end else begin
        mem_14 <= _GEN_1102;
      end
    end else begin
      mem_14 <= _GEN_1102;
    end
    if (io_writePorts_4_wen) begin // @[Regfile.scala 57:17]
      if (6'hf == io_writePorts_4_addr) begin // @[Regfile.scala 58:19]
        mem_15 <= io_writePorts_4_data; // @[Regfile.scala 58:19]
      end else begin
        mem_15 <= _GEN_1103;
      end
    end else begin
      mem_15 <= _GEN_1103;
    end
    if (io_writePorts_4_wen) begin // @[Regfile.scala 57:17]
      if (6'h10 == io_writePorts_4_addr) begin // @[Regfile.scala 58:19]
        mem_16 <= io_writePorts_4_data; // @[Regfile.scala 58:19]
      end else begin
        mem_16 <= _GEN_1104;
      end
    end else begin
      mem_16 <= _GEN_1104;
    end
    if (io_writePorts_4_wen) begin // @[Regfile.scala 57:17]
      if (6'h11 == io_writePorts_4_addr) begin // @[Regfile.scala 58:19]
        mem_17 <= io_writePorts_4_data; // @[Regfile.scala 58:19]
      end else begin
        mem_17 <= _GEN_1105;
      end
    end else begin
      mem_17 <= _GEN_1105;
    end
    if (io_writePorts_4_wen) begin // @[Regfile.scala 57:17]
      if (6'h12 == io_writePorts_4_addr) begin // @[Regfile.scala 58:19]
        mem_18 <= io_writePorts_4_data; // @[Regfile.scala 58:19]
      end else begin
        mem_18 <= _GEN_1106;
      end
    end else begin
      mem_18 <= _GEN_1106;
    end
    if (io_writePorts_4_wen) begin // @[Regfile.scala 57:17]
      if (6'h13 == io_writePorts_4_addr) begin // @[Regfile.scala 58:19]
        mem_19 <= io_writePorts_4_data; // @[Regfile.scala 58:19]
      end else begin
        mem_19 <= _GEN_1107;
      end
    end else begin
      mem_19 <= _GEN_1107;
    end
    if (io_writePorts_4_wen) begin // @[Regfile.scala 57:17]
      if (6'h14 == io_writePorts_4_addr) begin // @[Regfile.scala 58:19]
        mem_20 <= io_writePorts_4_data; // @[Regfile.scala 58:19]
      end else begin
        mem_20 <= _GEN_1108;
      end
    end else begin
      mem_20 <= _GEN_1108;
    end
    if (io_writePorts_4_wen) begin // @[Regfile.scala 57:17]
      if (6'h15 == io_writePorts_4_addr) begin // @[Regfile.scala 58:19]
        mem_21 <= io_writePorts_4_data; // @[Regfile.scala 58:19]
      end else begin
        mem_21 <= _GEN_1109;
      end
    end else begin
      mem_21 <= _GEN_1109;
    end
    if (io_writePorts_4_wen) begin // @[Regfile.scala 57:17]
      if (6'h16 == io_writePorts_4_addr) begin // @[Regfile.scala 58:19]
        mem_22 <= io_writePorts_4_data; // @[Regfile.scala 58:19]
      end else begin
        mem_22 <= _GEN_1110;
      end
    end else begin
      mem_22 <= _GEN_1110;
    end
    if (io_writePorts_4_wen) begin // @[Regfile.scala 57:17]
      if (6'h17 == io_writePorts_4_addr) begin // @[Regfile.scala 58:19]
        mem_23 <= io_writePorts_4_data; // @[Regfile.scala 58:19]
      end else begin
        mem_23 <= _GEN_1111;
      end
    end else begin
      mem_23 <= _GEN_1111;
    end
    if (io_writePorts_4_wen) begin // @[Regfile.scala 57:17]
      if (6'h18 == io_writePorts_4_addr) begin // @[Regfile.scala 58:19]
        mem_24 <= io_writePorts_4_data; // @[Regfile.scala 58:19]
      end else begin
        mem_24 <= _GEN_1112;
      end
    end else begin
      mem_24 <= _GEN_1112;
    end
    if (io_writePorts_4_wen) begin // @[Regfile.scala 57:17]
      if (6'h19 == io_writePorts_4_addr) begin // @[Regfile.scala 58:19]
        mem_25 <= io_writePorts_4_data; // @[Regfile.scala 58:19]
      end else begin
        mem_25 <= _GEN_1113;
      end
    end else begin
      mem_25 <= _GEN_1113;
    end
    if (io_writePorts_4_wen) begin // @[Regfile.scala 57:17]
      if (6'h1a == io_writePorts_4_addr) begin // @[Regfile.scala 58:19]
        mem_26 <= io_writePorts_4_data; // @[Regfile.scala 58:19]
      end else begin
        mem_26 <= _GEN_1114;
      end
    end else begin
      mem_26 <= _GEN_1114;
    end
    if (io_writePorts_4_wen) begin // @[Regfile.scala 57:17]
      if (6'h1b == io_writePorts_4_addr) begin // @[Regfile.scala 58:19]
        mem_27 <= io_writePorts_4_data; // @[Regfile.scala 58:19]
      end else begin
        mem_27 <= _GEN_1115;
      end
    end else begin
      mem_27 <= _GEN_1115;
    end
    if (io_writePorts_4_wen) begin // @[Regfile.scala 57:17]
      if (6'h1c == io_writePorts_4_addr) begin // @[Regfile.scala 58:19]
        mem_28 <= io_writePorts_4_data; // @[Regfile.scala 58:19]
      end else begin
        mem_28 <= _GEN_1116;
      end
    end else begin
      mem_28 <= _GEN_1116;
    end
    if (io_writePorts_4_wen) begin // @[Regfile.scala 57:17]
      if (6'h1d == io_writePorts_4_addr) begin // @[Regfile.scala 58:19]
        mem_29 <= io_writePorts_4_data; // @[Regfile.scala 58:19]
      end else begin
        mem_29 <= _GEN_1117;
      end
    end else begin
      mem_29 <= _GEN_1117;
    end
    if (io_writePorts_4_wen) begin // @[Regfile.scala 57:17]
      if (6'h1e == io_writePorts_4_addr) begin // @[Regfile.scala 58:19]
        mem_30 <= io_writePorts_4_data; // @[Regfile.scala 58:19]
      end else begin
        mem_30 <= _GEN_1118;
      end
    end else begin
      mem_30 <= _GEN_1118;
    end
    if (io_writePorts_4_wen) begin // @[Regfile.scala 57:17]
      if (6'h1f == io_writePorts_4_addr) begin // @[Regfile.scala 58:19]
        mem_31 <= io_writePorts_4_data; // @[Regfile.scala 58:19]
      end else begin
        mem_31 <= _GEN_1119;
      end
    end else begin
      mem_31 <= _GEN_1119;
    end
    if (io_writePorts_4_wen) begin // @[Regfile.scala 57:17]
      if (6'h20 == io_writePorts_4_addr) begin // @[Regfile.scala 58:19]
        mem_32 <= io_writePorts_4_data; // @[Regfile.scala 58:19]
      end else begin
        mem_32 <= _GEN_1120;
      end
    end else begin
      mem_32 <= _GEN_1120;
    end
    if (io_writePorts_4_wen) begin // @[Regfile.scala 57:17]
      if (6'h21 == io_writePorts_4_addr) begin // @[Regfile.scala 58:19]
        mem_33 <= io_writePorts_4_data; // @[Regfile.scala 58:19]
      end else begin
        mem_33 <= _GEN_1121;
      end
    end else begin
      mem_33 <= _GEN_1121;
    end
    if (io_writePorts_4_wen) begin // @[Regfile.scala 57:17]
      if (6'h22 == io_writePorts_4_addr) begin // @[Regfile.scala 58:19]
        mem_34 <= io_writePorts_4_data; // @[Regfile.scala 58:19]
      end else begin
        mem_34 <= _GEN_1122;
      end
    end else begin
      mem_34 <= _GEN_1122;
    end
    if (io_writePorts_4_wen) begin // @[Regfile.scala 57:17]
      if (6'h23 == io_writePorts_4_addr) begin // @[Regfile.scala 58:19]
        mem_35 <= io_writePorts_4_data; // @[Regfile.scala 58:19]
      end else begin
        mem_35 <= _GEN_1123;
      end
    end else begin
      mem_35 <= _GEN_1123;
    end
    if (io_writePorts_4_wen) begin // @[Regfile.scala 57:17]
      if (6'h24 == io_writePorts_4_addr) begin // @[Regfile.scala 58:19]
        mem_36 <= io_writePorts_4_data; // @[Regfile.scala 58:19]
      end else begin
        mem_36 <= _GEN_1124;
      end
    end else begin
      mem_36 <= _GEN_1124;
    end
    if (io_writePorts_4_wen) begin // @[Regfile.scala 57:17]
      if (6'h25 == io_writePorts_4_addr) begin // @[Regfile.scala 58:19]
        mem_37 <= io_writePorts_4_data; // @[Regfile.scala 58:19]
      end else begin
        mem_37 <= _GEN_1125;
      end
    end else begin
      mem_37 <= _GEN_1125;
    end
    if (io_writePorts_4_wen) begin // @[Regfile.scala 57:17]
      if (6'h26 == io_writePorts_4_addr) begin // @[Regfile.scala 58:19]
        mem_38 <= io_writePorts_4_data; // @[Regfile.scala 58:19]
      end else begin
        mem_38 <= _GEN_1126;
      end
    end else begin
      mem_38 <= _GEN_1126;
    end
    if (io_writePorts_4_wen) begin // @[Regfile.scala 57:17]
      if (6'h27 == io_writePorts_4_addr) begin // @[Regfile.scala 58:19]
        mem_39 <= io_writePorts_4_data; // @[Regfile.scala 58:19]
      end else begin
        mem_39 <= _GEN_1127;
      end
    end else begin
      mem_39 <= _GEN_1127;
    end
    if (io_writePorts_4_wen) begin // @[Regfile.scala 57:17]
      if (6'h28 == io_writePorts_4_addr) begin // @[Regfile.scala 58:19]
        mem_40 <= io_writePorts_4_data; // @[Regfile.scala 58:19]
      end else begin
        mem_40 <= _GEN_1128;
      end
    end else begin
      mem_40 <= _GEN_1128;
    end
    if (io_writePorts_4_wen) begin // @[Regfile.scala 57:17]
      if (6'h29 == io_writePorts_4_addr) begin // @[Regfile.scala 58:19]
        mem_41 <= io_writePorts_4_data; // @[Regfile.scala 58:19]
      end else begin
        mem_41 <= _GEN_1129;
      end
    end else begin
      mem_41 <= _GEN_1129;
    end
    if (io_writePorts_4_wen) begin // @[Regfile.scala 57:17]
      if (6'h2a == io_writePorts_4_addr) begin // @[Regfile.scala 58:19]
        mem_42 <= io_writePorts_4_data; // @[Regfile.scala 58:19]
      end else begin
        mem_42 <= _GEN_1130;
      end
    end else begin
      mem_42 <= _GEN_1130;
    end
    if (io_writePorts_4_wen) begin // @[Regfile.scala 57:17]
      if (6'h2b == io_writePorts_4_addr) begin // @[Regfile.scala 58:19]
        mem_43 <= io_writePorts_4_data; // @[Regfile.scala 58:19]
      end else begin
        mem_43 <= _GEN_1131;
      end
    end else begin
      mem_43 <= _GEN_1131;
    end
    if (io_writePorts_4_wen) begin // @[Regfile.scala 57:17]
      if (6'h2c == io_writePorts_4_addr) begin // @[Regfile.scala 58:19]
        mem_44 <= io_writePorts_4_data; // @[Regfile.scala 58:19]
      end else begin
        mem_44 <= _GEN_1132;
      end
    end else begin
      mem_44 <= _GEN_1132;
    end
    if (io_writePorts_4_wen) begin // @[Regfile.scala 57:17]
      if (6'h2d == io_writePorts_4_addr) begin // @[Regfile.scala 58:19]
        mem_45 <= io_writePorts_4_data; // @[Regfile.scala 58:19]
      end else begin
        mem_45 <= _GEN_1133;
      end
    end else begin
      mem_45 <= _GEN_1133;
    end
    if (io_writePorts_4_wen) begin // @[Regfile.scala 57:17]
      if (6'h2e == io_writePorts_4_addr) begin // @[Regfile.scala 58:19]
        mem_46 <= io_writePorts_4_data; // @[Regfile.scala 58:19]
      end else begin
        mem_46 <= _GEN_1134;
      end
    end else begin
      mem_46 <= _GEN_1134;
    end
    if (io_writePorts_4_wen) begin // @[Regfile.scala 57:17]
      if (6'h2f == io_writePorts_4_addr) begin // @[Regfile.scala 58:19]
        mem_47 <= io_writePorts_4_data; // @[Regfile.scala 58:19]
      end else begin
        mem_47 <= _GEN_1135;
      end
    end else begin
      mem_47 <= _GEN_1135;
    end
    if (io_writePorts_4_wen) begin // @[Regfile.scala 57:17]
      if (6'h30 == io_writePorts_4_addr) begin // @[Regfile.scala 58:19]
        mem_48 <= io_writePorts_4_data; // @[Regfile.scala 58:19]
      end else begin
        mem_48 <= _GEN_1136;
      end
    end else begin
      mem_48 <= _GEN_1136;
    end
    if (io_writePorts_4_wen) begin // @[Regfile.scala 57:17]
      if (6'h31 == io_writePorts_4_addr) begin // @[Regfile.scala 58:19]
        mem_49 <= io_writePorts_4_data; // @[Regfile.scala 58:19]
      end else begin
        mem_49 <= _GEN_1137;
      end
    end else begin
      mem_49 <= _GEN_1137;
    end
    if (io_writePorts_4_wen) begin // @[Regfile.scala 57:17]
      if (6'h32 == io_writePorts_4_addr) begin // @[Regfile.scala 58:19]
        mem_50 <= io_writePorts_4_data; // @[Regfile.scala 58:19]
      end else begin
        mem_50 <= _GEN_1138;
      end
    end else begin
      mem_50 <= _GEN_1138;
    end
    if (io_writePorts_4_wen) begin // @[Regfile.scala 57:17]
      if (6'h33 == io_writePorts_4_addr) begin // @[Regfile.scala 58:19]
        mem_51 <= io_writePorts_4_data; // @[Regfile.scala 58:19]
      end else begin
        mem_51 <= _GEN_1139;
      end
    end else begin
      mem_51 <= _GEN_1139;
    end
    if (io_writePorts_4_wen) begin // @[Regfile.scala 57:17]
      if (6'h34 == io_writePorts_4_addr) begin // @[Regfile.scala 58:19]
        mem_52 <= io_writePorts_4_data; // @[Regfile.scala 58:19]
      end else begin
        mem_52 <= _GEN_1140;
      end
    end else begin
      mem_52 <= _GEN_1140;
    end
    if (io_writePorts_4_wen) begin // @[Regfile.scala 57:17]
      if (6'h35 == io_writePorts_4_addr) begin // @[Regfile.scala 58:19]
        mem_53 <= io_writePorts_4_data; // @[Regfile.scala 58:19]
      end else begin
        mem_53 <= _GEN_1141;
      end
    end else begin
      mem_53 <= _GEN_1141;
    end
    if (io_writePorts_4_wen) begin // @[Regfile.scala 57:17]
      if (6'h36 == io_writePorts_4_addr) begin // @[Regfile.scala 58:19]
        mem_54 <= io_writePorts_4_data; // @[Regfile.scala 58:19]
      end else begin
        mem_54 <= _GEN_1142;
      end
    end else begin
      mem_54 <= _GEN_1142;
    end
    if (io_writePorts_4_wen) begin // @[Regfile.scala 57:17]
      if (6'h37 == io_writePorts_4_addr) begin // @[Regfile.scala 58:19]
        mem_55 <= io_writePorts_4_data; // @[Regfile.scala 58:19]
      end else begin
        mem_55 <= _GEN_1143;
      end
    end else begin
      mem_55 <= _GEN_1143;
    end
    if (io_writePorts_4_wen) begin // @[Regfile.scala 57:17]
      if (6'h38 == io_writePorts_4_addr) begin // @[Regfile.scala 58:19]
        mem_56 <= io_writePorts_4_data; // @[Regfile.scala 58:19]
      end else begin
        mem_56 <= _GEN_1144;
      end
    end else begin
      mem_56 <= _GEN_1144;
    end
    if (io_writePorts_4_wen) begin // @[Regfile.scala 57:17]
      if (6'h39 == io_writePorts_4_addr) begin // @[Regfile.scala 58:19]
        mem_57 <= io_writePorts_4_data; // @[Regfile.scala 58:19]
      end else begin
        mem_57 <= _GEN_1145;
      end
    end else begin
      mem_57 <= _GEN_1145;
    end
    if (io_writePorts_4_wen) begin // @[Regfile.scala 57:17]
      if (6'h3a == io_writePorts_4_addr) begin // @[Regfile.scala 58:19]
        mem_58 <= io_writePorts_4_data; // @[Regfile.scala 58:19]
      end else begin
        mem_58 <= _GEN_1146;
      end
    end else begin
      mem_58 <= _GEN_1146;
    end
    if (io_writePorts_4_wen) begin // @[Regfile.scala 57:17]
      if (6'h3b == io_writePorts_4_addr) begin // @[Regfile.scala 58:19]
        mem_59 <= io_writePorts_4_data; // @[Regfile.scala 58:19]
      end else begin
        mem_59 <= _GEN_1147;
      end
    end else begin
      mem_59 <= _GEN_1147;
    end
    if (io_writePorts_4_wen) begin // @[Regfile.scala 57:17]
      if (6'h3c == io_writePorts_4_addr) begin // @[Regfile.scala 58:19]
        mem_60 <= io_writePorts_4_data; // @[Regfile.scala 58:19]
      end else begin
        mem_60 <= _GEN_1148;
      end
    end else begin
      mem_60 <= _GEN_1148;
    end
    if (io_writePorts_4_wen) begin // @[Regfile.scala 57:17]
      if (6'h3d == io_writePorts_4_addr) begin // @[Regfile.scala 58:19]
        mem_61 <= io_writePorts_4_data; // @[Regfile.scala 58:19]
      end else begin
        mem_61 <= _GEN_1149;
      end
    end else begin
      mem_61 <= _GEN_1149;
    end
    if (io_writePorts_4_wen) begin // @[Regfile.scala 57:17]
      if (6'h3e == io_writePorts_4_addr) begin // @[Regfile.scala 58:19]
        mem_62 <= io_writePorts_4_data; // @[Regfile.scala 58:19]
      end else begin
        mem_62 <= _GEN_1150;
      end
    end else begin
      mem_62 <= _GEN_1150;
    end
    if (io_writePorts_4_wen) begin // @[Regfile.scala 57:17]
      if (6'h3f == io_writePorts_4_addr) begin // @[Regfile.scala 58:19]
        mem_63 <= io_writePorts_4_data; // @[Regfile.scala 58:19]
      end else begin
        mem_63 <= _GEN_1151;
      end
    end else begin
      mem_63 <= _GEN_1151;
    end
    if (io_readPorts_0_addr == 6'h0) begin // @[Regfile.scala 53:33]
      io_readPorts_0_data_REG <= 64'h0;
    end else if (6'h3f == io_readPorts_0_addr) begin // @[Regfile.scala 53:33]
      io_readPorts_0_data_REG <= mem_63; // @[Regfile.scala 53:33]
    end else if (6'h3e == io_readPorts_0_addr) begin // @[Regfile.scala 53:33]
      io_readPorts_0_data_REG <= mem_62; // @[Regfile.scala 53:33]
    end else if (6'h3d == io_readPorts_0_addr) begin // @[Regfile.scala 53:33]
      io_readPorts_0_data_REG <= mem_61; // @[Regfile.scala 53:33]
    end else begin
      io_readPorts_0_data_REG <= _GEN_60;
    end
    if (io_readPorts_1_addr == 6'h0) begin // @[Regfile.scala 53:33]
      io_readPorts_1_data_REG <= 64'h0;
    end else if (6'h3f == io_readPorts_1_addr) begin // @[Regfile.scala 53:33]
      io_readPorts_1_data_REG <= mem_63; // @[Regfile.scala 53:33]
    end else if (6'h3e == io_readPorts_1_addr) begin // @[Regfile.scala 53:33]
      io_readPorts_1_data_REG <= mem_62; // @[Regfile.scala 53:33]
    end else if (6'h3d == io_readPorts_1_addr) begin // @[Regfile.scala 53:33]
      io_readPorts_1_data_REG <= mem_61; // @[Regfile.scala 53:33]
    end else begin
      io_readPorts_1_data_REG <= _GEN_124;
    end
    if (io_readPorts_2_addr == 6'h0) begin // @[Regfile.scala 53:33]
      io_readPorts_2_data_REG <= 64'h0;
    end else if (6'h3f == io_readPorts_2_addr) begin // @[Regfile.scala 53:33]
      io_readPorts_2_data_REG <= mem_63; // @[Regfile.scala 53:33]
    end else if (6'h3e == io_readPorts_2_addr) begin // @[Regfile.scala 53:33]
      io_readPorts_2_data_REG <= mem_62; // @[Regfile.scala 53:33]
    end else if (6'h3d == io_readPorts_2_addr) begin // @[Regfile.scala 53:33]
      io_readPorts_2_data_REG <= mem_61; // @[Regfile.scala 53:33]
    end else begin
      io_readPorts_2_data_REG <= _GEN_188;
    end
    if (io_readPorts_3_addr == 6'h0) begin // @[Regfile.scala 53:33]
      io_readPorts_3_data_REG <= 64'h0;
    end else if (6'h3f == io_readPorts_3_addr) begin // @[Regfile.scala 53:33]
      io_readPorts_3_data_REG <= mem_63; // @[Regfile.scala 53:33]
    end else if (6'h3e == io_readPorts_3_addr) begin // @[Regfile.scala 53:33]
      io_readPorts_3_data_REG <= mem_62; // @[Regfile.scala 53:33]
    end else if (6'h3d == io_readPorts_3_addr) begin // @[Regfile.scala 53:33]
      io_readPorts_3_data_REG <= mem_61; // @[Regfile.scala 53:33]
    end else begin
      io_readPorts_3_data_REG <= _GEN_252;
    end
    if (io_readPorts_4_addr == 6'h0) begin // @[Regfile.scala 53:33]
      io_readPorts_4_data_REG <= 64'h0;
    end else if (6'h3f == io_readPorts_4_addr) begin // @[Regfile.scala 53:33]
      io_readPorts_4_data_REG <= mem_63; // @[Regfile.scala 53:33]
    end else if (6'h3e == io_readPorts_4_addr) begin // @[Regfile.scala 53:33]
      io_readPorts_4_data_REG <= mem_62; // @[Regfile.scala 53:33]
    end else if (6'h3d == io_readPorts_4_addr) begin // @[Regfile.scala 53:33]
      io_readPorts_4_data_REG <= mem_61; // @[Regfile.scala 53:33]
    end else begin
      io_readPorts_4_data_REG <= _GEN_316;
    end
    if (io_readPorts_5_addr == 6'h0) begin // @[Regfile.scala 53:33]
      io_readPorts_5_data_REG <= 64'h0;
    end else if (6'h3f == io_readPorts_5_addr) begin // @[Regfile.scala 53:33]
      io_readPorts_5_data_REG <= mem_63; // @[Regfile.scala 53:33]
    end else if (6'h3e == io_readPorts_5_addr) begin // @[Regfile.scala 53:33]
      io_readPorts_5_data_REG <= mem_62; // @[Regfile.scala 53:33]
    end else if (6'h3d == io_readPorts_5_addr) begin // @[Regfile.scala 53:33]
      io_readPorts_5_data_REG <= mem_61; // @[Regfile.scala 53:33]
    end else begin
      io_readPorts_5_data_REG <= _GEN_380;
    end
    if (io_readPorts_6_addr == 6'h0) begin // @[Regfile.scala 53:33]
      io_readPorts_6_data_REG <= 64'h0;
    end else if (6'h3f == io_readPorts_6_addr) begin // @[Regfile.scala 53:33]
      io_readPorts_6_data_REG <= mem_63; // @[Regfile.scala 53:33]
    end else if (6'h3e == io_readPorts_6_addr) begin // @[Regfile.scala 53:33]
      io_readPorts_6_data_REG <= mem_62; // @[Regfile.scala 53:33]
    end else if (6'h3d == io_readPorts_6_addr) begin // @[Regfile.scala 53:33]
      io_readPorts_6_data_REG <= mem_61; // @[Regfile.scala 53:33]
    end else begin
      io_readPorts_6_data_REG <= _GEN_444;
    end
    if (io_readPorts_7_addr == 6'h0) begin // @[Regfile.scala 53:33]
      io_readPorts_7_data_REG <= 64'h0;
    end else if (6'h3f == io_readPorts_7_addr) begin // @[Regfile.scala 53:33]
      io_readPorts_7_data_REG <= mem_63; // @[Regfile.scala 53:33]
    end else if (6'h3e == io_readPorts_7_addr) begin // @[Regfile.scala 53:33]
      io_readPorts_7_data_REG <= mem_62; // @[Regfile.scala 53:33]
    end else if (6'h3d == io_readPorts_7_addr) begin // @[Regfile.scala 53:33]
      io_readPorts_7_data_REG <= mem_61; // @[Regfile.scala 53:33]
    end else begin
      io_readPorts_7_data_REG <= _GEN_508;
    end
    if (io_readPorts_8_addr == 6'h0) begin // @[Regfile.scala 53:33]
      io_readPorts_8_data_REG <= 64'h0;
    end else if (6'h3f == io_readPorts_8_addr) begin // @[Regfile.scala 53:33]
      io_readPorts_8_data_REG <= mem_63; // @[Regfile.scala 53:33]
    end else if (6'h3e == io_readPorts_8_addr) begin // @[Regfile.scala 53:33]
      io_readPorts_8_data_REG <= mem_62; // @[Regfile.scala 53:33]
    end else if (6'h3d == io_readPorts_8_addr) begin // @[Regfile.scala 53:33]
      io_readPorts_8_data_REG <= mem_61; // @[Regfile.scala 53:33]
    end else begin
      io_readPorts_8_data_REG <= _GEN_572;
    end
    if (io_readPorts_9_addr == 6'h0) begin // @[Regfile.scala 53:33]
      io_readPorts_9_data_REG <= 64'h0;
    end else if (6'h3f == io_readPorts_9_addr) begin // @[Regfile.scala 53:33]
      io_readPorts_9_data_REG <= mem_63; // @[Regfile.scala 53:33]
    end else if (6'h3e == io_readPorts_9_addr) begin // @[Regfile.scala 53:33]
      io_readPorts_9_data_REG <= mem_62; // @[Regfile.scala 53:33]
    end else if (6'h3d == io_readPorts_9_addr) begin // @[Regfile.scala 53:33]
      io_readPorts_9_data_REG <= mem_61; // @[Regfile.scala 53:33]
    end else begin
      io_readPorts_9_data_REG <= _GEN_636;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  mem_0 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  mem_1 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  mem_2 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  mem_3 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  mem_4 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  mem_5 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  mem_6 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  mem_7 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  mem_8 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  mem_9 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  mem_10 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  mem_11 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  mem_12 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  mem_13 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  mem_14 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  mem_15 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  mem_16 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  mem_17 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  mem_18 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  mem_19 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  mem_20 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  mem_21 = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  mem_22 = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  mem_23 = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  mem_24 = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  mem_25 = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  mem_26 = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  mem_27 = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  mem_28 = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  mem_29 = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  mem_30 = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  mem_31 = _RAND_31[63:0];
  _RAND_32 = {2{`RANDOM}};
  mem_32 = _RAND_32[63:0];
  _RAND_33 = {2{`RANDOM}};
  mem_33 = _RAND_33[63:0];
  _RAND_34 = {2{`RANDOM}};
  mem_34 = _RAND_34[63:0];
  _RAND_35 = {2{`RANDOM}};
  mem_35 = _RAND_35[63:0];
  _RAND_36 = {2{`RANDOM}};
  mem_36 = _RAND_36[63:0];
  _RAND_37 = {2{`RANDOM}};
  mem_37 = _RAND_37[63:0];
  _RAND_38 = {2{`RANDOM}};
  mem_38 = _RAND_38[63:0];
  _RAND_39 = {2{`RANDOM}};
  mem_39 = _RAND_39[63:0];
  _RAND_40 = {2{`RANDOM}};
  mem_40 = _RAND_40[63:0];
  _RAND_41 = {2{`RANDOM}};
  mem_41 = _RAND_41[63:0];
  _RAND_42 = {2{`RANDOM}};
  mem_42 = _RAND_42[63:0];
  _RAND_43 = {2{`RANDOM}};
  mem_43 = _RAND_43[63:0];
  _RAND_44 = {2{`RANDOM}};
  mem_44 = _RAND_44[63:0];
  _RAND_45 = {2{`RANDOM}};
  mem_45 = _RAND_45[63:0];
  _RAND_46 = {2{`RANDOM}};
  mem_46 = _RAND_46[63:0];
  _RAND_47 = {2{`RANDOM}};
  mem_47 = _RAND_47[63:0];
  _RAND_48 = {2{`RANDOM}};
  mem_48 = _RAND_48[63:0];
  _RAND_49 = {2{`RANDOM}};
  mem_49 = _RAND_49[63:0];
  _RAND_50 = {2{`RANDOM}};
  mem_50 = _RAND_50[63:0];
  _RAND_51 = {2{`RANDOM}};
  mem_51 = _RAND_51[63:0];
  _RAND_52 = {2{`RANDOM}};
  mem_52 = _RAND_52[63:0];
  _RAND_53 = {2{`RANDOM}};
  mem_53 = _RAND_53[63:0];
  _RAND_54 = {2{`RANDOM}};
  mem_54 = _RAND_54[63:0];
  _RAND_55 = {2{`RANDOM}};
  mem_55 = _RAND_55[63:0];
  _RAND_56 = {2{`RANDOM}};
  mem_56 = _RAND_56[63:0];
  _RAND_57 = {2{`RANDOM}};
  mem_57 = _RAND_57[63:0];
  _RAND_58 = {2{`RANDOM}};
  mem_58 = _RAND_58[63:0];
  _RAND_59 = {2{`RANDOM}};
  mem_59 = _RAND_59[63:0];
  _RAND_60 = {2{`RANDOM}};
  mem_60 = _RAND_60[63:0];
  _RAND_61 = {2{`RANDOM}};
  mem_61 = _RAND_61[63:0];
  _RAND_62 = {2{`RANDOM}};
  mem_62 = _RAND_62[63:0];
  _RAND_63 = {2{`RANDOM}};
  mem_63 = _RAND_63[63:0];
  _RAND_64 = {2{`RANDOM}};
  io_readPorts_0_data_REG = _RAND_64[63:0];
  _RAND_65 = {2{`RANDOM}};
  io_readPorts_1_data_REG = _RAND_65[63:0];
  _RAND_66 = {2{`RANDOM}};
  io_readPorts_2_data_REG = _RAND_66[63:0];
  _RAND_67 = {2{`RANDOM}};
  io_readPorts_3_data_REG = _RAND_67[63:0];
  _RAND_68 = {2{`RANDOM}};
  io_readPorts_4_data_REG = _RAND_68[63:0];
  _RAND_69 = {2{`RANDOM}};
  io_readPorts_5_data_REG = _RAND_69[63:0];
  _RAND_70 = {2{`RANDOM}};
  io_readPorts_6_data_REG = _RAND_70[63:0];
  _RAND_71 = {2{`RANDOM}};
  io_readPorts_7_data_REG = _RAND_71[63:0];
  _RAND_72 = {2{`RANDOM}};
  io_readPorts_8_data_REG = _RAND_72[63:0];
  _RAND_73 = {2{`RANDOM}};
  io_readPorts_9_data_REG = _RAND_73[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule

