module DelayN_118(
  input  [38:0] io_in,
  output [38:0] io_out
);
  assign io_out = io_in; // @[Hold.scala 92:10]
endmodule

