module bosc_xsl2_ultiscan_top(
  output          xsl2_fscan_mode,
  output          xsl2_fscan_mode_atspeed,
  output          xsl2_fscan_state,
  output          xsl2_fscan_byplatrst_b,
  output          xsl2_fscan_byprst_b,
  output          xsl2_fscan_clkgenctrl,
  output          xsl2_fscan_clkgenctrlen,
  output          xsl2_fscan_clkungate,
  output          xsl2_fscan_clkungate_syn,
  output          xsl2_fscan_rstbypen,
  output          xsl2_fscan_shiften,
  output          xsl2_fscan_ram_bypsel,
  output          xsl2_fscan_ram_hold,
  output          xsl2_fscan_ram_init_en,
  output          xsl2_fscan_ram_init_val,
  output          xsl2_fscan_ram_mcp,
  output          xsl2_fscan_ram_odis_b,
  output          xsl2_fscan_ram_rddis_b,
  output          xsl2_fscan_ram_wrdis_b,
  input           xsl2_fdfx_powergood,
  input           xsl2_ijtag_capture,
  input           xsl2_ijtag_reset_b,
  input           xsl2_ijtag_select,
  input           xsl2_ijtag_shift,
  input           xsl2_ijtag_si,
  input           xsl2_ijtag_tck,
  input           xsl2_ijtag_update,
  output          xsl2_ijtag_so,
  input  [3397:0] xsl2_scanchains_so_end,
  output [3397:0] xsl2_scanchains_si_bgn,
  output          xsl2_dftclken,
  input           xsl2_core_clock_preclk,
  output          xsl2_core_clock_postclk,
  input           xsl2_uscan_state,
  input           xsl2_uscan_edt_update,
  input           xsl2_uscan_mode,
  input           xsl2_uscan_scanclk,
  input  [19:0]   xsl2_uscan_si,
  output [19:0]   xsl2_uscan_so
);
  ultiscan_xsl2_ult_scan_ctlr_wrap xsl2_ultiscan (
    .xsl2_fscan_mode(xsl2_fscan_mode),
    .xsl2_fscan_mode_atspeed(xsl2_fscan_mode_atspeed),
    .xsl2_fscan_state(xsl2_fscan_state),
    .xsl2_fscan_byplatrst_b(xsl2_fscan_byplatrst_b),
    .xsl2_fscan_byprst_b(xsl2_fscan_byprst_b),
    .xsl2_fscan_clkgenctrl(xsl2_fscan_clkgenctrl),
    .xsl2_fscan_clkgenctrlen(xsl2_fscan_clkgenctrlen),
    .xsl2_fscan_clkungate(xsl2_fscan_clkungate),
    .xsl2_fscan_clkungate_syn(xsl2_fscan_clkungate_syn),
    .xsl2_fscan_rstbypen(xsl2_fscan_rstbypen),
    .xsl2_fscan_shiften(xsl2_fscan_shiften),
    .xsl2_fscan_ram_bypsel(xsl2_fscan_ram_bypsel),
    .xsl2_fscan_ram_hold(xsl2_fscan_ram_hold),
    .xsl2_fscan_ram_init_en(xsl2_fscan_ram_init_en),
    .xsl2_fscan_ram_init_val(xsl2_fscan_ram_init_val),
    .xsl2_fscan_ram_mcp(xsl2_fscan_ram_mcp),
    .xsl2_fscan_ram_odis_b(xsl2_fscan_ram_odis_b),
    .xsl2_fscan_ram_rddis_b(xsl2_fscan_ram_rddis_b),
    .xsl2_fscan_ram_wrdis_b(xsl2_fscan_ram_wrdis_b),
    .xsl2_fdfx_powergood(xsl2_fdfx_powergood),
    .xsl2_ijtag_capture(xsl2_ijtag_capture),
    .xsl2_ijtag_reset_b(xsl2_ijtag_reset_b),
    .xsl2_ijtag_select(xsl2_ijtag_select),
    .xsl2_ijtag_shift(xsl2_ijtag_shift),
    .xsl2_ijtag_si(xsl2_ijtag_si),
    .xsl2_ijtag_tck(xsl2_ijtag_tck),
    .xsl2_ijtag_update(xsl2_ijtag_update),
    .xsl2_ijtag_so(xsl2_ijtag_so),
    .xsl2_scanchains_so_end(xsl2_scanchains_so_end),
    .xsl2_scanchains_si_bgn(xsl2_scanchains_si_bgn),
    .xsl2_dftclken(xsl2_dftclken),
    .xsl2_core_clock_preclk(xsl2_core_clock_preclk),
    .xsl2_core_clock_postclk(xsl2_core_clock_postclk),
    .xsl2_uscan_state(xsl2_uscan_state),
    .xsl2_uscan_edt_update(xsl2_uscan_edt_update),
    .xsl2_uscan_mode(xsl2_uscan_mode),
    .xsl2_uscan_scanclk(xsl2_uscan_scanclk),
    .xsl2_uscan_si(xsl2_uscan_si),
    .xsl2_uscan_so(xsl2_uscan_so)
  );
endmodule

