module AgeDetector(
  input         clock,
  input         reset,
  input  [15:0] io_enq_0,
  input  [15:0] io_enq_1,
  input  [15:0] io_deq,
  output [15:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
`endif // RANDOMIZE_REG_INIT
  reg  age_0_0; // @[SelectPolicy.scala 115:62]
  reg  age_0_1; // @[SelectPolicy.scala 115:62]
  reg  age_0_2; // @[SelectPolicy.scala 115:62]
  reg  age_0_3; // @[SelectPolicy.scala 115:62]
  reg  age_0_4; // @[SelectPolicy.scala 115:62]
  reg  age_0_5; // @[SelectPolicy.scala 115:62]
  reg  age_0_6; // @[SelectPolicy.scala 115:62]
  reg  age_0_7; // @[SelectPolicy.scala 115:62]
  reg  age_0_8; // @[SelectPolicy.scala 115:62]
  reg  age_0_9; // @[SelectPolicy.scala 115:62]
  reg  age_0_10; // @[SelectPolicy.scala 115:62]
  reg  age_0_11; // @[SelectPolicy.scala 115:62]
  reg  age_0_12; // @[SelectPolicy.scala 115:62]
  reg  age_0_13; // @[SelectPolicy.scala 115:62]
  reg  age_0_14; // @[SelectPolicy.scala 115:62]
  reg  age_0_15; // @[SelectPolicy.scala 115:62]
  reg  age_1_1; // @[SelectPolicy.scala 115:62]
  reg  age_1_2; // @[SelectPolicy.scala 115:62]
  reg  age_1_3; // @[SelectPolicy.scala 115:62]
  reg  age_1_4; // @[SelectPolicy.scala 115:62]
  reg  age_1_5; // @[SelectPolicy.scala 115:62]
  reg  age_1_6; // @[SelectPolicy.scala 115:62]
  reg  age_1_7; // @[SelectPolicy.scala 115:62]
  reg  age_1_8; // @[SelectPolicy.scala 115:62]
  reg  age_1_9; // @[SelectPolicy.scala 115:62]
  reg  age_1_10; // @[SelectPolicy.scala 115:62]
  reg  age_1_11; // @[SelectPolicy.scala 115:62]
  reg  age_1_12; // @[SelectPolicy.scala 115:62]
  reg  age_1_13; // @[SelectPolicy.scala 115:62]
  reg  age_1_14; // @[SelectPolicy.scala 115:62]
  reg  age_1_15; // @[SelectPolicy.scala 115:62]
  reg  age_2_2; // @[SelectPolicy.scala 115:62]
  reg  age_2_3; // @[SelectPolicy.scala 115:62]
  reg  age_2_4; // @[SelectPolicy.scala 115:62]
  reg  age_2_5; // @[SelectPolicy.scala 115:62]
  reg  age_2_6; // @[SelectPolicy.scala 115:62]
  reg  age_2_7; // @[SelectPolicy.scala 115:62]
  reg  age_2_8; // @[SelectPolicy.scala 115:62]
  reg  age_2_9; // @[SelectPolicy.scala 115:62]
  reg  age_2_10; // @[SelectPolicy.scala 115:62]
  reg  age_2_11; // @[SelectPolicy.scala 115:62]
  reg  age_2_12; // @[SelectPolicy.scala 115:62]
  reg  age_2_13; // @[SelectPolicy.scala 115:62]
  reg  age_2_14; // @[SelectPolicy.scala 115:62]
  reg  age_2_15; // @[SelectPolicy.scala 115:62]
  reg  age_3_3; // @[SelectPolicy.scala 115:62]
  reg  age_3_4; // @[SelectPolicy.scala 115:62]
  reg  age_3_5; // @[SelectPolicy.scala 115:62]
  reg  age_3_6; // @[SelectPolicy.scala 115:62]
  reg  age_3_7; // @[SelectPolicy.scala 115:62]
  reg  age_3_8; // @[SelectPolicy.scala 115:62]
  reg  age_3_9; // @[SelectPolicy.scala 115:62]
  reg  age_3_10; // @[SelectPolicy.scala 115:62]
  reg  age_3_11; // @[SelectPolicy.scala 115:62]
  reg  age_3_12; // @[SelectPolicy.scala 115:62]
  reg  age_3_13; // @[SelectPolicy.scala 115:62]
  reg  age_3_14; // @[SelectPolicy.scala 115:62]
  reg  age_3_15; // @[SelectPolicy.scala 115:62]
  reg  age_4_4; // @[SelectPolicy.scala 115:62]
  reg  age_4_5; // @[SelectPolicy.scala 115:62]
  reg  age_4_6; // @[SelectPolicy.scala 115:62]
  reg  age_4_7; // @[SelectPolicy.scala 115:62]
  reg  age_4_8; // @[SelectPolicy.scala 115:62]
  reg  age_4_9; // @[SelectPolicy.scala 115:62]
  reg  age_4_10; // @[SelectPolicy.scala 115:62]
  reg  age_4_11; // @[SelectPolicy.scala 115:62]
  reg  age_4_12; // @[SelectPolicy.scala 115:62]
  reg  age_4_13; // @[SelectPolicy.scala 115:62]
  reg  age_4_14; // @[SelectPolicy.scala 115:62]
  reg  age_4_15; // @[SelectPolicy.scala 115:62]
  reg  age_5_5; // @[SelectPolicy.scala 115:62]
  reg  age_5_6; // @[SelectPolicy.scala 115:62]
  reg  age_5_7; // @[SelectPolicy.scala 115:62]
  reg  age_5_8; // @[SelectPolicy.scala 115:62]
  reg  age_5_9; // @[SelectPolicy.scala 115:62]
  reg  age_5_10; // @[SelectPolicy.scala 115:62]
  reg  age_5_11; // @[SelectPolicy.scala 115:62]
  reg  age_5_12; // @[SelectPolicy.scala 115:62]
  reg  age_5_13; // @[SelectPolicy.scala 115:62]
  reg  age_5_14; // @[SelectPolicy.scala 115:62]
  reg  age_5_15; // @[SelectPolicy.scala 115:62]
  reg  age_6_6; // @[SelectPolicy.scala 115:62]
  reg  age_6_7; // @[SelectPolicy.scala 115:62]
  reg  age_6_8; // @[SelectPolicy.scala 115:62]
  reg  age_6_9; // @[SelectPolicy.scala 115:62]
  reg  age_6_10; // @[SelectPolicy.scala 115:62]
  reg  age_6_11; // @[SelectPolicy.scala 115:62]
  reg  age_6_12; // @[SelectPolicy.scala 115:62]
  reg  age_6_13; // @[SelectPolicy.scala 115:62]
  reg  age_6_14; // @[SelectPolicy.scala 115:62]
  reg  age_6_15; // @[SelectPolicy.scala 115:62]
  reg  age_7_7; // @[SelectPolicy.scala 115:62]
  reg  age_7_8; // @[SelectPolicy.scala 115:62]
  reg  age_7_9; // @[SelectPolicy.scala 115:62]
  reg  age_7_10; // @[SelectPolicy.scala 115:62]
  reg  age_7_11; // @[SelectPolicy.scala 115:62]
  reg  age_7_12; // @[SelectPolicy.scala 115:62]
  reg  age_7_13; // @[SelectPolicy.scala 115:62]
  reg  age_7_14; // @[SelectPolicy.scala 115:62]
  reg  age_7_15; // @[SelectPolicy.scala 115:62]
  reg  age_8_8; // @[SelectPolicy.scala 115:62]
  reg  age_8_9; // @[SelectPolicy.scala 115:62]
  reg  age_8_10; // @[SelectPolicy.scala 115:62]
  reg  age_8_11; // @[SelectPolicy.scala 115:62]
  reg  age_8_12; // @[SelectPolicy.scala 115:62]
  reg  age_8_13; // @[SelectPolicy.scala 115:62]
  reg  age_8_14; // @[SelectPolicy.scala 115:62]
  reg  age_8_15; // @[SelectPolicy.scala 115:62]
  reg  age_9_9; // @[SelectPolicy.scala 115:62]
  reg  age_9_10; // @[SelectPolicy.scala 115:62]
  reg  age_9_11; // @[SelectPolicy.scala 115:62]
  reg  age_9_12; // @[SelectPolicy.scala 115:62]
  reg  age_9_13; // @[SelectPolicy.scala 115:62]
  reg  age_9_14; // @[SelectPolicy.scala 115:62]
  reg  age_9_15; // @[SelectPolicy.scala 115:62]
  reg  age_10_10; // @[SelectPolicy.scala 115:62]
  reg  age_10_11; // @[SelectPolicy.scala 115:62]
  reg  age_10_12; // @[SelectPolicy.scala 115:62]
  reg  age_10_13; // @[SelectPolicy.scala 115:62]
  reg  age_10_14; // @[SelectPolicy.scala 115:62]
  reg  age_10_15; // @[SelectPolicy.scala 115:62]
  reg  age_11_11; // @[SelectPolicy.scala 115:62]
  reg  age_11_12; // @[SelectPolicy.scala 115:62]
  reg  age_11_13; // @[SelectPolicy.scala 115:62]
  reg  age_11_14; // @[SelectPolicy.scala 115:62]
  reg  age_11_15; // @[SelectPolicy.scala 115:62]
  reg  age_12_12; // @[SelectPolicy.scala 115:62]
  reg  age_12_13; // @[SelectPolicy.scala 115:62]
  reg  age_12_14; // @[SelectPolicy.scala 115:62]
  reg  age_12_15; // @[SelectPolicy.scala 115:62]
  reg  age_13_13; // @[SelectPolicy.scala 115:62]
  reg  age_13_14; // @[SelectPolicy.scala 115:62]
  reg  age_13_15; // @[SelectPolicy.scala 115:62]
  reg  age_14_14; // @[SelectPolicy.scala 115:62]
  reg  age_14_15; // @[SelectPolicy.scala 115:62]
  reg  age_15_15; // @[SelectPolicy.scala 115:62]
  wire [1:0] _thisValid_T_2 = {io_enq_1[0],io_enq_0[0]}; // @[SelectPolicy.scala 127:51]
  wire  _thisValid_T_5 = ~io_deq[0]; // @[SelectPolicy.scala 127:65]
  wire  _thisValid_T_6 = |_thisValid_T_2 & ~io_deq[0]; // @[SelectPolicy.scala 127:62]
  wire  thisValid = age_0_0 | _thisValid_T_6; // @[SelectPolicy.scala 132:35]
  wire  result_1 = io_enq_0[0] & _thisValid_T_5; // @[SelectPolicy.scala 126:32]
  wire  nextAge_0_0_xs_1 = io_enq_1[0] & result_1; // @[ParallelMux.scala 64:44]
  wire  _result_T_5 = ~io_deq[1]; // @[SelectPolicy.scala 126:35]
  wire  result_1_1 = io_enq_0[1] & ~io_deq[1]; // @[SelectPolicy.scala 126:32]
  wire  nextAge_0_1_xs_1 = io_enq_1[0] & result_1_1; // @[ParallelMux.scala 64:44]
  wire  _result_T_8 = ~io_deq[2]; // @[SelectPolicy.scala 126:35]
  wire  result_1_2 = io_enq_0[2] & ~io_deq[2]; // @[SelectPolicy.scala 126:32]
  wire  nextAge_0_2_xs_1 = io_enq_1[0] & result_1_2; // @[ParallelMux.scala 64:44]
  wire  _result_T_11 = ~io_deq[3]; // @[SelectPolicy.scala 126:35]
  wire  result_1_3 = io_enq_0[3] & ~io_deq[3]; // @[SelectPolicy.scala 126:32]
  wire  nextAge_0_3_xs_1 = io_enq_1[0] & result_1_3; // @[ParallelMux.scala 64:44]
  wire  _result_T_14 = ~io_deq[4]; // @[SelectPolicy.scala 126:35]
  wire  result_1_4 = io_enq_0[4] & ~io_deq[4]; // @[SelectPolicy.scala 126:32]
  wire  nextAge_0_4_xs_1 = io_enq_1[0] & result_1_4; // @[ParallelMux.scala 64:44]
  wire  _result_T_17 = ~io_deq[5]; // @[SelectPolicy.scala 126:35]
  wire  result_1_5 = io_enq_0[5] & ~io_deq[5]; // @[SelectPolicy.scala 126:32]
  wire  nextAge_0_5_xs_1 = io_enq_1[0] & result_1_5; // @[ParallelMux.scala 64:44]
  wire  _result_T_20 = ~io_deq[6]; // @[SelectPolicy.scala 126:35]
  wire  result_1_6 = io_enq_0[6] & ~io_deq[6]; // @[SelectPolicy.scala 126:32]
  wire  nextAge_0_6_xs_1 = io_enq_1[0] & result_1_6; // @[ParallelMux.scala 64:44]
  wire  _result_T_23 = ~io_deq[7]; // @[SelectPolicy.scala 126:35]
  wire  result_1_7 = io_enq_0[7] & ~io_deq[7]; // @[SelectPolicy.scala 126:32]
  wire  nextAge_0_7_xs_1 = io_enq_1[0] & result_1_7; // @[ParallelMux.scala 64:44]
  wire  _result_T_26 = ~io_deq[8]; // @[SelectPolicy.scala 126:35]
  wire  result_1_8 = io_enq_0[8] & ~io_deq[8]; // @[SelectPolicy.scala 126:32]
  wire  nextAge_0_8_xs_1 = io_enq_1[0] & result_1_8; // @[ParallelMux.scala 64:44]
  wire  _result_T_29 = ~io_deq[9]; // @[SelectPolicy.scala 126:35]
  wire  result_1_9 = io_enq_0[9] & ~io_deq[9]; // @[SelectPolicy.scala 126:32]
  wire  nextAge_0_9_xs_1 = io_enq_1[0] & result_1_9; // @[ParallelMux.scala 64:44]
  wire  _result_T_32 = ~io_deq[10]; // @[SelectPolicy.scala 126:35]
  wire  result_1_10 = io_enq_0[10] & ~io_deq[10]; // @[SelectPolicy.scala 126:32]
  wire  nextAge_0_10_xs_1 = io_enq_1[0] & result_1_10; // @[ParallelMux.scala 64:44]
  wire  _result_T_35 = ~io_deq[11]; // @[SelectPolicy.scala 126:35]
  wire  result_1_11 = io_enq_0[11] & ~io_deq[11]; // @[SelectPolicy.scala 126:32]
  wire  nextAge_0_11_xs_1 = io_enq_1[0] & result_1_11; // @[ParallelMux.scala 64:44]
  wire  _result_T_38 = ~io_deq[12]; // @[SelectPolicy.scala 126:35]
  wire  result_1_12 = io_enq_0[12] & ~io_deq[12]; // @[SelectPolicy.scala 126:32]
  wire  nextAge_0_12_xs_1 = io_enq_1[0] & result_1_12; // @[ParallelMux.scala 64:44]
  wire  _result_T_41 = ~io_deq[13]; // @[SelectPolicy.scala 126:35]
  wire  result_1_13 = io_enq_0[13] & ~io_deq[13]; // @[SelectPolicy.scala 126:32]
  wire  nextAge_0_13_xs_1 = io_enq_1[0] & result_1_13; // @[ParallelMux.scala 64:44]
  wire  _result_T_44 = ~io_deq[14]; // @[SelectPolicy.scala 126:35]
  wire  result_1_14 = io_enq_0[14] & ~io_deq[14]; // @[SelectPolicy.scala 126:32]
  wire  nextAge_0_14_xs_1 = io_enq_1[0] & result_1_14; // @[ParallelMux.scala 64:44]
  wire  _result_T_47 = ~io_deq[15]; // @[SelectPolicy.scala 126:35]
  wire  result_1_15 = io_enq_0[15] & ~io_deq[15]; // @[SelectPolicy.scala 126:32]
  wire  nextAge_0_15_xs_1 = io_enq_1[0] & result_1_15; // @[ParallelMux.scala 64:44]
  wire [1:0] _thisValid_T_9 = {io_enq_1[1],io_enq_0[1]}; // @[SelectPolicy.scala 127:51]
  wire  _thisValid_T_13 = |_thisValid_T_9 & _result_T_5; // @[SelectPolicy.scala 127:62]
  wire  thisValid_1 = age_1_1 | _thisValid_T_13; // @[SelectPolicy.scala 132:35]
  wire  _nextAge_1_0_T_4 = ~age_0_1; // @[SelectPolicy.scala 119:78]
  wire  nextAge_1_1_xs_1 = io_enq_1[1] & result_1_1; // @[ParallelMux.scala 64:44]
  wire  nextAge_1_2_xs_1 = io_enq_1[1] & result_1_2; // @[ParallelMux.scala 64:44]
  wire  nextAge_1_3_xs_1 = io_enq_1[1] & result_1_3; // @[ParallelMux.scala 64:44]
  wire  nextAge_1_4_xs_1 = io_enq_1[1] & result_1_4; // @[ParallelMux.scala 64:44]
  wire  nextAge_1_5_xs_1 = io_enq_1[1] & result_1_5; // @[ParallelMux.scala 64:44]
  wire  nextAge_1_6_xs_1 = io_enq_1[1] & result_1_6; // @[ParallelMux.scala 64:44]
  wire  nextAge_1_7_xs_1 = io_enq_1[1] & result_1_7; // @[ParallelMux.scala 64:44]
  wire  nextAge_1_8_xs_1 = io_enq_1[1] & result_1_8; // @[ParallelMux.scala 64:44]
  wire  nextAge_1_9_xs_1 = io_enq_1[1] & result_1_9; // @[ParallelMux.scala 64:44]
  wire  nextAge_1_10_xs_1 = io_enq_1[1] & result_1_10; // @[ParallelMux.scala 64:44]
  wire  nextAge_1_11_xs_1 = io_enq_1[1] & result_1_11; // @[ParallelMux.scala 64:44]
  wire  nextAge_1_12_xs_1 = io_enq_1[1] & result_1_12; // @[ParallelMux.scala 64:44]
  wire  nextAge_1_13_xs_1 = io_enq_1[1] & result_1_13; // @[ParallelMux.scala 64:44]
  wire  nextAge_1_14_xs_1 = io_enq_1[1] & result_1_14; // @[ParallelMux.scala 64:44]
  wire  nextAge_1_15_xs_1 = io_enq_1[1] & result_1_15; // @[ParallelMux.scala 64:44]
  wire [1:0] _thisValid_T_16 = {io_enq_1[2],io_enq_0[2]}; // @[SelectPolicy.scala 127:51]
  wire  _thisValid_T_20 = |_thisValid_T_16 & _result_T_8; // @[SelectPolicy.scala 127:62]
  wire  thisValid_2 = age_2_2 | _thisValid_T_20; // @[SelectPolicy.scala 132:35]
  wire  _nextAge_2_0_T_4 = ~age_0_2; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_2_1_T_4 = ~age_1_2; // @[SelectPolicy.scala 119:78]
  wire  nextAge_2_2_xs_1 = io_enq_1[2] & result_1_2; // @[ParallelMux.scala 64:44]
  wire  nextAge_2_3_xs_1 = io_enq_1[2] & result_1_3; // @[ParallelMux.scala 64:44]
  wire  nextAge_2_4_xs_1 = io_enq_1[2] & result_1_4; // @[ParallelMux.scala 64:44]
  wire  nextAge_2_5_xs_1 = io_enq_1[2] & result_1_5; // @[ParallelMux.scala 64:44]
  wire  nextAge_2_6_xs_1 = io_enq_1[2] & result_1_6; // @[ParallelMux.scala 64:44]
  wire  nextAge_2_7_xs_1 = io_enq_1[2] & result_1_7; // @[ParallelMux.scala 64:44]
  wire  nextAge_2_8_xs_1 = io_enq_1[2] & result_1_8; // @[ParallelMux.scala 64:44]
  wire  nextAge_2_9_xs_1 = io_enq_1[2] & result_1_9; // @[ParallelMux.scala 64:44]
  wire  nextAge_2_10_xs_1 = io_enq_1[2] & result_1_10; // @[ParallelMux.scala 64:44]
  wire  nextAge_2_11_xs_1 = io_enq_1[2] & result_1_11; // @[ParallelMux.scala 64:44]
  wire  nextAge_2_12_xs_1 = io_enq_1[2] & result_1_12; // @[ParallelMux.scala 64:44]
  wire  nextAge_2_13_xs_1 = io_enq_1[2] & result_1_13; // @[ParallelMux.scala 64:44]
  wire  nextAge_2_14_xs_1 = io_enq_1[2] & result_1_14; // @[ParallelMux.scala 64:44]
  wire  nextAge_2_15_xs_1 = io_enq_1[2] & result_1_15; // @[ParallelMux.scala 64:44]
  wire [1:0] _thisValid_T_23 = {io_enq_1[3],io_enq_0[3]}; // @[SelectPolicy.scala 127:51]
  wire  _thisValid_T_27 = |_thisValid_T_23 & _result_T_11; // @[SelectPolicy.scala 127:62]
  wire  thisValid_3 = age_3_3 | _thisValid_T_27; // @[SelectPolicy.scala 132:35]
  wire  _nextAge_3_0_T_4 = ~age_0_3; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_3_1_T_4 = ~age_1_3; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_3_2_T_4 = ~age_2_3; // @[SelectPolicy.scala 119:78]
  wire  nextAge_3_3_xs_1 = io_enq_1[3] & result_1_3; // @[ParallelMux.scala 64:44]
  wire  nextAge_3_4_xs_1 = io_enq_1[3] & result_1_4; // @[ParallelMux.scala 64:44]
  wire  nextAge_3_5_xs_1 = io_enq_1[3] & result_1_5; // @[ParallelMux.scala 64:44]
  wire  nextAge_3_6_xs_1 = io_enq_1[3] & result_1_6; // @[ParallelMux.scala 64:44]
  wire  nextAge_3_7_xs_1 = io_enq_1[3] & result_1_7; // @[ParallelMux.scala 64:44]
  wire  nextAge_3_8_xs_1 = io_enq_1[3] & result_1_8; // @[ParallelMux.scala 64:44]
  wire  nextAge_3_9_xs_1 = io_enq_1[3] & result_1_9; // @[ParallelMux.scala 64:44]
  wire  nextAge_3_10_xs_1 = io_enq_1[3] & result_1_10; // @[ParallelMux.scala 64:44]
  wire  nextAge_3_11_xs_1 = io_enq_1[3] & result_1_11; // @[ParallelMux.scala 64:44]
  wire  nextAge_3_12_xs_1 = io_enq_1[3] & result_1_12; // @[ParallelMux.scala 64:44]
  wire  nextAge_3_13_xs_1 = io_enq_1[3] & result_1_13; // @[ParallelMux.scala 64:44]
  wire  nextAge_3_14_xs_1 = io_enq_1[3] & result_1_14; // @[ParallelMux.scala 64:44]
  wire  nextAge_3_15_xs_1 = io_enq_1[3] & result_1_15; // @[ParallelMux.scala 64:44]
  wire [1:0] _thisValid_T_30 = {io_enq_1[4],io_enq_0[4]}; // @[SelectPolicy.scala 127:51]
  wire  _thisValid_T_34 = |_thisValid_T_30 & _result_T_14; // @[SelectPolicy.scala 127:62]
  wire  thisValid_4 = age_4_4 | _thisValid_T_34; // @[SelectPolicy.scala 132:35]
  wire  _nextAge_4_0_T_4 = ~age_0_4; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_4_1_T_4 = ~age_1_4; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_4_2_T_4 = ~age_2_4; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_4_3_T_4 = ~age_3_4; // @[SelectPolicy.scala 119:78]
  wire  nextAge_4_4_xs_1 = io_enq_1[4] & result_1_4; // @[ParallelMux.scala 64:44]
  wire  nextAge_4_5_xs_1 = io_enq_1[4] & result_1_5; // @[ParallelMux.scala 64:44]
  wire  nextAge_4_6_xs_1 = io_enq_1[4] & result_1_6; // @[ParallelMux.scala 64:44]
  wire  nextAge_4_7_xs_1 = io_enq_1[4] & result_1_7; // @[ParallelMux.scala 64:44]
  wire  nextAge_4_8_xs_1 = io_enq_1[4] & result_1_8; // @[ParallelMux.scala 64:44]
  wire  nextAge_4_9_xs_1 = io_enq_1[4] & result_1_9; // @[ParallelMux.scala 64:44]
  wire  nextAge_4_10_xs_1 = io_enq_1[4] & result_1_10; // @[ParallelMux.scala 64:44]
  wire  nextAge_4_11_xs_1 = io_enq_1[4] & result_1_11; // @[ParallelMux.scala 64:44]
  wire  nextAge_4_12_xs_1 = io_enq_1[4] & result_1_12; // @[ParallelMux.scala 64:44]
  wire  nextAge_4_13_xs_1 = io_enq_1[4] & result_1_13; // @[ParallelMux.scala 64:44]
  wire  nextAge_4_14_xs_1 = io_enq_1[4] & result_1_14; // @[ParallelMux.scala 64:44]
  wire  nextAge_4_15_xs_1 = io_enq_1[4] & result_1_15; // @[ParallelMux.scala 64:44]
  wire [1:0] _thisValid_T_37 = {io_enq_1[5],io_enq_0[5]}; // @[SelectPolicy.scala 127:51]
  wire  _thisValid_T_41 = |_thisValid_T_37 & _result_T_17; // @[SelectPolicy.scala 127:62]
  wire  thisValid_5 = age_5_5 | _thisValid_T_41; // @[SelectPolicy.scala 132:35]
  wire  _nextAge_5_0_T_4 = ~age_0_5; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_5_1_T_4 = ~age_1_5; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_5_2_T_4 = ~age_2_5; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_5_3_T_4 = ~age_3_5; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_5_4_T_4 = ~age_4_5; // @[SelectPolicy.scala 119:78]
  wire  nextAge_5_5_xs_1 = io_enq_1[5] & result_1_5; // @[ParallelMux.scala 64:44]
  wire  nextAge_5_6_xs_1 = io_enq_1[5] & result_1_6; // @[ParallelMux.scala 64:44]
  wire  nextAge_5_7_xs_1 = io_enq_1[5] & result_1_7; // @[ParallelMux.scala 64:44]
  wire  nextAge_5_8_xs_1 = io_enq_1[5] & result_1_8; // @[ParallelMux.scala 64:44]
  wire  nextAge_5_9_xs_1 = io_enq_1[5] & result_1_9; // @[ParallelMux.scala 64:44]
  wire  nextAge_5_10_xs_1 = io_enq_1[5] & result_1_10; // @[ParallelMux.scala 64:44]
  wire  nextAge_5_11_xs_1 = io_enq_1[5] & result_1_11; // @[ParallelMux.scala 64:44]
  wire  nextAge_5_12_xs_1 = io_enq_1[5] & result_1_12; // @[ParallelMux.scala 64:44]
  wire  nextAge_5_13_xs_1 = io_enq_1[5] & result_1_13; // @[ParallelMux.scala 64:44]
  wire  nextAge_5_14_xs_1 = io_enq_1[5] & result_1_14; // @[ParallelMux.scala 64:44]
  wire  nextAge_5_15_xs_1 = io_enq_1[5] & result_1_15; // @[ParallelMux.scala 64:44]
  wire [1:0] _thisValid_T_44 = {io_enq_1[6],io_enq_0[6]}; // @[SelectPolicy.scala 127:51]
  wire  _thisValid_T_48 = |_thisValid_T_44 & _result_T_20; // @[SelectPolicy.scala 127:62]
  wire  thisValid_6 = age_6_6 | _thisValid_T_48; // @[SelectPolicy.scala 132:35]
  wire  _nextAge_6_0_T_4 = ~age_0_6; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_6_1_T_4 = ~age_1_6; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_6_2_T_4 = ~age_2_6; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_6_3_T_4 = ~age_3_6; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_6_4_T_4 = ~age_4_6; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_6_5_T_4 = ~age_5_6; // @[SelectPolicy.scala 119:78]
  wire  nextAge_6_6_xs_1 = io_enq_1[6] & result_1_6; // @[ParallelMux.scala 64:44]
  wire  nextAge_6_7_xs_1 = io_enq_1[6] & result_1_7; // @[ParallelMux.scala 64:44]
  wire  nextAge_6_8_xs_1 = io_enq_1[6] & result_1_8; // @[ParallelMux.scala 64:44]
  wire  nextAge_6_9_xs_1 = io_enq_1[6] & result_1_9; // @[ParallelMux.scala 64:44]
  wire  nextAge_6_10_xs_1 = io_enq_1[6] & result_1_10; // @[ParallelMux.scala 64:44]
  wire  nextAge_6_11_xs_1 = io_enq_1[6] & result_1_11; // @[ParallelMux.scala 64:44]
  wire  nextAge_6_12_xs_1 = io_enq_1[6] & result_1_12; // @[ParallelMux.scala 64:44]
  wire  nextAge_6_13_xs_1 = io_enq_1[6] & result_1_13; // @[ParallelMux.scala 64:44]
  wire  nextAge_6_14_xs_1 = io_enq_1[6] & result_1_14; // @[ParallelMux.scala 64:44]
  wire  nextAge_6_15_xs_1 = io_enq_1[6] & result_1_15; // @[ParallelMux.scala 64:44]
  wire [1:0] _thisValid_T_51 = {io_enq_1[7],io_enq_0[7]}; // @[SelectPolicy.scala 127:51]
  wire  _thisValid_T_55 = |_thisValid_T_51 & _result_T_23; // @[SelectPolicy.scala 127:62]
  wire  thisValid_7 = age_7_7 | _thisValid_T_55; // @[SelectPolicy.scala 132:35]
  wire  _nextAge_7_0_T_4 = ~age_0_7; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_7_1_T_4 = ~age_1_7; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_7_2_T_4 = ~age_2_7; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_7_3_T_4 = ~age_3_7; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_7_4_T_4 = ~age_4_7; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_7_5_T_4 = ~age_5_7; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_7_6_T_4 = ~age_6_7; // @[SelectPolicy.scala 119:78]
  wire  nextAge_7_7_xs_1 = io_enq_1[7] & result_1_7; // @[ParallelMux.scala 64:44]
  wire  nextAge_7_8_xs_1 = io_enq_1[7] & result_1_8; // @[ParallelMux.scala 64:44]
  wire  nextAge_7_9_xs_1 = io_enq_1[7] & result_1_9; // @[ParallelMux.scala 64:44]
  wire  nextAge_7_10_xs_1 = io_enq_1[7] & result_1_10; // @[ParallelMux.scala 64:44]
  wire  nextAge_7_11_xs_1 = io_enq_1[7] & result_1_11; // @[ParallelMux.scala 64:44]
  wire  nextAge_7_12_xs_1 = io_enq_1[7] & result_1_12; // @[ParallelMux.scala 64:44]
  wire  nextAge_7_13_xs_1 = io_enq_1[7] & result_1_13; // @[ParallelMux.scala 64:44]
  wire  nextAge_7_14_xs_1 = io_enq_1[7] & result_1_14; // @[ParallelMux.scala 64:44]
  wire  nextAge_7_15_xs_1 = io_enq_1[7] & result_1_15; // @[ParallelMux.scala 64:44]
  wire [1:0] _thisValid_T_58 = {io_enq_1[8],io_enq_0[8]}; // @[SelectPolicy.scala 127:51]
  wire  _thisValid_T_62 = |_thisValid_T_58 & _result_T_26; // @[SelectPolicy.scala 127:62]
  wire  thisValid_8 = age_8_8 | _thisValid_T_62; // @[SelectPolicy.scala 132:35]
  wire  _nextAge_8_0_T_4 = ~age_0_8; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_8_1_T_4 = ~age_1_8; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_8_2_T_4 = ~age_2_8; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_8_3_T_4 = ~age_3_8; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_8_4_T_4 = ~age_4_8; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_8_5_T_4 = ~age_5_8; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_8_6_T_4 = ~age_6_8; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_8_7_T_4 = ~age_7_8; // @[SelectPolicy.scala 119:78]
  wire  nextAge_8_8_xs_1 = io_enq_1[8] & result_1_8; // @[ParallelMux.scala 64:44]
  wire  nextAge_8_9_xs_1 = io_enq_1[8] & result_1_9; // @[ParallelMux.scala 64:44]
  wire  nextAge_8_10_xs_1 = io_enq_1[8] & result_1_10; // @[ParallelMux.scala 64:44]
  wire  nextAge_8_11_xs_1 = io_enq_1[8] & result_1_11; // @[ParallelMux.scala 64:44]
  wire  nextAge_8_12_xs_1 = io_enq_1[8] & result_1_12; // @[ParallelMux.scala 64:44]
  wire  nextAge_8_13_xs_1 = io_enq_1[8] & result_1_13; // @[ParallelMux.scala 64:44]
  wire  nextAge_8_14_xs_1 = io_enq_1[8] & result_1_14; // @[ParallelMux.scala 64:44]
  wire  nextAge_8_15_xs_1 = io_enq_1[8] & result_1_15; // @[ParallelMux.scala 64:44]
  wire [1:0] _thisValid_T_65 = {io_enq_1[9],io_enq_0[9]}; // @[SelectPolicy.scala 127:51]
  wire  _thisValid_T_69 = |_thisValid_T_65 & _result_T_29; // @[SelectPolicy.scala 127:62]
  wire  thisValid_9 = age_9_9 | _thisValid_T_69; // @[SelectPolicy.scala 132:35]
  wire  _nextAge_9_0_T_4 = ~age_0_9; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_9_1_T_4 = ~age_1_9; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_9_2_T_4 = ~age_2_9; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_9_3_T_4 = ~age_3_9; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_9_4_T_4 = ~age_4_9; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_9_5_T_4 = ~age_5_9; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_9_6_T_4 = ~age_6_9; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_9_7_T_4 = ~age_7_9; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_9_8_T_4 = ~age_8_9; // @[SelectPolicy.scala 119:78]
  wire  nextAge_9_9_xs_1 = io_enq_1[9] & result_1_9; // @[ParallelMux.scala 64:44]
  wire  nextAge_9_10_xs_1 = io_enq_1[9] & result_1_10; // @[ParallelMux.scala 64:44]
  wire  nextAge_9_11_xs_1 = io_enq_1[9] & result_1_11; // @[ParallelMux.scala 64:44]
  wire  nextAge_9_12_xs_1 = io_enq_1[9] & result_1_12; // @[ParallelMux.scala 64:44]
  wire  nextAge_9_13_xs_1 = io_enq_1[9] & result_1_13; // @[ParallelMux.scala 64:44]
  wire  nextAge_9_14_xs_1 = io_enq_1[9] & result_1_14; // @[ParallelMux.scala 64:44]
  wire  nextAge_9_15_xs_1 = io_enq_1[9] & result_1_15; // @[ParallelMux.scala 64:44]
  wire [1:0] _thisValid_T_72 = {io_enq_1[10],io_enq_0[10]}; // @[SelectPolicy.scala 127:51]
  wire  _thisValid_T_76 = |_thisValid_T_72 & _result_T_32; // @[SelectPolicy.scala 127:62]
  wire  thisValid_10 = age_10_10 | _thisValid_T_76; // @[SelectPolicy.scala 132:35]
  wire  _nextAge_10_0_T_4 = ~age_0_10; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_10_1_T_4 = ~age_1_10; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_10_2_T_4 = ~age_2_10; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_10_3_T_4 = ~age_3_10; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_10_4_T_4 = ~age_4_10; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_10_5_T_4 = ~age_5_10; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_10_6_T_4 = ~age_6_10; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_10_7_T_4 = ~age_7_10; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_10_8_T_4 = ~age_8_10; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_10_9_T_4 = ~age_9_10; // @[SelectPolicy.scala 119:78]
  wire  nextAge_10_10_xs_1 = io_enq_1[10] & result_1_10; // @[ParallelMux.scala 64:44]
  wire  nextAge_10_11_xs_1 = io_enq_1[10] & result_1_11; // @[ParallelMux.scala 64:44]
  wire  nextAge_10_12_xs_1 = io_enq_1[10] & result_1_12; // @[ParallelMux.scala 64:44]
  wire  nextAge_10_13_xs_1 = io_enq_1[10] & result_1_13; // @[ParallelMux.scala 64:44]
  wire  nextAge_10_14_xs_1 = io_enq_1[10] & result_1_14; // @[ParallelMux.scala 64:44]
  wire  nextAge_10_15_xs_1 = io_enq_1[10] & result_1_15; // @[ParallelMux.scala 64:44]
  wire [1:0] _thisValid_T_79 = {io_enq_1[11],io_enq_0[11]}; // @[SelectPolicy.scala 127:51]
  wire  _thisValid_T_83 = |_thisValid_T_79 & _result_T_35; // @[SelectPolicy.scala 127:62]
  wire  thisValid_11 = age_11_11 | _thisValid_T_83; // @[SelectPolicy.scala 132:35]
  wire  _nextAge_11_0_T_4 = ~age_0_11; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_11_1_T_4 = ~age_1_11; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_11_2_T_4 = ~age_2_11; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_11_3_T_4 = ~age_3_11; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_11_4_T_4 = ~age_4_11; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_11_5_T_4 = ~age_5_11; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_11_6_T_4 = ~age_6_11; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_11_7_T_4 = ~age_7_11; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_11_8_T_4 = ~age_8_11; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_11_9_T_4 = ~age_9_11; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_11_10_T_4 = ~age_10_11; // @[SelectPolicy.scala 119:78]
  wire  nextAge_11_11_xs_1 = io_enq_1[11] & result_1_11; // @[ParallelMux.scala 64:44]
  wire  nextAge_11_12_xs_1 = io_enq_1[11] & result_1_12; // @[ParallelMux.scala 64:44]
  wire  nextAge_11_13_xs_1 = io_enq_1[11] & result_1_13; // @[ParallelMux.scala 64:44]
  wire  nextAge_11_14_xs_1 = io_enq_1[11] & result_1_14; // @[ParallelMux.scala 64:44]
  wire  nextAge_11_15_xs_1 = io_enq_1[11] & result_1_15; // @[ParallelMux.scala 64:44]
  wire [1:0] _thisValid_T_86 = {io_enq_1[12],io_enq_0[12]}; // @[SelectPolicy.scala 127:51]
  wire  _thisValid_T_90 = |_thisValid_T_86 & _result_T_38; // @[SelectPolicy.scala 127:62]
  wire  thisValid_12 = age_12_12 | _thisValid_T_90; // @[SelectPolicy.scala 132:35]
  wire  _nextAge_12_0_T_4 = ~age_0_12; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_12_1_T_4 = ~age_1_12; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_12_2_T_4 = ~age_2_12; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_12_3_T_4 = ~age_3_12; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_12_4_T_4 = ~age_4_12; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_12_5_T_4 = ~age_5_12; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_12_6_T_4 = ~age_6_12; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_12_7_T_4 = ~age_7_12; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_12_8_T_4 = ~age_8_12; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_12_9_T_4 = ~age_9_12; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_12_10_T_4 = ~age_10_12; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_12_11_T_4 = ~age_11_12; // @[SelectPolicy.scala 119:78]
  wire  nextAge_12_12_xs_1 = io_enq_1[12] & result_1_12; // @[ParallelMux.scala 64:44]
  wire  nextAge_12_13_xs_1 = io_enq_1[12] & result_1_13; // @[ParallelMux.scala 64:44]
  wire  nextAge_12_14_xs_1 = io_enq_1[12] & result_1_14; // @[ParallelMux.scala 64:44]
  wire  nextAge_12_15_xs_1 = io_enq_1[12] & result_1_15; // @[ParallelMux.scala 64:44]
  wire [1:0] _thisValid_T_93 = {io_enq_1[13],io_enq_0[13]}; // @[SelectPolicy.scala 127:51]
  wire  _thisValid_T_97 = |_thisValid_T_93 & _result_T_41; // @[SelectPolicy.scala 127:62]
  wire  thisValid_13 = age_13_13 | _thisValid_T_97; // @[SelectPolicy.scala 132:35]
  wire  _nextAge_13_0_T_4 = ~age_0_13; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_13_1_T_4 = ~age_1_13; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_13_2_T_4 = ~age_2_13; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_13_3_T_4 = ~age_3_13; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_13_4_T_4 = ~age_4_13; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_13_5_T_4 = ~age_5_13; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_13_6_T_4 = ~age_6_13; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_13_7_T_4 = ~age_7_13; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_13_8_T_4 = ~age_8_13; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_13_9_T_4 = ~age_9_13; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_13_10_T_4 = ~age_10_13; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_13_11_T_4 = ~age_11_13; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_13_12_T_4 = ~age_12_13; // @[SelectPolicy.scala 119:78]
  wire  nextAge_13_13_xs_1 = io_enq_1[13] & result_1_13; // @[ParallelMux.scala 64:44]
  wire  nextAge_13_14_xs_1 = io_enq_1[13] & result_1_14; // @[ParallelMux.scala 64:44]
  wire  nextAge_13_15_xs_1 = io_enq_1[13] & result_1_15; // @[ParallelMux.scala 64:44]
  wire [1:0] _thisValid_T_100 = {io_enq_1[14],io_enq_0[14]}; // @[SelectPolicy.scala 127:51]
  wire  _thisValid_T_104 = |_thisValid_T_100 & _result_T_44; // @[SelectPolicy.scala 127:62]
  wire  thisValid_14 = age_14_14 | _thisValid_T_104; // @[SelectPolicy.scala 132:35]
  wire  _nextAge_14_0_T_4 = ~age_0_14; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_14_1_T_4 = ~age_1_14; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_14_2_T_4 = ~age_2_14; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_14_3_T_4 = ~age_3_14; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_14_4_T_4 = ~age_4_14; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_14_5_T_4 = ~age_5_14; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_14_6_T_4 = ~age_6_14; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_14_7_T_4 = ~age_7_14; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_14_8_T_4 = ~age_8_14; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_14_9_T_4 = ~age_9_14; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_14_10_T_4 = ~age_10_14; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_14_11_T_4 = ~age_11_14; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_14_12_T_4 = ~age_12_14; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_14_13_T_4 = ~age_13_14; // @[SelectPolicy.scala 119:78]
  wire  nextAge_14_14_xs_1 = io_enq_1[14] & result_1_14; // @[ParallelMux.scala 64:44]
  wire  nextAge_14_15_xs_1 = io_enq_1[14] & result_1_15; // @[ParallelMux.scala 64:44]
  wire [1:0] _thisValid_T_107 = {io_enq_1[15],io_enq_0[15]}; // @[SelectPolicy.scala 127:51]
  wire  _thisValid_T_111 = |_thisValid_T_107 & _result_T_47; // @[SelectPolicy.scala 127:62]
  wire  thisValid_15 = age_15_15 | _thisValid_T_111; // @[SelectPolicy.scala 132:35]
  wire  _nextAge_15_0_T_4 = ~age_0_15; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_15_1_T_4 = ~age_1_15; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_15_2_T_4 = ~age_2_15; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_15_3_T_4 = ~age_3_15; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_15_4_T_4 = ~age_4_15; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_15_5_T_4 = ~age_5_15; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_15_6_T_4 = ~age_6_15; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_15_7_T_4 = ~age_7_15; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_15_8_T_4 = ~age_8_15; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_15_9_T_4 = ~age_9_15; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_15_10_T_4 = ~age_10_15; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_15_11_T_4 = ~age_11_15; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_15_12_T_4 = ~age_12_15; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_15_13_T_4 = ~age_13_15; // @[SelectPolicy.scala 119:78]
  wire  _nextAge_15_14_T_4 = ~age_14_15; // @[SelectPolicy.scala 119:78]
  wire  nextAge_15_15_xs_1 = io_enq_1[15] & result_1_15; // @[ParallelMux.scala 64:44]
  wire [7:0] best_lo = {age_0_7,age_0_6,age_0_5,age_0_4,age_0_3,age_0_2,age_0_1,age_0_0}; // @[SelectPolicy.scala 159:57]
  wire [15:0] _best_T = {age_0_15,age_0_14,age_0_13,age_0_12,age_0_11,age_0_10,age_0_9,age_0_8,best_lo}; // @[SelectPolicy.scala 159:57]
  wire  _best_T_1 = &_best_T; // @[SelectPolicy.scala 159:64]
  wire [7:0] best_lo_1 = {age_1_7,age_1_6,age_1_5,age_1_4,age_1_3,age_1_2,age_1_1,_nextAge_1_0_T_4}; // @[SelectPolicy.scala 159:57]
  wire [15:0] _best_T_3 = {age_1_15,age_1_14,age_1_13,age_1_12,age_1_11,age_1_10,age_1_9,age_1_8,best_lo_1}; // @[SelectPolicy.scala 159:57]
  wire  _best_T_4 = &_best_T_3; // @[SelectPolicy.scala 159:64]
  wire [7:0] best_lo_2 = {age_2_7,age_2_6,age_2_5,age_2_4,age_2_3,age_2_2,_nextAge_2_1_T_4,_nextAge_2_0_T_4}; // @[SelectPolicy.scala 159:57]
  wire [15:0] _best_T_7 = {age_2_15,age_2_14,age_2_13,age_2_12,age_2_11,age_2_10,age_2_9,age_2_8,best_lo_2}; // @[SelectPolicy.scala 159:57]
  wire  _best_T_8 = &_best_T_7; // @[SelectPolicy.scala 159:64]
  wire [7:0] best_lo_3 = {age_3_7,age_3_6,age_3_5,age_3_4,age_3_3,_nextAge_3_2_T_4,_nextAge_3_1_T_4,_nextAge_3_0_T_4}; // @[SelectPolicy.scala 159:57]
  wire [15:0] _best_T_12 = {age_3_15,age_3_14,age_3_13,age_3_12,age_3_11,age_3_10,age_3_9,age_3_8,best_lo_3}; // @[SelectPolicy.scala 159:57]
  wire  _best_T_13 = &_best_T_12; // @[SelectPolicy.scala 159:64]
  wire [7:0] best_lo_4 = {age_4_7,age_4_6,age_4_5,age_4_4,_nextAge_4_3_T_4,_nextAge_4_2_T_4,_nextAge_4_1_T_4,
    _nextAge_4_0_T_4}; // @[SelectPolicy.scala 159:57]
  wire [15:0] _best_T_18 = {age_4_15,age_4_14,age_4_13,age_4_12,age_4_11,age_4_10,age_4_9,age_4_8,best_lo_4}; // @[SelectPolicy.scala 159:57]
  wire  _best_T_19 = &_best_T_18; // @[SelectPolicy.scala 159:64]
  wire [7:0] best_lo_5 = {age_5_7,age_5_6,age_5_5,_nextAge_5_4_T_4,_nextAge_5_3_T_4,_nextAge_5_2_T_4,_nextAge_5_1_T_4,
    _nextAge_5_0_T_4}; // @[SelectPolicy.scala 159:57]
  wire [15:0] _best_T_25 = {age_5_15,age_5_14,age_5_13,age_5_12,age_5_11,age_5_10,age_5_9,age_5_8,best_lo_5}; // @[SelectPolicy.scala 159:57]
  wire  _best_T_26 = &_best_T_25; // @[SelectPolicy.scala 159:64]
  wire [7:0] best_lo_6 = {age_6_7,age_6_6,_nextAge_6_5_T_4,_nextAge_6_4_T_4,_nextAge_6_3_T_4,_nextAge_6_2_T_4,
    _nextAge_6_1_T_4,_nextAge_6_0_T_4}; // @[SelectPolicy.scala 159:57]
  wire [15:0] _best_T_33 = {age_6_15,age_6_14,age_6_13,age_6_12,age_6_11,age_6_10,age_6_9,age_6_8,best_lo_6}; // @[SelectPolicy.scala 159:57]
  wire  _best_T_34 = &_best_T_33; // @[SelectPolicy.scala 159:64]
  wire [7:0] best_lo_7 = {age_7_7,_nextAge_7_6_T_4,_nextAge_7_5_T_4,_nextAge_7_4_T_4,_nextAge_7_3_T_4,_nextAge_7_2_T_4,
    _nextAge_7_1_T_4,_nextAge_7_0_T_4}; // @[SelectPolicy.scala 159:57]
  wire [15:0] _best_T_42 = {age_7_15,age_7_14,age_7_13,age_7_12,age_7_11,age_7_10,age_7_9,age_7_8,best_lo_7}; // @[SelectPolicy.scala 159:57]
  wire  _best_T_43 = &_best_T_42; // @[SelectPolicy.scala 159:64]
  wire [7:0] best_lo_8 = {_nextAge_8_7_T_4,_nextAge_8_6_T_4,_nextAge_8_5_T_4,_nextAge_8_4_T_4,_nextAge_8_3_T_4,
    _nextAge_8_2_T_4,_nextAge_8_1_T_4,_nextAge_8_0_T_4}; // @[SelectPolicy.scala 159:57]
  wire [15:0] _best_T_52 = {age_8_15,age_8_14,age_8_13,age_8_12,age_8_11,age_8_10,age_8_9,age_8_8,best_lo_8}; // @[SelectPolicy.scala 159:57]
  wire  _best_T_53 = &_best_T_52; // @[SelectPolicy.scala 159:64]
  wire [7:0] best_lo_9 = {_nextAge_9_7_T_4,_nextAge_9_6_T_4,_nextAge_9_5_T_4,_nextAge_9_4_T_4,_nextAge_9_3_T_4,
    _nextAge_9_2_T_4,_nextAge_9_1_T_4,_nextAge_9_0_T_4}; // @[SelectPolicy.scala 159:57]
  wire [15:0] _best_T_63 = {age_9_15,age_9_14,age_9_13,age_9_12,age_9_11,age_9_10,age_9_9,_nextAge_9_8_T_4,best_lo_9}; // @[SelectPolicy.scala 159:57]
  wire  _best_T_64 = &_best_T_63; // @[SelectPolicy.scala 159:64]
  wire [7:0] best_lo_10 = {_nextAge_10_7_T_4,_nextAge_10_6_T_4,_nextAge_10_5_T_4,_nextAge_10_4_T_4,_nextAge_10_3_T_4,
    _nextAge_10_2_T_4,_nextAge_10_1_T_4,_nextAge_10_0_T_4}; // @[SelectPolicy.scala 159:57]
  wire [15:0] _best_T_75 = {age_10_15,age_10_14,age_10_13,age_10_12,age_10_11,age_10_10,_nextAge_10_9_T_4,
    _nextAge_10_8_T_4,best_lo_10}; // @[SelectPolicy.scala 159:57]
  wire  _best_T_76 = &_best_T_75; // @[SelectPolicy.scala 159:64]
  wire [7:0] best_lo_11 = {_nextAge_11_7_T_4,_nextAge_11_6_T_4,_nextAge_11_5_T_4,_nextAge_11_4_T_4,_nextAge_11_3_T_4,
    _nextAge_11_2_T_4,_nextAge_11_1_T_4,_nextAge_11_0_T_4}; // @[SelectPolicy.scala 159:57]
  wire [15:0] _best_T_88 = {age_11_15,age_11_14,age_11_13,age_11_12,age_11_11,_nextAge_11_10_T_4,_nextAge_11_9_T_4,
    _nextAge_11_8_T_4,best_lo_11}; // @[SelectPolicy.scala 159:57]
  wire  _best_T_89 = &_best_T_88; // @[SelectPolicy.scala 159:64]
  wire [7:0] best_lo_12 = {_nextAge_12_7_T_4,_nextAge_12_6_T_4,_nextAge_12_5_T_4,_nextAge_12_4_T_4,_nextAge_12_3_T_4,
    _nextAge_12_2_T_4,_nextAge_12_1_T_4,_nextAge_12_0_T_4}; // @[SelectPolicy.scala 159:57]
  wire [15:0] _best_T_102 = {age_12_15,age_12_14,age_12_13,age_12_12,_nextAge_12_11_T_4,_nextAge_12_10_T_4,
    _nextAge_12_9_T_4,_nextAge_12_8_T_4,best_lo_12}; // @[SelectPolicy.scala 159:57]
  wire  _best_T_103 = &_best_T_102; // @[SelectPolicy.scala 159:64]
  wire [7:0] best_lo_13 = {_nextAge_13_7_T_4,_nextAge_13_6_T_4,_nextAge_13_5_T_4,_nextAge_13_4_T_4,_nextAge_13_3_T_4,
    _nextAge_13_2_T_4,_nextAge_13_1_T_4,_nextAge_13_0_T_4}; // @[SelectPolicy.scala 159:57]
  wire [15:0] _best_T_117 = {age_13_15,age_13_14,age_13_13,_nextAge_13_12_T_4,_nextAge_13_11_T_4,_nextAge_13_10_T_4,
    _nextAge_13_9_T_4,_nextAge_13_8_T_4,best_lo_13}; // @[SelectPolicy.scala 159:57]
  wire  _best_T_118 = &_best_T_117; // @[SelectPolicy.scala 159:64]
  wire [7:0] best_lo_14 = {_nextAge_14_7_T_4,_nextAge_14_6_T_4,_nextAge_14_5_T_4,_nextAge_14_4_T_4,_nextAge_14_3_T_4,
    _nextAge_14_2_T_4,_nextAge_14_1_T_4,_nextAge_14_0_T_4}; // @[SelectPolicy.scala 159:57]
  wire [15:0] _best_T_133 = {age_14_15,age_14_14,_nextAge_14_13_T_4,_nextAge_14_12_T_4,_nextAge_14_11_T_4,
    _nextAge_14_10_T_4,_nextAge_14_9_T_4,_nextAge_14_8_T_4,best_lo_14}; // @[SelectPolicy.scala 159:57]
  wire  _best_T_134 = &_best_T_133; // @[SelectPolicy.scala 159:64]
  wire [7:0] best_lo_15 = {_nextAge_15_7_T_4,_nextAge_15_6_T_4,_nextAge_15_5_T_4,_nextAge_15_4_T_4,_nextAge_15_3_T_4,
    _nextAge_15_2_T_4,_nextAge_15_1_T_4,_nextAge_15_0_T_4}; // @[SelectPolicy.scala 159:57]
  wire [15:0] _best_T_150 = {age_15_15,_nextAge_15_14_T_4,_nextAge_15_13_T_4,_nextAge_15_12_T_4,_nextAge_15_11_T_4,
    _nextAge_15_10_T_4,_nextAge_15_9_T_4,_nextAge_15_8_T_4,best_lo_15}; // @[SelectPolicy.scala 159:57]
  wire  _best_T_151 = &_best_T_150; // @[SelectPolicy.scala 159:64]
  wire [7:0] best_lo_16 = {_best_T_43,_best_T_34,_best_T_26,_best_T_19,_best_T_13,_best_T_8,_best_T_4,_best_T_1}; // @[SelectPolicy.scala 160:9]
  wire [7:0] best_hi_16 = {_best_T_151,_best_T_134,_best_T_118,_best_T_103,_best_T_89,_best_T_76,_best_T_64,_best_T_53}; // @[SelectPolicy.scala 160:9]
  assign io_out = {best_hi_16,best_lo_16}; // @[SelectPolicy.scala 160:9]
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_0_0 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[0]) begin // @[SelectPolicy.scala 137:33]
      age_0_0 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[0]) begin // @[SelectPolicy.scala 140:34]
      age_0_0 <= thisValid; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_6) begin // @[SelectPolicy.scala 151:14]
      age_0_0 <= ~age_0_0 & ~nextAge_0_0_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_0_1 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[0]) begin // @[SelectPolicy.scala 137:33]
      age_0_1 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[1]) begin // @[SelectPolicy.scala 140:34]
      age_0_1 <= thisValid; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_6) begin // @[SelectPolicy.scala 151:14]
      age_0_1 <= ~age_1_1 & ~nextAge_0_1_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_0_2 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[0]) begin // @[SelectPolicy.scala 137:33]
      age_0_2 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[2]) begin // @[SelectPolicy.scala 140:34]
      age_0_2 <= thisValid; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_6) begin // @[SelectPolicy.scala 151:14]
      age_0_2 <= ~age_2_2 & ~nextAge_0_2_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_0_3 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[0]) begin // @[SelectPolicy.scala 137:33]
      age_0_3 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[3]) begin // @[SelectPolicy.scala 140:34]
      age_0_3 <= thisValid; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_6) begin // @[SelectPolicy.scala 151:14]
      age_0_3 <= ~age_3_3 & ~nextAge_0_3_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_0_4 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[0]) begin // @[SelectPolicy.scala 137:33]
      age_0_4 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[4]) begin // @[SelectPolicy.scala 140:34]
      age_0_4 <= thisValid; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_6) begin // @[SelectPolicy.scala 151:14]
      age_0_4 <= ~age_4_4 & ~nextAge_0_4_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_0_5 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[0]) begin // @[SelectPolicy.scala 137:33]
      age_0_5 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[5]) begin // @[SelectPolicy.scala 140:34]
      age_0_5 <= thisValid; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_6) begin // @[SelectPolicy.scala 151:14]
      age_0_5 <= ~age_5_5 & ~nextAge_0_5_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_0_6 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[0]) begin // @[SelectPolicy.scala 137:33]
      age_0_6 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[6]) begin // @[SelectPolicy.scala 140:34]
      age_0_6 <= thisValid; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_6) begin // @[SelectPolicy.scala 151:14]
      age_0_6 <= ~age_6_6 & ~nextAge_0_6_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_0_7 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[0]) begin // @[SelectPolicy.scala 137:33]
      age_0_7 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[7]) begin // @[SelectPolicy.scala 140:34]
      age_0_7 <= thisValid; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_6) begin // @[SelectPolicy.scala 151:14]
      age_0_7 <= ~age_7_7 & ~nextAge_0_7_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_0_8 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[0]) begin // @[SelectPolicy.scala 137:33]
      age_0_8 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[8]) begin // @[SelectPolicy.scala 140:34]
      age_0_8 <= thisValid; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_6) begin // @[SelectPolicy.scala 151:14]
      age_0_8 <= ~age_8_8 & ~nextAge_0_8_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_0_9 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[0]) begin // @[SelectPolicy.scala 137:33]
      age_0_9 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[9]) begin // @[SelectPolicy.scala 140:34]
      age_0_9 <= thisValid; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_6) begin // @[SelectPolicy.scala 151:14]
      age_0_9 <= ~age_9_9 & ~nextAge_0_9_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_0_10 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[0]) begin // @[SelectPolicy.scala 137:33]
      age_0_10 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[10]) begin // @[SelectPolicy.scala 140:34]
      age_0_10 <= thisValid; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_6) begin // @[SelectPolicy.scala 151:14]
      age_0_10 <= ~age_10_10 & ~nextAge_0_10_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_0_11 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[0]) begin // @[SelectPolicy.scala 137:33]
      age_0_11 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[11]) begin // @[SelectPolicy.scala 140:34]
      age_0_11 <= thisValid; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_6) begin // @[SelectPolicy.scala 151:14]
      age_0_11 <= ~age_11_11 & ~nextAge_0_11_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_0_12 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[0]) begin // @[SelectPolicy.scala 137:33]
      age_0_12 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[12]) begin // @[SelectPolicy.scala 140:34]
      age_0_12 <= thisValid; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_6) begin // @[SelectPolicy.scala 151:14]
      age_0_12 <= ~age_12_12 & ~nextAge_0_12_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_0_13 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[0]) begin // @[SelectPolicy.scala 137:33]
      age_0_13 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[13]) begin // @[SelectPolicy.scala 140:34]
      age_0_13 <= thisValid; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_6) begin // @[SelectPolicy.scala 151:14]
      age_0_13 <= ~age_13_13 & ~nextAge_0_13_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_0_14 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[0]) begin // @[SelectPolicy.scala 137:33]
      age_0_14 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[14]) begin // @[SelectPolicy.scala 140:34]
      age_0_14 <= thisValid; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_6) begin // @[SelectPolicy.scala 151:14]
      age_0_14 <= ~age_14_14 & ~nextAge_0_14_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_0_15 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[0]) begin // @[SelectPolicy.scala 137:33]
      age_0_15 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[15]) begin // @[SelectPolicy.scala 140:34]
      age_0_15 <= thisValid; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_6) begin // @[SelectPolicy.scala 151:14]
      age_0_15 <= ~age_15_15 & ~nextAge_0_15_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_1_1 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[1]) begin // @[SelectPolicy.scala 137:33]
      age_1_1 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[1]) begin // @[SelectPolicy.scala 140:34]
      age_1_1 <= thisValid_1; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_13) begin // @[SelectPolicy.scala 151:14]
      age_1_1 <= ~age_1_1 & ~nextAge_1_1_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_1_2 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[1]) begin // @[SelectPolicy.scala 137:33]
      age_1_2 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[2]) begin // @[SelectPolicy.scala 140:34]
      age_1_2 <= thisValid_1; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_13) begin // @[SelectPolicy.scala 151:14]
      age_1_2 <= ~age_2_2 & ~nextAge_1_2_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_1_3 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[1]) begin // @[SelectPolicy.scala 137:33]
      age_1_3 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[3]) begin // @[SelectPolicy.scala 140:34]
      age_1_3 <= thisValid_1; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_13) begin // @[SelectPolicy.scala 151:14]
      age_1_3 <= ~age_3_3 & ~nextAge_1_3_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_1_4 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[1]) begin // @[SelectPolicy.scala 137:33]
      age_1_4 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[4]) begin // @[SelectPolicy.scala 140:34]
      age_1_4 <= thisValid_1; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_13) begin // @[SelectPolicy.scala 151:14]
      age_1_4 <= ~age_4_4 & ~nextAge_1_4_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_1_5 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[1]) begin // @[SelectPolicy.scala 137:33]
      age_1_5 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[5]) begin // @[SelectPolicy.scala 140:34]
      age_1_5 <= thisValid_1; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_13) begin // @[SelectPolicy.scala 151:14]
      age_1_5 <= ~age_5_5 & ~nextAge_1_5_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_1_6 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[1]) begin // @[SelectPolicy.scala 137:33]
      age_1_6 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[6]) begin // @[SelectPolicy.scala 140:34]
      age_1_6 <= thisValid_1; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_13) begin // @[SelectPolicy.scala 151:14]
      age_1_6 <= ~age_6_6 & ~nextAge_1_6_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_1_7 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[1]) begin // @[SelectPolicy.scala 137:33]
      age_1_7 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[7]) begin // @[SelectPolicy.scala 140:34]
      age_1_7 <= thisValid_1; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_13) begin // @[SelectPolicy.scala 151:14]
      age_1_7 <= ~age_7_7 & ~nextAge_1_7_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_1_8 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[1]) begin // @[SelectPolicy.scala 137:33]
      age_1_8 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[8]) begin // @[SelectPolicy.scala 140:34]
      age_1_8 <= thisValid_1; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_13) begin // @[SelectPolicy.scala 151:14]
      age_1_8 <= ~age_8_8 & ~nextAge_1_8_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_1_9 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[1]) begin // @[SelectPolicy.scala 137:33]
      age_1_9 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[9]) begin // @[SelectPolicy.scala 140:34]
      age_1_9 <= thisValid_1; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_13) begin // @[SelectPolicy.scala 151:14]
      age_1_9 <= ~age_9_9 & ~nextAge_1_9_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_1_10 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[1]) begin // @[SelectPolicy.scala 137:33]
      age_1_10 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[10]) begin // @[SelectPolicy.scala 140:34]
      age_1_10 <= thisValid_1; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_13) begin // @[SelectPolicy.scala 151:14]
      age_1_10 <= ~age_10_10 & ~nextAge_1_10_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_1_11 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[1]) begin // @[SelectPolicy.scala 137:33]
      age_1_11 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[11]) begin // @[SelectPolicy.scala 140:34]
      age_1_11 <= thisValid_1; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_13) begin // @[SelectPolicy.scala 151:14]
      age_1_11 <= ~age_11_11 & ~nextAge_1_11_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_1_12 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[1]) begin // @[SelectPolicy.scala 137:33]
      age_1_12 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[12]) begin // @[SelectPolicy.scala 140:34]
      age_1_12 <= thisValid_1; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_13) begin // @[SelectPolicy.scala 151:14]
      age_1_12 <= ~age_12_12 & ~nextAge_1_12_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_1_13 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[1]) begin // @[SelectPolicy.scala 137:33]
      age_1_13 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[13]) begin // @[SelectPolicy.scala 140:34]
      age_1_13 <= thisValid_1; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_13) begin // @[SelectPolicy.scala 151:14]
      age_1_13 <= ~age_13_13 & ~nextAge_1_13_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_1_14 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[1]) begin // @[SelectPolicy.scala 137:33]
      age_1_14 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[14]) begin // @[SelectPolicy.scala 140:34]
      age_1_14 <= thisValid_1; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_13) begin // @[SelectPolicy.scala 151:14]
      age_1_14 <= ~age_14_14 & ~nextAge_1_14_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_1_15 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[1]) begin // @[SelectPolicy.scala 137:33]
      age_1_15 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[15]) begin // @[SelectPolicy.scala 140:34]
      age_1_15 <= thisValid_1; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_13) begin // @[SelectPolicy.scala 151:14]
      age_1_15 <= ~age_15_15 & ~nextAge_1_15_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_2_2 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[2]) begin // @[SelectPolicy.scala 137:33]
      age_2_2 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[2]) begin // @[SelectPolicy.scala 140:34]
      age_2_2 <= thisValid_2; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_20) begin // @[SelectPolicy.scala 151:14]
      age_2_2 <= ~age_2_2 & ~nextAge_2_2_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_2_3 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[2]) begin // @[SelectPolicy.scala 137:33]
      age_2_3 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[3]) begin // @[SelectPolicy.scala 140:34]
      age_2_3 <= thisValid_2; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_20) begin // @[SelectPolicy.scala 151:14]
      age_2_3 <= ~age_3_3 & ~nextAge_2_3_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_2_4 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[2]) begin // @[SelectPolicy.scala 137:33]
      age_2_4 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[4]) begin // @[SelectPolicy.scala 140:34]
      age_2_4 <= thisValid_2; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_20) begin // @[SelectPolicy.scala 151:14]
      age_2_4 <= ~age_4_4 & ~nextAge_2_4_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_2_5 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[2]) begin // @[SelectPolicy.scala 137:33]
      age_2_5 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[5]) begin // @[SelectPolicy.scala 140:34]
      age_2_5 <= thisValid_2; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_20) begin // @[SelectPolicy.scala 151:14]
      age_2_5 <= ~age_5_5 & ~nextAge_2_5_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_2_6 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[2]) begin // @[SelectPolicy.scala 137:33]
      age_2_6 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[6]) begin // @[SelectPolicy.scala 140:34]
      age_2_6 <= thisValid_2; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_20) begin // @[SelectPolicy.scala 151:14]
      age_2_6 <= ~age_6_6 & ~nextAge_2_6_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_2_7 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[2]) begin // @[SelectPolicy.scala 137:33]
      age_2_7 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[7]) begin // @[SelectPolicy.scala 140:34]
      age_2_7 <= thisValid_2; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_20) begin // @[SelectPolicy.scala 151:14]
      age_2_7 <= ~age_7_7 & ~nextAge_2_7_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_2_8 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[2]) begin // @[SelectPolicy.scala 137:33]
      age_2_8 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[8]) begin // @[SelectPolicy.scala 140:34]
      age_2_8 <= thisValid_2; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_20) begin // @[SelectPolicy.scala 151:14]
      age_2_8 <= ~age_8_8 & ~nextAge_2_8_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_2_9 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[2]) begin // @[SelectPolicy.scala 137:33]
      age_2_9 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[9]) begin // @[SelectPolicy.scala 140:34]
      age_2_9 <= thisValid_2; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_20) begin // @[SelectPolicy.scala 151:14]
      age_2_9 <= ~age_9_9 & ~nextAge_2_9_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_2_10 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[2]) begin // @[SelectPolicy.scala 137:33]
      age_2_10 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[10]) begin // @[SelectPolicy.scala 140:34]
      age_2_10 <= thisValid_2; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_20) begin // @[SelectPolicy.scala 151:14]
      age_2_10 <= ~age_10_10 & ~nextAge_2_10_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_2_11 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[2]) begin // @[SelectPolicy.scala 137:33]
      age_2_11 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[11]) begin // @[SelectPolicy.scala 140:34]
      age_2_11 <= thisValid_2; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_20) begin // @[SelectPolicy.scala 151:14]
      age_2_11 <= ~age_11_11 & ~nextAge_2_11_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_2_12 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[2]) begin // @[SelectPolicy.scala 137:33]
      age_2_12 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[12]) begin // @[SelectPolicy.scala 140:34]
      age_2_12 <= thisValid_2; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_20) begin // @[SelectPolicy.scala 151:14]
      age_2_12 <= ~age_12_12 & ~nextAge_2_12_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_2_13 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[2]) begin // @[SelectPolicy.scala 137:33]
      age_2_13 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[13]) begin // @[SelectPolicy.scala 140:34]
      age_2_13 <= thisValid_2; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_20) begin // @[SelectPolicy.scala 151:14]
      age_2_13 <= ~age_13_13 & ~nextAge_2_13_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_2_14 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[2]) begin // @[SelectPolicy.scala 137:33]
      age_2_14 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[14]) begin // @[SelectPolicy.scala 140:34]
      age_2_14 <= thisValid_2; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_20) begin // @[SelectPolicy.scala 151:14]
      age_2_14 <= ~age_14_14 & ~nextAge_2_14_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_2_15 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[2]) begin // @[SelectPolicy.scala 137:33]
      age_2_15 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[15]) begin // @[SelectPolicy.scala 140:34]
      age_2_15 <= thisValid_2; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_20) begin // @[SelectPolicy.scala 151:14]
      age_2_15 <= ~age_15_15 & ~nextAge_2_15_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_3_3 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[3]) begin // @[SelectPolicy.scala 137:33]
      age_3_3 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[3]) begin // @[SelectPolicy.scala 140:34]
      age_3_3 <= thisValid_3; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_27) begin // @[SelectPolicy.scala 151:14]
      age_3_3 <= ~age_3_3 & ~nextAge_3_3_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_3_4 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[3]) begin // @[SelectPolicy.scala 137:33]
      age_3_4 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[4]) begin // @[SelectPolicy.scala 140:34]
      age_3_4 <= thisValid_3; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_27) begin // @[SelectPolicy.scala 151:14]
      age_3_4 <= ~age_4_4 & ~nextAge_3_4_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_3_5 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[3]) begin // @[SelectPolicy.scala 137:33]
      age_3_5 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[5]) begin // @[SelectPolicy.scala 140:34]
      age_3_5 <= thisValid_3; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_27) begin // @[SelectPolicy.scala 151:14]
      age_3_5 <= ~age_5_5 & ~nextAge_3_5_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_3_6 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[3]) begin // @[SelectPolicy.scala 137:33]
      age_3_6 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[6]) begin // @[SelectPolicy.scala 140:34]
      age_3_6 <= thisValid_3; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_27) begin // @[SelectPolicy.scala 151:14]
      age_3_6 <= ~age_6_6 & ~nextAge_3_6_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_3_7 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[3]) begin // @[SelectPolicy.scala 137:33]
      age_3_7 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[7]) begin // @[SelectPolicy.scala 140:34]
      age_3_7 <= thisValid_3; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_27) begin // @[SelectPolicy.scala 151:14]
      age_3_7 <= ~age_7_7 & ~nextAge_3_7_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_3_8 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[3]) begin // @[SelectPolicy.scala 137:33]
      age_3_8 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[8]) begin // @[SelectPolicy.scala 140:34]
      age_3_8 <= thisValid_3; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_27) begin // @[SelectPolicy.scala 151:14]
      age_3_8 <= ~age_8_8 & ~nextAge_3_8_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_3_9 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[3]) begin // @[SelectPolicy.scala 137:33]
      age_3_9 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[9]) begin // @[SelectPolicy.scala 140:34]
      age_3_9 <= thisValid_3; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_27) begin // @[SelectPolicy.scala 151:14]
      age_3_9 <= ~age_9_9 & ~nextAge_3_9_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_3_10 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[3]) begin // @[SelectPolicy.scala 137:33]
      age_3_10 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[10]) begin // @[SelectPolicy.scala 140:34]
      age_3_10 <= thisValid_3; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_27) begin // @[SelectPolicy.scala 151:14]
      age_3_10 <= ~age_10_10 & ~nextAge_3_10_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_3_11 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[3]) begin // @[SelectPolicy.scala 137:33]
      age_3_11 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[11]) begin // @[SelectPolicy.scala 140:34]
      age_3_11 <= thisValid_3; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_27) begin // @[SelectPolicy.scala 151:14]
      age_3_11 <= ~age_11_11 & ~nextAge_3_11_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_3_12 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[3]) begin // @[SelectPolicy.scala 137:33]
      age_3_12 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[12]) begin // @[SelectPolicy.scala 140:34]
      age_3_12 <= thisValid_3; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_27) begin // @[SelectPolicy.scala 151:14]
      age_3_12 <= ~age_12_12 & ~nextAge_3_12_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_3_13 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[3]) begin // @[SelectPolicy.scala 137:33]
      age_3_13 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[13]) begin // @[SelectPolicy.scala 140:34]
      age_3_13 <= thisValid_3; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_27) begin // @[SelectPolicy.scala 151:14]
      age_3_13 <= ~age_13_13 & ~nextAge_3_13_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_3_14 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[3]) begin // @[SelectPolicy.scala 137:33]
      age_3_14 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[14]) begin // @[SelectPolicy.scala 140:34]
      age_3_14 <= thisValid_3; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_27) begin // @[SelectPolicy.scala 151:14]
      age_3_14 <= ~age_14_14 & ~nextAge_3_14_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_3_15 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[3]) begin // @[SelectPolicy.scala 137:33]
      age_3_15 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[15]) begin // @[SelectPolicy.scala 140:34]
      age_3_15 <= thisValid_3; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_27) begin // @[SelectPolicy.scala 151:14]
      age_3_15 <= ~age_15_15 & ~nextAge_3_15_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_4_4 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[4]) begin // @[SelectPolicy.scala 137:33]
      age_4_4 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[4]) begin // @[SelectPolicy.scala 140:34]
      age_4_4 <= thisValid_4; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_34) begin // @[SelectPolicy.scala 151:14]
      age_4_4 <= ~age_4_4 & ~nextAge_4_4_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_4_5 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[4]) begin // @[SelectPolicy.scala 137:33]
      age_4_5 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[5]) begin // @[SelectPolicy.scala 140:34]
      age_4_5 <= thisValid_4; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_34) begin // @[SelectPolicy.scala 151:14]
      age_4_5 <= ~age_5_5 & ~nextAge_4_5_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_4_6 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[4]) begin // @[SelectPolicy.scala 137:33]
      age_4_6 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[6]) begin // @[SelectPolicy.scala 140:34]
      age_4_6 <= thisValid_4; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_34) begin // @[SelectPolicy.scala 151:14]
      age_4_6 <= ~age_6_6 & ~nextAge_4_6_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_4_7 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[4]) begin // @[SelectPolicy.scala 137:33]
      age_4_7 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[7]) begin // @[SelectPolicy.scala 140:34]
      age_4_7 <= thisValid_4; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_34) begin // @[SelectPolicy.scala 151:14]
      age_4_7 <= ~age_7_7 & ~nextAge_4_7_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_4_8 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[4]) begin // @[SelectPolicy.scala 137:33]
      age_4_8 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[8]) begin // @[SelectPolicy.scala 140:34]
      age_4_8 <= thisValid_4; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_34) begin // @[SelectPolicy.scala 151:14]
      age_4_8 <= ~age_8_8 & ~nextAge_4_8_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_4_9 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[4]) begin // @[SelectPolicy.scala 137:33]
      age_4_9 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[9]) begin // @[SelectPolicy.scala 140:34]
      age_4_9 <= thisValid_4; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_34) begin // @[SelectPolicy.scala 151:14]
      age_4_9 <= ~age_9_9 & ~nextAge_4_9_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_4_10 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[4]) begin // @[SelectPolicy.scala 137:33]
      age_4_10 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[10]) begin // @[SelectPolicy.scala 140:34]
      age_4_10 <= thisValid_4; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_34) begin // @[SelectPolicy.scala 151:14]
      age_4_10 <= ~age_10_10 & ~nextAge_4_10_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_4_11 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[4]) begin // @[SelectPolicy.scala 137:33]
      age_4_11 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[11]) begin // @[SelectPolicy.scala 140:34]
      age_4_11 <= thisValid_4; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_34) begin // @[SelectPolicy.scala 151:14]
      age_4_11 <= ~age_11_11 & ~nextAge_4_11_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_4_12 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[4]) begin // @[SelectPolicy.scala 137:33]
      age_4_12 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[12]) begin // @[SelectPolicy.scala 140:34]
      age_4_12 <= thisValid_4; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_34) begin // @[SelectPolicy.scala 151:14]
      age_4_12 <= ~age_12_12 & ~nextAge_4_12_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_4_13 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[4]) begin // @[SelectPolicy.scala 137:33]
      age_4_13 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[13]) begin // @[SelectPolicy.scala 140:34]
      age_4_13 <= thisValid_4; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_34) begin // @[SelectPolicy.scala 151:14]
      age_4_13 <= ~age_13_13 & ~nextAge_4_13_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_4_14 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[4]) begin // @[SelectPolicy.scala 137:33]
      age_4_14 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[14]) begin // @[SelectPolicy.scala 140:34]
      age_4_14 <= thisValid_4; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_34) begin // @[SelectPolicy.scala 151:14]
      age_4_14 <= ~age_14_14 & ~nextAge_4_14_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_4_15 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[4]) begin // @[SelectPolicy.scala 137:33]
      age_4_15 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[15]) begin // @[SelectPolicy.scala 140:34]
      age_4_15 <= thisValid_4; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_34) begin // @[SelectPolicy.scala 151:14]
      age_4_15 <= ~age_15_15 & ~nextAge_4_15_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_5_5 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[5]) begin // @[SelectPolicy.scala 137:33]
      age_5_5 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[5]) begin // @[SelectPolicy.scala 140:34]
      age_5_5 <= thisValid_5; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_41) begin // @[SelectPolicy.scala 151:14]
      age_5_5 <= ~age_5_5 & ~nextAge_5_5_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_5_6 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[5]) begin // @[SelectPolicy.scala 137:33]
      age_5_6 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[6]) begin // @[SelectPolicy.scala 140:34]
      age_5_6 <= thisValid_5; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_41) begin // @[SelectPolicy.scala 151:14]
      age_5_6 <= ~age_6_6 & ~nextAge_5_6_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_5_7 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[5]) begin // @[SelectPolicy.scala 137:33]
      age_5_7 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[7]) begin // @[SelectPolicy.scala 140:34]
      age_5_7 <= thisValid_5; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_41) begin // @[SelectPolicy.scala 151:14]
      age_5_7 <= ~age_7_7 & ~nextAge_5_7_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_5_8 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[5]) begin // @[SelectPolicy.scala 137:33]
      age_5_8 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[8]) begin // @[SelectPolicy.scala 140:34]
      age_5_8 <= thisValid_5; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_41) begin // @[SelectPolicy.scala 151:14]
      age_5_8 <= ~age_8_8 & ~nextAge_5_8_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_5_9 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[5]) begin // @[SelectPolicy.scala 137:33]
      age_5_9 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[9]) begin // @[SelectPolicy.scala 140:34]
      age_5_9 <= thisValid_5; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_41) begin // @[SelectPolicy.scala 151:14]
      age_5_9 <= ~age_9_9 & ~nextAge_5_9_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_5_10 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[5]) begin // @[SelectPolicy.scala 137:33]
      age_5_10 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[10]) begin // @[SelectPolicy.scala 140:34]
      age_5_10 <= thisValid_5; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_41) begin // @[SelectPolicy.scala 151:14]
      age_5_10 <= ~age_10_10 & ~nextAge_5_10_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_5_11 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[5]) begin // @[SelectPolicy.scala 137:33]
      age_5_11 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[11]) begin // @[SelectPolicy.scala 140:34]
      age_5_11 <= thisValid_5; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_41) begin // @[SelectPolicy.scala 151:14]
      age_5_11 <= ~age_11_11 & ~nextAge_5_11_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_5_12 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[5]) begin // @[SelectPolicy.scala 137:33]
      age_5_12 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[12]) begin // @[SelectPolicy.scala 140:34]
      age_5_12 <= thisValid_5; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_41) begin // @[SelectPolicy.scala 151:14]
      age_5_12 <= ~age_12_12 & ~nextAge_5_12_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_5_13 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[5]) begin // @[SelectPolicy.scala 137:33]
      age_5_13 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[13]) begin // @[SelectPolicy.scala 140:34]
      age_5_13 <= thisValid_5; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_41) begin // @[SelectPolicy.scala 151:14]
      age_5_13 <= ~age_13_13 & ~nextAge_5_13_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_5_14 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[5]) begin // @[SelectPolicy.scala 137:33]
      age_5_14 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[14]) begin // @[SelectPolicy.scala 140:34]
      age_5_14 <= thisValid_5; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_41) begin // @[SelectPolicy.scala 151:14]
      age_5_14 <= ~age_14_14 & ~nextAge_5_14_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_5_15 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[5]) begin // @[SelectPolicy.scala 137:33]
      age_5_15 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[15]) begin // @[SelectPolicy.scala 140:34]
      age_5_15 <= thisValid_5; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_41) begin // @[SelectPolicy.scala 151:14]
      age_5_15 <= ~age_15_15 & ~nextAge_5_15_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_6_6 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[6]) begin // @[SelectPolicy.scala 137:33]
      age_6_6 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[6]) begin // @[SelectPolicy.scala 140:34]
      age_6_6 <= thisValid_6; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_48) begin // @[SelectPolicy.scala 151:14]
      age_6_6 <= ~age_6_6 & ~nextAge_6_6_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_6_7 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[6]) begin // @[SelectPolicy.scala 137:33]
      age_6_7 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[7]) begin // @[SelectPolicy.scala 140:34]
      age_6_7 <= thisValid_6; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_48) begin // @[SelectPolicy.scala 151:14]
      age_6_7 <= ~age_7_7 & ~nextAge_6_7_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_6_8 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[6]) begin // @[SelectPolicy.scala 137:33]
      age_6_8 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[8]) begin // @[SelectPolicy.scala 140:34]
      age_6_8 <= thisValid_6; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_48) begin // @[SelectPolicy.scala 151:14]
      age_6_8 <= ~age_8_8 & ~nextAge_6_8_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_6_9 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[6]) begin // @[SelectPolicy.scala 137:33]
      age_6_9 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[9]) begin // @[SelectPolicy.scala 140:34]
      age_6_9 <= thisValid_6; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_48) begin // @[SelectPolicy.scala 151:14]
      age_6_9 <= ~age_9_9 & ~nextAge_6_9_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_6_10 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[6]) begin // @[SelectPolicy.scala 137:33]
      age_6_10 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[10]) begin // @[SelectPolicy.scala 140:34]
      age_6_10 <= thisValid_6; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_48) begin // @[SelectPolicy.scala 151:14]
      age_6_10 <= ~age_10_10 & ~nextAge_6_10_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_6_11 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[6]) begin // @[SelectPolicy.scala 137:33]
      age_6_11 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[11]) begin // @[SelectPolicy.scala 140:34]
      age_6_11 <= thisValid_6; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_48) begin // @[SelectPolicy.scala 151:14]
      age_6_11 <= ~age_11_11 & ~nextAge_6_11_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_6_12 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[6]) begin // @[SelectPolicy.scala 137:33]
      age_6_12 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[12]) begin // @[SelectPolicy.scala 140:34]
      age_6_12 <= thisValid_6; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_48) begin // @[SelectPolicy.scala 151:14]
      age_6_12 <= ~age_12_12 & ~nextAge_6_12_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_6_13 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[6]) begin // @[SelectPolicy.scala 137:33]
      age_6_13 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[13]) begin // @[SelectPolicy.scala 140:34]
      age_6_13 <= thisValid_6; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_48) begin // @[SelectPolicy.scala 151:14]
      age_6_13 <= ~age_13_13 & ~nextAge_6_13_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_6_14 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[6]) begin // @[SelectPolicy.scala 137:33]
      age_6_14 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[14]) begin // @[SelectPolicy.scala 140:34]
      age_6_14 <= thisValid_6; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_48) begin // @[SelectPolicy.scala 151:14]
      age_6_14 <= ~age_14_14 & ~nextAge_6_14_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_6_15 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[6]) begin // @[SelectPolicy.scala 137:33]
      age_6_15 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[15]) begin // @[SelectPolicy.scala 140:34]
      age_6_15 <= thisValid_6; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_48) begin // @[SelectPolicy.scala 151:14]
      age_6_15 <= ~age_15_15 & ~nextAge_6_15_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_7_7 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[7]) begin // @[SelectPolicy.scala 137:33]
      age_7_7 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[7]) begin // @[SelectPolicy.scala 140:34]
      age_7_7 <= thisValid_7; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_55) begin // @[SelectPolicy.scala 151:14]
      age_7_7 <= ~age_7_7 & ~nextAge_7_7_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_7_8 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[7]) begin // @[SelectPolicy.scala 137:33]
      age_7_8 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[8]) begin // @[SelectPolicy.scala 140:34]
      age_7_8 <= thisValid_7; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_55) begin // @[SelectPolicy.scala 151:14]
      age_7_8 <= ~age_8_8 & ~nextAge_7_8_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_7_9 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[7]) begin // @[SelectPolicy.scala 137:33]
      age_7_9 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[9]) begin // @[SelectPolicy.scala 140:34]
      age_7_9 <= thisValid_7; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_55) begin // @[SelectPolicy.scala 151:14]
      age_7_9 <= ~age_9_9 & ~nextAge_7_9_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_7_10 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[7]) begin // @[SelectPolicy.scala 137:33]
      age_7_10 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[10]) begin // @[SelectPolicy.scala 140:34]
      age_7_10 <= thisValid_7; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_55) begin // @[SelectPolicy.scala 151:14]
      age_7_10 <= ~age_10_10 & ~nextAge_7_10_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_7_11 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[7]) begin // @[SelectPolicy.scala 137:33]
      age_7_11 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[11]) begin // @[SelectPolicy.scala 140:34]
      age_7_11 <= thisValid_7; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_55) begin // @[SelectPolicy.scala 151:14]
      age_7_11 <= ~age_11_11 & ~nextAge_7_11_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_7_12 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[7]) begin // @[SelectPolicy.scala 137:33]
      age_7_12 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[12]) begin // @[SelectPolicy.scala 140:34]
      age_7_12 <= thisValid_7; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_55) begin // @[SelectPolicy.scala 151:14]
      age_7_12 <= ~age_12_12 & ~nextAge_7_12_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_7_13 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[7]) begin // @[SelectPolicy.scala 137:33]
      age_7_13 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[13]) begin // @[SelectPolicy.scala 140:34]
      age_7_13 <= thisValid_7; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_55) begin // @[SelectPolicy.scala 151:14]
      age_7_13 <= ~age_13_13 & ~nextAge_7_13_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_7_14 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[7]) begin // @[SelectPolicy.scala 137:33]
      age_7_14 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[14]) begin // @[SelectPolicy.scala 140:34]
      age_7_14 <= thisValid_7; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_55) begin // @[SelectPolicy.scala 151:14]
      age_7_14 <= ~age_14_14 & ~nextAge_7_14_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_7_15 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[7]) begin // @[SelectPolicy.scala 137:33]
      age_7_15 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[15]) begin // @[SelectPolicy.scala 140:34]
      age_7_15 <= thisValid_7; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_55) begin // @[SelectPolicy.scala 151:14]
      age_7_15 <= ~age_15_15 & ~nextAge_7_15_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_8_8 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[8]) begin // @[SelectPolicy.scala 137:33]
      age_8_8 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[8]) begin // @[SelectPolicy.scala 140:34]
      age_8_8 <= thisValid_8; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_62) begin // @[SelectPolicy.scala 151:14]
      age_8_8 <= ~age_8_8 & ~nextAge_8_8_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_8_9 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[8]) begin // @[SelectPolicy.scala 137:33]
      age_8_9 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[9]) begin // @[SelectPolicy.scala 140:34]
      age_8_9 <= thisValid_8; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_62) begin // @[SelectPolicy.scala 151:14]
      age_8_9 <= ~age_9_9 & ~nextAge_8_9_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_8_10 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[8]) begin // @[SelectPolicy.scala 137:33]
      age_8_10 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[10]) begin // @[SelectPolicy.scala 140:34]
      age_8_10 <= thisValid_8; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_62) begin // @[SelectPolicy.scala 151:14]
      age_8_10 <= ~age_10_10 & ~nextAge_8_10_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_8_11 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[8]) begin // @[SelectPolicy.scala 137:33]
      age_8_11 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[11]) begin // @[SelectPolicy.scala 140:34]
      age_8_11 <= thisValid_8; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_62) begin // @[SelectPolicy.scala 151:14]
      age_8_11 <= ~age_11_11 & ~nextAge_8_11_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_8_12 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[8]) begin // @[SelectPolicy.scala 137:33]
      age_8_12 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[12]) begin // @[SelectPolicy.scala 140:34]
      age_8_12 <= thisValid_8; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_62) begin // @[SelectPolicy.scala 151:14]
      age_8_12 <= ~age_12_12 & ~nextAge_8_12_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_8_13 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[8]) begin // @[SelectPolicy.scala 137:33]
      age_8_13 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[13]) begin // @[SelectPolicy.scala 140:34]
      age_8_13 <= thisValid_8; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_62) begin // @[SelectPolicy.scala 151:14]
      age_8_13 <= ~age_13_13 & ~nextAge_8_13_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_8_14 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[8]) begin // @[SelectPolicy.scala 137:33]
      age_8_14 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[14]) begin // @[SelectPolicy.scala 140:34]
      age_8_14 <= thisValid_8; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_62) begin // @[SelectPolicy.scala 151:14]
      age_8_14 <= ~age_14_14 & ~nextAge_8_14_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_8_15 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[8]) begin // @[SelectPolicy.scala 137:33]
      age_8_15 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[15]) begin // @[SelectPolicy.scala 140:34]
      age_8_15 <= thisValid_8; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_62) begin // @[SelectPolicy.scala 151:14]
      age_8_15 <= ~age_15_15 & ~nextAge_8_15_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_9_9 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[9]) begin // @[SelectPolicy.scala 137:33]
      age_9_9 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[9]) begin // @[SelectPolicy.scala 140:34]
      age_9_9 <= thisValid_9; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_69) begin // @[SelectPolicy.scala 151:14]
      age_9_9 <= ~age_9_9 & ~nextAge_9_9_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_9_10 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[9]) begin // @[SelectPolicy.scala 137:33]
      age_9_10 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[10]) begin // @[SelectPolicy.scala 140:34]
      age_9_10 <= thisValid_9; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_69) begin // @[SelectPolicy.scala 151:14]
      age_9_10 <= ~age_10_10 & ~nextAge_9_10_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_9_11 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[9]) begin // @[SelectPolicy.scala 137:33]
      age_9_11 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[11]) begin // @[SelectPolicy.scala 140:34]
      age_9_11 <= thisValid_9; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_69) begin // @[SelectPolicy.scala 151:14]
      age_9_11 <= ~age_11_11 & ~nextAge_9_11_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_9_12 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[9]) begin // @[SelectPolicy.scala 137:33]
      age_9_12 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[12]) begin // @[SelectPolicy.scala 140:34]
      age_9_12 <= thisValid_9; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_69) begin // @[SelectPolicy.scala 151:14]
      age_9_12 <= ~age_12_12 & ~nextAge_9_12_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_9_13 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[9]) begin // @[SelectPolicy.scala 137:33]
      age_9_13 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[13]) begin // @[SelectPolicy.scala 140:34]
      age_9_13 <= thisValid_9; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_69) begin // @[SelectPolicy.scala 151:14]
      age_9_13 <= ~age_13_13 & ~nextAge_9_13_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_9_14 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[9]) begin // @[SelectPolicy.scala 137:33]
      age_9_14 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[14]) begin // @[SelectPolicy.scala 140:34]
      age_9_14 <= thisValid_9; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_69) begin // @[SelectPolicy.scala 151:14]
      age_9_14 <= ~age_14_14 & ~nextAge_9_14_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_9_15 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[9]) begin // @[SelectPolicy.scala 137:33]
      age_9_15 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[15]) begin // @[SelectPolicy.scala 140:34]
      age_9_15 <= thisValid_9; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_69) begin // @[SelectPolicy.scala 151:14]
      age_9_15 <= ~age_15_15 & ~nextAge_9_15_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_10_10 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[10]) begin // @[SelectPolicy.scala 137:33]
      age_10_10 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[10]) begin // @[SelectPolicy.scala 140:34]
      age_10_10 <= thisValid_10; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_76) begin // @[SelectPolicy.scala 151:14]
      age_10_10 <= ~age_10_10 & ~nextAge_10_10_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_10_11 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[10]) begin // @[SelectPolicy.scala 137:33]
      age_10_11 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[11]) begin // @[SelectPolicy.scala 140:34]
      age_10_11 <= thisValid_10; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_76) begin // @[SelectPolicy.scala 151:14]
      age_10_11 <= ~age_11_11 & ~nextAge_10_11_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_10_12 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[10]) begin // @[SelectPolicy.scala 137:33]
      age_10_12 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[12]) begin // @[SelectPolicy.scala 140:34]
      age_10_12 <= thisValid_10; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_76) begin // @[SelectPolicy.scala 151:14]
      age_10_12 <= ~age_12_12 & ~nextAge_10_12_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_10_13 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[10]) begin // @[SelectPolicy.scala 137:33]
      age_10_13 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[13]) begin // @[SelectPolicy.scala 140:34]
      age_10_13 <= thisValid_10; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_76) begin // @[SelectPolicy.scala 151:14]
      age_10_13 <= ~age_13_13 & ~nextAge_10_13_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_10_14 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[10]) begin // @[SelectPolicy.scala 137:33]
      age_10_14 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[14]) begin // @[SelectPolicy.scala 140:34]
      age_10_14 <= thisValid_10; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_76) begin // @[SelectPolicy.scala 151:14]
      age_10_14 <= ~age_14_14 & ~nextAge_10_14_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_10_15 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[10]) begin // @[SelectPolicy.scala 137:33]
      age_10_15 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[15]) begin // @[SelectPolicy.scala 140:34]
      age_10_15 <= thisValid_10; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_76) begin // @[SelectPolicy.scala 151:14]
      age_10_15 <= ~age_15_15 & ~nextAge_10_15_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_11_11 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[11]) begin // @[SelectPolicy.scala 137:33]
      age_11_11 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[11]) begin // @[SelectPolicy.scala 140:34]
      age_11_11 <= thisValid_11; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_83) begin // @[SelectPolicy.scala 151:14]
      age_11_11 <= ~age_11_11 & ~nextAge_11_11_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_11_12 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[11]) begin // @[SelectPolicy.scala 137:33]
      age_11_12 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[12]) begin // @[SelectPolicy.scala 140:34]
      age_11_12 <= thisValid_11; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_83) begin // @[SelectPolicy.scala 151:14]
      age_11_12 <= ~age_12_12 & ~nextAge_11_12_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_11_13 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[11]) begin // @[SelectPolicy.scala 137:33]
      age_11_13 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[13]) begin // @[SelectPolicy.scala 140:34]
      age_11_13 <= thisValid_11; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_83) begin // @[SelectPolicy.scala 151:14]
      age_11_13 <= ~age_13_13 & ~nextAge_11_13_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_11_14 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[11]) begin // @[SelectPolicy.scala 137:33]
      age_11_14 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[14]) begin // @[SelectPolicy.scala 140:34]
      age_11_14 <= thisValid_11; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_83) begin // @[SelectPolicy.scala 151:14]
      age_11_14 <= ~age_14_14 & ~nextAge_11_14_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_11_15 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[11]) begin // @[SelectPolicy.scala 137:33]
      age_11_15 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[15]) begin // @[SelectPolicy.scala 140:34]
      age_11_15 <= thisValid_11; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_83) begin // @[SelectPolicy.scala 151:14]
      age_11_15 <= ~age_15_15 & ~nextAge_11_15_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_12_12 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[12]) begin // @[SelectPolicy.scala 137:33]
      age_12_12 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[12]) begin // @[SelectPolicy.scala 140:34]
      age_12_12 <= thisValid_12; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_90) begin // @[SelectPolicy.scala 151:14]
      age_12_12 <= ~age_12_12 & ~nextAge_12_12_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_12_13 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[12]) begin // @[SelectPolicy.scala 137:33]
      age_12_13 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[13]) begin // @[SelectPolicy.scala 140:34]
      age_12_13 <= thisValid_12; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_90) begin // @[SelectPolicy.scala 151:14]
      age_12_13 <= ~age_13_13 & ~nextAge_12_13_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_12_14 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[12]) begin // @[SelectPolicy.scala 137:33]
      age_12_14 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[14]) begin // @[SelectPolicy.scala 140:34]
      age_12_14 <= thisValid_12; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_90) begin // @[SelectPolicy.scala 151:14]
      age_12_14 <= ~age_14_14 & ~nextAge_12_14_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_12_15 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[12]) begin // @[SelectPolicy.scala 137:33]
      age_12_15 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[15]) begin // @[SelectPolicy.scala 140:34]
      age_12_15 <= thisValid_12; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_90) begin // @[SelectPolicy.scala 151:14]
      age_12_15 <= ~age_15_15 & ~nextAge_12_15_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_13_13 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[13]) begin // @[SelectPolicy.scala 137:33]
      age_13_13 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[13]) begin // @[SelectPolicy.scala 140:34]
      age_13_13 <= thisValid_13; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_97) begin // @[SelectPolicy.scala 151:14]
      age_13_13 <= ~age_13_13 & ~nextAge_13_13_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_13_14 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[13]) begin // @[SelectPolicy.scala 137:33]
      age_13_14 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[14]) begin // @[SelectPolicy.scala 140:34]
      age_13_14 <= thisValid_13; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_97) begin // @[SelectPolicy.scala 151:14]
      age_13_14 <= ~age_14_14 & ~nextAge_13_14_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_13_15 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[13]) begin // @[SelectPolicy.scala 137:33]
      age_13_15 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[15]) begin // @[SelectPolicy.scala 140:34]
      age_13_15 <= thisValid_13; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_97) begin // @[SelectPolicy.scala 151:14]
      age_13_15 <= ~age_15_15 & ~nextAge_13_15_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_14_14 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[14]) begin // @[SelectPolicy.scala 137:33]
      age_14_14 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[14]) begin // @[SelectPolicy.scala 140:34]
      age_14_14 <= thisValid_14; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_104) begin // @[SelectPolicy.scala 151:14]
      age_14_14 <= ~age_14_14 & ~nextAge_14_14_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_14_15 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[14]) begin // @[SelectPolicy.scala 137:33]
      age_14_15 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[15]) begin // @[SelectPolicy.scala 140:34]
      age_14_15 <= thisValid_14; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_104) begin // @[SelectPolicy.scala 151:14]
      age_14_15 <= ~age_15_15 & ~nextAge_14_15_xs_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SelectPolicy.scala 134:27]
      age_15_15 <= 1'h0; // @[SelectPolicy.scala 136:14]
    end else if (io_deq[15]) begin // @[SelectPolicy.scala 137:33]
      age_15_15 <= 1'h0; // @[SelectPolicy.scala 139:14]
    end else if (io_deq[15]) begin // @[SelectPolicy.scala 140:34]
      age_15_15 <= thisValid_15; // @[SelectPolicy.scala 148:14]
    end else if (_thisValid_T_111) begin // @[SelectPolicy.scala 151:14]
      age_15_15 <= ~age_15_15 & ~nextAge_15_15_xs_1;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  age_0_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  age_0_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  age_0_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  age_0_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  age_0_4 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  age_0_5 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  age_0_6 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  age_0_7 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  age_0_8 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  age_0_9 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  age_0_10 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  age_0_11 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  age_0_12 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  age_0_13 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  age_0_14 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  age_0_15 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  age_1_1 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  age_1_2 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  age_1_3 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  age_1_4 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  age_1_5 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  age_1_6 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  age_1_7 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  age_1_8 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  age_1_9 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  age_1_10 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  age_1_11 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  age_1_12 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  age_1_13 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  age_1_14 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  age_1_15 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  age_2_2 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  age_2_3 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  age_2_4 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  age_2_5 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  age_2_6 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  age_2_7 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  age_2_8 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  age_2_9 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  age_2_10 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  age_2_11 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  age_2_12 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  age_2_13 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  age_2_14 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  age_2_15 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  age_3_3 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  age_3_4 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  age_3_5 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  age_3_6 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  age_3_7 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  age_3_8 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  age_3_9 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  age_3_10 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  age_3_11 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  age_3_12 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  age_3_13 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  age_3_14 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  age_3_15 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  age_4_4 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  age_4_5 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  age_4_6 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  age_4_7 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  age_4_8 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  age_4_9 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  age_4_10 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  age_4_11 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  age_4_12 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  age_4_13 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  age_4_14 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  age_4_15 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  age_5_5 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  age_5_6 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  age_5_7 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  age_5_8 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  age_5_9 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  age_5_10 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  age_5_11 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  age_5_12 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  age_5_13 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  age_5_14 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  age_5_15 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  age_6_6 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  age_6_7 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  age_6_8 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  age_6_9 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  age_6_10 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  age_6_11 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  age_6_12 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  age_6_13 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  age_6_14 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  age_6_15 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  age_7_7 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  age_7_8 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  age_7_9 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  age_7_10 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  age_7_11 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  age_7_12 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  age_7_13 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  age_7_14 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  age_7_15 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  age_8_8 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  age_8_9 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  age_8_10 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  age_8_11 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  age_8_12 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  age_8_13 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  age_8_14 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  age_8_15 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  age_9_9 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  age_9_10 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  age_9_11 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  age_9_12 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  age_9_13 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  age_9_14 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  age_9_15 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  age_10_10 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  age_10_11 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  age_10_12 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  age_10_13 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  age_10_14 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  age_10_15 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  age_11_11 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  age_11_12 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  age_11_13 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  age_11_14 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  age_11_15 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  age_12_12 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  age_12_13 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  age_12_14 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  age_12_15 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  age_13_13 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  age_13_14 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  age_13_15 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  age_14_14 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  age_14_15 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  age_15_15 = _RAND_135[0:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    age_0_0 = 1'h0;
  end
  if (reset) begin
    age_0_1 = 1'h0;
  end
  if (reset) begin
    age_0_2 = 1'h0;
  end
  if (reset) begin
    age_0_3 = 1'h0;
  end
  if (reset) begin
    age_0_4 = 1'h0;
  end
  if (reset) begin
    age_0_5 = 1'h0;
  end
  if (reset) begin
    age_0_6 = 1'h0;
  end
  if (reset) begin
    age_0_7 = 1'h0;
  end
  if (reset) begin
    age_0_8 = 1'h0;
  end
  if (reset) begin
    age_0_9 = 1'h0;
  end
  if (reset) begin
    age_0_10 = 1'h0;
  end
  if (reset) begin
    age_0_11 = 1'h0;
  end
  if (reset) begin
    age_0_12 = 1'h0;
  end
  if (reset) begin
    age_0_13 = 1'h0;
  end
  if (reset) begin
    age_0_14 = 1'h0;
  end
  if (reset) begin
    age_0_15 = 1'h0;
  end
  if (reset) begin
    age_1_1 = 1'h0;
  end
  if (reset) begin
    age_1_2 = 1'h0;
  end
  if (reset) begin
    age_1_3 = 1'h0;
  end
  if (reset) begin
    age_1_4 = 1'h0;
  end
  if (reset) begin
    age_1_5 = 1'h0;
  end
  if (reset) begin
    age_1_6 = 1'h0;
  end
  if (reset) begin
    age_1_7 = 1'h0;
  end
  if (reset) begin
    age_1_8 = 1'h0;
  end
  if (reset) begin
    age_1_9 = 1'h0;
  end
  if (reset) begin
    age_1_10 = 1'h0;
  end
  if (reset) begin
    age_1_11 = 1'h0;
  end
  if (reset) begin
    age_1_12 = 1'h0;
  end
  if (reset) begin
    age_1_13 = 1'h0;
  end
  if (reset) begin
    age_1_14 = 1'h0;
  end
  if (reset) begin
    age_1_15 = 1'h0;
  end
  if (reset) begin
    age_2_2 = 1'h0;
  end
  if (reset) begin
    age_2_3 = 1'h0;
  end
  if (reset) begin
    age_2_4 = 1'h0;
  end
  if (reset) begin
    age_2_5 = 1'h0;
  end
  if (reset) begin
    age_2_6 = 1'h0;
  end
  if (reset) begin
    age_2_7 = 1'h0;
  end
  if (reset) begin
    age_2_8 = 1'h0;
  end
  if (reset) begin
    age_2_9 = 1'h0;
  end
  if (reset) begin
    age_2_10 = 1'h0;
  end
  if (reset) begin
    age_2_11 = 1'h0;
  end
  if (reset) begin
    age_2_12 = 1'h0;
  end
  if (reset) begin
    age_2_13 = 1'h0;
  end
  if (reset) begin
    age_2_14 = 1'h0;
  end
  if (reset) begin
    age_2_15 = 1'h0;
  end
  if (reset) begin
    age_3_3 = 1'h0;
  end
  if (reset) begin
    age_3_4 = 1'h0;
  end
  if (reset) begin
    age_3_5 = 1'h0;
  end
  if (reset) begin
    age_3_6 = 1'h0;
  end
  if (reset) begin
    age_3_7 = 1'h0;
  end
  if (reset) begin
    age_3_8 = 1'h0;
  end
  if (reset) begin
    age_3_9 = 1'h0;
  end
  if (reset) begin
    age_3_10 = 1'h0;
  end
  if (reset) begin
    age_3_11 = 1'h0;
  end
  if (reset) begin
    age_3_12 = 1'h0;
  end
  if (reset) begin
    age_3_13 = 1'h0;
  end
  if (reset) begin
    age_3_14 = 1'h0;
  end
  if (reset) begin
    age_3_15 = 1'h0;
  end
  if (reset) begin
    age_4_4 = 1'h0;
  end
  if (reset) begin
    age_4_5 = 1'h0;
  end
  if (reset) begin
    age_4_6 = 1'h0;
  end
  if (reset) begin
    age_4_7 = 1'h0;
  end
  if (reset) begin
    age_4_8 = 1'h0;
  end
  if (reset) begin
    age_4_9 = 1'h0;
  end
  if (reset) begin
    age_4_10 = 1'h0;
  end
  if (reset) begin
    age_4_11 = 1'h0;
  end
  if (reset) begin
    age_4_12 = 1'h0;
  end
  if (reset) begin
    age_4_13 = 1'h0;
  end
  if (reset) begin
    age_4_14 = 1'h0;
  end
  if (reset) begin
    age_4_15 = 1'h0;
  end
  if (reset) begin
    age_5_5 = 1'h0;
  end
  if (reset) begin
    age_5_6 = 1'h0;
  end
  if (reset) begin
    age_5_7 = 1'h0;
  end
  if (reset) begin
    age_5_8 = 1'h0;
  end
  if (reset) begin
    age_5_9 = 1'h0;
  end
  if (reset) begin
    age_5_10 = 1'h0;
  end
  if (reset) begin
    age_5_11 = 1'h0;
  end
  if (reset) begin
    age_5_12 = 1'h0;
  end
  if (reset) begin
    age_5_13 = 1'h0;
  end
  if (reset) begin
    age_5_14 = 1'h0;
  end
  if (reset) begin
    age_5_15 = 1'h0;
  end
  if (reset) begin
    age_6_6 = 1'h0;
  end
  if (reset) begin
    age_6_7 = 1'h0;
  end
  if (reset) begin
    age_6_8 = 1'h0;
  end
  if (reset) begin
    age_6_9 = 1'h0;
  end
  if (reset) begin
    age_6_10 = 1'h0;
  end
  if (reset) begin
    age_6_11 = 1'h0;
  end
  if (reset) begin
    age_6_12 = 1'h0;
  end
  if (reset) begin
    age_6_13 = 1'h0;
  end
  if (reset) begin
    age_6_14 = 1'h0;
  end
  if (reset) begin
    age_6_15 = 1'h0;
  end
  if (reset) begin
    age_7_7 = 1'h0;
  end
  if (reset) begin
    age_7_8 = 1'h0;
  end
  if (reset) begin
    age_7_9 = 1'h0;
  end
  if (reset) begin
    age_7_10 = 1'h0;
  end
  if (reset) begin
    age_7_11 = 1'h0;
  end
  if (reset) begin
    age_7_12 = 1'h0;
  end
  if (reset) begin
    age_7_13 = 1'h0;
  end
  if (reset) begin
    age_7_14 = 1'h0;
  end
  if (reset) begin
    age_7_15 = 1'h0;
  end
  if (reset) begin
    age_8_8 = 1'h0;
  end
  if (reset) begin
    age_8_9 = 1'h0;
  end
  if (reset) begin
    age_8_10 = 1'h0;
  end
  if (reset) begin
    age_8_11 = 1'h0;
  end
  if (reset) begin
    age_8_12 = 1'h0;
  end
  if (reset) begin
    age_8_13 = 1'h0;
  end
  if (reset) begin
    age_8_14 = 1'h0;
  end
  if (reset) begin
    age_8_15 = 1'h0;
  end
  if (reset) begin
    age_9_9 = 1'h0;
  end
  if (reset) begin
    age_9_10 = 1'h0;
  end
  if (reset) begin
    age_9_11 = 1'h0;
  end
  if (reset) begin
    age_9_12 = 1'h0;
  end
  if (reset) begin
    age_9_13 = 1'h0;
  end
  if (reset) begin
    age_9_14 = 1'h0;
  end
  if (reset) begin
    age_9_15 = 1'h0;
  end
  if (reset) begin
    age_10_10 = 1'h0;
  end
  if (reset) begin
    age_10_11 = 1'h0;
  end
  if (reset) begin
    age_10_12 = 1'h0;
  end
  if (reset) begin
    age_10_13 = 1'h0;
  end
  if (reset) begin
    age_10_14 = 1'h0;
  end
  if (reset) begin
    age_10_15 = 1'h0;
  end
  if (reset) begin
    age_11_11 = 1'h0;
  end
  if (reset) begin
    age_11_12 = 1'h0;
  end
  if (reset) begin
    age_11_13 = 1'h0;
  end
  if (reset) begin
    age_11_14 = 1'h0;
  end
  if (reset) begin
    age_11_15 = 1'h0;
  end
  if (reset) begin
    age_12_12 = 1'h0;
  end
  if (reset) begin
    age_12_13 = 1'h0;
  end
  if (reset) begin
    age_12_14 = 1'h0;
  end
  if (reset) begin
    age_12_15 = 1'h0;
  end
  if (reset) begin
    age_13_13 = 1'h0;
  end
  if (reset) begin
    age_13_14 = 1'h0;
  end
  if (reset) begin
    age_13_15 = 1'h0;
  end
  if (reset) begin
    age_14_14 = 1'h0;
  end
  if (reset) begin
    age_14_15 = 1'h0;
  end
  if (reset) begin
    age_15_15 = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule

