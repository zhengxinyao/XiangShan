module NegedgeDataModule__64entry_32(
  input        clock,
  input  [5:0] io_raddr_0,
  input  [5:0] io_raddr_1,
  output [4:0] io_rdata_0_ssid,
  output       io_rdata_0_strict,
  output [4:0] io_rdata_1_ssid,
  output       io_rdata_1_strict,
  input        io_wen_0,
  input        io_wen_1,
  input  [5:0] io_waddr_0,
  input  [5:0] io_waddr_1,
  input  [4:0] io_wdata_0_ssid,
  input        io_wdata_0_strict,
  input  [4:0] io_wdata_1_ssid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
`endif // RANDOMIZE_REG_INIT
  reg [4:0] data_0_ssid; // @[DataModuleTemplate.scala 168:17]
  reg  data_0_strict; // @[DataModuleTemplate.scala 168:17]
  reg [4:0] data_1_ssid; // @[DataModuleTemplate.scala 168:17]
  reg  data_1_strict; // @[DataModuleTemplate.scala 168:17]
  reg [4:0] data_2_ssid; // @[DataModuleTemplate.scala 168:17]
  reg  data_2_strict; // @[DataModuleTemplate.scala 168:17]
  reg [4:0] data_3_ssid; // @[DataModuleTemplate.scala 168:17]
  reg  data_3_strict; // @[DataModuleTemplate.scala 168:17]
  reg [4:0] data_4_ssid; // @[DataModuleTemplate.scala 168:17]
  reg  data_4_strict; // @[DataModuleTemplate.scala 168:17]
  reg [4:0] data_5_ssid; // @[DataModuleTemplate.scala 168:17]
  reg  data_5_strict; // @[DataModuleTemplate.scala 168:17]
  reg [4:0] data_6_ssid; // @[DataModuleTemplate.scala 168:17]
  reg  data_6_strict; // @[DataModuleTemplate.scala 168:17]
  reg [4:0] data_7_ssid; // @[DataModuleTemplate.scala 168:17]
  reg  data_7_strict; // @[DataModuleTemplate.scala 168:17]
  reg [4:0] data_8_ssid; // @[DataModuleTemplate.scala 168:17]
  reg  data_8_strict; // @[DataModuleTemplate.scala 168:17]
  reg [4:0] data_9_ssid; // @[DataModuleTemplate.scala 168:17]
  reg  data_9_strict; // @[DataModuleTemplate.scala 168:17]
  reg [4:0] data_10_ssid; // @[DataModuleTemplate.scala 168:17]
  reg  data_10_strict; // @[DataModuleTemplate.scala 168:17]
  reg [4:0] data_11_ssid; // @[DataModuleTemplate.scala 168:17]
  reg  data_11_strict; // @[DataModuleTemplate.scala 168:17]
  reg [4:0] data_12_ssid; // @[DataModuleTemplate.scala 168:17]
  reg  data_12_strict; // @[DataModuleTemplate.scala 168:17]
  reg [4:0] data_13_ssid; // @[DataModuleTemplate.scala 168:17]
  reg  data_13_strict; // @[DataModuleTemplate.scala 168:17]
  reg [4:0] data_14_ssid; // @[DataModuleTemplate.scala 168:17]
  reg  data_14_strict; // @[DataModuleTemplate.scala 168:17]
  reg [4:0] data_15_ssid; // @[DataModuleTemplate.scala 168:17]
  reg  data_15_strict; // @[DataModuleTemplate.scala 168:17]
  reg [4:0] data_16_ssid; // @[DataModuleTemplate.scala 168:17]
  reg  data_16_strict; // @[DataModuleTemplate.scala 168:17]
  reg [4:0] data_17_ssid; // @[DataModuleTemplate.scala 168:17]
  reg  data_17_strict; // @[DataModuleTemplate.scala 168:17]
  reg [4:0] data_18_ssid; // @[DataModuleTemplate.scala 168:17]
  reg  data_18_strict; // @[DataModuleTemplate.scala 168:17]
  reg [4:0] data_19_ssid; // @[DataModuleTemplate.scala 168:17]
  reg  data_19_strict; // @[DataModuleTemplate.scala 168:17]
  reg [4:0] data_20_ssid; // @[DataModuleTemplate.scala 168:17]
  reg  data_20_strict; // @[DataModuleTemplate.scala 168:17]
  reg [4:0] data_21_ssid; // @[DataModuleTemplate.scala 168:17]
  reg  data_21_strict; // @[DataModuleTemplate.scala 168:17]
  reg [4:0] data_22_ssid; // @[DataModuleTemplate.scala 168:17]
  reg  data_22_strict; // @[DataModuleTemplate.scala 168:17]
  reg [4:0] data_23_ssid; // @[DataModuleTemplate.scala 168:17]
  reg  data_23_strict; // @[DataModuleTemplate.scala 168:17]
  reg [4:0] data_24_ssid; // @[DataModuleTemplate.scala 168:17]
  reg  data_24_strict; // @[DataModuleTemplate.scala 168:17]
  reg [4:0] data_25_ssid; // @[DataModuleTemplate.scala 168:17]
  reg  data_25_strict; // @[DataModuleTemplate.scala 168:17]
  reg [4:0] data_26_ssid; // @[DataModuleTemplate.scala 168:17]
  reg  data_26_strict; // @[DataModuleTemplate.scala 168:17]
  reg [4:0] data_27_ssid; // @[DataModuleTemplate.scala 168:17]
  reg  data_27_strict; // @[DataModuleTemplate.scala 168:17]
  reg [4:0] data_28_ssid; // @[DataModuleTemplate.scala 168:17]
  reg  data_28_strict; // @[DataModuleTemplate.scala 168:17]
  reg [4:0] data_29_ssid; // @[DataModuleTemplate.scala 168:17]
  reg  data_29_strict; // @[DataModuleTemplate.scala 168:17]
  reg [4:0] data_30_ssid; // @[DataModuleTemplate.scala 168:17]
  reg  data_30_strict; // @[DataModuleTemplate.scala 168:17]
  reg [4:0] data_31_ssid; // @[DataModuleTemplate.scala 168:17]
  reg  data_31_strict; // @[DataModuleTemplate.scala 168:17]
  reg [4:0] data_32_ssid; // @[DataModuleTemplate.scala 168:17]
  reg  data_32_strict; // @[DataModuleTemplate.scala 168:17]
  reg [4:0] data_33_ssid; // @[DataModuleTemplate.scala 168:17]
  reg  data_33_strict; // @[DataModuleTemplate.scala 168:17]
  reg [4:0] data_34_ssid; // @[DataModuleTemplate.scala 168:17]
  reg  data_34_strict; // @[DataModuleTemplate.scala 168:17]
  reg [4:0] data_35_ssid; // @[DataModuleTemplate.scala 168:17]
  reg  data_35_strict; // @[DataModuleTemplate.scala 168:17]
  reg [4:0] data_36_ssid; // @[DataModuleTemplate.scala 168:17]
  reg  data_36_strict; // @[DataModuleTemplate.scala 168:17]
  reg [4:0] data_37_ssid; // @[DataModuleTemplate.scala 168:17]
  reg  data_37_strict; // @[DataModuleTemplate.scala 168:17]
  reg [4:0] data_38_ssid; // @[DataModuleTemplate.scala 168:17]
  reg  data_38_strict; // @[DataModuleTemplate.scala 168:17]
  reg [4:0] data_39_ssid; // @[DataModuleTemplate.scala 168:17]
  reg  data_39_strict; // @[DataModuleTemplate.scala 168:17]
  reg [4:0] data_40_ssid; // @[DataModuleTemplate.scala 168:17]
  reg  data_40_strict; // @[DataModuleTemplate.scala 168:17]
  reg [4:0] data_41_ssid; // @[DataModuleTemplate.scala 168:17]
  reg  data_41_strict; // @[DataModuleTemplate.scala 168:17]
  reg [4:0] data_42_ssid; // @[DataModuleTemplate.scala 168:17]
  reg  data_42_strict; // @[DataModuleTemplate.scala 168:17]
  reg [4:0] data_43_ssid; // @[DataModuleTemplate.scala 168:17]
  reg  data_43_strict; // @[DataModuleTemplate.scala 168:17]
  reg [4:0] data_44_ssid; // @[DataModuleTemplate.scala 168:17]
  reg  data_44_strict; // @[DataModuleTemplate.scala 168:17]
  reg [4:0] data_45_ssid; // @[DataModuleTemplate.scala 168:17]
  reg  data_45_strict; // @[DataModuleTemplate.scala 168:17]
  reg [4:0] data_46_ssid; // @[DataModuleTemplate.scala 168:17]
  reg  data_46_strict; // @[DataModuleTemplate.scala 168:17]
  reg [4:0] data_47_ssid; // @[DataModuleTemplate.scala 168:17]
  reg  data_47_strict; // @[DataModuleTemplate.scala 168:17]
  reg [4:0] data_48_ssid; // @[DataModuleTemplate.scala 168:17]
  reg  data_48_strict; // @[DataModuleTemplate.scala 168:17]
  reg [4:0] data_49_ssid; // @[DataModuleTemplate.scala 168:17]
  reg  data_49_strict; // @[DataModuleTemplate.scala 168:17]
  reg [4:0] data_50_ssid; // @[DataModuleTemplate.scala 168:17]
  reg  data_50_strict; // @[DataModuleTemplate.scala 168:17]
  reg [4:0] data_51_ssid; // @[DataModuleTemplate.scala 168:17]
  reg  data_51_strict; // @[DataModuleTemplate.scala 168:17]
  reg [4:0] data_52_ssid; // @[DataModuleTemplate.scala 168:17]
  reg  data_52_strict; // @[DataModuleTemplate.scala 168:17]
  reg [4:0] data_53_ssid; // @[DataModuleTemplate.scala 168:17]
  reg  data_53_strict; // @[DataModuleTemplate.scala 168:17]
  reg [4:0] data_54_ssid; // @[DataModuleTemplate.scala 168:17]
  reg  data_54_strict; // @[DataModuleTemplate.scala 168:17]
  reg [4:0] data_55_ssid; // @[DataModuleTemplate.scala 168:17]
  reg  data_55_strict; // @[DataModuleTemplate.scala 168:17]
  reg [4:0] data_56_ssid; // @[DataModuleTemplate.scala 168:17]
  reg  data_56_strict; // @[DataModuleTemplate.scala 168:17]
  reg [4:0] data_57_ssid; // @[DataModuleTemplate.scala 168:17]
  reg  data_57_strict; // @[DataModuleTemplate.scala 168:17]
  reg [4:0] data_58_ssid; // @[DataModuleTemplate.scala 168:17]
  reg  data_58_strict; // @[DataModuleTemplate.scala 168:17]
  reg [4:0] data_59_ssid; // @[DataModuleTemplate.scala 168:17]
  reg  data_59_strict; // @[DataModuleTemplate.scala 168:17]
  reg [4:0] data_60_ssid; // @[DataModuleTemplate.scala 168:17]
  reg  data_60_strict; // @[DataModuleTemplate.scala 168:17]
  reg [4:0] data_61_ssid; // @[DataModuleTemplate.scala 168:17]
  reg  data_61_strict; // @[DataModuleTemplate.scala 168:17]
  reg [4:0] data_62_ssid; // @[DataModuleTemplate.scala 168:17]
  reg  data_62_strict; // @[DataModuleTemplate.scala 168:17]
  reg [4:0] data_63_ssid; // @[DataModuleTemplate.scala 168:17]
  reg  data_63_strict; // @[DataModuleTemplate.scala 168:17]
  wire  read_by_0 = io_wen_0 & io_waddr_0 == io_raddr_0; // @[DataModuleTemplate.scala 176:54]
  wire  read_by_1 = io_wen_1 & io_waddr_1 == io_raddr_0; // @[DataModuleTemplate.scala 176:54]
  wire [63:0] addr_dec = 64'h1 << io_raddr_0; // @[OneHot.scala 64:12]
  wire [1:0] _T = {read_by_1,read_by_0}; // @[DataModuleTemplate.scala 178:28]
  wire  _io_rdata_0_T = read_by_0 & io_wdata_0_strict; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_3 = read_by_0 ? io_wdata_0_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_4 = read_by_1 ? io_wdata_1_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_5 = _io_rdata_0_T_3 | _io_rdata_0_T_4; // @[Mux.scala 27:73]
  wire  _io_rdata_0_T_85 = addr_dec[15] & data_15_strict; // @[Mux.scala 27:73]
  wire  _io_rdata_0_T_148 = addr_dec[0] & data_0_strict | addr_dec[1] & data_1_strict | addr_dec[2] & data_2_strict |
    addr_dec[3] & data_3_strict | addr_dec[4] & data_4_strict | addr_dec[5] & data_5_strict | addr_dec[6] &
    data_6_strict | addr_dec[7] & data_7_strict | addr_dec[8] & data_8_strict | addr_dec[9] & data_9_strict | addr_dec[
    10] & data_10_strict | addr_dec[11] & data_11_strict | addr_dec[12] & data_12_strict | addr_dec[13] & data_13_strict
     | addr_dec[14] & data_14_strict | _io_rdata_0_T_85; // @[Mux.scala 27:73]
  wire  _io_rdata_0_T_163 = _io_rdata_0_T_148 | addr_dec[16] & data_16_strict | addr_dec[17] & data_17_strict | addr_dec
    [18] & data_18_strict | addr_dec[19] & data_19_strict | addr_dec[20] & data_20_strict | addr_dec[21] &
    data_21_strict | addr_dec[22] & data_22_strict | addr_dec[23] & data_23_strict | addr_dec[24] & data_24_strict |
    addr_dec[25] & data_25_strict | addr_dec[26] & data_26_strict | addr_dec[27] & data_27_strict | addr_dec[28] &
    data_28_strict | addr_dec[29] & data_29_strict | addr_dec[30] & data_30_strict; // @[Mux.scala 27:73]
  wire  _io_rdata_0_T_178 = _io_rdata_0_T_163 | addr_dec[31] & data_31_strict | addr_dec[32] & data_32_strict | addr_dec
    [33] & data_33_strict | addr_dec[34] & data_34_strict | addr_dec[35] & data_35_strict | addr_dec[36] &
    data_36_strict | addr_dec[37] & data_37_strict | addr_dec[38] & data_38_strict | addr_dec[39] & data_39_strict |
    addr_dec[40] & data_40_strict | addr_dec[41] & data_41_strict | addr_dec[42] & data_42_strict | addr_dec[43] &
    data_43_strict | addr_dec[44] & data_44_strict | addr_dec[45] & data_45_strict; // @[Mux.scala 27:73]
  wire  _io_rdata_0_T_193 = _io_rdata_0_T_178 | addr_dec[46] & data_46_strict | addr_dec[47] & data_47_strict | addr_dec
    [48] & data_48_strict | addr_dec[49] & data_49_strict | addr_dec[50] & data_50_strict | addr_dec[51] &
    data_51_strict | addr_dec[52] & data_52_strict | addr_dec[53] & data_53_strict | addr_dec[54] & data_54_strict |
    addr_dec[55] & data_55_strict | addr_dec[56] & data_56_strict | addr_dec[57] & data_57_strict | addr_dec[58] &
    data_58_strict | addr_dec[59] & data_59_strict | addr_dec[60] & data_60_strict; // @[Mux.scala 27:73]
  wire  _io_rdata_0_T_196 = _io_rdata_0_T_193 | addr_dec[61] & data_61_strict | addr_dec[62] & data_62_strict | addr_dec
    [63] & data_63_strict; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_197 = addr_dec[0] ? data_0_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_198 = addr_dec[1] ? data_1_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_199 = addr_dec[2] ? data_2_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_200 = addr_dec[3] ? data_3_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_201 = addr_dec[4] ? data_4_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_202 = addr_dec[5] ? data_5_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_203 = addr_dec[6] ? data_6_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_204 = addr_dec[7] ? data_7_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_205 = addr_dec[8] ? data_8_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_206 = addr_dec[9] ? data_9_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_207 = addr_dec[10] ? data_10_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_208 = addr_dec[11] ? data_11_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_209 = addr_dec[12] ? data_12_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_210 = addr_dec[13] ? data_13_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_211 = addr_dec[14] ? data_14_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_212 = addr_dec[15] ? data_15_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_213 = addr_dec[16] ? data_16_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_214 = addr_dec[17] ? data_17_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_215 = addr_dec[18] ? data_18_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_216 = addr_dec[19] ? data_19_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_217 = addr_dec[20] ? data_20_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_218 = addr_dec[21] ? data_21_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_219 = addr_dec[22] ? data_22_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_220 = addr_dec[23] ? data_23_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_221 = addr_dec[24] ? data_24_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_222 = addr_dec[25] ? data_25_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_223 = addr_dec[26] ? data_26_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_224 = addr_dec[27] ? data_27_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_225 = addr_dec[28] ? data_28_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_226 = addr_dec[29] ? data_29_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_227 = addr_dec[30] ? data_30_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_228 = addr_dec[31] ? data_31_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_229 = addr_dec[32] ? data_32_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_230 = addr_dec[33] ? data_33_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_231 = addr_dec[34] ? data_34_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_232 = addr_dec[35] ? data_35_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_233 = addr_dec[36] ? data_36_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_234 = addr_dec[37] ? data_37_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_235 = addr_dec[38] ? data_38_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_236 = addr_dec[39] ? data_39_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_237 = addr_dec[40] ? data_40_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_238 = addr_dec[41] ? data_41_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_239 = addr_dec[42] ? data_42_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_240 = addr_dec[43] ? data_43_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_241 = addr_dec[44] ? data_44_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_242 = addr_dec[45] ? data_45_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_243 = addr_dec[46] ? data_46_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_244 = addr_dec[47] ? data_47_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_245 = addr_dec[48] ? data_48_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_246 = addr_dec[49] ? data_49_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_247 = addr_dec[50] ? data_50_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_248 = addr_dec[51] ? data_51_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_249 = addr_dec[52] ? data_52_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_250 = addr_dec[53] ? data_53_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_251 = addr_dec[54] ? data_54_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_252 = addr_dec[55] ? data_55_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_253 = addr_dec[56] ? data_56_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_254 = addr_dec[57] ? data_57_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_255 = addr_dec[58] ? data_58_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_256 = addr_dec[59] ? data_59_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_257 = addr_dec[60] ? data_60_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_258 = addr_dec[61] ? data_61_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_259 = addr_dec[62] ? data_62_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_260 = addr_dec[63] ? data_63_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_261 = _io_rdata_0_T_197 | _io_rdata_0_T_198; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_262 = _io_rdata_0_T_261 | _io_rdata_0_T_199; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_263 = _io_rdata_0_T_262 | _io_rdata_0_T_200; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_264 = _io_rdata_0_T_263 | _io_rdata_0_T_201; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_265 = _io_rdata_0_T_264 | _io_rdata_0_T_202; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_266 = _io_rdata_0_T_265 | _io_rdata_0_T_203; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_267 = _io_rdata_0_T_266 | _io_rdata_0_T_204; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_268 = _io_rdata_0_T_267 | _io_rdata_0_T_205; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_269 = _io_rdata_0_T_268 | _io_rdata_0_T_206; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_270 = _io_rdata_0_T_269 | _io_rdata_0_T_207; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_271 = _io_rdata_0_T_270 | _io_rdata_0_T_208; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_272 = _io_rdata_0_T_271 | _io_rdata_0_T_209; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_273 = _io_rdata_0_T_272 | _io_rdata_0_T_210; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_274 = _io_rdata_0_T_273 | _io_rdata_0_T_211; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_275 = _io_rdata_0_T_274 | _io_rdata_0_T_212; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_276 = _io_rdata_0_T_275 | _io_rdata_0_T_213; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_277 = _io_rdata_0_T_276 | _io_rdata_0_T_214; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_278 = _io_rdata_0_T_277 | _io_rdata_0_T_215; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_279 = _io_rdata_0_T_278 | _io_rdata_0_T_216; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_280 = _io_rdata_0_T_279 | _io_rdata_0_T_217; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_281 = _io_rdata_0_T_280 | _io_rdata_0_T_218; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_282 = _io_rdata_0_T_281 | _io_rdata_0_T_219; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_283 = _io_rdata_0_T_282 | _io_rdata_0_T_220; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_284 = _io_rdata_0_T_283 | _io_rdata_0_T_221; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_285 = _io_rdata_0_T_284 | _io_rdata_0_T_222; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_286 = _io_rdata_0_T_285 | _io_rdata_0_T_223; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_287 = _io_rdata_0_T_286 | _io_rdata_0_T_224; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_288 = _io_rdata_0_T_287 | _io_rdata_0_T_225; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_289 = _io_rdata_0_T_288 | _io_rdata_0_T_226; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_290 = _io_rdata_0_T_289 | _io_rdata_0_T_227; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_291 = _io_rdata_0_T_290 | _io_rdata_0_T_228; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_292 = _io_rdata_0_T_291 | _io_rdata_0_T_229; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_293 = _io_rdata_0_T_292 | _io_rdata_0_T_230; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_294 = _io_rdata_0_T_293 | _io_rdata_0_T_231; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_295 = _io_rdata_0_T_294 | _io_rdata_0_T_232; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_296 = _io_rdata_0_T_295 | _io_rdata_0_T_233; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_297 = _io_rdata_0_T_296 | _io_rdata_0_T_234; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_298 = _io_rdata_0_T_297 | _io_rdata_0_T_235; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_299 = _io_rdata_0_T_298 | _io_rdata_0_T_236; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_300 = _io_rdata_0_T_299 | _io_rdata_0_T_237; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_301 = _io_rdata_0_T_300 | _io_rdata_0_T_238; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_302 = _io_rdata_0_T_301 | _io_rdata_0_T_239; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_303 = _io_rdata_0_T_302 | _io_rdata_0_T_240; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_304 = _io_rdata_0_T_303 | _io_rdata_0_T_241; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_305 = _io_rdata_0_T_304 | _io_rdata_0_T_242; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_306 = _io_rdata_0_T_305 | _io_rdata_0_T_243; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_307 = _io_rdata_0_T_306 | _io_rdata_0_T_244; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_308 = _io_rdata_0_T_307 | _io_rdata_0_T_245; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_309 = _io_rdata_0_T_308 | _io_rdata_0_T_246; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_310 = _io_rdata_0_T_309 | _io_rdata_0_T_247; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_311 = _io_rdata_0_T_310 | _io_rdata_0_T_248; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_312 = _io_rdata_0_T_311 | _io_rdata_0_T_249; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_313 = _io_rdata_0_T_312 | _io_rdata_0_T_250; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_314 = _io_rdata_0_T_313 | _io_rdata_0_T_251; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_315 = _io_rdata_0_T_314 | _io_rdata_0_T_252; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_316 = _io_rdata_0_T_315 | _io_rdata_0_T_253; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_317 = _io_rdata_0_T_316 | _io_rdata_0_T_254; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_318 = _io_rdata_0_T_317 | _io_rdata_0_T_255; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_319 = _io_rdata_0_T_318 | _io_rdata_0_T_256; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_320 = _io_rdata_0_T_319 | _io_rdata_0_T_257; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_321 = _io_rdata_0_T_320 | _io_rdata_0_T_258; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_322 = _io_rdata_0_T_321 | _io_rdata_0_T_259; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_0_T_323 = _io_rdata_0_T_322 | _io_rdata_0_T_260; // @[Mux.scala 27:73]
  wire  read_by_0_1 = io_wen_0 & io_waddr_0 == io_raddr_1; // @[DataModuleTemplate.scala 176:54]
  wire  read_by_1_1 = io_wen_1 & io_waddr_1 == io_raddr_1; // @[DataModuleTemplate.scala 176:54]
  wire [63:0] addr_dec_1 = 64'h1 << io_raddr_1; // @[OneHot.scala 64:12]
  wire [1:0] _T_2 = {read_by_1_1,read_by_0_1}; // @[DataModuleTemplate.scala 178:28]
  wire  _io_rdata_1_T = read_by_0_1 & io_wdata_0_strict; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_3 = read_by_0_1 ? io_wdata_0_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_4 = read_by_1_1 ? io_wdata_1_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_5 = _io_rdata_1_T_3 | _io_rdata_1_T_4; // @[Mux.scala 27:73]
  wire  _io_rdata_1_T_85 = addr_dec_1[15] & data_15_strict; // @[Mux.scala 27:73]
  wire  _io_rdata_1_T_148 = addr_dec_1[0] & data_0_strict | addr_dec_1[1] & data_1_strict | addr_dec_1[2] &
    data_2_strict | addr_dec_1[3] & data_3_strict | addr_dec_1[4] & data_4_strict | addr_dec_1[5] & data_5_strict |
    addr_dec_1[6] & data_6_strict | addr_dec_1[7] & data_7_strict | addr_dec_1[8] & data_8_strict | addr_dec_1[9] &
    data_9_strict | addr_dec_1[10] & data_10_strict | addr_dec_1[11] & data_11_strict | addr_dec_1[12] & data_12_strict
     | addr_dec_1[13] & data_13_strict | addr_dec_1[14] & data_14_strict | _io_rdata_1_T_85; // @[Mux.scala 27:73]
  wire  _io_rdata_1_T_163 = _io_rdata_1_T_148 | addr_dec_1[16] & data_16_strict | addr_dec_1[17] & data_17_strict |
    addr_dec_1[18] & data_18_strict | addr_dec_1[19] & data_19_strict | addr_dec_1[20] & data_20_strict | addr_dec_1[21]
     & data_21_strict | addr_dec_1[22] & data_22_strict | addr_dec_1[23] & data_23_strict | addr_dec_1[24] &
    data_24_strict | addr_dec_1[25] & data_25_strict | addr_dec_1[26] & data_26_strict | addr_dec_1[27] & data_27_strict
     | addr_dec_1[28] & data_28_strict | addr_dec_1[29] & data_29_strict | addr_dec_1[30] & data_30_strict; // @[Mux.scala 27:73]
  wire  _io_rdata_1_T_178 = _io_rdata_1_T_163 | addr_dec_1[31] & data_31_strict | addr_dec_1[32] & data_32_strict |
    addr_dec_1[33] & data_33_strict | addr_dec_1[34] & data_34_strict | addr_dec_1[35] & data_35_strict | addr_dec_1[36]
     & data_36_strict | addr_dec_1[37] & data_37_strict | addr_dec_1[38] & data_38_strict | addr_dec_1[39] &
    data_39_strict | addr_dec_1[40] & data_40_strict | addr_dec_1[41] & data_41_strict | addr_dec_1[42] & data_42_strict
     | addr_dec_1[43] & data_43_strict | addr_dec_1[44] & data_44_strict | addr_dec_1[45] & data_45_strict; // @[Mux.scala 27:73]
  wire  _io_rdata_1_T_193 = _io_rdata_1_T_178 | addr_dec_1[46] & data_46_strict | addr_dec_1[47] & data_47_strict |
    addr_dec_1[48] & data_48_strict | addr_dec_1[49] & data_49_strict | addr_dec_1[50] & data_50_strict | addr_dec_1[51]
     & data_51_strict | addr_dec_1[52] & data_52_strict | addr_dec_1[53] & data_53_strict | addr_dec_1[54] &
    data_54_strict | addr_dec_1[55] & data_55_strict | addr_dec_1[56] & data_56_strict | addr_dec_1[57] & data_57_strict
     | addr_dec_1[58] & data_58_strict | addr_dec_1[59] & data_59_strict | addr_dec_1[60] & data_60_strict; // @[Mux.scala 27:73]
  wire  _io_rdata_1_T_196 = _io_rdata_1_T_193 | addr_dec_1[61] & data_61_strict | addr_dec_1[62] & data_62_strict |
    addr_dec_1[63] & data_63_strict; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_197 = addr_dec_1[0] ? data_0_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_198 = addr_dec_1[1] ? data_1_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_199 = addr_dec_1[2] ? data_2_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_200 = addr_dec_1[3] ? data_3_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_201 = addr_dec_1[4] ? data_4_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_202 = addr_dec_1[5] ? data_5_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_203 = addr_dec_1[6] ? data_6_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_204 = addr_dec_1[7] ? data_7_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_205 = addr_dec_1[8] ? data_8_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_206 = addr_dec_1[9] ? data_9_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_207 = addr_dec_1[10] ? data_10_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_208 = addr_dec_1[11] ? data_11_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_209 = addr_dec_1[12] ? data_12_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_210 = addr_dec_1[13] ? data_13_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_211 = addr_dec_1[14] ? data_14_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_212 = addr_dec_1[15] ? data_15_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_213 = addr_dec_1[16] ? data_16_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_214 = addr_dec_1[17] ? data_17_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_215 = addr_dec_1[18] ? data_18_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_216 = addr_dec_1[19] ? data_19_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_217 = addr_dec_1[20] ? data_20_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_218 = addr_dec_1[21] ? data_21_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_219 = addr_dec_1[22] ? data_22_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_220 = addr_dec_1[23] ? data_23_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_221 = addr_dec_1[24] ? data_24_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_222 = addr_dec_1[25] ? data_25_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_223 = addr_dec_1[26] ? data_26_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_224 = addr_dec_1[27] ? data_27_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_225 = addr_dec_1[28] ? data_28_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_226 = addr_dec_1[29] ? data_29_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_227 = addr_dec_1[30] ? data_30_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_228 = addr_dec_1[31] ? data_31_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_229 = addr_dec_1[32] ? data_32_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_230 = addr_dec_1[33] ? data_33_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_231 = addr_dec_1[34] ? data_34_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_232 = addr_dec_1[35] ? data_35_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_233 = addr_dec_1[36] ? data_36_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_234 = addr_dec_1[37] ? data_37_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_235 = addr_dec_1[38] ? data_38_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_236 = addr_dec_1[39] ? data_39_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_237 = addr_dec_1[40] ? data_40_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_238 = addr_dec_1[41] ? data_41_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_239 = addr_dec_1[42] ? data_42_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_240 = addr_dec_1[43] ? data_43_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_241 = addr_dec_1[44] ? data_44_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_242 = addr_dec_1[45] ? data_45_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_243 = addr_dec_1[46] ? data_46_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_244 = addr_dec_1[47] ? data_47_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_245 = addr_dec_1[48] ? data_48_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_246 = addr_dec_1[49] ? data_49_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_247 = addr_dec_1[50] ? data_50_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_248 = addr_dec_1[51] ? data_51_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_249 = addr_dec_1[52] ? data_52_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_250 = addr_dec_1[53] ? data_53_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_251 = addr_dec_1[54] ? data_54_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_252 = addr_dec_1[55] ? data_55_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_253 = addr_dec_1[56] ? data_56_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_254 = addr_dec_1[57] ? data_57_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_255 = addr_dec_1[58] ? data_58_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_256 = addr_dec_1[59] ? data_59_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_257 = addr_dec_1[60] ? data_60_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_258 = addr_dec_1[61] ? data_61_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_259 = addr_dec_1[62] ? data_62_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_260 = addr_dec_1[63] ? data_63_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_261 = _io_rdata_1_T_197 | _io_rdata_1_T_198; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_262 = _io_rdata_1_T_261 | _io_rdata_1_T_199; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_263 = _io_rdata_1_T_262 | _io_rdata_1_T_200; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_264 = _io_rdata_1_T_263 | _io_rdata_1_T_201; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_265 = _io_rdata_1_T_264 | _io_rdata_1_T_202; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_266 = _io_rdata_1_T_265 | _io_rdata_1_T_203; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_267 = _io_rdata_1_T_266 | _io_rdata_1_T_204; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_268 = _io_rdata_1_T_267 | _io_rdata_1_T_205; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_269 = _io_rdata_1_T_268 | _io_rdata_1_T_206; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_270 = _io_rdata_1_T_269 | _io_rdata_1_T_207; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_271 = _io_rdata_1_T_270 | _io_rdata_1_T_208; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_272 = _io_rdata_1_T_271 | _io_rdata_1_T_209; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_273 = _io_rdata_1_T_272 | _io_rdata_1_T_210; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_274 = _io_rdata_1_T_273 | _io_rdata_1_T_211; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_275 = _io_rdata_1_T_274 | _io_rdata_1_T_212; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_276 = _io_rdata_1_T_275 | _io_rdata_1_T_213; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_277 = _io_rdata_1_T_276 | _io_rdata_1_T_214; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_278 = _io_rdata_1_T_277 | _io_rdata_1_T_215; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_279 = _io_rdata_1_T_278 | _io_rdata_1_T_216; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_280 = _io_rdata_1_T_279 | _io_rdata_1_T_217; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_281 = _io_rdata_1_T_280 | _io_rdata_1_T_218; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_282 = _io_rdata_1_T_281 | _io_rdata_1_T_219; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_283 = _io_rdata_1_T_282 | _io_rdata_1_T_220; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_284 = _io_rdata_1_T_283 | _io_rdata_1_T_221; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_285 = _io_rdata_1_T_284 | _io_rdata_1_T_222; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_286 = _io_rdata_1_T_285 | _io_rdata_1_T_223; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_287 = _io_rdata_1_T_286 | _io_rdata_1_T_224; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_288 = _io_rdata_1_T_287 | _io_rdata_1_T_225; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_289 = _io_rdata_1_T_288 | _io_rdata_1_T_226; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_290 = _io_rdata_1_T_289 | _io_rdata_1_T_227; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_291 = _io_rdata_1_T_290 | _io_rdata_1_T_228; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_292 = _io_rdata_1_T_291 | _io_rdata_1_T_229; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_293 = _io_rdata_1_T_292 | _io_rdata_1_T_230; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_294 = _io_rdata_1_T_293 | _io_rdata_1_T_231; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_295 = _io_rdata_1_T_294 | _io_rdata_1_T_232; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_296 = _io_rdata_1_T_295 | _io_rdata_1_T_233; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_297 = _io_rdata_1_T_296 | _io_rdata_1_T_234; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_298 = _io_rdata_1_T_297 | _io_rdata_1_T_235; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_299 = _io_rdata_1_T_298 | _io_rdata_1_T_236; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_300 = _io_rdata_1_T_299 | _io_rdata_1_T_237; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_301 = _io_rdata_1_T_300 | _io_rdata_1_T_238; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_302 = _io_rdata_1_T_301 | _io_rdata_1_T_239; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_303 = _io_rdata_1_T_302 | _io_rdata_1_T_240; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_304 = _io_rdata_1_T_303 | _io_rdata_1_T_241; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_305 = _io_rdata_1_T_304 | _io_rdata_1_T_242; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_306 = _io_rdata_1_T_305 | _io_rdata_1_T_243; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_307 = _io_rdata_1_T_306 | _io_rdata_1_T_244; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_308 = _io_rdata_1_T_307 | _io_rdata_1_T_245; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_309 = _io_rdata_1_T_308 | _io_rdata_1_T_246; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_310 = _io_rdata_1_T_309 | _io_rdata_1_T_247; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_311 = _io_rdata_1_T_310 | _io_rdata_1_T_248; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_312 = _io_rdata_1_T_311 | _io_rdata_1_T_249; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_313 = _io_rdata_1_T_312 | _io_rdata_1_T_250; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_314 = _io_rdata_1_T_313 | _io_rdata_1_T_251; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_315 = _io_rdata_1_T_314 | _io_rdata_1_T_252; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_316 = _io_rdata_1_T_315 | _io_rdata_1_T_253; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_317 = _io_rdata_1_T_316 | _io_rdata_1_T_254; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_318 = _io_rdata_1_T_317 | _io_rdata_1_T_255; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_319 = _io_rdata_1_T_318 | _io_rdata_1_T_256; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_320 = _io_rdata_1_T_319 | _io_rdata_1_T_257; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_321 = _io_rdata_1_T_320 | _io_rdata_1_T_258; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_322 = _io_rdata_1_T_321 | _io_rdata_1_T_259; // @[Mux.scala 27:73]
  wire [4:0] _io_rdata_1_T_323 = _io_rdata_1_T_322 | _io_rdata_1_T_260; // @[Mux.scala 27:73]
  wire [63:0] waddr_dec_0 = 64'h1 << io_waddr_0; // @[OneHot.scala 57:35]
  wire [63:0] waddr_dec_1 = 64'h1 << io_waddr_1; // @[OneHot.scala 57:35]
  wire  write_wen_0 = io_wen_0 & waddr_dec_0[0]; // @[DataModuleTemplate.scala 188:57]
  wire  write_wen_1 = io_wen_1 & waddr_dec_1[0]; // @[DataModuleTemplate.scala 188:57]
  wire [1:0] _T_4 = {write_wen_1,write_wen_0}; // @[DataModuleTemplate.scala 189:30]
  wire  _data_0_T = write_wen_0 & io_wdata_0_strict; // @[Mux.scala 27:73]
  wire [4:0] _data_0_T_3 = write_wen_0 ? io_wdata_0_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_0_T_4 = write_wen_1 ? io_wdata_1_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_0_T_5 = _data_0_T_3 | _data_0_T_4; // @[Mux.scala 27:73]
  wire  write_wen_0_1 = io_wen_0 & waddr_dec_0[1]; // @[DataModuleTemplate.scala 188:57]
  wire  write_wen_1_1 = io_wen_1 & waddr_dec_1[1]; // @[DataModuleTemplate.scala 188:57]
  wire [1:0] _T_6 = {write_wen_1_1,write_wen_0_1}; // @[DataModuleTemplate.scala 189:30]
  wire  _data_1_T = write_wen_0_1 & io_wdata_0_strict; // @[Mux.scala 27:73]
  wire [4:0] _data_1_T_3 = write_wen_0_1 ? io_wdata_0_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_1_T_4 = write_wen_1_1 ? io_wdata_1_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_1_T_5 = _data_1_T_3 | _data_1_T_4; // @[Mux.scala 27:73]
  wire  write_wen_0_2 = io_wen_0 & waddr_dec_0[2]; // @[DataModuleTemplate.scala 188:57]
  wire  write_wen_1_2 = io_wen_1 & waddr_dec_1[2]; // @[DataModuleTemplate.scala 188:57]
  wire [1:0] _T_8 = {write_wen_1_2,write_wen_0_2}; // @[DataModuleTemplate.scala 189:30]
  wire  _data_2_T = write_wen_0_2 & io_wdata_0_strict; // @[Mux.scala 27:73]
  wire [4:0] _data_2_T_3 = write_wen_0_2 ? io_wdata_0_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_2_T_4 = write_wen_1_2 ? io_wdata_1_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_2_T_5 = _data_2_T_3 | _data_2_T_4; // @[Mux.scala 27:73]
  wire  write_wen_0_3 = io_wen_0 & waddr_dec_0[3]; // @[DataModuleTemplate.scala 188:57]
  wire  write_wen_1_3 = io_wen_1 & waddr_dec_1[3]; // @[DataModuleTemplate.scala 188:57]
  wire [1:0] _T_10 = {write_wen_1_3,write_wen_0_3}; // @[DataModuleTemplate.scala 189:30]
  wire  _data_3_T = write_wen_0_3 & io_wdata_0_strict; // @[Mux.scala 27:73]
  wire [4:0] _data_3_T_3 = write_wen_0_3 ? io_wdata_0_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_3_T_4 = write_wen_1_3 ? io_wdata_1_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_3_T_5 = _data_3_T_3 | _data_3_T_4; // @[Mux.scala 27:73]
  wire  write_wen_0_4 = io_wen_0 & waddr_dec_0[4]; // @[DataModuleTemplate.scala 188:57]
  wire  write_wen_1_4 = io_wen_1 & waddr_dec_1[4]; // @[DataModuleTemplate.scala 188:57]
  wire [1:0] _T_12 = {write_wen_1_4,write_wen_0_4}; // @[DataModuleTemplate.scala 189:30]
  wire  _data_4_T = write_wen_0_4 & io_wdata_0_strict; // @[Mux.scala 27:73]
  wire [4:0] _data_4_T_3 = write_wen_0_4 ? io_wdata_0_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_4_T_4 = write_wen_1_4 ? io_wdata_1_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_4_T_5 = _data_4_T_3 | _data_4_T_4; // @[Mux.scala 27:73]
  wire  write_wen_0_5 = io_wen_0 & waddr_dec_0[5]; // @[DataModuleTemplate.scala 188:57]
  wire  write_wen_1_5 = io_wen_1 & waddr_dec_1[5]; // @[DataModuleTemplate.scala 188:57]
  wire [1:0] _T_14 = {write_wen_1_5,write_wen_0_5}; // @[DataModuleTemplate.scala 189:30]
  wire  _data_5_T = write_wen_0_5 & io_wdata_0_strict; // @[Mux.scala 27:73]
  wire [4:0] _data_5_T_3 = write_wen_0_5 ? io_wdata_0_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_5_T_4 = write_wen_1_5 ? io_wdata_1_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_5_T_5 = _data_5_T_3 | _data_5_T_4; // @[Mux.scala 27:73]
  wire  write_wen_0_6 = io_wen_0 & waddr_dec_0[6]; // @[DataModuleTemplate.scala 188:57]
  wire  write_wen_1_6 = io_wen_1 & waddr_dec_1[6]; // @[DataModuleTemplate.scala 188:57]
  wire [1:0] _T_16 = {write_wen_1_6,write_wen_0_6}; // @[DataModuleTemplate.scala 189:30]
  wire  _data_6_T = write_wen_0_6 & io_wdata_0_strict; // @[Mux.scala 27:73]
  wire [4:0] _data_6_T_3 = write_wen_0_6 ? io_wdata_0_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_6_T_4 = write_wen_1_6 ? io_wdata_1_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_6_T_5 = _data_6_T_3 | _data_6_T_4; // @[Mux.scala 27:73]
  wire  write_wen_0_7 = io_wen_0 & waddr_dec_0[7]; // @[DataModuleTemplate.scala 188:57]
  wire  write_wen_1_7 = io_wen_1 & waddr_dec_1[7]; // @[DataModuleTemplate.scala 188:57]
  wire [1:0] _T_18 = {write_wen_1_7,write_wen_0_7}; // @[DataModuleTemplate.scala 189:30]
  wire  _data_7_T = write_wen_0_7 & io_wdata_0_strict; // @[Mux.scala 27:73]
  wire [4:0] _data_7_T_3 = write_wen_0_7 ? io_wdata_0_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_7_T_4 = write_wen_1_7 ? io_wdata_1_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_7_T_5 = _data_7_T_3 | _data_7_T_4; // @[Mux.scala 27:73]
  wire  write_wen_0_8 = io_wen_0 & waddr_dec_0[8]; // @[DataModuleTemplate.scala 188:57]
  wire  write_wen_1_8 = io_wen_1 & waddr_dec_1[8]; // @[DataModuleTemplate.scala 188:57]
  wire [1:0] _T_20 = {write_wen_1_8,write_wen_0_8}; // @[DataModuleTemplate.scala 189:30]
  wire  _data_8_T = write_wen_0_8 & io_wdata_0_strict; // @[Mux.scala 27:73]
  wire [4:0] _data_8_T_3 = write_wen_0_8 ? io_wdata_0_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_8_T_4 = write_wen_1_8 ? io_wdata_1_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_8_T_5 = _data_8_T_3 | _data_8_T_4; // @[Mux.scala 27:73]
  wire  write_wen_0_9 = io_wen_0 & waddr_dec_0[9]; // @[DataModuleTemplate.scala 188:57]
  wire  write_wen_1_9 = io_wen_1 & waddr_dec_1[9]; // @[DataModuleTemplate.scala 188:57]
  wire [1:0] _T_22 = {write_wen_1_9,write_wen_0_9}; // @[DataModuleTemplate.scala 189:30]
  wire  _data_9_T = write_wen_0_9 & io_wdata_0_strict; // @[Mux.scala 27:73]
  wire [4:0] _data_9_T_3 = write_wen_0_9 ? io_wdata_0_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_9_T_4 = write_wen_1_9 ? io_wdata_1_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_9_T_5 = _data_9_T_3 | _data_9_T_4; // @[Mux.scala 27:73]
  wire  write_wen_0_10 = io_wen_0 & waddr_dec_0[10]; // @[DataModuleTemplate.scala 188:57]
  wire  write_wen_1_10 = io_wen_1 & waddr_dec_1[10]; // @[DataModuleTemplate.scala 188:57]
  wire [1:0] _T_24 = {write_wen_1_10,write_wen_0_10}; // @[DataModuleTemplate.scala 189:30]
  wire  _data_10_T = write_wen_0_10 & io_wdata_0_strict; // @[Mux.scala 27:73]
  wire [4:0] _data_10_T_3 = write_wen_0_10 ? io_wdata_0_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_10_T_4 = write_wen_1_10 ? io_wdata_1_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_10_T_5 = _data_10_T_3 | _data_10_T_4; // @[Mux.scala 27:73]
  wire  write_wen_0_11 = io_wen_0 & waddr_dec_0[11]; // @[DataModuleTemplate.scala 188:57]
  wire  write_wen_1_11 = io_wen_1 & waddr_dec_1[11]; // @[DataModuleTemplate.scala 188:57]
  wire [1:0] _T_26 = {write_wen_1_11,write_wen_0_11}; // @[DataModuleTemplate.scala 189:30]
  wire  _data_11_T = write_wen_0_11 & io_wdata_0_strict; // @[Mux.scala 27:73]
  wire [4:0] _data_11_T_3 = write_wen_0_11 ? io_wdata_0_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_11_T_4 = write_wen_1_11 ? io_wdata_1_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_11_T_5 = _data_11_T_3 | _data_11_T_4; // @[Mux.scala 27:73]
  wire  write_wen_0_12 = io_wen_0 & waddr_dec_0[12]; // @[DataModuleTemplate.scala 188:57]
  wire  write_wen_1_12 = io_wen_1 & waddr_dec_1[12]; // @[DataModuleTemplate.scala 188:57]
  wire [1:0] _T_28 = {write_wen_1_12,write_wen_0_12}; // @[DataModuleTemplate.scala 189:30]
  wire  _data_12_T = write_wen_0_12 & io_wdata_0_strict; // @[Mux.scala 27:73]
  wire [4:0] _data_12_T_3 = write_wen_0_12 ? io_wdata_0_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_12_T_4 = write_wen_1_12 ? io_wdata_1_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_12_T_5 = _data_12_T_3 | _data_12_T_4; // @[Mux.scala 27:73]
  wire  write_wen_0_13 = io_wen_0 & waddr_dec_0[13]; // @[DataModuleTemplate.scala 188:57]
  wire  write_wen_1_13 = io_wen_1 & waddr_dec_1[13]; // @[DataModuleTemplate.scala 188:57]
  wire [1:0] _T_30 = {write_wen_1_13,write_wen_0_13}; // @[DataModuleTemplate.scala 189:30]
  wire  _data_13_T = write_wen_0_13 & io_wdata_0_strict; // @[Mux.scala 27:73]
  wire [4:0] _data_13_T_3 = write_wen_0_13 ? io_wdata_0_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_13_T_4 = write_wen_1_13 ? io_wdata_1_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_13_T_5 = _data_13_T_3 | _data_13_T_4; // @[Mux.scala 27:73]
  wire  write_wen_0_14 = io_wen_0 & waddr_dec_0[14]; // @[DataModuleTemplate.scala 188:57]
  wire  write_wen_1_14 = io_wen_1 & waddr_dec_1[14]; // @[DataModuleTemplate.scala 188:57]
  wire [1:0] _T_32 = {write_wen_1_14,write_wen_0_14}; // @[DataModuleTemplate.scala 189:30]
  wire  _data_14_T = write_wen_0_14 & io_wdata_0_strict; // @[Mux.scala 27:73]
  wire [4:0] _data_14_T_3 = write_wen_0_14 ? io_wdata_0_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_14_T_4 = write_wen_1_14 ? io_wdata_1_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_14_T_5 = _data_14_T_3 | _data_14_T_4; // @[Mux.scala 27:73]
  wire  write_wen_0_15 = io_wen_0 & waddr_dec_0[15]; // @[DataModuleTemplate.scala 188:57]
  wire  write_wen_1_15 = io_wen_1 & waddr_dec_1[15]; // @[DataModuleTemplate.scala 188:57]
  wire [1:0] _T_34 = {write_wen_1_15,write_wen_0_15}; // @[DataModuleTemplate.scala 189:30]
  wire  _data_15_T = write_wen_0_15 & io_wdata_0_strict; // @[Mux.scala 27:73]
  wire [4:0] _data_15_T_3 = write_wen_0_15 ? io_wdata_0_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_15_T_4 = write_wen_1_15 ? io_wdata_1_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_15_T_5 = _data_15_T_3 | _data_15_T_4; // @[Mux.scala 27:73]
  wire  write_wen_0_16 = io_wen_0 & waddr_dec_0[16]; // @[DataModuleTemplate.scala 188:57]
  wire  write_wen_1_16 = io_wen_1 & waddr_dec_1[16]; // @[DataModuleTemplate.scala 188:57]
  wire [1:0] _T_36 = {write_wen_1_16,write_wen_0_16}; // @[DataModuleTemplate.scala 189:30]
  wire  _data_16_T = write_wen_0_16 & io_wdata_0_strict; // @[Mux.scala 27:73]
  wire [4:0] _data_16_T_3 = write_wen_0_16 ? io_wdata_0_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_16_T_4 = write_wen_1_16 ? io_wdata_1_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_16_T_5 = _data_16_T_3 | _data_16_T_4; // @[Mux.scala 27:73]
  wire  write_wen_0_17 = io_wen_0 & waddr_dec_0[17]; // @[DataModuleTemplate.scala 188:57]
  wire  write_wen_1_17 = io_wen_1 & waddr_dec_1[17]; // @[DataModuleTemplate.scala 188:57]
  wire [1:0] _T_38 = {write_wen_1_17,write_wen_0_17}; // @[DataModuleTemplate.scala 189:30]
  wire  _data_17_T = write_wen_0_17 & io_wdata_0_strict; // @[Mux.scala 27:73]
  wire [4:0] _data_17_T_3 = write_wen_0_17 ? io_wdata_0_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_17_T_4 = write_wen_1_17 ? io_wdata_1_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_17_T_5 = _data_17_T_3 | _data_17_T_4; // @[Mux.scala 27:73]
  wire  write_wen_0_18 = io_wen_0 & waddr_dec_0[18]; // @[DataModuleTemplate.scala 188:57]
  wire  write_wen_1_18 = io_wen_1 & waddr_dec_1[18]; // @[DataModuleTemplate.scala 188:57]
  wire [1:0] _T_40 = {write_wen_1_18,write_wen_0_18}; // @[DataModuleTemplate.scala 189:30]
  wire  _data_18_T = write_wen_0_18 & io_wdata_0_strict; // @[Mux.scala 27:73]
  wire [4:0] _data_18_T_3 = write_wen_0_18 ? io_wdata_0_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_18_T_4 = write_wen_1_18 ? io_wdata_1_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_18_T_5 = _data_18_T_3 | _data_18_T_4; // @[Mux.scala 27:73]
  wire  write_wen_0_19 = io_wen_0 & waddr_dec_0[19]; // @[DataModuleTemplate.scala 188:57]
  wire  write_wen_1_19 = io_wen_1 & waddr_dec_1[19]; // @[DataModuleTemplate.scala 188:57]
  wire [1:0] _T_42 = {write_wen_1_19,write_wen_0_19}; // @[DataModuleTemplate.scala 189:30]
  wire  _data_19_T = write_wen_0_19 & io_wdata_0_strict; // @[Mux.scala 27:73]
  wire [4:0] _data_19_T_3 = write_wen_0_19 ? io_wdata_0_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_19_T_4 = write_wen_1_19 ? io_wdata_1_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_19_T_5 = _data_19_T_3 | _data_19_T_4; // @[Mux.scala 27:73]
  wire  write_wen_0_20 = io_wen_0 & waddr_dec_0[20]; // @[DataModuleTemplate.scala 188:57]
  wire  write_wen_1_20 = io_wen_1 & waddr_dec_1[20]; // @[DataModuleTemplate.scala 188:57]
  wire [1:0] _T_44 = {write_wen_1_20,write_wen_0_20}; // @[DataModuleTemplate.scala 189:30]
  wire  _data_20_T = write_wen_0_20 & io_wdata_0_strict; // @[Mux.scala 27:73]
  wire [4:0] _data_20_T_3 = write_wen_0_20 ? io_wdata_0_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_20_T_4 = write_wen_1_20 ? io_wdata_1_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_20_T_5 = _data_20_T_3 | _data_20_T_4; // @[Mux.scala 27:73]
  wire  write_wen_0_21 = io_wen_0 & waddr_dec_0[21]; // @[DataModuleTemplate.scala 188:57]
  wire  write_wen_1_21 = io_wen_1 & waddr_dec_1[21]; // @[DataModuleTemplate.scala 188:57]
  wire [1:0] _T_46 = {write_wen_1_21,write_wen_0_21}; // @[DataModuleTemplate.scala 189:30]
  wire  _data_21_T = write_wen_0_21 & io_wdata_0_strict; // @[Mux.scala 27:73]
  wire [4:0] _data_21_T_3 = write_wen_0_21 ? io_wdata_0_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_21_T_4 = write_wen_1_21 ? io_wdata_1_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_21_T_5 = _data_21_T_3 | _data_21_T_4; // @[Mux.scala 27:73]
  wire  write_wen_0_22 = io_wen_0 & waddr_dec_0[22]; // @[DataModuleTemplate.scala 188:57]
  wire  write_wen_1_22 = io_wen_1 & waddr_dec_1[22]; // @[DataModuleTemplate.scala 188:57]
  wire [1:0] _T_48 = {write_wen_1_22,write_wen_0_22}; // @[DataModuleTemplate.scala 189:30]
  wire  _data_22_T = write_wen_0_22 & io_wdata_0_strict; // @[Mux.scala 27:73]
  wire [4:0] _data_22_T_3 = write_wen_0_22 ? io_wdata_0_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_22_T_4 = write_wen_1_22 ? io_wdata_1_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_22_T_5 = _data_22_T_3 | _data_22_T_4; // @[Mux.scala 27:73]
  wire  write_wen_0_23 = io_wen_0 & waddr_dec_0[23]; // @[DataModuleTemplate.scala 188:57]
  wire  write_wen_1_23 = io_wen_1 & waddr_dec_1[23]; // @[DataModuleTemplate.scala 188:57]
  wire [1:0] _T_50 = {write_wen_1_23,write_wen_0_23}; // @[DataModuleTemplate.scala 189:30]
  wire  _data_23_T = write_wen_0_23 & io_wdata_0_strict; // @[Mux.scala 27:73]
  wire [4:0] _data_23_T_3 = write_wen_0_23 ? io_wdata_0_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_23_T_4 = write_wen_1_23 ? io_wdata_1_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_23_T_5 = _data_23_T_3 | _data_23_T_4; // @[Mux.scala 27:73]
  wire  write_wen_0_24 = io_wen_0 & waddr_dec_0[24]; // @[DataModuleTemplate.scala 188:57]
  wire  write_wen_1_24 = io_wen_1 & waddr_dec_1[24]; // @[DataModuleTemplate.scala 188:57]
  wire [1:0] _T_52 = {write_wen_1_24,write_wen_0_24}; // @[DataModuleTemplate.scala 189:30]
  wire  _data_24_T = write_wen_0_24 & io_wdata_0_strict; // @[Mux.scala 27:73]
  wire [4:0] _data_24_T_3 = write_wen_0_24 ? io_wdata_0_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_24_T_4 = write_wen_1_24 ? io_wdata_1_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_24_T_5 = _data_24_T_3 | _data_24_T_4; // @[Mux.scala 27:73]
  wire  write_wen_0_25 = io_wen_0 & waddr_dec_0[25]; // @[DataModuleTemplate.scala 188:57]
  wire  write_wen_1_25 = io_wen_1 & waddr_dec_1[25]; // @[DataModuleTemplate.scala 188:57]
  wire [1:0] _T_54 = {write_wen_1_25,write_wen_0_25}; // @[DataModuleTemplate.scala 189:30]
  wire  _data_25_T = write_wen_0_25 & io_wdata_0_strict; // @[Mux.scala 27:73]
  wire [4:0] _data_25_T_3 = write_wen_0_25 ? io_wdata_0_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_25_T_4 = write_wen_1_25 ? io_wdata_1_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_25_T_5 = _data_25_T_3 | _data_25_T_4; // @[Mux.scala 27:73]
  wire  write_wen_0_26 = io_wen_0 & waddr_dec_0[26]; // @[DataModuleTemplate.scala 188:57]
  wire  write_wen_1_26 = io_wen_1 & waddr_dec_1[26]; // @[DataModuleTemplate.scala 188:57]
  wire [1:0] _T_56 = {write_wen_1_26,write_wen_0_26}; // @[DataModuleTemplate.scala 189:30]
  wire  _data_26_T = write_wen_0_26 & io_wdata_0_strict; // @[Mux.scala 27:73]
  wire [4:0] _data_26_T_3 = write_wen_0_26 ? io_wdata_0_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_26_T_4 = write_wen_1_26 ? io_wdata_1_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_26_T_5 = _data_26_T_3 | _data_26_T_4; // @[Mux.scala 27:73]
  wire  write_wen_0_27 = io_wen_0 & waddr_dec_0[27]; // @[DataModuleTemplate.scala 188:57]
  wire  write_wen_1_27 = io_wen_1 & waddr_dec_1[27]; // @[DataModuleTemplate.scala 188:57]
  wire [1:0] _T_58 = {write_wen_1_27,write_wen_0_27}; // @[DataModuleTemplate.scala 189:30]
  wire  _data_27_T = write_wen_0_27 & io_wdata_0_strict; // @[Mux.scala 27:73]
  wire [4:0] _data_27_T_3 = write_wen_0_27 ? io_wdata_0_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_27_T_4 = write_wen_1_27 ? io_wdata_1_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_27_T_5 = _data_27_T_3 | _data_27_T_4; // @[Mux.scala 27:73]
  wire  write_wen_0_28 = io_wen_0 & waddr_dec_0[28]; // @[DataModuleTemplate.scala 188:57]
  wire  write_wen_1_28 = io_wen_1 & waddr_dec_1[28]; // @[DataModuleTemplate.scala 188:57]
  wire [1:0] _T_60 = {write_wen_1_28,write_wen_0_28}; // @[DataModuleTemplate.scala 189:30]
  wire  _data_28_T = write_wen_0_28 & io_wdata_0_strict; // @[Mux.scala 27:73]
  wire [4:0] _data_28_T_3 = write_wen_0_28 ? io_wdata_0_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_28_T_4 = write_wen_1_28 ? io_wdata_1_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_28_T_5 = _data_28_T_3 | _data_28_T_4; // @[Mux.scala 27:73]
  wire  write_wen_0_29 = io_wen_0 & waddr_dec_0[29]; // @[DataModuleTemplate.scala 188:57]
  wire  write_wen_1_29 = io_wen_1 & waddr_dec_1[29]; // @[DataModuleTemplate.scala 188:57]
  wire [1:0] _T_62 = {write_wen_1_29,write_wen_0_29}; // @[DataModuleTemplate.scala 189:30]
  wire  _data_29_T = write_wen_0_29 & io_wdata_0_strict; // @[Mux.scala 27:73]
  wire [4:0] _data_29_T_3 = write_wen_0_29 ? io_wdata_0_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_29_T_4 = write_wen_1_29 ? io_wdata_1_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_29_T_5 = _data_29_T_3 | _data_29_T_4; // @[Mux.scala 27:73]
  wire  write_wen_0_30 = io_wen_0 & waddr_dec_0[30]; // @[DataModuleTemplate.scala 188:57]
  wire  write_wen_1_30 = io_wen_1 & waddr_dec_1[30]; // @[DataModuleTemplate.scala 188:57]
  wire [1:0] _T_64 = {write_wen_1_30,write_wen_0_30}; // @[DataModuleTemplate.scala 189:30]
  wire  _data_30_T = write_wen_0_30 & io_wdata_0_strict; // @[Mux.scala 27:73]
  wire [4:0] _data_30_T_3 = write_wen_0_30 ? io_wdata_0_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_30_T_4 = write_wen_1_30 ? io_wdata_1_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_30_T_5 = _data_30_T_3 | _data_30_T_4; // @[Mux.scala 27:73]
  wire  write_wen_0_31 = io_wen_0 & waddr_dec_0[31]; // @[DataModuleTemplate.scala 188:57]
  wire  write_wen_1_31 = io_wen_1 & waddr_dec_1[31]; // @[DataModuleTemplate.scala 188:57]
  wire [1:0] _T_66 = {write_wen_1_31,write_wen_0_31}; // @[DataModuleTemplate.scala 189:30]
  wire  _data_31_T = write_wen_0_31 & io_wdata_0_strict; // @[Mux.scala 27:73]
  wire [4:0] _data_31_T_3 = write_wen_0_31 ? io_wdata_0_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_31_T_4 = write_wen_1_31 ? io_wdata_1_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_31_T_5 = _data_31_T_3 | _data_31_T_4; // @[Mux.scala 27:73]
  wire  write_wen_0_32 = io_wen_0 & waddr_dec_0[32]; // @[DataModuleTemplate.scala 188:57]
  wire  write_wen_1_32 = io_wen_1 & waddr_dec_1[32]; // @[DataModuleTemplate.scala 188:57]
  wire [1:0] _T_68 = {write_wen_1_32,write_wen_0_32}; // @[DataModuleTemplate.scala 189:30]
  wire  _data_32_T = write_wen_0_32 & io_wdata_0_strict; // @[Mux.scala 27:73]
  wire [4:0] _data_32_T_3 = write_wen_0_32 ? io_wdata_0_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_32_T_4 = write_wen_1_32 ? io_wdata_1_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_32_T_5 = _data_32_T_3 | _data_32_T_4; // @[Mux.scala 27:73]
  wire  write_wen_0_33 = io_wen_0 & waddr_dec_0[33]; // @[DataModuleTemplate.scala 188:57]
  wire  write_wen_1_33 = io_wen_1 & waddr_dec_1[33]; // @[DataModuleTemplate.scala 188:57]
  wire [1:0] _T_70 = {write_wen_1_33,write_wen_0_33}; // @[DataModuleTemplate.scala 189:30]
  wire  _data_33_T = write_wen_0_33 & io_wdata_0_strict; // @[Mux.scala 27:73]
  wire [4:0] _data_33_T_3 = write_wen_0_33 ? io_wdata_0_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_33_T_4 = write_wen_1_33 ? io_wdata_1_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_33_T_5 = _data_33_T_3 | _data_33_T_4; // @[Mux.scala 27:73]
  wire  write_wen_0_34 = io_wen_0 & waddr_dec_0[34]; // @[DataModuleTemplate.scala 188:57]
  wire  write_wen_1_34 = io_wen_1 & waddr_dec_1[34]; // @[DataModuleTemplate.scala 188:57]
  wire [1:0] _T_72 = {write_wen_1_34,write_wen_0_34}; // @[DataModuleTemplate.scala 189:30]
  wire  _data_34_T = write_wen_0_34 & io_wdata_0_strict; // @[Mux.scala 27:73]
  wire [4:0] _data_34_T_3 = write_wen_0_34 ? io_wdata_0_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_34_T_4 = write_wen_1_34 ? io_wdata_1_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_34_T_5 = _data_34_T_3 | _data_34_T_4; // @[Mux.scala 27:73]
  wire  write_wen_0_35 = io_wen_0 & waddr_dec_0[35]; // @[DataModuleTemplate.scala 188:57]
  wire  write_wen_1_35 = io_wen_1 & waddr_dec_1[35]; // @[DataModuleTemplate.scala 188:57]
  wire [1:0] _T_74 = {write_wen_1_35,write_wen_0_35}; // @[DataModuleTemplate.scala 189:30]
  wire  _data_35_T = write_wen_0_35 & io_wdata_0_strict; // @[Mux.scala 27:73]
  wire [4:0] _data_35_T_3 = write_wen_0_35 ? io_wdata_0_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_35_T_4 = write_wen_1_35 ? io_wdata_1_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_35_T_5 = _data_35_T_3 | _data_35_T_4; // @[Mux.scala 27:73]
  wire  write_wen_0_36 = io_wen_0 & waddr_dec_0[36]; // @[DataModuleTemplate.scala 188:57]
  wire  write_wen_1_36 = io_wen_1 & waddr_dec_1[36]; // @[DataModuleTemplate.scala 188:57]
  wire [1:0] _T_76 = {write_wen_1_36,write_wen_0_36}; // @[DataModuleTemplate.scala 189:30]
  wire  _data_36_T = write_wen_0_36 & io_wdata_0_strict; // @[Mux.scala 27:73]
  wire [4:0] _data_36_T_3 = write_wen_0_36 ? io_wdata_0_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_36_T_4 = write_wen_1_36 ? io_wdata_1_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_36_T_5 = _data_36_T_3 | _data_36_T_4; // @[Mux.scala 27:73]
  wire  write_wen_0_37 = io_wen_0 & waddr_dec_0[37]; // @[DataModuleTemplate.scala 188:57]
  wire  write_wen_1_37 = io_wen_1 & waddr_dec_1[37]; // @[DataModuleTemplate.scala 188:57]
  wire [1:0] _T_78 = {write_wen_1_37,write_wen_0_37}; // @[DataModuleTemplate.scala 189:30]
  wire  _data_37_T = write_wen_0_37 & io_wdata_0_strict; // @[Mux.scala 27:73]
  wire [4:0] _data_37_T_3 = write_wen_0_37 ? io_wdata_0_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_37_T_4 = write_wen_1_37 ? io_wdata_1_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_37_T_5 = _data_37_T_3 | _data_37_T_4; // @[Mux.scala 27:73]
  wire  write_wen_0_38 = io_wen_0 & waddr_dec_0[38]; // @[DataModuleTemplate.scala 188:57]
  wire  write_wen_1_38 = io_wen_1 & waddr_dec_1[38]; // @[DataModuleTemplate.scala 188:57]
  wire [1:0] _T_80 = {write_wen_1_38,write_wen_0_38}; // @[DataModuleTemplate.scala 189:30]
  wire  _data_38_T = write_wen_0_38 & io_wdata_0_strict; // @[Mux.scala 27:73]
  wire [4:0] _data_38_T_3 = write_wen_0_38 ? io_wdata_0_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_38_T_4 = write_wen_1_38 ? io_wdata_1_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_38_T_5 = _data_38_T_3 | _data_38_T_4; // @[Mux.scala 27:73]
  wire  write_wen_0_39 = io_wen_0 & waddr_dec_0[39]; // @[DataModuleTemplate.scala 188:57]
  wire  write_wen_1_39 = io_wen_1 & waddr_dec_1[39]; // @[DataModuleTemplate.scala 188:57]
  wire [1:0] _T_82 = {write_wen_1_39,write_wen_0_39}; // @[DataModuleTemplate.scala 189:30]
  wire  _data_39_T = write_wen_0_39 & io_wdata_0_strict; // @[Mux.scala 27:73]
  wire [4:0] _data_39_T_3 = write_wen_0_39 ? io_wdata_0_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_39_T_4 = write_wen_1_39 ? io_wdata_1_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_39_T_5 = _data_39_T_3 | _data_39_T_4; // @[Mux.scala 27:73]
  wire  write_wen_0_40 = io_wen_0 & waddr_dec_0[40]; // @[DataModuleTemplate.scala 188:57]
  wire  write_wen_1_40 = io_wen_1 & waddr_dec_1[40]; // @[DataModuleTemplate.scala 188:57]
  wire [1:0] _T_84 = {write_wen_1_40,write_wen_0_40}; // @[DataModuleTemplate.scala 189:30]
  wire  _data_40_T = write_wen_0_40 & io_wdata_0_strict; // @[Mux.scala 27:73]
  wire [4:0] _data_40_T_3 = write_wen_0_40 ? io_wdata_0_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_40_T_4 = write_wen_1_40 ? io_wdata_1_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_40_T_5 = _data_40_T_3 | _data_40_T_4; // @[Mux.scala 27:73]
  wire  write_wen_0_41 = io_wen_0 & waddr_dec_0[41]; // @[DataModuleTemplate.scala 188:57]
  wire  write_wen_1_41 = io_wen_1 & waddr_dec_1[41]; // @[DataModuleTemplate.scala 188:57]
  wire [1:0] _T_86 = {write_wen_1_41,write_wen_0_41}; // @[DataModuleTemplate.scala 189:30]
  wire  _data_41_T = write_wen_0_41 & io_wdata_0_strict; // @[Mux.scala 27:73]
  wire [4:0] _data_41_T_3 = write_wen_0_41 ? io_wdata_0_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_41_T_4 = write_wen_1_41 ? io_wdata_1_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_41_T_5 = _data_41_T_3 | _data_41_T_4; // @[Mux.scala 27:73]
  wire  write_wen_0_42 = io_wen_0 & waddr_dec_0[42]; // @[DataModuleTemplate.scala 188:57]
  wire  write_wen_1_42 = io_wen_1 & waddr_dec_1[42]; // @[DataModuleTemplate.scala 188:57]
  wire [1:0] _T_88 = {write_wen_1_42,write_wen_0_42}; // @[DataModuleTemplate.scala 189:30]
  wire  _data_42_T = write_wen_0_42 & io_wdata_0_strict; // @[Mux.scala 27:73]
  wire [4:0] _data_42_T_3 = write_wen_0_42 ? io_wdata_0_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_42_T_4 = write_wen_1_42 ? io_wdata_1_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_42_T_5 = _data_42_T_3 | _data_42_T_4; // @[Mux.scala 27:73]
  wire  write_wen_0_43 = io_wen_0 & waddr_dec_0[43]; // @[DataModuleTemplate.scala 188:57]
  wire  write_wen_1_43 = io_wen_1 & waddr_dec_1[43]; // @[DataModuleTemplate.scala 188:57]
  wire [1:0] _T_90 = {write_wen_1_43,write_wen_0_43}; // @[DataModuleTemplate.scala 189:30]
  wire  _data_43_T = write_wen_0_43 & io_wdata_0_strict; // @[Mux.scala 27:73]
  wire [4:0] _data_43_T_3 = write_wen_0_43 ? io_wdata_0_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_43_T_4 = write_wen_1_43 ? io_wdata_1_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_43_T_5 = _data_43_T_3 | _data_43_T_4; // @[Mux.scala 27:73]
  wire  write_wen_0_44 = io_wen_0 & waddr_dec_0[44]; // @[DataModuleTemplate.scala 188:57]
  wire  write_wen_1_44 = io_wen_1 & waddr_dec_1[44]; // @[DataModuleTemplate.scala 188:57]
  wire [1:0] _T_92 = {write_wen_1_44,write_wen_0_44}; // @[DataModuleTemplate.scala 189:30]
  wire  _data_44_T = write_wen_0_44 & io_wdata_0_strict; // @[Mux.scala 27:73]
  wire [4:0] _data_44_T_3 = write_wen_0_44 ? io_wdata_0_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_44_T_4 = write_wen_1_44 ? io_wdata_1_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_44_T_5 = _data_44_T_3 | _data_44_T_4; // @[Mux.scala 27:73]
  wire  write_wen_0_45 = io_wen_0 & waddr_dec_0[45]; // @[DataModuleTemplate.scala 188:57]
  wire  write_wen_1_45 = io_wen_1 & waddr_dec_1[45]; // @[DataModuleTemplate.scala 188:57]
  wire [1:0] _T_94 = {write_wen_1_45,write_wen_0_45}; // @[DataModuleTemplate.scala 189:30]
  wire  _data_45_T = write_wen_0_45 & io_wdata_0_strict; // @[Mux.scala 27:73]
  wire [4:0] _data_45_T_3 = write_wen_0_45 ? io_wdata_0_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_45_T_4 = write_wen_1_45 ? io_wdata_1_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_45_T_5 = _data_45_T_3 | _data_45_T_4; // @[Mux.scala 27:73]
  wire  write_wen_0_46 = io_wen_0 & waddr_dec_0[46]; // @[DataModuleTemplate.scala 188:57]
  wire  write_wen_1_46 = io_wen_1 & waddr_dec_1[46]; // @[DataModuleTemplate.scala 188:57]
  wire [1:0] _T_96 = {write_wen_1_46,write_wen_0_46}; // @[DataModuleTemplate.scala 189:30]
  wire  _data_46_T = write_wen_0_46 & io_wdata_0_strict; // @[Mux.scala 27:73]
  wire [4:0] _data_46_T_3 = write_wen_0_46 ? io_wdata_0_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_46_T_4 = write_wen_1_46 ? io_wdata_1_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_46_T_5 = _data_46_T_3 | _data_46_T_4; // @[Mux.scala 27:73]
  wire  write_wen_0_47 = io_wen_0 & waddr_dec_0[47]; // @[DataModuleTemplate.scala 188:57]
  wire  write_wen_1_47 = io_wen_1 & waddr_dec_1[47]; // @[DataModuleTemplate.scala 188:57]
  wire [1:0] _T_98 = {write_wen_1_47,write_wen_0_47}; // @[DataModuleTemplate.scala 189:30]
  wire  _data_47_T = write_wen_0_47 & io_wdata_0_strict; // @[Mux.scala 27:73]
  wire [4:0] _data_47_T_3 = write_wen_0_47 ? io_wdata_0_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_47_T_4 = write_wen_1_47 ? io_wdata_1_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_47_T_5 = _data_47_T_3 | _data_47_T_4; // @[Mux.scala 27:73]
  wire  write_wen_0_48 = io_wen_0 & waddr_dec_0[48]; // @[DataModuleTemplate.scala 188:57]
  wire  write_wen_1_48 = io_wen_1 & waddr_dec_1[48]; // @[DataModuleTemplate.scala 188:57]
  wire [1:0] _T_100 = {write_wen_1_48,write_wen_0_48}; // @[DataModuleTemplate.scala 189:30]
  wire  _data_48_T = write_wen_0_48 & io_wdata_0_strict; // @[Mux.scala 27:73]
  wire [4:0] _data_48_T_3 = write_wen_0_48 ? io_wdata_0_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_48_T_4 = write_wen_1_48 ? io_wdata_1_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_48_T_5 = _data_48_T_3 | _data_48_T_4; // @[Mux.scala 27:73]
  wire  write_wen_0_49 = io_wen_0 & waddr_dec_0[49]; // @[DataModuleTemplate.scala 188:57]
  wire  write_wen_1_49 = io_wen_1 & waddr_dec_1[49]; // @[DataModuleTemplate.scala 188:57]
  wire [1:0] _T_102 = {write_wen_1_49,write_wen_0_49}; // @[DataModuleTemplate.scala 189:30]
  wire  _data_49_T = write_wen_0_49 & io_wdata_0_strict; // @[Mux.scala 27:73]
  wire [4:0] _data_49_T_3 = write_wen_0_49 ? io_wdata_0_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_49_T_4 = write_wen_1_49 ? io_wdata_1_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_49_T_5 = _data_49_T_3 | _data_49_T_4; // @[Mux.scala 27:73]
  wire  write_wen_0_50 = io_wen_0 & waddr_dec_0[50]; // @[DataModuleTemplate.scala 188:57]
  wire  write_wen_1_50 = io_wen_1 & waddr_dec_1[50]; // @[DataModuleTemplate.scala 188:57]
  wire [1:0] _T_104 = {write_wen_1_50,write_wen_0_50}; // @[DataModuleTemplate.scala 189:30]
  wire  _data_50_T = write_wen_0_50 & io_wdata_0_strict; // @[Mux.scala 27:73]
  wire [4:0] _data_50_T_3 = write_wen_0_50 ? io_wdata_0_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_50_T_4 = write_wen_1_50 ? io_wdata_1_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_50_T_5 = _data_50_T_3 | _data_50_T_4; // @[Mux.scala 27:73]
  wire  write_wen_0_51 = io_wen_0 & waddr_dec_0[51]; // @[DataModuleTemplate.scala 188:57]
  wire  write_wen_1_51 = io_wen_1 & waddr_dec_1[51]; // @[DataModuleTemplate.scala 188:57]
  wire [1:0] _T_106 = {write_wen_1_51,write_wen_0_51}; // @[DataModuleTemplate.scala 189:30]
  wire  _data_51_T = write_wen_0_51 & io_wdata_0_strict; // @[Mux.scala 27:73]
  wire [4:0] _data_51_T_3 = write_wen_0_51 ? io_wdata_0_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_51_T_4 = write_wen_1_51 ? io_wdata_1_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_51_T_5 = _data_51_T_3 | _data_51_T_4; // @[Mux.scala 27:73]
  wire  write_wen_0_52 = io_wen_0 & waddr_dec_0[52]; // @[DataModuleTemplate.scala 188:57]
  wire  write_wen_1_52 = io_wen_1 & waddr_dec_1[52]; // @[DataModuleTemplate.scala 188:57]
  wire [1:0] _T_108 = {write_wen_1_52,write_wen_0_52}; // @[DataModuleTemplate.scala 189:30]
  wire  _data_52_T = write_wen_0_52 & io_wdata_0_strict; // @[Mux.scala 27:73]
  wire [4:0] _data_52_T_3 = write_wen_0_52 ? io_wdata_0_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_52_T_4 = write_wen_1_52 ? io_wdata_1_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_52_T_5 = _data_52_T_3 | _data_52_T_4; // @[Mux.scala 27:73]
  wire  write_wen_0_53 = io_wen_0 & waddr_dec_0[53]; // @[DataModuleTemplate.scala 188:57]
  wire  write_wen_1_53 = io_wen_1 & waddr_dec_1[53]; // @[DataModuleTemplate.scala 188:57]
  wire [1:0] _T_110 = {write_wen_1_53,write_wen_0_53}; // @[DataModuleTemplate.scala 189:30]
  wire  _data_53_T = write_wen_0_53 & io_wdata_0_strict; // @[Mux.scala 27:73]
  wire [4:0] _data_53_T_3 = write_wen_0_53 ? io_wdata_0_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_53_T_4 = write_wen_1_53 ? io_wdata_1_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_53_T_5 = _data_53_T_3 | _data_53_T_4; // @[Mux.scala 27:73]
  wire  write_wen_0_54 = io_wen_0 & waddr_dec_0[54]; // @[DataModuleTemplate.scala 188:57]
  wire  write_wen_1_54 = io_wen_1 & waddr_dec_1[54]; // @[DataModuleTemplate.scala 188:57]
  wire [1:0] _T_112 = {write_wen_1_54,write_wen_0_54}; // @[DataModuleTemplate.scala 189:30]
  wire  _data_54_T = write_wen_0_54 & io_wdata_0_strict; // @[Mux.scala 27:73]
  wire [4:0] _data_54_T_3 = write_wen_0_54 ? io_wdata_0_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_54_T_4 = write_wen_1_54 ? io_wdata_1_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_54_T_5 = _data_54_T_3 | _data_54_T_4; // @[Mux.scala 27:73]
  wire  write_wen_0_55 = io_wen_0 & waddr_dec_0[55]; // @[DataModuleTemplate.scala 188:57]
  wire  write_wen_1_55 = io_wen_1 & waddr_dec_1[55]; // @[DataModuleTemplate.scala 188:57]
  wire [1:0] _T_114 = {write_wen_1_55,write_wen_0_55}; // @[DataModuleTemplate.scala 189:30]
  wire  _data_55_T = write_wen_0_55 & io_wdata_0_strict; // @[Mux.scala 27:73]
  wire [4:0] _data_55_T_3 = write_wen_0_55 ? io_wdata_0_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_55_T_4 = write_wen_1_55 ? io_wdata_1_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_55_T_5 = _data_55_T_3 | _data_55_T_4; // @[Mux.scala 27:73]
  wire  write_wen_0_56 = io_wen_0 & waddr_dec_0[56]; // @[DataModuleTemplate.scala 188:57]
  wire  write_wen_1_56 = io_wen_1 & waddr_dec_1[56]; // @[DataModuleTemplate.scala 188:57]
  wire [1:0] _T_116 = {write_wen_1_56,write_wen_0_56}; // @[DataModuleTemplate.scala 189:30]
  wire  _data_56_T = write_wen_0_56 & io_wdata_0_strict; // @[Mux.scala 27:73]
  wire [4:0] _data_56_T_3 = write_wen_0_56 ? io_wdata_0_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_56_T_4 = write_wen_1_56 ? io_wdata_1_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_56_T_5 = _data_56_T_3 | _data_56_T_4; // @[Mux.scala 27:73]
  wire  write_wen_0_57 = io_wen_0 & waddr_dec_0[57]; // @[DataModuleTemplate.scala 188:57]
  wire  write_wen_1_57 = io_wen_1 & waddr_dec_1[57]; // @[DataModuleTemplate.scala 188:57]
  wire [1:0] _T_118 = {write_wen_1_57,write_wen_0_57}; // @[DataModuleTemplate.scala 189:30]
  wire  _data_57_T = write_wen_0_57 & io_wdata_0_strict; // @[Mux.scala 27:73]
  wire [4:0] _data_57_T_3 = write_wen_0_57 ? io_wdata_0_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_57_T_4 = write_wen_1_57 ? io_wdata_1_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_57_T_5 = _data_57_T_3 | _data_57_T_4; // @[Mux.scala 27:73]
  wire  write_wen_0_58 = io_wen_0 & waddr_dec_0[58]; // @[DataModuleTemplate.scala 188:57]
  wire  write_wen_1_58 = io_wen_1 & waddr_dec_1[58]; // @[DataModuleTemplate.scala 188:57]
  wire [1:0] _T_120 = {write_wen_1_58,write_wen_0_58}; // @[DataModuleTemplate.scala 189:30]
  wire  _data_58_T = write_wen_0_58 & io_wdata_0_strict; // @[Mux.scala 27:73]
  wire [4:0] _data_58_T_3 = write_wen_0_58 ? io_wdata_0_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_58_T_4 = write_wen_1_58 ? io_wdata_1_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_58_T_5 = _data_58_T_3 | _data_58_T_4; // @[Mux.scala 27:73]
  wire  write_wen_0_59 = io_wen_0 & waddr_dec_0[59]; // @[DataModuleTemplate.scala 188:57]
  wire  write_wen_1_59 = io_wen_1 & waddr_dec_1[59]; // @[DataModuleTemplate.scala 188:57]
  wire [1:0] _T_122 = {write_wen_1_59,write_wen_0_59}; // @[DataModuleTemplate.scala 189:30]
  wire  _data_59_T = write_wen_0_59 & io_wdata_0_strict; // @[Mux.scala 27:73]
  wire [4:0] _data_59_T_3 = write_wen_0_59 ? io_wdata_0_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_59_T_4 = write_wen_1_59 ? io_wdata_1_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_59_T_5 = _data_59_T_3 | _data_59_T_4; // @[Mux.scala 27:73]
  wire  write_wen_0_60 = io_wen_0 & waddr_dec_0[60]; // @[DataModuleTemplate.scala 188:57]
  wire  write_wen_1_60 = io_wen_1 & waddr_dec_1[60]; // @[DataModuleTemplate.scala 188:57]
  wire [1:0] _T_124 = {write_wen_1_60,write_wen_0_60}; // @[DataModuleTemplate.scala 189:30]
  wire  _data_60_T = write_wen_0_60 & io_wdata_0_strict; // @[Mux.scala 27:73]
  wire [4:0] _data_60_T_3 = write_wen_0_60 ? io_wdata_0_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_60_T_4 = write_wen_1_60 ? io_wdata_1_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_60_T_5 = _data_60_T_3 | _data_60_T_4; // @[Mux.scala 27:73]
  wire  write_wen_0_61 = io_wen_0 & waddr_dec_0[61]; // @[DataModuleTemplate.scala 188:57]
  wire  write_wen_1_61 = io_wen_1 & waddr_dec_1[61]; // @[DataModuleTemplate.scala 188:57]
  wire [1:0] _T_126 = {write_wen_1_61,write_wen_0_61}; // @[DataModuleTemplate.scala 189:30]
  wire  _data_61_T = write_wen_0_61 & io_wdata_0_strict; // @[Mux.scala 27:73]
  wire [4:0] _data_61_T_3 = write_wen_0_61 ? io_wdata_0_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_61_T_4 = write_wen_1_61 ? io_wdata_1_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_61_T_5 = _data_61_T_3 | _data_61_T_4; // @[Mux.scala 27:73]
  wire  write_wen_0_62 = io_wen_0 & waddr_dec_0[62]; // @[DataModuleTemplate.scala 188:57]
  wire  write_wen_1_62 = io_wen_1 & waddr_dec_1[62]; // @[DataModuleTemplate.scala 188:57]
  wire [1:0] _T_128 = {write_wen_1_62,write_wen_0_62}; // @[DataModuleTemplate.scala 189:30]
  wire  _data_62_T = write_wen_0_62 & io_wdata_0_strict; // @[Mux.scala 27:73]
  wire [4:0] _data_62_T_3 = write_wen_0_62 ? io_wdata_0_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_62_T_4 = write_wen_1_62 ? io_wdata_1_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_62_T_5 = _data_62_T_3 | _data_62_T_4; // @[Mux.scala 27:73]
  wire  write_wen_0_63 = io_wen_0 & waddr_dec_0[63]; // @[DataModuleTemplate.scala 188:57]
  wire  write_wen_1_63 = io_wen_1 & waddr_dec_1[63]; // @[DataModuleTemplate.scala 188:57]
  wire [1:0] _T_130 = {write_wen_1_63,write_wen_0_63}; // @[DataModuleTemplate.scala 189:30]
  wire  _data_63_T = write_wen_0_63 & io_wdata_0_strict; // @[Mux.scala 27:73]
  wire [4:0] _data_63_T_3 = write_wen_0_63 ? io_wdata_0_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_63_T_4 = write_wen_1_63 ? io_wdata_1_ssid : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _data_63_T_5 = _data_63_T_3 | _data_63_T_4; // @[Mux.scala 27:73]
  assign io_rdata_0_ssid = |_T ? _io_rdata_0_T_5 : _io_rdata_0_T_323; // @[DataModuleTemplate.scala 178:40 179:19 181:19]
  assign io_rdata_0_strict = |_T ? _io_rdata_0_T : _io_rdata_0_T_196; // @[DataModuleTemplate.scala 178:40 179:19 181:19]
  assign io_rdata_1_ssid = |_T_2 ? _io_rdata_1_T_5 : _io_rdata_1_T_323; // @[DataModuleTemplate.scala 178:40 179:19 181:19]
  assign io_rdata_1_strict = |_T_2 ? _io_rdata_1_T : _io_rdata_1_T_196; // @[DataModuleTemplate.scala 178:40 179:19 181:19]
  always @(negedge clock) begin
    if (|_T_4) begin // @[DataModuleTemplate.scala 189:42]
      data_0_ssid <= _data_0_T_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_4) begin // @[DataModuleTemplate.scala 189:42]
      data_0_strict <= _data_0_T; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_6) begin // @[DataModuleTemplate.scala 189:42]
      data_1_ssid <= _data_1_T_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_6) begin // @[DataModuleTemplate.scala 189:42]
      data_1_strict <= _data_1_T; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_8) begin // @[DataModuleTemplate.scala 189:42]
      data_2_ssid <= _data_2_T_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_8) begin // @[DataModuleTemplate.scala 189:42]
      data_2_strict <= _data_2_T; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_10) begin // @[DataModuleTemplate.scala 189:42]
      data_3_ssid <= _data_3_T_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_10) begin // @[DataModuleTemplate.scala 189:42]
      data_3_strict <= _data_3_T; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_12) begin // @[DataModuleTemplate.scala 189:42]
      data_4_ssid <= _data_4_T_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_12) begin // @[DataModuleTemplate.scala 189:42]
      data_4_strict <= _data_4_T; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_14) begin // @[DataModuleTemplate.scala 189:42]
      data_5_ssid <= _data_5_T_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_14) begin // @[DataModuleTemplate.scala 189:42]
      data_5_strict <= _data_5_T; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_16) begin // @[DataModuleTemplate.scala 189:42]
      data_6_ssid <= _data_6_T_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_16) begin // @[DataModuleTemplate.scala 189:42]
      data_6_strict <= _data_6_T; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_18) begin // @[DataModuleTemplate.scala 189:42]
      data_7_ssid <= _data_7_T_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_18) begin // @[DataModuleTemplate.scala 189:42]
      data_7_strict <= _data_7_T; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_20) begin // @[DataModuleTemplate.scala 189:42]
      data_8_ssid <= _data_8_T_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_20) begin // @[DataModuleTemplate.scala 189:42]
      data_8_strict <= _data_8_T; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_22) begin // @[DataModuleTemplate.scala 189:42]
      data_9_ssid <= _data_9_T_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_22) begin // @[DataModuleTemplate.scala 189:42]
      data_9_strict <= _data_9_T; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_24) begin // @[DataModuleTemplate.scala 189:42]
      data_10_ssid <= _data_10_T_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_24) begin // @[DataModuleTemplate.scala 189:42]
      data_10_strict <= _data_10_T; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_26) begin // @[DataModuleTemplate.scala 189:42]
      data_11_ssid <= _data_11_T_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_26) begin // @[DataModuleTemplate.scala 189:42]
      data_11_strict <= _data_11_T; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_28) begin // @[DataModuleTemplate.scala 189:42]
      data_12_ssid <= _data_12_T_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_28) begin // @[DataModuleTemplate.scala 189:42]
      data_12_strict <= _data_12_T; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_30) begin // @[DataModuleTemplate.scala 189:42]
      data_13_ssid <= _data_13_T_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_30) begin // @[DataModuleTemplate.scala 189:42]
      data_13_strict <= _data_13_T; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_32) begin // @[DataModuleTemplate.scala 189:42]
      data_14_ssid <= _data_14_T_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_32) begin // @[DataModuleTemplate.scala 189:42]
      data_14_strict <= _data_14_T; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_34) begin // @[DataModuleTemplate.scala 189:42]
      data_15_ssid <= _data_15_T_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_34) begin // @[DataModuleTemplate.scala 189:42]
      data_15_strict <= _data_15_T; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_36) begin // @[DataModuleTemplate.scala 189:42]
      data_16_ssid <= _data_16_T_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_36) begin // @[DataModuleTemplate.scala 189:42]
      data_16_strict <= _data_16_T; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_38) begin // @[DataModuleTemplate.scala 189:42]
      data_17_ssid <= _data_17_T_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_38) begin // @[DataModuleTemplate.scala 189:42]
      data_17_strict <= _data_17_T; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_40) begin // @[DataModuleTemplate.scala 189:42]
      data_18_ssid <= _data_18_T_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_40) begin // @[DataModuleTemplate.scala 189:42]
      data_18_strict <= _data_18_T; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_42) begin // @[DataModuleTemplate.scala 189:42]
      data_19_ssid <= _data_19_T_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_42) begin // @[DataModuleTemplate.scala 189:42]
      data_19_strict <= _data_19_T; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_44) begin // @[DataModuleTemplate.scala 189:42]
      data_20_ssid <= _data_20_T_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_44) begin // @[DataModuleTemplate.scala 189:42]
      data_20_strict <= _data_20_T; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_46) begin // @[DataModuleTemplate.scala 189:42]
      data_21_ssid <= _data_21_T_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_46) begin // @[DataModuleTemplate.scala 189:42]
      data_21_strict <= _data_21_T; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_48) begin // @[DataModuleTemplate.scala 189:42]
      data_22_ssid <= _data_22_T_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_48) begin // @[DataModuleTemplate.scala 189:42]
      data_22_strict <= _data_22_T; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_50) begin // @[DataModuleTemplate.scala 189:42]
      data_23_ssid <= _data_23_T_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_50) begin // @[DataModuleTemplate.scala 189:42]
      data_23_strict <= _data_23_T; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_52) begin // @[DataModuleTemplate.scala 189:42]
      data_24_ssid <= _data_24_T_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_52) begin // @[DataModuleTemplate.scala 189:42]
      data_24_strict <= _data_24_T; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_54) begin // @[DataModuleTemplate.scala 189:42]
      data_25_ssid <= _data_25_T_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_54) begin // @[DataModuleTemplate.scala 189:42]
      data_25_strict <= _data_25_T; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_56) begin // @[DataModuleTemplate.scala 189:42]
      data_26_ssid <= _data_26_T_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_56) begin // @[DataModuleTemplate.scala 189:42]
      data_26_strict <= _data_26_T; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_58) begin // @[DataModuleTemplate.scala 189:42]
      data_27_ssid <= _data_27_T_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_58) begin // @[DataModuleTemplate.scala 189:42]
      data_27_strict <= _data_27_T; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_60) begin // @[DataModuleTemplate.scala 189:42]
      data_28_ssid <= _data_28_T_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_60) begin // @[DataModuleTemplate.scala 189:42]
      data_28_strict <= _data_28_T; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_62) begin // @[DataModuleTemplate.scala 189:42]
      data_29_ssid <= _data_29_T_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_62) begin // @[DataModuleTemplate.scala 189:42]
      data_29_strict <= _data_29_T; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_64) begin // @[DataModuleTemplate.scala 189:42]
      data_30_ssid <= _data_30_T_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_64) begin // @[DataModuleTemplate.scala 189:42]
      data_30_strict <= _data_30_T; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_66) begin // @[DataModuleTemplate.scala 189:42]
      data_31_ssid <= _data_31_T_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_66) begin // @[DataModuleTemplate.scala 189:42]
      data_31_strict <= _data_31_T; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_68) begin // @[DataModuleTemplate.scala 189:42]
      data_32_ssid <= _data_32_T_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_68) begin // @[DataModuleTemplate.scala 189:42]
      data_32_strict <= _data_32_T; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_70) begin // @[DataModuleTemplate.scala 189:42]
      data_33_ssid <= _data_33_T_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_70) begin // @[DataModuleTemplate.scala 189:42]
      data_33_strict <= _data_33_T; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_72) begin // @[DataModuleTemplate.scala 189:42]
      data_34_ssid <= _data_34_T_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_72) begin // @[DataModuleTemplate.scala 189:42]
      data_34_strict <= _data_34_T; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_74) begin // @[DataModuleTemplate.scala 189:42]
      data_35_ssid <= _data_35_T_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_74) begin // @[DataModuleTemplate.scala 189:42]
      data_35_strict <= _data_35_T; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_76) begin // @[DataModuleTemplate.scala 189:42]
      data_36_ssid <= _data_36_T_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_76) begin // @[DataModuleTemplate.scala 189:42]
      data_36_strict <= _data_36_T; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_78) begin // @[DataModuleTemplate.scala 189:42]
      data_37_ssid <= _data_37_T_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_78) begin // @[DataModuleTemplate.scala 189:42]
      data_37_strict <= _data_37_T; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_80) begin // @[DataModuleTemplate.scala 189:42]
      data_38_ssid <= _data_38_T_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_80) begin // @[DataModuleTemplate.scala 189:42]
      data_38_strict <= _data_38_T; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_82) begin // @[DataModuleTemplate.scala 189:42]
      data_39_ssid <= _data_39_T_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_82) begin // @[DataModuleTemplate.scala 189:42]
      data_39_strict <= _data_39_T; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_84) begin // @[DataModuleTemplate.scala 189:42]
      data_40_ssid <= _data_40_T_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_84) begin // @[DataModuleTemplate.scala 189:42]
      data_40_strict <= _data_40_T; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_86) begin // @[DataModuleTemplate.scala 189:42]
      data_41_ssid <= _data_41_T_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_86) begin // @[DataModuleTemplate.scala 189:42]
      data_41_strict <= _data_41_T; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_88) begin // @[DataModuleTemplate.scala 189:42]
      data_42_ssid <= _data_42_T_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_88) begin // @[DataModuleTemplate.scala 189:42]
      data_42_strict <= _data_42_T; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_90) begin // @[DataModuleTemplate.scala 189:42]
      data_43_ssid <= _data_43_T_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_90) begin // @[DataModuleTemplate.scala 189:42]
      data_43_strict <= _data_43_T; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_92) begin // @[DataModuleTemplate.scala 189:42]
      data_44_ssid <= _data_44_T_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_92) begin // @[DataModuleTemplate.scala 189:42]
      data_44_strict <= _data_44_T; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_94) begin // @[DataModuleTemplate.scala 189:42]
      data_45_ssid <= _data_45_T_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_94) begin // @[DataModuleTemplate.scala 189:42]
      data_45_strict <= _data_45_T; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_96) begin // @[DataModuleTemplate.scala 189:42]
      data_46_ssid <= _data_46_T_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_96) begin // @[DataModuleTemplate.scala 189:42]
      data_46_strict <= _data_46_T; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_98) begin // @[DataModuleTemplate.scala 189:42]
      data_47_ssid <= _data_47_T_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_98) begin // @[DataModuleTemplate.scala 189:42]
      data_47_strict <= _data_47_T; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_100) begin // @[DataModuleTemplate.scala 189:42]
      data_48_ssid <= _data_48_T_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_100) begin // @[DataModuleTemplate.scala 189:42]
      data_48_strict <= _data_48_T; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_102) begin // @[DataModuleTemplate.scala 189:42]
      data_49_ssid <= _data_49_T_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_102) begin // @[DataModuleTemplate.scala 189:42]
      data_49_strict <= _data_49_T; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_104) begin // @[DataModuleTemplate.scala 189:42]
      data_50_ssid <= _data_50_T_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_104) begin // @[DataModuleTemplate.scala 189:42]
      data_50_strict <= _data_50_T; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_106) begin // @[DataModuleTemplate.scala 189:42]
      data_51_ssid <= _data_51_T_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_106) begin // @[DataModuleTemplate.scala 189:42]
      data_51_strict <= _data_51_T; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_108) begin // @[DataModuleTemplate.scala 189:42]
      data_52_ssid <= _data_52_T_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_108) begin // @[DataModuleTemplate.scala 189:42]
      data_52_strict <= _data_52_T; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_110) begin // @[DataModuleTemplate.scala 189:42]
      data_53_ssid <= _data_53_T_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_110) begin // @[DataModuleTemplate.scala 189:42]
      data_53_strict <= _data_53_T; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_112) begin // @[DataModuleTemplate.scala 189:42]
      data_54_ssid <= _data_54_T_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_112) begin // @[DataModuleTemplate.scala 189:42]
      data_54_strict <= _data_54_T; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_114) begin // @[DataModuleTemplate.scala 189:42]
      data_55_ssid <= _data_55_T_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_114) begin // @[DataModuleTemplate.scala 189:42]
      data_55_strict <= _data_55_T; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_116) begin // @[DataModuleTemplate.scala 189:42]
      data_56_ssid <= _data_56_T_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_116) begin // @[DataModuleTemplate.scala 189:42]
      data_56_strict <= _data_56_T; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_118) begin // @[DataModuleTemplate.scala 189:42]
      data_57_ssid <= _data_57_T_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_118) begin // @[DataModuleTemplate.scala 189:42]
      data_57_strict <= _data_57_T; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_120) begin // @[DataModuleTemplate.scala 189:42]
      data_58_ssid <= _data_58_T_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_120) begin // @[DataModuleTemplate.scala 189:42]
      data_58_strict <= _data_58_T; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_122) begin // @[DataModuleTemplate.scala 189:42]
      data_59_ssid <= _data_59_T_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_122) begin // @[DataModuleTemplate.scala 189:42]
      data_59_strict <= _data_59_T; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_124) begin // @[DataModuleTemplate.scala 189:42]
      data_60_ssid <= _data_60_T_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_124) begin // @[DataModuleTemplate.scala 189:42]
      data_60_strict <= _data_60_T; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_126) begin // @[DataModuleTemplate.scala 189:42]
      data_61_ssid <= _data_61_T_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_126) begin // @[DataModuleTemplate.scala 189:42]
      data_61_strict <= _data_61_T; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_128) begin // @[DataModuleTemplate.scala 189:42]
      data_62_ssid <= _data_62_T_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_128) begin // @[DataModuleTemplate.scala 189:42]
      data_62_strict <= _data_62_T; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_130) begin // @[DataModuleTemplate.scala 189:42]
      data_63_ssid <= _data_63_T_5; // @[DataModuleTemplate.scala 190:15]
    end
    if (|_T_130) begin // @[DataModuleTemplate.scala 189:42]
      data_63_strict <= _data_63_T; // @[DataModuleTemplate.scala 190:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  data_0_ssid = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  data_0_strict = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  data_1_ssid = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  data_1_strict = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  data_2_ssid = _RAND_4[4:0];
  _RAND_5 = {1{`RANDOM}};
  data_2_strict = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  data_3_ssid = _RAND_6[4:0];
  _RAND_7 = {1{`RANDOM}};
  data_3_strict = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  data_4_ssid = _RAND_8[4:0];
  _RAND_9 = {1{`RANDOM}};
  data_4_strict = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  data_5_ssid = _RAND_10[4:0];
  _RAND_11 = {1{`RANDOM}};
  data_5_strict = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  data_6_ssid = _RAND_12[4:0];
  _RAND_13 = {1{`RANDOM}};
  data_6_strict = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  data_7_ssid = _RAND_14[4:0];
  _RAND_15 = {1{`RANDOM}};
  data_7_strict = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  data_8_ssid = _RAND_16[4:0];
  _RAND_17 = {1{`RANDOM}};
  data_8_strict = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  data_9_ssid = _RAND_18[4:0];
  _RAND_19 = {1{`RANDOM}};
  data_9_strict = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  data_10_ssid = _RAND_20[4:0];
  _RAND_21 = {1{`RANDOM}};
  data_10_strict = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  data_11_ssid = _RAND_22[4:0];
  _RAND_23 = {1{`RANDOM}};
  data_11_strict = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  data_12_ssid = _RAND_24[4:0];
  _RAND_25 = {1{`RANDOM}};
  data_12_strict = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  data_13_ssid = _RAND_26[4:0];
  _RAND_27 = {1{`RANDOM}};
  data_13_strict = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  data_14_ssid = _RAND_28[4:0];
  _RAND_29 = {1{`RANDOM}};
  data_14_strict = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  data_15_ssid = _RAND_30[4:0];
  _RAND_31 = {1{`RANDOM}};
  data_15_strict = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  data_16_ssid = _RAND_32[4:0];
  _RAND_33 = {1{`RANDOM}};
  data_16_strict = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  data_17_ssid = _RAND_34[4:0];
  _RAND_35 = {1{`RANDOM}};
  data_17_strict = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  data_18_ssid = _RAND_36[4:0];
  _RAND_37 = {1{`RANDOM}};
  data_18_strict = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  data_19_ssid = _RAND_38[4:0];
  _RAND_39 = {1{`RANDOM}};
  data_19_strict = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  data_20_ssid = _RAND_40[4:0];
  _RAND_41 = {1{`RANDOM}};
  data_20_strict = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  data_21_ssid = _RAND_42[4:0];
  _RAND_43 = {1{`RANDOM}};
  data_21_strict = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  data_22_ssid = _RAND_44[4:0];
  _RAND_45 = {1{`RANDOM}};
  data_22_strict = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  data_23_ssid = _RAND_46[4:0];
  _RAND_47 = {1{`RANDOM}};
  data_23_strict = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  data_24_ssid = _RAND_48[4:0];
  _RAND_49 = {1{`RANDOM}};
  data_24_strict = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  data_25_ssid = _RAND_50[4:0];
  _RAND_51 = {1{`RANDOM}};
  data_25_strict = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  data_26_ssid = _RAND_52[4:0];
  _RAND_53 = {1{`RANDOM}};
  data_26_strict = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  data_27_ssid = _RAND_54[4:0];
  _RAND_55 = {1{`RANDOM}};
  data_27_strict = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  data_28_ssid = _RAND_56[4:0];
  _RAND_57 = {1{`RANDOM}};
  data_28_strict = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  data_29_ssid = _RAND_58[4:0];
  _RAND_59 = {1{`RANDOM}};
  data_29_strict = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  data_30_ssid = _RAND_60[4:0];
  _RAND_61 = {1{`RANDOM}};
  data_30_strict = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  data_31_ssid = _RAND_62[4:0];
  _RAND_63 = {1{`RANDOM}};
  data_31_strict = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  data_32_ssid = _RAND_64[4:0];
  _RAND_65 = {1{`RANDOM}};
  data_32_strict = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  data_33_ssid = _RAND_66[4:0];
  _RAND_67 = {1{`RANDOM}};
  data_33_strict = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  data_34_ssid = _RAND_68[4:0];
  _RAND_69 = {1{`RANDOM}};
  data_34_strict = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  data_35_ssid = _RAND_70[4:0];
  _RAND_71 = {1{`RANDOM}};
  data_35_strict = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  data_36_ssid = _RAND_72[4:0];
  _RAND_73 = {1{`RANDOM}};
  data_36_strict = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  data_37_ssid = _RAND_74[4:0];
  _RAND_75 = {1{`RANDOM}};
  data_37_strict = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  data_38_ssid = _RAND_76[4:0];
  _RAND_77 = {1{`RANDOM}};
  data_38_strict = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  data_39_ssid = _RAND_78[4:0];
  _RAND_79 = {1{`RANDOM}};
  data_39_strict = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  data_40_ssid = _RAND_80[4:0];
  _RAND_81 = {1{`RANDOM}};
  data_40_strict = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  data_41_ssid = _RAND_82[4:0];
  _RAND_83 = {1{`RANDOM}};
  data_41_strict = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  data_42_ssid = _RAND_84[4:0];
  _RAND_85 = {1{`RANDOM}};
  data_42_strict = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  data_43_ssid = _RAND_86[4:0];
  _RAND_87 = {1{`RANDOM}};
  data_43_strict = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  data_44_ssid = _RAND_88[4:0];
  _RAND_89 = {1{`RANDOM}};
  data_44_strict = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  data_45_ssid = _RAND_90[4:0];
  _RAND_91 = {1{`RANDOM}};
  data_45_strict = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  data_46_ssid = _RAND_92[4:0];
  _RAND_93 = {1{`RANDOM}};
  data_46_strict = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  data_47_ssid = _RAND_94[4:0];
  _RAND_95 = {1{`RANDOM}};
  data_47_strict = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  data_48_ssid = _RAND_96[4:0];
  _RAND_97 = {1{`RANDOM}};
  data_48_strict = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  data_49_ssid = _RAND_98[4:0];
  _RAND_99 = {1{`RANDOM}};
  data_49_strict = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  data_50_ssid = _RAND_100[4:0];
  _RAND_101 = {1{`RANDOM}};
  data_50_strict = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  data_51_ssid = _RAND_102[4:0];
  _RAND_103 = {1{`RANDOM}};
  data_51_strict = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  data_52_ssid = _RAND_104[4:0];
  _RAND_105 = {1{`RANDOM}};
  data_52_strict = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  data_53_ssid = _RAND_106[4:0];
  _RAND_107 = {1{`RANDOM}};
  data_53_strict = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  data_54_ssid = _RAND_108[4:0];
  _RAND_109 = {1{`RANDOM}};
  data_54_strict = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  data_55_ssid = _RAND_110[4:0];
  _RAND_111 = {1{`RANDOM}};
  data_55_strict = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  data_56_ssid = _RAND_112[4:0];
  _RAND_113 = {1{`RANDOM}};
  data_56_strict = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  data_57_ssid = _RAND_114[4:0];
  _RAND_115 = {1{`RANDOM}};
  data_57_strict = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  data_58_ssid = _RAND_116[4:0];
  _RAND_117 = {1{`RANDOM}};
  data_58_strict = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  data_59_ssid = _RAND_118[4:0];
  _RAND_119 = {1{`RANDOM}};
  data_59_strict = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  data_60_ssid = _RAND_120[4:0];
  _RAND_121 = {1{`RANDOM}};
  data_60_strict = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  data_61_ssid = _RAND_122[4:0];
  _RAND_123 = {1{`RANDOM}};
  data_61_strict = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  data_62_ssid = _RAND_124[4:0];
  _RAND_125 = {1{`RANDOM}};
  data_62_strict = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  data_63_ssid = _RAND_126[4:0];
  _RAND_127 = {1{`RANDOM}};
  data_63_strict = _RAND_127[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule

