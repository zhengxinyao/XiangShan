module MaxPeriodFibonacciLFSR(
  input   clock,
  input   reset,
  input   io_increment,
  output  io_out_0,
  output  io_out_1,
  output  io_out_2,
  output  io_out_3,
  output  io_out_4,
  output  io_out_5,
  output  io_out_6,
  output  io_out_7,
  output  io_out_8,
  output  io_out_9,
  output  io_out_10,
  output  io_out_11,
  output  io_out_12,
  output  io_out_13,
  output  io_out_14,
  output  io_out_15
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
`endif // RANDOMIZE_REG_INIT
  reg  state_0; // @[PRNG.scala 55:49]
  reg  state_1; // @[PRNG.scala 55:49]
  reg  state_2; // @[PRNG.scala 55:49]
  reg  state_3; // @[PRNG.scala 55:49]
  reg  state_4; // @[PRNG.scala 55:49]
  reg  state_5; // @[PRNG.scala 55:49]
  reg  state_6; // @[PRNG.scala 55:49]
  reg  state_7; // @[PRNG.scala 55:49]
  reg  state_8; // @[PRNG.scala 55:49]
  reg  state_9; // @[PRNG.scala 55:49]
  reg  state_10; // @[PRNG.scala 55:49]
  reg  state_11; // @[PRNG.scala 55:49]
  reg  state_12; // @[PRNG.scala 55:49]
  reg  state_13; // @[PRNG.scala 55:49]
  reg  state_14; // @[PRNG.scala 55:49]
  reg  state_15; // @[PRNG.scala 55:49]
  wire  _T_2 = state_15 ^ state_13 ^ state_12 ^ state_10; // @[LFSR.scala 15:41]
  assign io_out_0 = state_0; // @[PRNG.scala 78:10]
  assign io_out_1 = state_1; // @[PRNG.scala 78:10]
  assign io_out_2 = state_2; // @[PRNG.scala 78:10]
  assign io_out_3 = state_3; // @[PRNG.scala 78:10]
  assign io_out_4 = state_4; // @[PRNG.scala 78:10]
  assign io_out_5 = state_5; // @[PRNG.scala 78:10]
  assign io_out_6 = state_6; // @[PRNG.scala 78:10]
  assign io_out_7 = state_7; // @[PRNG.scala 78:10]
  assign io_out_8 = state_8; // @[PRNG.scala 78:10]
  assign io_out_9 = state_9; // @[PRNG.scala 78:10]
  assign io_out_10 = state_10; // @[PRNG.scala 78:10]
  assign io_out_11 = state_11; // @[PRNG.scala 78:10]
  assign io_out_12 = state_12; // @[PRNG.scala 78:10]
  assign io_out_13 = state_13; // @[PRNG.scala 78:10]
  assign io_out_14 = state_14; // @[PRNG.scala 78:10]
  assign io_out_15 = state_15; // @[PRNG.scala 78:10]
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PRNG.scala 69:22]
      state_0 <= 1'h1; // @[PRNG.scala 70:11]
    end else if (io_increment) begin // @[PRNG.scala 55:49]
      state_0 <= _T_2;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PRNG.scala 69:22]
      state_1 <= 1'h0; // @[PRNG.scala 70:11]
    end else if (io_increment) begin // @[PRNG.scala 55:49]
      state_1 <= state_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PRNG.scala 69:22]
      state_2 <= 1'h0; // @[PRNG.scala 70:11]
    end else if (io_increment) begin // @[PRNG.scala 55:49]
      state_2 <= state_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PRNG.scala 69:22]
      state_3 <= 1'h0; // @[PRNG.scala 70:11]
    end else if (io_increment) begin // @[PRNG.scala 55:49]
      state_3 <= state_2;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PRNG.scala 69:22]
      state_4 <= 1'h0; // @[PRNG.scala 70:11]
    end else if (io_increment) begin // @[PRNG.scala 55:49]
      state_4 <= state_3;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PRNG.scala 69:22]
      state_5 <= 1'h0; // @[PRNG.scala 70:11]
    end else if (io_increment) begin // @[PRNG.scala 55:49]
      state_5 <= state_4;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PRNG.scala 69:22]
      state_6 <= 1'h0; // @[PRNG.scala 70:11]
    end else if (io_increment) begin // @[PRNG.scala 55:49]
      state_6 <= state_5;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PRNG.scala 69:22]
      state_7 <= 1'h0; // @[PRNG.scala 70:11]
    end else if (io_increment) begin // @[PRNG.scala 55:49]
      state_7 <= state_6;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PRNG.scala 69:22]
      state_8 <= 1'h0; // @[PRNG.scala 70:11]
    end else if (io_increment) begin // @[PRNG.scala 55:49]
      state_8 <= state_7;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PRNG.scala 69:22]
      state_9 <= 1'h0; // @[PRNG.scala 70:11]
    end else if (io_increment) begin // @[PRNG.scala 55:49]
      state_9 <= state_8;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PRNG.scala 69:22]
      state_10 <= 1'h0; // @[PRNG.scala 70:11]
    end else if (io_increment) begin // @[PRNG.scala 55:49]
      state_10 <= state_9;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PRNG.scala 69:22]
      state_11 <= 1'h0; // @[PRNG.scala 70:11]
    end else if (io_increment) begin // @[PRNG.scala 55:49]
      state_11 <= state_10;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PRNG.scala 69:22]
      state_12 <= 1'h0; // @[PRNG.scala 70:11]
    end else if (io_increment) begin // @[PRNG.scala 55:49]
      state_12 <= state_11;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PRNG.scala 69:22]
      state_13 <= 1'h0; // @[PRNG.scala 70:11]
    end else if (io_increment) begin // @[PRNG.scala 55:49]
      state_13 <= state_12;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PRNG.scala 69:22]
      state_14 <= 1'h0; // @[PRNG.scala 70:11]
    end else if (io_increment) begin // @[PRNG.scala 55:49]
      state_14 <= state_13;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PRNG.scala 69:22]
      state_15 <= 1'h0; // @[PRNG.scala 70:11]
    end else if (io_increment) begin // @[PRNG.scala 55:49]
      state_15 <= state_14;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  state_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  state_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  state_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  state_4 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  state_5 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  state_6 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  state_7 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  state_8 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  state_9 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  state_10 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  state_11 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  state_12 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  state_13 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  state_14 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  state_15 = _RAND_15[0:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    state_0 = 1'h1;
  end
  if (reset) begin
    state_1 = 1'h0;
  end
  if (reset) begin
    state_2 = 1'h0;
  end
  if (reset) begin
    state_3 = 1'h0;
  end
  if (reset) begin
    state_4 = 1'h0;
  end
  if (reset) begin
    state_5 = 1'h0;
  end
  if (reset) begin
    state_6 = 1'h0;
  end
  if (reset) begin
    state_7 = 1'h0;
  end
  if (reset) begin
    state_8 = 1'h0;
  end
  if (reset) begin
    state_9 = 1'h0;
  end
  if (reset) begin
    state_10 = 1'h0;
  end
  if (reset) begin
    state_11 = 1'h0;
  end
  if (reset) begin
    state_12 = 1'h0;
  end
  if (reset) begin
    state_13 = 1'h0;
  end
  if (reset) begin
    state_14 = 1'h0;
  end
  if (reset) begin
    state_15 = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule

