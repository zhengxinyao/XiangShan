module LZA(
  input  [63:0] io_b,
  output [63:0] io_f
);
  wire  p_0 = io_b[0]; // @[LZA.scala 18:21]
  wire  k_0 = ~p_0; // @[LZA.scala 19:24]
  wire  p_1 = io_b[1]; // @[LZA.scala 18:21]
  wire  k_1 = ~p_1; // @[LZA.scala 19:24]
  wire  f_1 = p_1 ^ ~k_0; // @[LZA.scala 23:20]
  wire  p_2 = io_b[2]; // @[LZA.scala 18:21]
  wire  k_2 = ~p_2; // @[LZA.scala 19:24]
  wire  f_2 = p_2 ^ ~k_1; // @[LZA.scala 23:20]
  wire  p_3 = io_b[3]; // @[LZA.scala 18:21]
  wire  k_3 = ~p_3; // @[LZA.scala 19:24]
  wire  f_3 = p_3 ^ ~k_2; // @[LZA.scala 23:20]
  wire  p_4 = io_b[4]; // @[LZA.scala 18:21]
  wire  k_4 = ~p_4; // @[LZA.scala 19:24]
  wire  f_4 = p_4 ^ ~k_3; // @[LZA.scala 23:20]
  wire  p_5 = io_b[5]; // @[LZA.scala 18:21]
  wire  k_5 = ~p_5; // @[LZA.scala 19:24]
  wire  f_5 = p_5 ^ ~k_4; // @[LZA.scala 23:20]
  wire  p_6 = io_b[6]; // @[LZA.scala 18:21]
  wire  k_6 = ~p_6; // @[LZA.scala 19:24]
  wire  f_6 = p_6 ^ ~k_5; // @[LZA.scala 23:20]
  wire  p_7 = io_b[7]; // @[LZA.scala 18:21]
  wire  k_7 = ~p_7; // @[LZA.scala 19:24]
  wire  f_7 = p_7 ^ ~k_6; // @[LZA.scala 23:20]
  wire  p_8 = io_b[8]; // @[LZA.scala 18:21]
  wire  k_8 = ~p_8; // @[LZA.scala 19:24]
  wire  f_8 = p_8 ^ ~k_7; // @[LZA.scala 23:20]
  wire  p_9 = io_b[9]; // @[LZA.scala 18:21]
  wire  k_9 = ~p_9; // @[LZA.scala 19:24]
  wire  f_9 = p_9 ^ ~k_8; // @[LZA.scala 23:20]
  wire  p_10 = io_b[10]; // @[LZA.scala 18:21]
  wire  k_10 = ~p_10; // @[LZA.scala 19:24]
  wire  f_10 = p_10 ^ ~k_9; // @[LZA.scala 23:20]
  wire  p_11 = io_b[11]; // @[LZA.scala 18:21]
  wire  k_11 = ~p_11; // @[LZA.scala 19:24]
  wire  f_11 = p_11 ^ ~k_10; // @[LZA.scala 23:20]
  wire  p_12 = io_b[12]; // @[LZA.scala 18:21]
  wire  k_12 = ~p_12; // @[LZA.scala 19:24]
  wire  f_12 = p_12 ^ ~k_11; // @[LZA.scala 23:20]
  wire  p_13 = io_b[13]; // @[LZA.scala 18:21]
  wire  k_13 = ~p_13; // @[LZA.scala 19:24]
  wire  f_13 = p_13 ^ ~k_12; // @[LZA.scala 23:20]
  wire  p_14 = io_b[14]; // @[LZA.scala 18:21]
  wire  k_14 = ~p_14; // @[LZA.scala 19:24]
  wire  f_14 = p_14 ^ ~k_13; // @[LZA.scala 23:20]
  wire  p_15 = io_b[15]; // @[LZA.scala 18:21]
  wire  k_15 = ~p_15; // @[LZA.scala 19:24]
  wire  f_15 = p_15 ^ ~k_14; // @[LZA.scala 23:20]
  wire  p_16 = io_b[16]; // @[LZA.scala 18:21]
  wire  k_16 = ~p_16; // @[LZA.scala 19:24]
  wire  f_16 = p_16 ^ ~k_15; // @[LZA.scala 23:20]
  wire  p_17 = io_b[17]; // @[LZA.scala 18:21]
  wire  k_17 = ~p_17; // @[LZA.scala 19:24]
  wire  f_17 = p_17 ^ ~k_16; // @[LZA.scala 23:20]
  wire  p_18 = io_b[18]; // @[LZA.scala 18:21]
  wire  k_18 = ~p_18; // @[LZA.scala 19:24]
  wire  f_18 = p_18 ^ ~k_17; // @[LZA.scala 23:20]
  wire  p_19 = io_b[19]; // @[LZA.scala 18:21]
  wire  k_19 = ~p_19; // @[LZA.scala 19:24]
  wire  f_19 = p_19 ^ ~k_18; // @[LZA.scala 23:20]
  wire  p_20 = io_b[20]; // @[LZA.scala 18:21]
  wire  k_20 = ~p_20; // @[LZA.scala 19:24]
  wire  f_20 = p_20 ^ ~k_19; // @[LZA.scala 23:20]
  wire  p_21 = io_b[21]; // @[LZA.scala 18:21]
  wire  k_21 = ~p_21; // @[LZA.scala 19:24]
  wire  f_21 = p_21 ^ ~k_20; // @[LZA.scala 23:20]
  wire  p_22 = io_b[22]; // @[LZA.scala 18:21]
  wire  k_22 = ~p_22; // @[LZA.scala 19:24]
  wire  f_22 = p_22 ^ ~k_21; // @[LZA.scala 23:20]
  wire  p_23 = io_b[23]; // @[LZA.scala 18:21]
  wire  k_23 = ~p_23; // @[LZA.scala 19:24]
  wire  f_23 = p_23 ^ ~k_22; // @[LZA.scala 23:20]
  wire  p_24 = io_b[24]; // @[LZA.scala 18:21]
  wire  k_24 = ~p_24; // @[LZA.scala 19:24]
  wire  f_24 = p_24 ^ ~k_23; // @[LZA.scala 23:20]
  wire  p_25 = io_b[25]; // @[LZA.scala 18:21]
  wire  k_25 = ~p_25; // @[LZA.scala 19:24]
  wire  f_25 = p_25 ^ ~k_24; // @[LZA.scala 23:20]
  wire  p_26 = io_b[26]; // @[LZA.scala 18:21]
  wire  k_26 = ~p_26; // @[LZA.scala 19:24]
  wire  f_26 = p_26 ^ ~k_25; // @[LZA.scala 23:20]
  wire  p_27 = io_b[27]; // @[LZA.scala 18:21]
  wire  k_27 = ~p_27; // @[LZA.scala 19:24]
  wire  f_27 = p_27 ^ ~k_26; // @[LZA.scala 23:20]
  wire  p_28 = io_b[28]; // @[LZA.scala 18:21]
  wire  k_28 = ~p_28; // @[LZA.scala 19:24]
  wire  f_28 = p_28 ^ ~k_27; // @[LZA.scala 23:20]
  wire  p_29 = io_b[29]; // @[LZA.scala 18:21]
  wire  k_29 = ~p_29; // @[LZA.scala 19:24]
  wire  f_29 = p_29 ^ ~k_28; // @[LZA.scala 23:20]
  wire  p_30 = io_b[30]; // @[LZA.scala 18:21]
  wire  k_30 = ~p_30; // @[LZA.scala 19:24]
  wire  f_30 = p_30 ^ ~k_29; // @[LZA.scala 23:20]
  wire  p_31 = io_b[31]; // @[LZA.scala 18:21]
  wire  k_31 = ~p_31; // @[LZA.scala 19:24]
  wire  f_31 = p_31 ^ ~k_30; // @[LZA.scala 23:20]
  wire  p_32 = io_b[32]; // @[LZA.scala 18:21]
  wire  k_32 = ~p_32; // @[LZA.scala 19:24]
  wire  f_32 = p_32 ^ ~k_31; // @[LZA.scala 23:20]
  wire  p_33 = io_b[33]; // @[LZA.scala 18:21]
  wire  k_33 = ~p_33; // @[LZA.scala 19:24]
  wire  f_33 = p_33 ^ ~k_32; // @[LZA.scala 23:20]
  wire  p_34 = io_b[34]; // @[LZA.scala 18:21]
  wire  k_34 = ~p_34; // @[LZA.scala 19:24]
  wire  f_34 = p_34 ^ ~k_33; // @[LZA.scala 23:20]
  wire  p_35 = io_b[35]; // @[LZA.scala 18:21]
  wire  k_35 = ~p_35; // @[LZA.scala 19:24]
  wire  f_35 = p_35 ^ ~k_34; // @[LZA.scala 23:20]
  wire  p_36 = io_b[36]; // @[LZA.scala 18:21]
  wire  k_36 = ~p_36; // @[LZA.scala 19:24]
  wire  f_36 = p_36 ^ ~k_35; // @[LZA.scala 23:20]
  wire  p_37 = io_b[37]; // @[LZA.scala 18:21]
  wire  k_37 = ~p_37; // @[LZA.scala 19:24]
  wire  f_37 = p_37 ^ ~k_36; // @[LZA.scala 23:20]
  wire  p_38 = io_b[38]; // @[LZA.scala 18:21]
  wire  k_38 = ~p_38; // @[LZA.scala 19:24]
  wire  f_38 = p_38 ^ ~k_37; // @[LZA.scala 23:20]
  wire  p_39 = io_b[39]; // @[LZA.scala 18:21]
  wire  k_39 = ~p_39; // @[LZA.scala 19:24]
  wire  f_39 = p_39 ^ ~k_38; // @[LZA.scala 23:20]
  wire  p_40 = io_b[40]; // @[LZA.scala 18:21]
  wire  k_40 = ~p_40; // @[LZA.scala 19:24]
  wire  f_40 = p_40 ^ ~k_39; // @[LZA.scala 23:20]
  wire  p_41 = io_b[41]; // @[LZA.scala 18:21]
  wire  k_41 = ~p_41; // @[LZA.scala 19:24]
  wire  f_41 = p_41 ^ ~k_40; // @[LZA.scala 23:20]
  wire  p_42 = io_b[42]; // @[LZA.scala 18:21]
  wire  k_42 = ~p_42; // @[LZA.scala 19:24]
  wire  f_42 = p_42 ^ ~k_41; // @[LZA.scala 23:20]
  wire  p_43 = io_b[43]; // @[LZA.scala 18:21]
  wire  k_43 = ~p_43; // @[LZA.scala 19:24]
  wire  f_43 = p_43 ^ ~k_42; // @[LZA.scala 23:20]
  wire  p_44 = io_b[44]; // @[LZA.scala 18:21]
  wire  k_44 = ~p_44; // @[LZA.scala 19:24]
  wire  f_44 = p_44 ^ ~k_43; // @[LZA.scala 23:20]
  wire  p_45 = io_b[45]; // @[LZA.scala 18:21]
  wire  k_45 = ~p_45; // @[LZA.scala 19:24]
  wire  f_45 = p_45 ^ ~k_44; // @[LZA.scala 23:20]
  wire  p_46 = io_b[46]; // @[LZA.scala 18:21]
  wire  k_46 = ~p_46; // @[LZA.scala 19:24]
  wire  f_46 = p_46 ^ ~k_45; // @[LZA.scala 23:20]
  wire  p_47 = io_b[47]; // @[LZA.scala 18:21]
  wire  k_47 = ~p_47; // @[LZA.scala 19:24]
  wire  f_47 = p_47 ^ ~k_46; // @[LZA.scala 23:20]
  wire  p_48 = io_b[48]; // @[LZA.scala 18:21]
  wire  k_48 = ~p_48; // @[LZA.scala 19:24]
  wire  f_48 = p_48 ^ ~k_47; // @[LZA.scala 23:20]
  wire  p_49 = io_b[49]; // @[LZA.scala 18:21]
  wire  k_49 = ~p_49; // @[LZA.scala 19:24]
  wire  f_49 = p_49 ^ ~k_48; // @[LZA.scala 23:20]
  wire  p_50 = io_b[50]; // @[LZA.scala 18:21]
  wire  k_50 = ~p_50; // @[LZA.scala 19:24]
  wire  f_50 = p_50 ^ ~k_49; // @[LZA.scala 23:20]
  wire  p_51 = io_b[51]; // @[LZA.scala 18:21]
  wire  k_51 = ~p_51; // @[LZA.scala 19:24]
  wire  f_51 = p_51 ^ ~k_50; // @[LZA.scala 23:20]
  wire  p_52 = io_b[52]; // @[LZA.scala 18:21]
  wire  k_52 = ~p_52; // @[LZA.scala 19:24]
  wire  f_52 = p_52 ^ ~k_51; // @[LZA.scala 23:20]
  wire  p_53 = io_b[53]; // @[LZA.scala 18:21]
  wire  k_53 = ~p_53; // @[LZA.scala 19:24]
  wire  f_53 = p_53 ^ ~k_52; // @[LZA.scala 23:20]
  wire  p_54 = io_b[54]; // @[LZA.scala 18:21]
  wire  k_54 = ~p_54; // @[LZA.scala 19:24]
  wire  f_54 = p_54 ^ ~k_53; // @[LZA.scala 23:20]
  wire  p_55 = io_b[55]; // @[LZA.scala 18:21]
  wire  k_55 = ~p_55; // @[LZA.scala 19:24]
  wire  f_55 = p_55 ^ ~k_54; // @[LZA.scala 23:20]
  wire  p_56 = io_b[56]; // @[LZA.scala 18:21]
  wire  k_56 = ~p_56; // @[LZA.scala 19:24]
  wire  f_56 = p_56 ^ ~k_55; // @[LZA.scala 23:20]
  wire  p_57 = io_b[57]; // @[LZA.scala 18:21]
  wire  k_57 = ~p_57; // @[LZA.scala 19:24]
  wire  f_57 = p_57 ^ ~k_56; // @[LZA.scala 23:20]
  wire  p_58 = io_b[58]; // @[LZA.scala 18:21]
  wire  k_58 = ~p_58; // @[LZA.scala 19:24]
  wire  f_58 = p_58 ^ ~k_57; // @[LZA.scala 23:20]
  wire  p_59 = io_b[59]; // @[LZA.scala 18:21]
  wire  k_59 = ~p_59; // @[LZA.scala 19:24]
  wire  f_59 = p_59 ^ ~k_58; // @[LZA.scala 23:20]
  wire  p_60 = io_b[60]; // @[LZA.scala 18:21]
  wire  k_60 = ~p_60; // @[LZA.scala 19:24]
  wire  f_60 = p_60 ^ ~k_59; // @[LZA.scala 23:20]
  wire  p_61 = io_b[61]; // @[LZA.scala 18:21]
  wire  k_61 = ~p_61; // @[LZA.scala 19:24]
  wire  f_61 = p_61 ^ ~k_60; // @[LZA.scala 23:20]
  wire  p_62 = io_b[62]; // @[LZA.scala 18:21]
  wire  k_62 = ~p_62; // @[LZA.scala 19:24]
  wire  f_62 = p_62 ^ ~k_61; // @[LZA.scala 23:20]
  wire  p_63 = io_b[63]; // @[LZA.scala 18:21]
  wire  f_63 = p_63 ^ ~k_62; // @[LZA.scala 23:20]
  wire [7:0] io_f_lo_lo_lo = {f_7,f_6,f_5,f_4,f_3,f_2,f_1,1'h0}; // @[Cat.scala 31:58]
  wire [15:0] io_f_lo_lo = {f_15,f_14,f_13,f_12,f_11,f_10,f_9,f_8,io_f_lo_lo_lo}; // @[Cat.scala 31:58]
  wire [7:0] io_f_lo_hi_lo = {f_23,f_22,f_21,f_20,f_19,f_18,f_17,f_16}; // @[Cat.scala 31:58]
  wire [31:0] io_f_lo = {f_31,f_30,f_29,f_28,f_27,f_26,f_25,f_24,io_f_lo_hi_lo,io_f_lo_lo}; // @[Cat.scala 31:58]
  wire [7:0] io_f_hi_lo_lo = {f_39,f_38,f_37,f_36,f_35,f_34,f_33,f_32}; // @[Cat.scala 31:58]
  wire [15:0] io_f_hi_lo = {f_47,f_46,f_45,f_44,f_43,f_42,f_41,f_40,io_f_hi_lo_lo}; // @[Cat.scala 31:58]
  wire [7:0] io_f_hi_hi_lo = {f_55,f_54,f_53,f_52,f_51,f_50,f_49,f_48}; // @[Cat.scala 31:58]
  wire [31:0] io_f_hi = {f_63,f_62,f_61,f_60,f_59,f_58,f_57,f_56,io_f_hi_hi_lo,io_f_hi_lo}; // @[Cat.scala 31:58]
  assign io_f = {io_f_hi,io_f_lo}; // @[Cat.scala 31:58]
endmodule

