module CSA3_2_3362(
  input  [26:0] io_in_0,
  input  [26:0] io_in_1,
  input  [26:0] io_in_2,
  output [26:0] io_out_0,
  output [26:0] io_out_1
);
  wire  a = io_in_0[0]; // @[FDIV.scala 677:32]
  wire  b = io_in_1[0]; // @[FDIV.scala 677:45]
  wire  cin = io_in_2[0]; // @[FDIV.scala 677:58]
  wire  a_xor_b = a ^ b; // @[FDIV.scala 678:21]
  wire  a_and_b = a & b; // @[FDIV.scala 679:21]
  wire  sum = a_xor_b ^ cin; // @[FDIV.scala 680:23]
  wire  cout = a_and_b | a_xor_b & cin; // @[FDIV.scala 681:24]
  wire [1:0] temp_0 = {cout,sum}; // @[Cat.scala 31:58]
  wire  a_1 = io_in_0[1]; // @[FDIV.scala 677:32]
  wire  b_1 = io_in_1[1]; // @[FDIV.scala 677:45]
  wire  cin_1 = io_in_2[1]; // @[FDIV.scala 677:58]
  wire  a_xor_b1 = a_1 ^ b_1; // @[FDIV.scala 678:21]
  wire  a_and_b1 = a_1 & b_1; // @[FDIV.scala 679:21]
  wire  sum_1 = a_xor_b1 ^ cin_1; // @[FDIV.scala 680:23]
  wire  cout_1 = a_and_b1 | a_xor_b1 & cin_1; // @[FDIV.scala 681:24]
  wire [1:0] temp_1 = {cout_1,sum_1}; // @[Cat.scala 31:58]
  wire  a_2 = io_in_0[2]; // @[FDIV.scala 677:32]
  wire  b_2 = io_in_1[2]; // @[FDIV.scala 677:45]
  wire  cin_2 = io_in_2[2]; // @[FDIV.scala 677:58]
  wire  a_xor_b2 = a_2 ^ b_2; // @[FDIV.scala 678:21]
  wire  a_and_b2 = a_2 & b_2; // @[FDIV.scala 679:21]
  wire  sum_2 = a_xor_b2 ^ cin_2; // @[FDIV.scala 680:23]
  wire  cout_2 = a_and_b2 | a_xor_b2 & cin_2; // @[FDIV.scala 681:24]
  wire [1:0] temp_2 = {cout_2,sum_2}; // @[Cat.scala 31:58]
  wire  a_3 = io_in_0[3]; // @[FDIV.scala 677:32]
  wire  b_3 = io_in_1[3]; // @[FDIV.scala 677:45]
  wire  cin_3 = io_in_2[3]; // @[FDIV.scala 677:58]
  wire  a_xor_b3 = a_3 ^ b_3; // @[FDIV.scala 678:21]
  wire  a_and_b3 = a_3 & b_3; // @[FDIV.scala 679:21]
  wire  sum_3 = a_xor_b3 ^ cin_3; // @[FDIV.scala 680:23]
  wire  cout_3 = a_and_b3 | a_xor_b3 & cin_3; // @[FDIV.scala 681:24]
  wire [1:0] temp_3 = {cout_3,sum_3}; // @[Cat.scala 31:58]
  wire  a_4 = io_in_0[4]; // @[FDIV.scala 677:32]
  wire  b_4 = io_in_1[4]; // @[FDIV.scala 677:45]
  wire  cin_4 = io_in_2[4]; // @[FDIV.scala 677:58]
  wire  a_xor_b4 = a_4 ^ b_4; // @[FDIV.scala 678:21]
  wire  a_and_b4 = a_4 & b_4; // @[FDIV.scala 679:21]
  wire  sum_4 = a_xor_b4 ^ cin_4; // @[FDIV.scala 680:23]
  wire  cout_4 = a_and_b4 | a_xor_b4 & cin_4; // @[FDIV.scala 681:24]
  wire [1:0] temp_4 = {cout_4,sum_4}; // @[Cat.scala 31:58]
  wire  a_5 = io_in_0[5]; // @[FDIV.scala 677:32]
  wire  b_5 = io_in_1[5]; // @[FDIV.scala 677:45]
  wire  cin_5 = io_in_2[5]; // @[FDIV.scala 677:58]
  wire  a_xor_b5 = a_5 ^ b_5; // @[FDIV.scala 678:21]
  wire  a_and_b5 = a_5 & b_5; // @[FDIV.scala 679:21]
  wire  sum_5 = a_xor_b5 ^ cin_5; // @[FDIV.scala 680:23]
  wire  cout_5 = a_and_b5 | a_xor_b5 & cin_5; // @[FDIV.scala 681:24]
  wire [1:0] temp_5 = {cout_5,sum_5}; // @[Cat.scala 31:58]
  wire  a_6 = io_in_0[6]; // @[FDIV.scala 677:32]
  wire  b_6 = io_in_1[6]; // @[FDIV.scala 677:45]
  wire  cin_6 = io_in_2[6]; // @[FDIV.scala 677:58]
  wire  a_xor_b6 = a_6 ^ b_6; // @[FDIV.scala 678:21]
  wire  a_and_b6 = a_6 & b_6; // @[FDIV.scala 679:21]
  wire  sum_6 = a_xor_b6 ^ cin_6; // @[FDIV.scala 680:23]
  wire  cout_6 = a_and_b6 | a_xor_b6 & cin_6; // @[FDIV.scala 681:24]
  wire [1:0] temp_6 = {cout_6,sum_6}; // @[Cat.scala 31:58]
  wire  a_7 = io_in_0[7]; // @[FDIV.scala 677:32]
  wire  b_7 = io_in_1[7]; // @[FDIV.scala 677:45]
  wire  cin_7 = io_in_2[7]; // @[FDIV.scala 677:58]
  wire  a_xor_b7 = a_7 ^ b_7; // @[FDIV.scala 678:21]
  wire  a_and_b7 = a_7 & b_7; // @[FDIV.scala 679:21]
  wire  sum_7 = a_xor_b7 ^ cin_7; // @[FDIV.scala 680:23]
  wire  cout_7 = a_and_b7 | a_xor_b7 & cin_7; // @[FDIV.scala 681:24]
  wire [1:0] temp_7 = {cout_7,sum_7}; // @[Cat.scala 31:58]
  wire  a_8 = io_in_0[8]; // @[FDIV.scala 677:32]
  wire  b_8 = io_in_1[8]; // @[FDIV.scala 677:45]
  wire  cin_8 = io_in_2[8]; // @[FDIV.scala 677:58]
  wire  a_xor_b8 = a_8 ^ b_8; // @[FDIV.scala 678:21]
  wire  a_and_b8 = a_8 & b_8; // @[FDIV.scala 679:21]
  wire  sum_8 = a_xor_b8 ^ cin_8; // @[FDIV.scala 680:23]
  wire  cout_8 = a_and_b8 | a_xor_b8 & cin_8; // @[FDIV.scala 681:24]
  wire [1:0] temp_8 = {cout_8,sum_8}; // @[Cat.scala 31:58]
  wire  a_9 = io_in_0[9]; // @[FDIV.scala 677:32]
  wire  b_9 = io_in_1[9]; // @[FDIV.scala 677:45]
  wire  cin_9 = io_in_2[9]; // @[FDIV.scala 677:58]
  wire  a_xor_b9 = a_9 ^ b_9; // @[FDIV.scala 678:21]
  wire  a_and_b9 = a_9 & b_9; // @[FDIV.scala 679:21]
  wire  sum_9 = a_xor_b9 ^ cin_9; // @[FDIV.scala 680:23]
  wire  cout_9 = a_and_b9 | a_xor_b9 & cin_9; // @[FDIV.scala 681:24]
  wire [1:0] temp_9 = {cout_9,sum_9}; // @[Cat.scala 31:58]
  wire  a_10 = io_in_0[10]; // @[FDIV.scala 677:32]
  wire  b_10 = io_in_1[10]; // @[FDIV.scala 677:45]
  wire  cin_10 = io_in_2[10]; // @[FDIV.scala 677:58]
  wire  a_xor_b10 = a_10 ^ b_10; // @[FDIV.scala 678:21]
  wire  a_and_b10 = a_10 & b_10; // @[FDIV.scala 679:21]
  wire  sum_10 = a_xor_b10 ^ cin_10; // @[FDIV.scala 680:23]
  wire  cout_10 = a_and_b10 | a_xor_b10 & cin_10; // @[FDIV.scala 681:24]
  wire [1:0] temp_10 = {cout_10,sum_10}; // @[Cat.scala 31:58]
  wire  a_11 = io_in_0[11]; // @[FDIV.scala 677:32]
  wire  b_11 = io_in_1[11]; // @[FDIV.scala 677:45]
  wire  cin_11 = io_in_2[11]; // @[FDIV.scala 677:58]
  wire  a_xor_b11 = a_11 ^ b_11; // @[FDIV.scala 678:21]
  wire  a_and_b11 = a_11 & b_11; // @[FDIV.scala 679:21]
  wire  sum_11 = a_xor_b11 ^ cin_11; // @[FDIV.scala 680:23]
  wire  cout_11 = a_and_b11 | a_xor_b11 & cin_11; // @[FDIV.scala 681:24]
  wire [1:0] temp_11 = {cout_11,sum_11}; // @[Cat.scala 31:58]
  wire  a_12 = io_in_0[12]; // @[FDIV.scala 677:32]
  wire  b_12 = io_in_1[12]; // @[FDIV.scala 677:45]
  wire  cin_12 = io_in_2[12]; // @[FDIV.scala 677:58]
  wire  a_xor_b12 = a_12 ^ b_12; // @[FDIV.scala 678:21]
  wire  a_and_b12 = a_12 & b_12; // @[FDIV.scala 679:21]
  wire  sum_12 = a_xor_b12 ^ cin_12; // @[FDIV.scala 680:23]
  wire  cout_12 = a_and_b12 | a_xor_b12 & cin_12; // @[FDIV.scala 681:24]
  wire [1:0] temp_12 = {cout_12,sum_12}; // @[Cat.scala 31:58]
  wire  a_13 = io_in_0[13]; // @[FDIV.scala 677:32]
  wire  b_13 = io_in_1[13]; // @[FDIV.scala 677:45]
  wire  cin_13 = io_in_2[13]; // @[FDIV.scala 677:58]
  wire  a_xor_b13 = a_13 ^ b_13; // @[FDIV.scala 678:21]
  wire  a_and_b13 = a_13 & b_13; // @[FDIV.scala 679:21]
  wire  sum_13 = a_xor_b13 ^ cin_13; // @[FDIV.scala 680:23]
  wire  cout_13 = a_and_b13 | a_xor_b13 & cin_13; // @[FDIV.scala 681:24]
  wire [1:0] temp_13 = {cout_13,sum_13}; // @[Cat.scala 31:58]
  wire  a_14 = io_in_0[14]; // @[FDIV.scala 677:32]
  wire  b_14 = io_in_1[14]; // @[FDIV.scala 677:45]
  wire  cin_14 = io_in_2[14]; // @[FDIV.scala 677:58]
  wire  a_xor_b14 = a_14 ^ b_14; // @[FDIV.scala 678:21]
  wire  a_and_b14 = a_14 & b_14; // @[FDIV.scala 679:21]
  wire  sum_14 = a_xor_b14 ^ cin_14; // @[FDIV.scala 680:23]
  wire  cout_14 = a_and_b14 | a_xor_b14 & cin_14; // @[FDIV.scala 681:24]
  wire [1:0] temp_14 = {cout_14,sum_14}; // @[Cat.scala 31:58]
  wire  a_15 = io_in_0[15]; // @[FDIV.scala 677:32]
  wire  b_15 = io_in_1[15]; // @[FDIV.scala 677:45]
  wire  cin_15 = io_in_2[15]; // @[FDIV.scala 677:58]
  wire  a_xor_b15 = a_15 ^ b_15; // @[FDIV.scala 678:21]
  wire  a_and_b15 = a_15 & b_15; // @[FDIV.scala 679:21]
  wire  sum_15 = a_xor_b15 ^ cin_15; // @[FDIV.scala 680:23]
  wire  cout_15 = a_and_b15 | a_xor_b15 & cin_15; // @[FDIV.scala 681:24]
  wire [1:0] temp_15 = {cout_15,sum_15}; // @[Cat.scala 31:58]
  wire  a_16 = io_in_0[16]; // @[FDIV.scala 677:32]
  wire  b_16 = io_in_1[16]; // @[FDIV.scala 677:45]
  wire  cin_16 = io_in_2[16]; // @[FDIV.scala 677:58]
  wire  a_xor_b16 = a_16 ^ b_16; // @[FDIV.scala 678:21]
  wire  a_and_b16 = a_16 & b_16; // @[FDIV.scala 679:21]
  wire  sum_16 = a_xor_b16 ^ cin_16; // @[FDIV.scala 680:23]
  wire  cout_16 = a_and_b16 | a_xor_b16 & cin_16; // @[FDIV.scala 681:24]
  wire [1:0] temp_16 = {cout_16,sum_16}; // @[Cat.scala 31:58]
  wire  a_17 = io_in_0[17]; // @[FDIV.scala 677:32]
  wire  b_17 = io_in_1[17]; // @[FDIV.scala 677:45]
  wire  cin_17 = io_in_2[17]; // @[FDIV.scala 677:58]
  wire  a_xor_b17 = a_17 ^ b_17; // @[FDIV.scala 678:21]
  wire  a_and_b17 = a_17 & b_17; // @[FDIV.scala 679:21]
  wire  sum_17 = a_xor_b17 ^ cin_17; // @[FDIV.scala 680:23]
  wire  cout_17 = a_and_b17 | a_xor_b17 & cin_17; // @[FDIV.scala 681:24]
  wire [1:0] temp_17 = {cout_17,sum_17}; // @[Cat.scala 31:58]
  wire  a_18 = io_in_0[18]; // @[FDIV.scala 677:32]
  wire  b_18 = io_in_1[18]; // @[FDIV.scala 677:45]
  wire  cin_18 = io_in_2[18]; // @[FDIV.scala 677:58]
  wire  a_xor_b18 = a_18 ^ b_18; // @[FDIV.scala 678:21]
  wire  a_and_b18 = a_18 & b_18; // @[FDIV.scala 679:21]
  wire  sum_18 = a_xor_b18 ^ cin_18; // @[FDIV.scala 680:23]
  wire  cout_18 = a_and_b18 | a_xor_b18 & cin_18; // @[FDIV.scala 681:24]
  wire [1:0] temp_18 = {cout_18,sum_18}; // @[Cat.scala 31:58]
  wire  a_19 = io_in_0[19]; // @[FDIV.scala 677:32]
  wire  b_19 = io_in_1[19]; // @[FDIV.scala 677:45]
  wire  cin_19 = io_in_2[19]; // @[FDIV.scala 677:58]
  wire  a_xor_b19 = a_19 ^ b_19; // @[FDIV.scala 678:21]
  wire  a_and_b19 = a_19 & b_19; // @[FDIV.scala 679:21]
  wire  sum_19 = a_xor_b19 ^ cin_19; // @[FDIV.scala 680:23]
  wire  cout_19 = a_and_b19 | a_xor_b19 & cin_19; // @[FDIV.scala 681:24]
  wire [1:0] temp_19 = {cout_19,sum_19}; // @[Cat.scala 31:58]
  wire  a_20 = io_in_0[20]; // @[FDIV.scala 677:32]
  wire  b_20 = io_in_1[20]; // @[FDIV.scala 677:45]
  wire  cin_20 = io_in_2[20]; // @[FDIV.scala 677:58]
  wire  a_xor_b20 = a_20 ^ b_20; // @[FDIV.scala 678:21]
  wire  a_and_b20 = a_20 & b_20; // @[FDIV.scala 679:21]
  wire  sum_20 = a_xor_b20 ^ cin_20; // @[FDIV.scala 680:23]
  wire  cout_20 = a_and_b20 | a_xor_b20 & cin_20; // @[FDIV.scala 681:24]
  wire [1:0] temp_20 = {cout_20,sum_20}; // @[Cat.scala 31:58]
  wire  a_21 = io_in_0[21]; // @[FDIV.scala 677:32]
  wire  b_21 = io_in_1[21]; // @[FDIV.scala 677:45]
  wire  cin_21 = io_in_2[21]; // @[FDIV.scala 677:58]
  wire  a_xor_b21 = a_21 ^ b_21; // @[FDIV.scala 678:21]
  wire  a_and_b21 = a_21 & b_21; // @[FDIV.scala 679:21]
  wire  sum_21 = a_xor_b21 ^ cin_21; // @[FDIV.scala 680:23]
  wire  cout_21 = a_and_b21 | a_xor_b21 & cin_21; // @[FDIV.scala 681:24]
  wire [1:0] temp_21 = {cout_21,sum_21}; // @[Cat.scala 31:58]
  wire  a_22 = io_in_0[22]; // @[FDIV.scala 677:32]
  wire  b_22 = io_in_1[22]; // @[FDIV.scala 677:45]
  wire  cin_22 = io_in_2[22]; // @[FDIV.scala 677:58]
  wire  a_xor_b22 = a_22 ^ b_22; // @[FDIV.scala 678:21]
  wire  a_and_b22 = a_22 & b_22; // @[FDIV.scala 679:21]
  wire  sum_22 = a_xor_b22 ^ cin_22; // @[FDIV.scala 680:23]
  wire  cout_22 = a_and_b22 | a_xor_b22 & cin_22; // @[FDIV.scala 681:24]
  wire [1:0] temp_22 = {cout_22,sum_22}; // @[Cat.scala 31:58]
  wire  a_23 = io_in_0[23]; // @[FDIV.scala 677:32]
  wire  b_23 = io_in_1[23]; // @[FDIV.scala 677:45]
  wire  cin_23 = io_in_2[23]; // @[FDIV.scala 677:58]
  wire  a_xor_b23 = a_23 ^ b_23; // @[FDIV.scala 678:21]
  wire  a_and_b23 = a_23 & b_23; // @[FDIV.scala 679:21]
  wire  sum_23 = a_xor_b23 ^ cin_23; // @[FDIV.scala 680:23]
  wire  cout_23 = a_and_b23 | a_xor_b23 & cin_23; // @[FDIV.scala 681:24]
  wire [1:0] temp_23 = {cout_23,sum_23}; // @[Cat.scala 31:58]
  wire  a_24 = io_in_0[24]; // @[FDIV.scala 677:32]
  wire  b_24 = io_in_1[24]; // @[FDIV.scala 677:45]
  wire  cin_24 = io_in_2[24]; // @[FDIV.scala 677:58]
  wire  a_xor_b24 = a_24 ^ b_24; // @[FDIV.scala 678:21]
  wire  a_and_b24 = a_24 & b_24; // @[FDIV.scala 679:21]
  wire  sum_24 = a_xor_b24 ^ cin_24; // @[FDIV.scala 680:23]
  wire  cout_24 = a_and_b24 | a_xor_b24 & cin_24; // @[FDIV.scala 681:24]
  wire [1:0] temp_24 = {cout_24,sum_24}; // @[Cat.scala 31:58]
  wire  a_25 = io_in_0[25]; // @[FDIV.scala 677:32]
  wire  b_25 = io_in_1[25]; // @[FDIV.scala 677:45]
  wire  cin_25 = io_in_2[25]; // @[FDIV.scala 677:58]
  wire  a_xor_b25 = a_25 ^ b_25; // @[FDIV.scala 678:21]
  wire  a_and_b25 = a_25 & b_25; // @[FDIV.scala 679:21]
  wire  sum_25 = a_xor_b25 ^ cin_25; // @[FDIV.scala 680:23]
  wire  cout_25 = a_and_b25 | a_xor_b25 & cin_25; // @[FDIV.scala 681:24]
  wire [1:0] temp_25 = {cout_25,sum_25}; // @[Cat.scala 31:58]
  wire  a_26 = io_in_0[26]; // @[FDIV.scala 677:32]
  wire  b_26 = io_in_1[26]; // @[FDIV.scala 677:45]
  wire  cin_26 = io_in_2[26]; // @[FDIV.scala 677:58]
  wire  a_xor_b26 = a_26 ^ b_26; // @[FDIV.scala 678:21]
  wire  a_and_b26 = a_26 & b_26; // @[FDIV.scala 679:21]
  wire  sum_26 = a_xor_b26 ^ cin_26; // @[FDIV.scala 680:23]
  wire  cout_26 = a_and_b26 | a_xor_b26 & cin_26; // @[FDIV.scala 681:24]
  wire [1:0] temp_26 = {cout_26,sum_26}; // @[Cat.scala 31:58]
  wire [5:0] io_out_0_lo_lo = {temp_5[0],temp_4[0],temp_3[0],temp_2[0],temp_1[0],temp_0[0]}; // @[Cat.scala 31:58]
  wire [12:0] io_out_0_lo = {temp_12[0],temp_11[0],temp_10[0],temp_9[0],temp_8[0],temp_7[0],temp_6[0],io_out_0_lo_lo}; // @[Cat.scala 31:58]
  wire [6:0] io_out_0_hi_lo = {temp_19[0],temp_18[0],temp_17[0],temp_16[0],temp_15[0],temp_14[0],temp_13[0]}; // @[Cat.scala 31:58]
  wire [13:0] io_out_0_hi = {temp_26[0],temp_25[0],temp_24[0],temp_23[0],temp_22[0],temp_21[0],temp_20[0],io_out_0_hi_lo
    }; // @[Cat.scala 31:58]
  wire [5:0] io_out_1_lo_lo = {temp_5[1],temp_4[1],temp_3[1],temp_2[1],temp_1[1],temp_0[1]}; // @[Cat.scala 31:58]
  wire [12:0] io_out_1_lo = {temp_12[1],temp_11[1],temp_10[1],temp_9[1],temp_8[1],temp_7[1],temp_6[1],io_out_1_lo_lo}; // @[Cat.scala 31:58]
  wire [6:0] io_out_1_hi_lo = {temp_19[1],temp_18[1],temp_17[1],temp_16[1],temp_15[1],temp_14[1],temp_13[1]}; // @[Cat.scala 31:58]
  wire [13:0] io_out_1_hi = {temp_26[1],temp_25[1],temp_24[1],temp_23[1],temp_22[1],temp_21[1],temp_20[1],io_out_1_hi_lo
    }; // @[Cat.scala 31:58]
  assign io_out_0 = {io_out_0_hi,io_out_0_lo}; // @[Cat.scala 31:58]
  assign io_out_1 = {io_out_1_hi,io_out_1_lo}; // @[Cat.scala 31:58]
endmodule

