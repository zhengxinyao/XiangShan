module Predictor(
  input          clock,
  input          reset,
  input          io_bpu_to_ftq_resp_ready,
  output         io_bpu_to_ftq_resp_valid,
  output [38:0]  io_bpu_to_ftq_resp_bits_s1_pc,
  output         io_bpu_to_ftq_resp_bits_s1_full_pred_br_taken_mask_0,
  output         io_bpu_to_ftq_resp_bits_s1_full_pred_br_taken_mask_1,
  output         io_bpu_to_ftq_resp_bits_s1_full_pred_slot_valids_0,
  output         io_bpu_to_ftq_resp_bits_s1_full_pred_slot_valids_1,
  output [38:0]  io_bpu_to_ftq_resp_bits_s1_full_pred_targets_0,
  output [38:0]  io_bpu_to_ftq_resp_bits_s1_full_pred_targets_1,
  output [2:0]   io_bpu_to_ftq_resp_bits_s1_full_pred_offsets_0,
  output [2:0]   io_bpu_to_ftq_resp_bits_s1_full_pred_offsets_1,
  output [38:0]  io_bpu_to_ftq_resp_bits_s1_full_pred_fallThroughAddr,
  output         io_bpu_to_ftq_resp_bits_s1_full_pred_fallThroughErr,
  output         io_bpu_to_ftq_resp_bits_s1_full_pred_is_br_sharing,
  output         io_bpu_to_ftq_resp_bits_s1_full_pred_hit,
  output [38:0]  io_bpu_to_ftq_resp_bits_s2_pc,
  output         io_bpu_to_ftq_resp_bits_s2_valid,
  output         io_bpu_to_ftq_resp_bits_s2_hasRedirect,
  output         io_bpu_to_ftq_resp_bits_s2_ftq_idx_flag,
  output [2:0]   io_bpu_to_ftq_resp_bits_s2_ftq_idx_value,
  output         io_bpu_to_ftq_resp_bits_s2_full_pred_br_taken_mask_0,
  output         io_bpu_to_ftq_resp_bits_s2_full_pred_br_taken_mask_1,
  output         io_bpu_to_ftq_resp_bits_s2_full_pred_slot_valids_0,
  output         io_bpu_to_ftq_resp_bits_s2_full_pred_slot_valids_1,
  output [38:0]  io_bpu_to_ftq_resp_bits_s2_full_pred_targets_0,
  output [38:0]  io_bpu_to_ftq_resp_bits_s2_full_pred_targets_1,
  output [2:0]   io_bpu_to_ftq_resp_bits_s2_full_pred_offsets_0,
  output [2:0]   io_bpu_to_ftq_resp_bits_s2_full_pred_offsets_1,
  output [38:0]  io_bpu_to_ftq_resp_bits_s2_full_pred_fallThroughAddr,
  output         io_bpu_to_ftq_resp_bits_s2_full_pred_fallThroughErr,
  output         io_bpu_to_ftq_resp_bits_s2_full_pred_is_br_sharing,
  output         io_bpu_to_ftq_resp_bits_s2_full_pred_hit,
  output [38:0]  io_bpu_to_ftq_resp_bits_s3_pc,
  output         io_bpu_to_ftq_resp_bits_s3_valid,
  output         io_bpu_to_ftq_resp_bits_s3_hasRedirect,
  output         io_bpu_to_ftq_resp_bits_s3_ftq_idx_flag,
  output [2:0]   io_bpu_to_ftq_resp_bits_s3_ftq_idx_value,
  output         io_bpu_to_ftq_resp_bits_s3_full_pred_br_taken_mask_0,
  output         io_bpu_to_ftq_resp_bits_s3_full_pred_br_taken_mask_1,
  output         io_bpu_to_ftq_resp_bits_s3_full_pred_slot_valids_0,
  output         io_bpu_to_ftq_resp_bits_s3_full_pred_slot_valids_1,
  output [38:0]  io_bpu_to_ftq_resp_bits_s3_full_pred_targets_0,
  output [38:0]  io_bpu_to_ftq_resp_bits_s3_full_pred_targets_1,
  output [2:0]   io_bpu_to_ftq_resp_bits_s3_full_pred_offsets_0,
  output [2:0]   io_bpu_to_ftq_resp_bits_s3_full_pred_offsets_1,
  output [38:0]  io_bpu_to_ftq_resp_bits_s3_full_pred_fallThroughAddr,
  output         io_bpu_to_ftq_resp_bits_s3_full_pred_fallThroughErr,
  output         io_bpu_to_ftq_resp_bits_s3_full_pred_is_br_sharing,
  output         io_bpu_to_ftq_resp_bits_s3_full_pred_hit,
  output [255:0] io_bpu_to_ftq_resp_bits_last_stage_meta,
  output [7:0]   io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_17_folded_hist,
  output [7:0]   io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_16_folded_hist,
  output [10:0]  io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_15_folded_hist,
  output [6:0]   io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_14_folded_hist,
  output [6:0]   io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_13_folded_hist,
  output [6:0]   io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_12_folded_hist,
  output [7:0]   io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_11_folded_hist,
  output [8:0]   io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_10_folded_hist,
  output [6:0]   io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_9_folded_hist,
  output [7:0]   io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_8_folded_hist,
  output [8:0]   io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_7_folded_hist,
  output [8:0]   io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_6_folded_hist,
  output [10:0]  io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_5_folded_hist,
  output [3:0]   io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_4_folded_hist,
  output [10:0]  io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_3_folded_hist,
  output [7:0]   io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_2_folded_hist,
  output [7:0]   io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_1_folded_hist,
  output [7:0]   io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_0_folded_hist,
  output         io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_5_bits_0,
  output         io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_5_bits_1,
  output         io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_5_bits_2,
  output         io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_5_bits_3,
  output         io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_4_bits_0,
  output         io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_4_bits_1,
  output         io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_4_bits_2,
  output         io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_4_bits_3,
  output         io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_3_bits_0,
  output         io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_3_bits_1,
  output         io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_3_bits_2,
  output         io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_3_bits_3,
  output         io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_2_bits_0,
  output         io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_2_bits_1,
  output         io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_2_bits_2,
  output         io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_2_bits_3,
  output         io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_1_bits_0,
  output         io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_1_bits_1,
  output         io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_1_bits_2,
  output         io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_1_bits_3,
  output         io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_0_bits_0,
  output         io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_0_bits_1,
  output         io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_0_bits_2,
  output         io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_0_bits_3,
  output [2:0]   io_bpu_to_ftq_resp_bits_last_stage_spec_info_lastBrNumOH,
  output         io_bpu_to_ftq_resp_bits_last_stage_spec_info_histPtr_flag,
  output [7:0]   io_bpu_to_ftq_resp_bits_last_stage_spec_info_histPtr_value,
  output [4:0]   io_bpu_to_ftq_resp_bits_last_stage_spec_info_rasSp,
  output [38:0]  io_bpu_to_ftq_resp_bits_last_stage_spec_info_rasTop_retAddr,
  output [7:0]   io_bpu_to_ftq_resp_bits_last_stage_spec_info_rasTop_ctr,
  output         io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_valid,
  output [2:0]   io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_brSlots_0_offset,
  output [11:0]  io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_brSlots_0_lower,
  output [1:0]   io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_brSlots_0_tarStat,
  output         io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_brSlots_0_sharing,
  output         io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_brSlots_0_valid,
  output [2:0]   io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_tailSlot_offset,
  output [19:0]  io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_tailSlot_lower,
  output [1:0]   io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_tailSlot_tarStat,
  output         io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_tailSlot_sharing,
  output         io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_tailSlot_valid,
  output [2:0]   io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_pftAddr,
  output         io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_carry,
  output         io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_isCall,
  output         io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_isRet,
  output         io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_isJalr,
  output         io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_last_may_be_rvi_call,
  output         io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_always_taken_0,
  output         io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_always_taken_1,
  input          io_ftq_to_bpu_redirect_valid,
  input          io_ftq_to_bpu_redirect_bits_level,
  input  [38:0]  io_ftq_to_bpu_redirect_bits_cfiUpdate_pc,
  input          io_ftq_to_bpu_redirect_bits_cfiUpdate_pd_isRVC,
  input          io_ftq_to_bpu_redirect_bits_cfiUpdate_pd_isCall,
  input          io_ftq_to_bpu_redirect_bits_cfiUpdate_pd_isRet,
  input  [4:0]   io_ftq_to_bpu_redirect_bits_cfiUpdate_rasSp,
  input  [38:0]  io_ftq_to_bpu_redirect_bits_cfiUpdate_rasEntry_retAddr,
  input  [7:0]   io_ftq_to_bpu_redirect_bits_cfiUpdate_rasEntry_ctr,
  input  [7:0]   io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_17_folded_hist,
  input  [7:0]   io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_16_folded_hist,
  input  [10:0]  io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_15_folded_hist,
  input  [6:0]   io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_14_folded_hist,
  input  [6:0]   io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_13_folded_hist,
  input  [6:0]   io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_12_folded_hist,
  input  [7:0]   io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_11_folded_hist,
  input  [8:0]   io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_10_folded_hist,
  input  [6:0]   io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_9_folded_hist,
  input  [7:0]   io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_8_folded_hist,
  input  [8:0]   io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_7_folded_hist,
  input  [8:0]   io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_6_folded_hist,
  input  [10:0]  io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_5_folded_hist,
  input  [3:0]   io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_4_folded_hist,
  input  [10:0]  io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_3_folded_hist,
  input  [7:0]   io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_2_folded_hist,
  input  [7:0]   io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_1_folded_hist,
  input  [7:0]   io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_0_folded_hist,
  input          io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_5_bits_0,
  input          io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_5_bits_1,
  input          io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_5_bits_2,
  input          io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_5_bits_3,
  input          io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_4_bits_0,
  input          io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_4_bits_1,
  input          io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_4_bits_2,
  input          io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_3_bits_0,
  input          io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_3_bits_1,
  input          io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_3_bits_2,
  input          io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_3_bits_3,
  input          io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_2_bits_0,
  input          io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_2_bits_1,
  input          io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_2_bits_2,
  input          io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_2_bits_3,
  input          io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_1_bits_0,
  input          io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_1_bits_1,
  input          io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_1_bits_2,
  input          io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_1_bits_3,
  input          io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_0_bits_0,
  input          io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_0_bits_1,
  input          io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_0_bits_2,
  input          io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_0_bits_3,
  input  [2:0]   io_ftq_to_bpu_redirect_bits_cfiUpdate_lastBrNumOH,
  input          io_ftq_to_bpu_redirect_bits_cfiUpdate_histPtr_flag,
  input  [7:0]   io_ftq_to_bpu_redirect_bits_cfiUpdate_histPtr_value,
  input  [38:0]  io_ftq_to_bpu_redirect_bits_cfiUpdate_target,
  input          io_ftq_to_bpu_redirect_bits_cfiUpdate_taken,
  input  [1:0]   io_ftq_to_bpu_redirect_bits_cfiUpdate_shift,
  input          io_ftq_to_bpu_redirect_bits_cfiUpdate_addIntoHist,
  input          io_ftq_to_bpu_update_valid,
  input  [38:0]  io_ftq_to_bpu_update_bits_pc,
  input  [7:0]   io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_17_folded_hist,
  input  [7:0]   io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_16_folded_hist,
  input  [10:0]  io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_15_folded_hist,
  input  [6:0]   io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_14_folded_hist,
  input  [6:0]   io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_13_folded_hist,
  input  [6:0]   io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_12_folded_hist,
  input  [8:0]   io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_10_folded_hist,
  input  [6:0]   io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_9_folded_hist,
  input  [7:0]   io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_8_folded_hist,
  input  [8:0]   io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_7_folded_hist,
  input  [8:0]   io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_6_folded_hist,
  input  [10:0]  io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_5_folded_hist,
  input  [3:0]   io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_4_folded_hist,
  input  [10:0]  io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_3_folded_hist,
  input  [7:0]   io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_2_folded_hist,
  input  [7:0]   io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_1_folded_hist,
  input  [7:0]   io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_0_folded_hist,
  input          io_ftq_to_bpu_update_bits_ftb_entry_valid,
  input  [2:0]   io_ftq_to_bpu_update_bits_ftb_entry_brSlots_0_offset,
  input  [11:0]  io_ftq_to_bpu_update_bits_ftb_entry_brSlots_0_lower,
  input  [1:0]   io_ftq_to_bpu_update_bits_ftb_entry_brSlots_0_tarStat,
  input          io_ftq_to_bpu_update_bits_ftb_entry_brSlots_0_sharing,
  input          io_ftq_to_bpu_update_bits_ftb_entry_brSlots_0_valid,
  input  [2:0]   io_ftq_to_bpu_update_bits_ftb_entry_tailSlot_offset,
  input  [19:0]  io_ftq_to_bpu_update_bits_ftb_entry_tailSlot_lower,
  input  [1:0]   io_ftq_to_bpu_update_bits_ftb_entry_tailSlot_tarStat,
  input          io_ftq_to_bpu_update_bits_ftb_entry_tailSlot_sharing,
  input          io_ftq_to_bpu_update_bits_ftb_entry_tailSlot_valid,
  input  [2:0]   io_ftq_to_bpu_update_bits_ftb_entry_pftAddr,
  input          io_ftq_to_bpu_update_bits_ftb_entry_carry,
  input          io_ftq_to_bpu_update_bits_ftb_entry_isCall,
  input          io_ftq_to_bpu_update_bits_ftb_entry_isRet,
  input          io_ftq_to_bpu_update_bits_ftb_entry_isJalr,
  input          io_ftq_to_bpu_update_bits_ftb_entry_last_may_be_rvi_call,
  input          io_ftq_to_bpu_update_bits_ftb_entry_always_taken_0,
  input          io_ftq_to_bpu_update_bits_ftb_entry_always_taken_1,
  input          io_ftq_to_bpu_update_bits_br_taken_mask_0,
  input          io_ftq_to_bpu_update_bits_br_taken_mask_1,
  input          io_ftq_to_bpu_update_bits_jmp_taken,
  input          io_ftq_to_bpu_update_bits_mispred_mask_0,
  input          io_ftq_to_bpu_update_bits_mispred_mask_1,
  input          io_ftq_to_bpu_update_bits_mispred_mask_2,
  input          io_ftq_to_bpu_update_bits_old_entry,
  input  [255:0] io_ftq_to_bpu_update_bits_meta,
  input  [38:0]  io_ftq_to_bpu_update_bits_full_target,
  input          io_ftq_to_bpu_enq_ptr_flag,
  input  [2:0]   io_ftq_to_bpu_enq_ptr_value,
  input          io_ctrl_ubtb_enable,
  input          io_ctrl_btb_enable,
  input          io_ctrl_tage_enable,
  input          io_ctrl_sc_enable,
  input          io_ctrl_ras_enable,
  input  [35:0]  io_reset_vector,
  output [5:0]   io_perf_0_value,
  output [5:0]   io_perf_1_value,
  output [5:0]   io_perf_2_value,
  output [5:0]   io_perf_3_value,
  output [5:0]   io_perf_4_value,
  output [5:0]   io_perf_5_value,
  output [5:0]   io_perf_6_value
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [63:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [63:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [63:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [63:0] _RAND_393;
  reg [63:0] _RAND_394;
  reg [63:0] _RAND_395;
  reg [63:0] _RAND_396;
  reg [63:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [63:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [255:0] _RAND_450;
  reg [63:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
`endif // RANDOMIZE_REG_INIT
  wire  ctrl_delay_clock; // @[Hold.scala 97:23]
  wire  ctrl_delay_io_in_ubtb_enable; // @[Hold.scala 97:23]
  wire  ctrl_delay_io_in_btb_enable; // @[Hold.scala 97:23]
  wire  ctrl_delay_io_in_tage_enable; // @[Hold.scala 97:23]
  wire  ctrl_delay_io_in_sc_enable; // @[Hold.scala 97:23]
  wire  ctrl_delay_io_in_ras_enable; // @[Hold.scala 97:23]
  wire  ctrl_delay_io_out_ubtb_enable; // @[Hold.scala 97:23]
  wire  ctrl_delay_io_out_btb_enable; // @[Hold.scala 97:23]
  wire  ctrl_delay_io_out_tage_enable; // @[Hold.scala 97:23]
  wire  ctrl_delay_io_out_sc_enable; // @[Hold.scala 97:23]
  wire  ctrl_delay_io_out_ras_enable; // @[Hold.scala 97:23]
  wire  predictors_clock; // @[BPU.scala 245:26]
  wire  predictors_reset; // @[BPU.scala 245:26]
  wire [35:0] predictors_io_reset_vector; // @[BPU.scala 245:26]
  wire [38:0] predictors_io_in_bits_s0_pc; // @[BPU.scala 245:26]
  wire [7:0] predictors_io_in_bits_folded_hist_hist_17_folded_hist; // @[BPU.scala 245:26]
  wire [7:0] predictors_io_in_bits_folded_hist_hist_16_folded_hist; // @[BPU.scala 245:26]
  wire [10:0] predictors_io_in_bits_folded_hist_hist_15_folded_hist; // @[BPU.scala 245:26]
  wire [6:0] predictors_io_in_bits_folded_hist_hist_14_folded_hist; // @[BPU.scala 245:26]
  wire [6:0] predictors_io_in_bits_folded_hist_hist_13_folded_hist; // @[BPU.scala 245:26]
  wire [6:0] predictors_io_in_bits_folded_hist_hist_12_folded_hist; // @[BPU.scala 245:26]
  wire [8:0] predictors_io_in_bits_folded_hist_hist_10_folded_hist; // @[BPU.scala 245:26]
  wire [6:0] predictors_io_in_bits_folded_hist_hist_9_folded_hist; // @[BPU.scala 245:26]
  wire [7:0] predictors_io_in_bits_folded_hist_hist_8_folded_hist; // @[BPU.scala 245:26]
  wire [8:0] predictors_io_in_bits_folded_hist_hist_7_folded_hist; // @[BPU.scala 245:26]
  wire [8:0] predictors_io_in_bits_folded_hist_hist_6_folded_hist; // @[BPU.scala 245:26]
  wire [10:0] predictors_io_in_bits_folded_hist_hist_5_folded_hist; // @[BPU.scala 245:26]
  wire [3:0] predictors_io_in_bits_folded_hist_hist_4_folded_hist; // @[BPU.scala 245:26]
  wire [10:0] predictors_io_in_bits_folded_hist_hist_3_folded_hist; // @[BPU.scala 245:26]
  wire [7:0] predictors_io_in_bits_folded_hist_hist_2_folded_hist; // @[BPU.scala 245:26]
  wire [7:0] predictors_io_in_bits_folded_hist_hist_1_folded_hist; // @[BPU.scala 245:26]
  wire [7:0] predictors_io_in_bits_folded_hist_hist_0_folded_hist; // @[BPU.scala 245:26]
  wire [38:0] predictors_io_out_s1_pc; // @[BPU.scala 245:26]
  wire  predictors_io_out_s1_full_pred_br_taken_mask_0; // @[BPU.scala 245:26]
  wire  predictors_io_out_s1_full_pred_br_taken_mask_1; // @[BPU.scala 245:26]
  wire  predictors_io_out_s1_full_pred_slot_valids_0; // @[BPU.scala 245:26]
  wire  predictors_io_out_s1_full_pred_slot_valids_1; // @[BPU.scala 245:26]
  wire [38:0] predictors_io_out_s1_full_pred_targets_0; // @[BPU.scala 245:26]
  wire [38:0] predictors_io_out_s1_full_pred_targets_1; // @[BPU.scala 245:26]
  wire [2:0] predictors_io_out_s1_full_pred_offsets_0; // @[BPU.scala 245:26]
  wire [2:0] predictors_io_out_s1_full_pred_offsets_1; // @[BPU.scala 245:26]
  wire [38:0] predictors_io_out_s1_full_pred_fallThroughAddr; // @[BPU.scala 245:26]
  wire  predictors_io_out_s1_full_pred_fallThroughErr; // @[BPU.scala 245:26]
  wire  predictors_io_out_s1_full_pred_is_br_sharing; // @[BPU.scala 245:26]
  wire  predictors_io_out_s1_full_pred_hit; // @[BPU.scala 245:26]
  wire [38:0] predictors_io_out_s2_pc; // @[BPU.scala 245:26]
  wire  predictors_io_out_s2_full_pred_br_taken_mask_0; // @[BPU.scala 245:26]
  wire  predictors_io_out_s2_full_pred_br_taken_mask_1; // @[BPU.scala 245:26]
  wire  predictors_io_out_s2_full_pred_slot_valids_0; // @[BPU.scala 245:26]
  wire  predictors_io_out_s2_full_pred_slot_valids_1; // @[BPU.scala 245:26]
  wire [38:0] predictors_io_out_s2_full_pred_targets_0; // @[BPU.scala 245:26]
  wire [38:0] predictors_io_out_s2_full_pred_targets_1; // @[BPU.scala 245:26]
  wire [2:0] predictors_io_out_s2_full_pred_offsets_0; // @[BPU.scala 245:26]
  wire [2:0] predictors_io_out_s2_full_pred_offsets_1; // @[BPU.scala 245:26]
  wire [38:0] predictors_io_out_s2_full_pred_fallThroughAddr; // @[BPU.scala 245:26]
  wire  predictors_io_out_s2_full_pred_fallThroughErr; // @[BPU.scala 245:26]
  wire  predictors_io_out_s2_full_pred_is_br_sharing; // @[BPU.scala 245:26]
  wire  predictors_io_out_s2_full_pred_hit; // @[BPU.scala 245:26]
  wire [38:0] predictors_io_out_s3_pc; // @[BPU.scala 245:26]
  wire  predictors_io_out_s3_full_pred_br_taken_mask_0; // @[BPU.scala 245:26]
  wire  predictors_io_out_s3_full_pred_br_taken_mask_1; // @[BPU.scala 245:26]
  wire  predictors_io_out_s3_full_pred_slot_valids_0; // @[BPU.scala 245:26]
  wire  predictors_io_out_s3_full_pred_slot_valids_1; // @[BPU.scala 245:26]
  wire [38:0] predictors_io_out_s3_full_pred_targets_0; // @[BPU.scala 245:26]
  wire [38:0] predictors_io_out_s3_full_pred_targets_1; // @[BPU.scala 245:26]
  wire [2:0] predictors_io_out_s3_full_pred_offsets_0; // @[BPU.scala 245:26]
  wire [2:0] predictors_io_out_s3_full_pred_offsets_1; // @[BPU.scala 245:26]
  wire [38:0] predictors_io_out_s3_full_pred_fallThroughAddr; // @[BPU.scala 245:26]
  wire  predictors_io_out_s3_full_pred_fallThroughErr; // @[BPU.scala 245:26]
  wire  predictors_io_out_s3_full_pred_is_br_sharing; // @[BPU.scala 245:26]
  wire  predictors_io_out_s3_full_pred_hit; // @[BPU.scala 245:26]
  wire [255:0] predictors_io_out_last_stage_meta; // @[BPU.scala 245:26]
  wire [4:0] predictors_io_out_last_stage_spec_info_rasSp; // @[BPU.scala 245:26]
  wire [38:0] predictors_io_out_last_stage_spec_info_rasTop_retAddr; // @[BPU.scala 245:26]
  wire [7:0] predictors_io_out_last_stage_spec_info_rasTop_ctr; // @[BPU.scala 245:26]
  wire  predictors_io_out_last_stage_ftb_entry_valid; // @[BPU.scala 245:26]
  wire [2:0] predictors_io_out_last_stage_ftb_entry_brSlots_0_offset; // @[BPU.scala 245:26]
  wire [11:0] predictors_io_out_last_stage_ftb_entry_brSlots_0_lower; // @[BPU.scala 245:26]
  wire [1:0] predictors_io_out_last_stage_ftb_entry_brSlots_0_tarStat; // @[BPU.scala 245:26]
  wire  predictors_io_out_last_stage_ftb_entry_brSlots_0_sharing; // @[BPU.scala 245:26]
  wire  predictors_io_out_last_stage_ftb_entry_brSlots_0_valid; // @[BPU.scala 245:26]
  wire [2:0] predictors_io_out_last_stage_ftb_entry_tailSlot_offset; // @[BPU.scala 245:26]
  wire [19:0] predictors_io_out_last_stage_ftb_entry_tailSlot_lower; // @[BPU.scala 245:26]
  wire [1:0] predictors_io_out_last_stage_ftb_entry_tailSlot_tarStat; // @[BPU.scala 245:26]
  wire  predictors_io_out_last_stage_ftb_entry_tailSlot_sharing; // @[BPU.scala 245:26]
  wire  predictors_io_out_last_stage_ftb_entry_tailSlot_valid; // @[BPU.scala 245:26]
  wire [2:0] predictors_io_out_last_stage_ftb_entry_pftAddr; // @[BPU.scala 245:26]
  wire  predictors_io_out_last_stage_ftb_entry_carry; // @[BPU.scala 245:26]
  wire  predictors_io_out_last_stage_ftb_entry_isCall; // @[BPU.scala 245:26]
  wire  predictors_io_out_last_stage_ftb_entry_isRet; // @[BPU.scala 245:26]
  wire  predictors_io_out_last_stage_ftb_entry_isJalr; // @[BPU.scala 245:26]
  wire  predictors_io_out_last_stage_ftb_entry_last_may_be_rvi_call; // @[BPU.scala 245:26]
  wire  predictors_io_out_last_stage_ftb_entry_always_taken_0; // @[BPU.scala 245:26]
  wire  predictors_io_out_last_stage_ftb_entry_always_taken_1; // @[BPU.scala 245:26]
  wire  predictors_io_ctrl_ubtb_enable; // @[BPU.scala 245:26]
  wire  predictors_io_ctrl_btb_enable; // @[BPU.scala 245:26]
  wire  predictors_io_ctrl_tage_enable; // @[BPU.scala 245:26]
  wire  predictors_io_ctrl_sc_enable; // @[BPU.scala 245:26]
  wire  predictors_io_ctrl_ras_enable; // @[BPU.scala 245:26]
  wire  predictors_io_s0_fire; // @[BPU.scala 245:26]
  wire  predictors_io_s1_fire; // @[BPU.scala 245:26]
  wire  predictors_io_s2_fire; // @[BPU.scala 245:26]
  wire  predictors_io_s3_fire; // @[BPU.scala 245:26]
  wire  predictors_io_s3_redirect; // @[BPU.scala 245:26]
  wire  predictors_io_s1_ready; // @[BPU.scala 245:26]
  wire  predictors_io_update_valid; // @[BPU.scala 245:26]
  wire [38:0] predictors_io_update_bits_pc; // @[BPU.scala 245:26]
  wire [7:0] predictors_io_update_bits_spec_info_folded_hist_hist_17_folded_hist; // @[BPU.scala 245:26]
  wire [7:0] predictors_io_update_bits_spec_info_folded_hist_hist_16_folded_hist; // @[BPU.scala 245:26]
  wire [10:0] predictors_io_update_bits_spec_info_folded_hist_hist_15_folded_hist; // @[BPU.scala 245:26]
  wire [6:0] predictors_io_update_bits_spec_info_folded_hist_hist_14_folded_hist; // @[BPU.scala 245:26]
  wire [6:0] predictors_io_update_bits_spec_info_folded_hist_hist_13_folded_hist; // @[BPU.scala 245:26]
  wire [6:0] predictors_io_update_bits_spec_info_folded_hist_hist_12_folded_hist; // @[BPU.scala 245:26]
  wire [8:0] predictors_io_update_bits_spec_info_folded_hist_hist_10_folded_hist; // @[BPU.scala 245:26]
  wire [6:0] predictors_io_update_bits_spec_info_folded_hist_hist_9_folded_hist; // @[BPU.scala 245:26]
  wire [7:0] predictors_io_update_bits_spec_info_folded_hist_hist_8_folded_hist; // @[BPU.scala 245:26]
  wire [8:0] predictors_io_update_bits_spec_info_folded_hist_hist_7_folded_hist; // @[BPU.scala 245:26]
  wire [8:0] predictors_io_update_bits_spec_info_folded_hist_hist_6_folded_hist; // @[BPU.scala 245:26]
  wire [10:0] predictors_io_update_bits_spec_info_folded_hist_hist_5_folded_hist; // @[BPU.scala 245:26]
  wire [3:0] predictors_io_update_bits_spec_info_folded_hist_hist_4_folded_hist; // @[BPU.scala 245:26]
  wire [10:0] predictors_io_update_bits_spec_info_folded_hist_hist_3_folded_hist; // @[BPU.scala 245:26]
  wire [7:0] predictors_io_update_bits_spec_info_folded_hist_hist_2_folded_hist; // @[BPU.scala 245:26]
  wire [7:0] predictors_io_update_bits_spec_info_folded_hist_hist_1_folded_hist; // @[BPU.scala 245:26]
  wire [7:0] predictors_io_update_bits_spec_info_folded_hist_hist_0_folded_hist; // @[BPU.scala 245:26]
  wire  predictors_io_update_bits_ftb_entry_valid; // @[BPU.scala 245:26]
  wire [2:0] predictors_io_update_bits_ftb_entry_brSlots_0_offset; // @[BPU.scala 245:26]
  wire [11:0] predictors_io_update_bits_ftb_entry_brSlots_0_lower; // @[BPU.scala 245:26]
  wire [1:0] predictors_io_update_bits_ftb_entry_brSlots_0_tarStat; // @[BPU.scala 245:26]
  wire  predictors_io_update_bits_ftb_entry_brSlots_0_sharing; // @[BPU.scala 245:26]
  wire  predictors_io_update_bits_ftb_entry_brSlots_0_valid; // @[BPU.scala 245:26]
  wire [2:0] predictors_io_update_bits_ftb_entry_tailSlot_offset; // @[BPU.scala 245:26]
  wire [19:0] predictors_io_update_bits_ftb_entry_tailSlot_lower; // @[BPU.scala 245:26]
  wire [1:0] predictors_io_update_bits_ftb_entry_tailSlot_tarStat; // @[BPU.scala 245:26]
  wire  predictors_io_update_bits_ftb_entry_tailSlot_sharing; // @[BPU.scala 245:26]
  wire  predictors_io_update_bits_ftb_entry_tailSlot_valid; // @[BPU.scala 245:26]
  wire [2:0] predictors_io_update_bits_ftb_entry_pftAddr; // @[BPU.scala 245:26]
  wire  predictors_io_update_bits_ftb_entry_carry; // @[BPU.scala 245:26]
  wire  predictors_io_update_bits_ftb_entry_isCall; // @[BPU.scala 245:26]
  wire  predictors_io_update_bits_ftb_entry_isRet; // @[BPU.scala 245:26]
  wire  predictors_io_update_bits_ftb_entry_isJalr; // @[BPU.scala 245:26]
  wire  predictors_io_update_bits_ftb_entry_last_may_be_rvi_call; // @[BPU.scala 245:26]
  wire  predictors_io_update_bits_ftb_entry_always_taken_0; // @[BPU.scala 245:26]
  wire  predictors_io_update_bits_ftb_entry_always_taken_1; // @[BPU.scala 245:26]
  wire  predictors_io_update_bits_br_taken_mask_0; // @[BPU.scala 245:26]
  wire  predictors_io_update_bits_br_taken_mask_1; // @[BPU.scala 245:26]
  wire  predictors_io_update_bits_jmp_taken; // @[BPU.scala 245:26]
  wire  predictors_io_update_bits_mispred_mask_0; // @[BPU.scala 245:26]
  wire  predictors_io_update_bits_mispred_mask_1; // @[BPU.scala 245:26]
  wire  predictors_io_update_bits_mispred_mask_2; // @[BPU.scala 245:26]
  wire  predictors_io_update_bits_old_entry; // @[BPU.scala 245:26]
  wire [255:0] predictors_io_update_bits_meta; // @[BPU.scala 245:26]
  wire [38:0] predictors_io_update_bits_full_target; // @[BPU.scala 245:26]
  wire  predictors_io_redirect_valid; // @[BPU.scala 245:26]
  wire  predictors_io_redirect_bits_level; // @[BPU.scala 245:26]
  wire [38:0] predictors_io_redirect_bits_cfiUpdate_pc; // @[BPU.scala 245:26]
  wire  predictors_io_redirect_bits_cfiUpdate_pd_isRVC; // @[BPU.scala 245:26]
  wire  predictors_io_redirect_bits_cfiUpdate_pd_isCall; // @[BPU.scala 245:26]
  wire  predictors_io_redirect_bits_cfiUpdate_pd_isRet; // @[BPU.scala 245:26]
  wire [4:0] predictors_io_redirect_bits_cfiUpdate_rasSp; // @[BPU.scala 245:26]
  wire [38:0] predictors_io_redirect_bits_cfiUpdate_rasEntry_retAddr; // @[BPU.scala 245:26]
  wire [7:0] predictors_io_redirect_bits_cfiUpdate_rasEntry_ctr; // @[BPU.scala 245:26]
  wire [5:0] predictors_io_perf_0_value; // @[BPU.scala 245:26]
  wire [5:0] predictors_io_perf_1_value; // @[BPU.scala 245:26]
  wire [5:0] predictors_io_perf_2_value; // @[BPU.scala 245:26]
  wire [5:0] predictors_io_perf_3_value; // @[BPU.scala 245:26]
  wire [5:0] predictors_io_perf_4_value; // @[BPU.scala 245:26]
  wire [5:0] predictors_io_perf_5_value; // @[BPU.scala 245:26]
  wire [5:0] predictors_io_perf_6_value; // @[BPU.scala 245:26]
  wire  reset_vector_delay_clock; // @[Hold.scala 97:23]
  wire [35:0] reset_vector_delay_io_in; // @[Hold.scala 97:23]
  wire [35:0] reset_vector_delay_io_out; // @[Hold.scala 97:23]
  wire  s0_pc_ppm_s2_target_sel; // @[PriorityMuxGen.scala 136:25]
  wire [38:0] s0_pc_ppm_s2_target_src; // @[PriorityMuxGen.scala 136:25]
  wire  s0_pc_ppm_s1_target_sel; // @[PriorityMuxGen.scala 136:25]
  wire [38:0] s0_pc_ppm_s1_target_src; // @[PriorityMuxGen.scala 136:25]
  wire  s0_pc_ppm_s3_target_sel; // @[PriorityMuxGen.scala 136:25]
  wire [38:0] s0_pc_ppm_s3_target_src; // @[PriorityMuxGen.scala 136:25]
  wire  s0_pc_ppm_redirect_target_sel; // @[PriorityMuxGen.scala 136:25]
  wire [38:0] s0_pc_ppm_redirect_target_src; // @[PriorityMuxGen.scala 136:25]
  wire [38:0] s0_pc_ppm_stallPC_src; // @[PriorityMuxGen.scala 136:25]
  wire [38:0] s0_pc_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  s0_folded_gh_ppm_s2_FGH_sel; // @[PriorityMuxGen.scala 136:25]
  wire [7:0] s0_folded_gh_ppm_s2_FGH_src_hist_17_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [7:0] s0_folded_gh_ppm_s2_FGH_src_hist_16_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [10:0] s0_folded_gh_ppm_s2_FGH_src_hist_15_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [6:0] s0_folded_gh_ppm_s2_FGH_src_hist_14_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [6:0] s0_folded_gh_ppm_s2_FGH_src_hist_13_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [6:0] s0_folded_gh_ppm_s2_FGH_src_hist_12_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [7:0] s0_folded_gh_ppm_s2_FGH_src_hist_11_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [8:0] s0_folded_gh_ppm_s2_FGH_src_hist_10_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [6:0] s0_folded_gh_ppm_s2_FGH_src_hist_9_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [7:0] s0_folded_gh_ppm_s2_FGH_src_hist_8_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [8:0] s0_folded_gh_ppm_s2_FGH_src_hist_7_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [8:0] s0_folded_gh_ppm_s2_FGH_src_hist_6_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [10:0] s0_folded_gh_ppm_s2_FGH_src_hist_5_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [3:0] s0_folded_gh_ppm_s2_FGH_src_hist_4_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [10:0] s0_folded_gh_ppm_s2_FGH_src_hist_3_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [7:0] s0_folded_gh_ppm_s2_FGH_src_hist_2_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [7:0] s0_folded_gh_ppm_s2_FGH_src_hist_1_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [7:0] s0_folded_gh_ppm_s2_FGH_src_hist_0_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire  s0_folded_gh_ppm_s1_FGH_sel; // @[PriorityMuxGen.scala 136:25]
  wire [7:0] s0_folded_gh_ppm_s1_FGH_src_hist_17_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [7:0] s0_folded_gh_ppm_s1_FGH_src_hist_16_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [10:0] s0_folded_gh_ppm_s1_FGH_src_hist_15_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [6:0] s0_folded_gh_ppm_s1_FGH_src_hist_14_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [6:0] s0_folded_gh_ppm_s1_FGH_src_hist_13_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [6:0] s0_folded_gh_ppm_s1_FGH_src_hist_12_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [7:0] s0_folded_gh_ppm_s1_FGH_src_hist_11_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [8:0] s0_folded_gh_ppm_s1_FGH_src_hist_10_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [6:0] s0_folded_gh_ppm_s1_FGH_src_hist_9_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [7:0] s0_folded_gh_ppm_s1_FGH_src_hist_8_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [8:0] s0_folded_gh_ppm_s1_FGH_src_hist_7_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [8:0] s0_folded_gh_ppm_s1_FGH_src_hist_6_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [10:0] s0_folded_gh_ppm_s1_FGH_src_hist_5_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [3:0] s0_folded_gh_ppm_s1_FGH_src_hist_4_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [10:0] s0_folded_gh_ppm_s1_FGH_src_hist_3_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [7:0] s0_folded_gh_ppm_s1_FGH_src_hist_2_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [7:0] s0_folded_gh_ppm_s1_FGH_src_hist_1_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [7:0] s0_folded_gh_ppm_s1_FGH_src_hist_0_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire  s0_folded_gh_ppm_s3_FGH_sel; // @[PriorityMuxGen.scala 136:25]
  wire [7:0] s0_folded_gh_ppm_s3_FGH_src_hist_17_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [7:0] s0_folded_gh_ppm_s3_FGH_src_hist_16_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [10:0] s0_folded_gh_ppm_s3_FGH_src_hist_15_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [6:0] s0_folded_gh_ppm_s3_FGH_src_hist_14_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [6:0] s0_folded_gh_ppm_s3_FGH_src_hist_13_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [6:0] s0_folded_gh_ppm_s3_FGH_src_hist_12_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [7:0] s0_folded_gh_ppm_s3_FGH_src_hist_11_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [8:0] s0_folded_gh_ppm_s3_FGH_src_hist_10_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [6:0] s0_folded_gh_ppm_s3_FGH_src_hist_9_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [7:0] s0_folded_gh_ppm_s3_FGH_src_hist_8_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [8:0] s0_folded_gh_ppm_s3_FGH_src_hist_7_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [8:0] s0_folded_gh_ppm_s3_FGH_src_hist_6_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [10:0] s0_folded_gh_ppm_s3_FGH_src_hist_5_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [3:0] s0_folded_gh_ppm_s3_FGH_src_hist_4_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [10:0] s0_folded_gh_ppm_s3_FGH_src_hist_3_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [7:0] s0_folded_gh_ppm_s3_FGH_src_hist_2_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [7:0] s0_folded_gh_ppm_s3_FGH_src_hist_1_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [7:0] s0_folded_gh_ppm_s3_FGH_src_hist_0_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire  s0_folded_gh_ppm_redirect_FGHT_sel; // @[PriorityMuxGen.scala 136:25]
  wire [7:0] s0_folded_gh_ppm_redirect_FGHT_src_hist_17_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [7:0] s0_folded_gh_ppm_redirect_FGHT_src_hist_16_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [10:0] s0_folded_gh_ppm_redirect_FGHT_src_hist_15_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [6:0] s0_folded_gh_ppm_redirect_FGHT_src_hist_14_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [6:0] s0_folded_gh_ppm_redirect_FGHT_src_hist_13_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [6:0] s0_folded_gh_ppm_redirect_FGHT_src_hist_12_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [7:0] s0_folded_gh_ppm_redirect_FGHT_src_hist_11_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [8:0] s0_folded_gh_ppm_redirect_FGHT_src_hist_10_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [6:0] s0_folded_gh_ppm_redirect_FGHT_src_hist_9_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [7:0] s0_folded_gh_ppm_redirect_FGHT_src_hist_8_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [8:0] s0_folded_gh_ppm_redirect_FGHT_src_hist_7_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [8:0] s0_folded_gh_ppm_redirect_FGHT_src_hist_6_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [10:0] s0_folded_gh_ppm_redirect_FGHT_src_hist_5_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [3:0] s0_folded_gh_ppm_redirect_FGHT_src_hist_4_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [10:0] s0_folded_gh_ppm_redirect_FGHT_src_hist_3_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [7:0] s0_folded_gh_ppm_redirect_FGHT_src_hist_2_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [7:0] s0_folded_gh_ppm_redirect_FGHT_src_hist_1_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [7:0] s0_folded_gh_ppm_redirect_FGHT_src_hist_0_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [7:0] s0_folded_gh_ppm_stallFGH_src_hist_17_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [7:0] s0_folded_gh_ppm_stallFGH_src_hist_16_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [10:0] s0_folded_gh_ppm_stallFGH_src_hist_15_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [6:0] s0_folded_gh_ppm_stallFGH_src_hist_14_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [6:0] s0_folded_gh_ppm_stallFGH_src_hist_13_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [6:0] s0_folded_gh_ppm_stallFGH_src_hist_12_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [7:0] s0_folded_gh_ppm_stallFGH_src_hist_11_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [8:0] s0_folded_gh_ppm_stallFGH_src_hist_10_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [6:0] s0_folded_gh_ppm_stallFGH_src_hist_9_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [7:0] s0_folded_gh_ppm_stallFGH_src_hist_8_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [8:0] s0_folded_gh_ppm_stallFGH_src_hist_7_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [8:0] s0_folded_gh_ppm_stallFGH_src_hist_6_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [10:0] s0_folded_gh_ppm_stallFGH_src_hist_5_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [3:0] s0_folded_gh_ppm_stallFGH_src_hist_4_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [10:0] s0_folded_gh_ppm_stallFGH_src_hist_3_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [7:0] s0_folded_gh_ppm_stallFGH_src_hist_2_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [7:0] s0_folded_gh_ppm_stallFGH_src_hist_1_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [7:0] s0_folded_gh_ppm_stallFGH_src_hist_0_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [7:0] s0_folded_gh_ppm_out_res_hist_17_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [7:0] s0_folded_gh_ppm_out_res_hist_16_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [10:0] s0_folded_gh_ppm_out_res_hist_15_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [6:0] s0_folded_gh_ppm_out_res_hist_14_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [6:0] s0_folded_gh_ppm_out_res_hist_13_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [6:0] s0_folded_gh_ppm_out_res_hist_12_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [7:0] s0_folded_gh_ppm_out_res_hist_11_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [8:0] s0_folded_gh_ppm_out_res_hist_10_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [6:0] s0_folded_gh_ppm_out_res_hist_9_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [7:0] s0_folded_gh_ppm_out_res_hist_8_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [8:0] s0_folded_gh_ppm_out_res_hist_7_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [8:0] s0_folded_gh_ppm_out_res_hist_6_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [10:0] s0_folded_gh_ppm_out_res_hist_5_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [3:0] s0_folded_gh_ppm_out_res_hist_4_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [10:0] s0_folded_gh_ppm_out_res_hist_3_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [7:0] s0_folded_gh_ppm_out_res_hist_2_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [7:0] s0_folded_gh_ppm_out_res_hist_1_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire [7:0] s0_folded_gh_ppm_out_res_hist_0_folded_hist; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ghist_ptr_ppm_s2_GHPtr_sel; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ghist_ptr_ppm_s2_GHPtr_src_flag; // @[PriorityMuxGen.scala 136:25]
  wire [7:0] s0_ghist_ptr_ppm_s2_GHPtr_src_value; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ghist_ptr_ppm_s1_GHPtr_sel; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ghist_ptr_ppm_s1_GHPtr_src_flag; // @[PriorityMuxGen.scala 136:25]
  wire [7:0] s0_ghist_ptr_ppm_s1_GHPtr_src_value; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ghist_ptr_ppm_s3_GHPtr_sel; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ghist_ptr_ppm_s3_GHPtr_src_flag; // @[PriorityMuxGen.scala 136:25]
  wire [7:0] s0_ghist_ptr_ppm_s3_GHPtr_src_value; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ghist_ptr_ppm_redirect_GHPtr_sel; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ghist_ptr_ppm_redirect_GHPtr_src_flag; // @[PriorityMuxGen.scala 136:25]
  wire [7:0] s0_ghist_ptr_ppm_redirect_GHPtr_src_value; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ghist_ptr_ppm_stallGHPtr_src_flag; // @[PriorityMuxGen.scala 136:25]
  wire [7:0] s0_ghist_ptr_ppm_stallGHPtr_src_value; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ghist_ptr_ppm_out_res_flag; // @[PriorityMuxGen.scala 136:25]
  wire [7:0] s0_ghist_ptr_ppm_out_res_value; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_sel; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_src_afhob_5_bits_0; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_src_afhob_5_bits_1; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_src_afhob_5_bits_2; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_src_afhob_5_bits_3; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_src_afhob_4_bits_0; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_src_afhob_4_bits_1; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_src_afhob_4_bits_2; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_src_afhob_4_bits_3; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_src_afhob_3_bits_0; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_src_afhob_3_bits_1; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_src_afhob_3_bits_2; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_src_afhob_3_bits_3; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_src_afhob_2_bits_0; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_src_afhob_2_bits_1; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_src_afhob_2_bits_2; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_src_afhob_2_bits_3; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_src_afhob_1_bits_0; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_src_afhob_1_bits_1; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_src_afhob_1_bits_2; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_src_afhob_1_bits_3; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_src_afhob_0_bits_0; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_src_afhob_0_bits_1; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_src_afhob_0_bits_2; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_src_afhob_0_bits_3; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_sel; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_src_afhob_5_bits_0; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_src_afhob_5_bits_1; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_src_afhob_5_bits_2; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_src_afhob_5_bits_3; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_src_afhob_4_bits_0; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_src_afhob_4_bits_1; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_src_afhob_4_bits_2; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_src_afhob_4_bits_3; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_src_afhob_3_bits_0; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_src_afhob_3_bits_1; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_src_afhob_3_bits_2; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_src_afhob_3_bits_3; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_src_afhob_2_bits_0; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_src_afhob_2_bits_1; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_src_afhob_2_bits_2; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_src_afhob_2_bits_3; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_src_afhob_1_bits_0; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_src_afhob_1_bits_1; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_src_afhob_1_bits_2; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_src_afhob_1_bits_3; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_src_afhob_0_bits_0; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_src_afhob_0_bits_1; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_src_afhob_0_bits_2; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_src_afhob_0_bits_3; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_sel; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_src_afhob_5_bits_0; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_src_afhob_5_bits_1; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_src_afhob_5_bits_2; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_src_afhob_5_bits_3; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_src_afhob_4_bits_0; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_src_afhob_4_bits_1; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_src_afhob_4_bits_2; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_src_afhob_4_bits_3; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_src_afhob_3_bits_0; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_src_afhob_3_bits_1; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_src_afhob_3_bits_2; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_src_afhob_3_bits_3; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_src_afhob_2_bits_0; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_src_afhob_2_bits_1; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_src_afhob_2_bits_2; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_src_afhob_2_bits_3; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_src_afhob_1_bits_0; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_src_afhob_1_bits_1; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_src_afhob_1_bits_2; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_src_afhob_1_bits_3; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_src_afhob_0_bits_0; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_src_afhob_0_bits_1; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_src_afhob_0_bits_2; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_src_afhob_0_bits_3; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_sel; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_src_afhob_5_bits_0; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_src_afhob_5_bits_1; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_src_afhob_5_bits_2; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_src_afhob_5_bits_3; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_src_afhob_4_bits_0; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_src_afhob_4_bits_1; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_src_afhob_4_bits_2; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_src_afhob_4_bits_3; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_src_afhob_3_bits_0; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_src_afhob_3_bits_1; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_src_afhob_3_bits_2; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_src_afhob_3_bits_3; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_src_afhob_2_bits_0; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_src_afhob_2_bits_1; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_src_afhob_2_bits_2; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_src_afhob_2_bits_3; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_src_afhob_1_bits_0; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_src_afhob_1_bits_1; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_src_afhob_1_bits_2; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_src_afhob_1_bits_3; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_src_afhob_0_bits_0; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_src_afhob_0_bits_1; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_src_afhob_0_bits_2; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_src_afhob_0_bits_3; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_stallAFHOB_src_afhob_5_bits_0; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_stallAFHOB_src_afhob_5_bits_1; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_stallAFHOB_src_afhob_5_bits_2; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_stallAFHOB_src_afhob_5_bits_3; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_stallAFHOB_src_afhob_4_bits_0; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_stallAFHOB_src_afhob_4_bits_1; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_stallAFHOB_src_afhob_4_bits_2; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_stallAFHOB_src_afhob_4_bits_3; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_stallAFHOB_src_afhob_3_bits_0; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_stallAFHOB_src_afhob_3_bits_1; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_stallAFHOB_src_afhob_3_bits_2; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_stallAFHOB_src_afhob_3_bits_3; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_stallAFHOB_src_afhob_2_bits_0; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_stallAFHOB_src_afhob_2_bits_1; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_stallAFHOB_src_afhob_2_bits_2; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_stallAFHOB_src_afhob_2_bits_3; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_stallAFHOB_src_afhob_1_bits_0; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_stallAFHOB_src_afhob_1_bits_1; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_stallAFHOB_src_afhob_1_bits_2; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_stallAFHOB_src_afhob_1_bits_3; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_stallAFHOB_src_afhob_0_bits_0; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_stallAFHOB_src_afhob_0_bits_1; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_stallAFHOB_src_afhob_0_bits_2; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_stallAFHOB_src_afhob_0_bits_3; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_out_res_afhob_5_bits_0; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_out_res_afhob_5_bits_1; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_out_res_afhob_5_bits_2; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_out_res_afhob_5_bits_3; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_out_res_afhob_4_bits_0; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_out_res_afhob_4_bits_1; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_out_res_afhob_4_bits_2; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_out_res_afhob_4_bits_3; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_out_res_afhob_3_bits_0; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_out_res_afhob_3_bits_1; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_out_res_afhob_3_bits_2; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_out_res_afhob_3_bits_3; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_out_res_afhob_2_bits_0; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_out_res_afhob_2_bits_1; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_out_res_afhob_2_bits_2; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_out_res_afhob_2_bits_3; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_out_res_afhob_1_bits_0; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_out_res_afhob_1_bits_1; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_out_res_afhob_1_bits_2; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_out_res_afhob_1_bits_3; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_out_res_afhob_0_bits_0; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_out_res_afhob_0_bits_1; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_out_res_afhob_0_bits_2; // @[PriorityMuxGen.scala 136:25]
  wire  s0_ahead_fh_oldest_bits_ppm_out_res_afhob_0_bits_3; // @[PriorityMuxGen.scala 136:25]
  wire  s0_last_br_num_oh_ppm_s2_BrNumOH_sel; // @[PriorityMuxGen.scala 136:25]
  wire [2:0] s0_last_br_num_oh_ppm_s2_BrNumOH_src; // @[PriorityMuxGen.scala 136:25]
  wire  s0_last_br_num_oh_ppm_s1_BrNumOH_sel; // @[PriorityMuxGen.scala 136:25]
  wire [2:0] s0_last_br_num_oh_ppm_s1_BrNumOH_src; // @[PriorityMuxGen.scala 136:25]
  wire  s0_last_br_num_oh_ppm_s3_BrNumOH_sel; // @[PriorityMuxGen.scala 136:25]
  wire [2:0] s0_last_br_num_oh_ppm_s3_BrNumOH_src; // @[PriorityMuxGen.scala 136:25]
  wire  s0_last_br_num_oh_ppm_redirect_BrNumOH_sel; // @[PriorityMuxGen.scala 136:25]
  wire [2:0] s0_last_br_num_oh_ppm_redirect_BrNumOH_src; // @[PriorityMuxGen.scala 136:25]
  wire [2:0] s0_last_br_num_oh_ppm_stallBrNumOH_src; // @[PriorityMuxGen.scala 136:25]
  wire [2:0] s0_last_br_num_oh_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_0_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_0_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_0_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_0_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_0_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_0_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_0_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_0_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_1_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_1_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_1_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_1_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_1_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_1_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_1_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_1_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_2_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_2_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_2_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_2_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_2_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_2_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_2_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_2_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_3_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_3_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_3_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_3_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_3_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_3_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_3_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_3_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_4_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_4_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_4_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_4_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_4_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_4_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_4_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_4_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_5_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_5_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_5_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_5_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_5_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_5_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_5_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_5_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_6_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_6_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_6_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_6_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_6_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_6_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_6_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_6_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_7_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_7_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_7_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_7_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_7_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_7_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_7_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_7_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_8_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_8_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_8_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_8_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_8_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_8_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_8_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_8_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_9_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_9_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_9_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_9_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_9_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_9_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_9_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_9_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_10_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_10_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_10_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_10_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_10_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_10_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_10_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_10_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_11_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_11_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_11_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_11_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_11_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_11_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_11_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_11_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_12_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_12_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_12_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_12_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_12_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_12_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_12_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_12_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_13_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_13_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_13_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_13_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_13_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_13_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_13_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_13_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_14_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_14_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_14_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_14_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_14_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_14_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_14_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_14_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_15_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_15_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_15_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_15_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_15_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_15_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_15_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_15_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_16_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_16_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_16_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_16_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_16_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_16_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_16_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_16_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_17_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_17_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_17_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_17_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_17_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_17_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_17_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_17_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_18_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_18_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_18_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_18_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_18_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_18_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_18_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_18_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_19_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_19_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_19_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_19_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_19_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_19_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_19_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_19_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_20_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_20_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_20_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_20_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_20_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_20_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_20_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_20_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_21_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_21_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_21_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_21_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_21_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_21_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_21_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_21_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_22_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_22_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_22_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_22_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_22_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_22_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_22_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_22_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_23_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_23_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_23_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_23_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_23_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_23_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_23_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_23_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_24_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_24_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_24_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_24_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_24_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_24_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_24_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_24_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_25_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_25_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_25_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_25_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_25_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_25_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_25_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_25_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_26_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_26_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_26_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_26_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_26_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_26_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_26_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_26_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_27_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_27_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_27_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_27_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_27_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_27_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_27_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_27_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_28_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_28_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_28_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_28_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_28_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_28_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_28_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_28_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_29_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_29_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_29_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_29_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_29_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_29_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_29_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_29_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_30_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_30_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_30_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_30_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_30_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_30_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_30_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_30_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_31_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_31_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_31_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_31_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_31_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_31_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_31_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_31_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_32_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_32_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_32_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_32_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_32_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_32_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_32_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_32_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_33_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_33_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_33_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_33_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_33_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_33_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_33_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_33_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_34_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_34_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_34_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_34_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_34_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_34_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_34_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_34_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_35_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_35_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_35_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_35_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_35_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_35_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_35_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_35_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_36_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_36_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_36_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_36_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_36_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_36_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_36_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_36_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_37_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_37_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_37_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_37_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_37_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_37_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_37_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_37_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_38_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_38_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_38_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_38_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_38_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_38_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_38_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_38_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_39_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_39_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_39_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_39_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_39_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_39_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_39_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_39_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_40_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_40_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_40_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_40_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_40_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_40_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_40_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_40_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_41_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_41_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_41_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_41_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_41_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_41_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_41_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_41_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_42_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_42_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_42_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_42_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_42_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_42_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_42_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_42_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_43_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_43_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_43_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_43_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_43_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_43_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_43_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_43_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_44_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_44_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_44_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_44_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_44_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_44_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_44_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_44_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_45_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_45_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_45_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_45_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_45_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_45_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_45_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_45_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_46_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_46_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_46_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_46_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_46_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_46_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_46_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_46_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_47_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_47_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_47_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_47_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_47_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_47_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_47_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_47_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_48_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_48_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_48_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_48_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_48_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_48_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_48_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_48_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_49_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_49_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_49_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_49_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_49_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_49_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_49_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_49_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_50_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_50_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_50_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_50_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_50_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_50_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_50_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_50_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_51_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_51_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_51_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_51_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_51_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_51_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_51_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_51_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_52_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_52_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_52_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_52_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_52_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_52_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_52_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_52_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_53_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_53_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_53_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_53_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_53_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_53_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_53_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_53_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_54_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_54_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_54_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_54_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_54_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_54_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_54_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_54_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_55_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_55_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_55_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_55_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_55_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_55_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_55_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_55_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_56_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_56_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_56_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_56_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_56_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_56_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_56_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_56_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_57_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_57_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_57_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_57_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_57_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_57_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_57_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_57_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_58_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_58_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_58_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_58_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_58_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_58_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_58_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_58_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_59_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_59_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_59_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_59_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_59_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_59_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_59_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_59_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_60_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_60_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_60_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_60_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_60_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_60_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_60_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_60_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_61_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_61_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_61_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_61_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_61_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_61_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_61_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_61_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_62_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_62_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_62_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_62_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_62_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_62_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_62_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_62_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_63_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_63_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_63_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_63_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_63_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_63_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_63_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_63_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_64_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_64_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_64_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_64_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_64_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_64_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_64_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_64_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_65_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_65_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_65_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_65_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_65_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_65_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_65_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_65_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_66_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_66_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_66_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_66_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_66_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_66_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_66_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_66_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_67_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_67_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_67_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_67_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_67_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_67_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_67_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_67_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_68_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_68_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_68_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_68_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_68_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_68_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_68_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_68_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_69_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_69_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_69_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_69_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_69_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_69_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_69_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_69_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_70_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_70_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_70_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_70_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_70_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_70_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_70_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_70_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_71_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_71_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_71_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_71_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_71_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_71_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_71_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_71_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_72_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_72_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_72_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_72_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_72_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_72_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_72_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_72_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_73_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_73_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_73_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_73_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_73_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_73_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_73_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_73_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_74_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_74_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_74_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_74_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_74_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_74_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_74_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_74_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_75_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_75_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_75_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_75_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_75_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_75_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_75_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_75_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_76_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_76_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_76_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_76_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_76_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_76_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_76_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_76_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_77_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_77_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_77_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_77_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_77_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_77_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_77_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_77_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_78_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_78_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_78_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_78_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_78_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_78_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_78_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_78_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_79_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_79_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_79_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_79_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_79_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_79_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_79_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_79_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_80_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_80_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_80_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_80_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_80_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_80_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_80_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_80_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_81_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_81_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_81_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_81_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_81_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_81_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_81_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_81_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_82_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_82_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_82_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_82_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_82_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_82_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_82_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_82_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_83_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_83_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_83_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_83_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_83_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_83_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_83_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_83_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_84_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_84_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_84_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_84_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_84_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_84_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_84_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_84_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_85_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_85_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_85_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_85_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_85_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_85_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_85_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_85_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_86_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_86_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_86_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_86_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_86_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_86_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_86_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_86_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_87_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_87_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_87_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_87_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_87_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_87_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_87_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_87_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_88_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_88_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_88_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_88_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_88_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_88_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_88_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_88_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_89_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_89_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_89_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_89_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_89_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_89_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_89_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_89_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_90_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_90_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_90_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_90_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_90_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_90_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_90_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_90_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_91_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_91_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_91_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_91_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_91_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_91_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_91_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_91_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_92_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_92_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_92_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_92_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_92_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_92_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_92_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_92_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_93_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_93_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_93_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_93_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_93_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_93_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_93_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_93_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_94_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_94_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_94_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_94_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_94_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_94_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_94_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_94_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_95_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_95_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_95_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_95_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_95_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_95_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_95_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_95_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_96_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_96_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_96_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_96_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_96_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_96_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_96_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_96_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_97_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_97_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_97_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_97_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_97_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_97_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_97_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_97_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_98_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_98_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_98_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_98_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_98_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_98_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_98_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_98_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_99_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_99_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_99_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_99_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_99_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_99_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_99_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_99_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_100_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_100_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_100_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_100_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_100_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_100_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_100_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_100_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_101_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_101_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_101_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_101_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_101_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_101_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_101_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_101_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_102_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_102_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_102_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_102_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_102_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_102_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_102_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_102_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_103_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_103_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_103_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_103_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_103_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_103_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_103_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_103_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_104_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_104_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_104_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_104_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_104_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_104_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_104_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_104_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_105_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_105_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_105_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_105_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_105_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_105_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_105_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_105_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_106_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_106_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_106_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_106_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_106_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_106_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_106_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_106_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_107_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_107_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_107_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_107_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_107_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_107_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_107_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_107_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_108_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_108_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_108_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_108_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_108_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_108_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_108_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_108_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_109_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_109_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_109_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_109_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_109_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_109_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_109_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_109_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_110_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_110_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_110_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_110_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_110_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_110_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_110_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_110_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_111_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_111_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_111_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_111_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_111_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_111_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_111_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_111_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_112_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_112_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_112_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_112_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_112_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_112_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_112_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_112_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_113_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_113_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_113_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_113_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_113_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_113_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_113_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_113_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_114_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_114_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_114_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_114_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_114_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_114_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_114_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_114_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_115_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_115_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_115_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_115_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_115_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_115_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_115_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_115_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_116_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_116_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_116_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_116_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_116_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_116_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_116_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_116_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_117_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_117_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_117_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_117_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_117_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_117_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_117_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_117_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_118_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_118_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_118_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_118_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_118_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_118_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_118_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_118_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_119_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_119_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_119_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_119_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_119_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_119_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_119_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_119_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_120_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_120_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_120_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_120_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_120_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_120_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_120_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_120_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_121_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_121_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_121_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_121_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_121_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_121_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_121_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_121_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_122_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_122_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_122_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_122_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_122_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_122_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_122_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_122_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_123_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_123_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_123_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_123_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_123_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_123_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_123_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_123_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_124_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_124_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_124_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_124_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_124_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_124_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_124_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_124_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_125_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_125_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_125_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_125_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_125_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_125_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_125_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_125_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_126_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_126_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_126_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_126_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_126_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_126_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_126_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_126_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_127_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_127_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_127_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_127_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_127_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_127_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_127_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_127_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_128_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_128_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_128_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_128_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_128_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_128_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_128_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_128_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_129_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_129_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_129_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_129_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_129_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_129_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_129_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_129_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_130_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_130_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_130_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_130_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_130_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_130_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_130_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_130_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_131_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_131_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_131_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_131_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_131_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_131_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_131_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_131_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_132_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_132_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_132_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_132_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_132_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_132_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_132_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_132_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_133_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_133_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_133_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_133_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_133_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_133_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_133_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_133_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_134_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_134_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_134_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_134_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_134_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_134_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_134_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_134_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_135_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_135_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_135_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_135_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_135_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_135_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_135_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_135_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_136_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_136_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_136_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_136_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_136_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_136_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_136_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_136_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_137_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_137_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_137_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_137_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_137_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_137_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_137_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_137_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_138_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_138_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_138_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_138_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_138_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_138_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_138_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_138_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_139_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_139_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_139_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_139_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_139_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_139_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_139_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_139_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_140_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_140_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_140_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_140_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_140_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_140_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_140_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_140_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_141_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_141_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_141_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_141_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_141_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_141_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_141_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_141_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_142_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_142_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_142_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_142_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_142_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_142_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_142_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_142_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_143_ppm_s2_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_143_ppm_s2_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_143_ppm_s1_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_143_ppm_s1_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_143_ppm_s3_new_bit_0_sel; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_143_ppm_s3_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_143_ppm_redirect_new_bit_0_src; // @[PriorityMuxGen.scala 136:25]
  wire  ghv_write_datas_143_ppm_out_res; // @[PriorityMuxGen.scala 136:25]
  reg  s1_valid; // @[BPU.scala 252:45]
  reg  s2_valid; // @[BPU.scala 252:45]
  reg  s3_valid; // @[BPU.scala 252:45]
  reg [38:0] s0_pc_reg; // @[BPU.scala 258:26]
  reg  REG; // @[BPU.scala 259:24]
  reg  REG_1; // @[BPU.scala 259:16]
  wire [38:0] s0_pc = s0_pc_ppm_out_res; // @[BPU.scala 257:19 667:17]
  wire  s1_components_ready = predictors_io_s1_ready; // @[BPU.scala 254:75 342:23]
  wire  s2_ready = s2_valid | ~s2_valid; // @[BPU.scala 348:23]
  wire  _s1_fire_T_1 = s1_valid & s2_ready; // @[BPU.scala 349:46]
  wire  s1_fire = s1_valid & s2_ready & io_bpu_to_ftq_resp_ready; // @[BPU.scala 349:58]
  wire  s1_ready = s1_fire | ~s1_valid; // @[BPU.scala 343:23]
  wire  s0_fire = s1_components_ready & s1_ready; // @[BPU.scala 344:34]
  reg [7:0] s0_folded_gh_reg_hist_17_folded_hist; // @[BPU.scala 267:33]
  reg [7:0] s0_folded_gh_reg_hist_16_folded_hist; // @[BPU.scala 267:33]
  reg [10:0] s0_folded_gh_reg_hist_15_folded_hist; // @[BPU.scala 267:33]
  reg [6:0] s0_folded_gh_reg_hist_14_folded_hist; // @[BPU.scala 267:33]
  reg [6:0] s0_folded_gh_reg_hist_13_folded_hist; // @[BPU.scala 267:33]
  reg [6:0] s0_folded_gh_reg_hist_12_folded_hist; // @[BPU.scala 267:33]
  reg [7:0] s0_folded_gh_reg_hist_11_folded_hist; // @[BPU.scala 267:33]
  reg [8:0] s0_folded_gh_reg_hist_10_folded_hist; // @[BPU.scala 267:33]
  reg [6:0] s0_folded_gh_reg_hist_9_folded_hist; // @[BPU.scala 267:33]
  reg [7:0] s0_folded_gh_reg_hist_8_folded_hist; // @[BPU.scala 267:33]
  reg [8:0] s0_folded_gh_reg_hist_7_folded_hist; // @[BPU.scala 267:33]
  reg [8:0] s0_folded_gh_reg_hist_6_folded_hist; // @[BPU.scala 267:33]
  reg [10:0] s0_folded_gh_reg_hist_5_folded_hist; // @[BPU.scala 267:33]
  reg [3:0] s0_folded_gh_reg_hist_4_folded_hist; // @[BPU.scala 267:33]
  reg [10:0] s0_folded_gh_reg_hist_3_folded_hist; // @[BPU.scala 267:33]
  reg [7:0] s0_folded_gh_reg_hist_2_folded_hist; // @[BPU.scala 267:33]
  reg [7:0] s0_folded_gh_reg_hist_1_folded_hist; // @[BPU.scala 267:33]
  reg [7:0] s0_folded_gh_reg_hist_0_folded_hist; // @[BPU.scala 267:33]
  reg [7:0] s1_folded_gh_hist_17_folded_hist; // @[Reg.scala 28:20]
  reg [7:0] s1_folded_gh_hist_16_folded_hist; // @[Reg.scala 28:20]
  reg [10:0] s1_folded_gh_hist_15_folded_hist; // @[Reg.scala 28:20]
  reg [6:0] s1_folded_gh_hist_14_folded_hist; // @[Reg.scala 28:20]
  reg [6:0] s1_folded_gh_hist_13_folded_hist; // @[Reg.scala 28:20]
  reg [6:0] s1_folded_gh_hist_12_folded_hist; // @[Reg.scala 28:20]
  reg [7:0] s1_folded_gh_hist_11_folded_hist; // @[Reg.scala 28:20]
  reg [8:0] s1_folded_gh_hist_10_folded_hist; // @[Reg.scala 28:20]
  reg [6:0] s1_folded_gh_hist_9_folded_hist; // @[Reg.scala 28:20]
  reg [7:0] s1_folded_gh_hist_8_folded_hist; // @[Reg.scala 28:20]
  reg [8:0] s1_folded_gh_hist_7_folded_hist; // @[Reg.scala 28:20]
  reg [8:0] s1_folded_gh_hist_6_folded_hist; // @[Reg.scala 28:20]
  reg [10:0] s1_folded_gh_hist_5_folded_hist; // @[Reg.scala 28:20]
  reg [3:0] s1_folded_gh_hist_4_folded_hist; // @[Reg.scala 28:20]
  reg [10:0] s1_folded_gh_hist_3_folded_hist; // @[Reg.scala 28:20]
  reg [7:0] s1_folded_gh_hist_2_folded_hist; // @[Reg.scala 28:20]
  reg [7:0] s1_folded_gh_hist_1_folded_hist; // @[Reg.scala 28:20]
  reg [7:0] s1_folded_gh_hist_0_folded_hist; // @[Reg.scala 28:20]
  wire [7:0] s0_folded_gh_hist_17_folded_hist = s0_folded_gh_ppm_out_res_hist_17_folded_hist; // @[BPU.scala 266:26 668:17]
  wire [7:0] s0_folded_gh_hist_16_folded_hist = s0_folded_gh_ppm_out_res_hist_16_folded_hist; // @[BPU.scala 266:26 668:17]
  wire [10:0] s0_folded_gh_hist_15_folded_hist = s0_folded_gh_ppm_out_res_hist_15_folded_hist; // @[BPU.scala 266:26 668:17]
  wire [6:0] s0_folded_gh_hist_14_folded_hist = s0_folded_gh_ppm_out_res_hist_14_folded_hist; // @[BPU.scala 266:26 668:17]
  wire [6:0] s0_folded_gh_hist_13_folded_hist = s0_folded_gh_ppm_out_res_hist_13_folded_hist; // @[BPU.scala 266:26 668:17]
  wire [6:0] s0_folded_gh_hist_12_folded_hist = s0_folded_gh_ppm_out_res_hist_12_folded_hist; // @[BPU.scala 266:26 668:17]
  wire [7:0] s0_folded_gh_hist_11_folded_hist = s0_folded_gh_ppm_out_res_hist_11_folded_hist; // @[BPU.scala 266:26 668:17]
  wire [8:0] s0_folded_gh_hist_10_folded_hist = s0_folded_gh_ppm_out_res_hist_10_folded_hist; // @[BPU.scala 266:26 668:17]
  wire [6:0] s0_folded_gh_hist_9_folded_hist = s0_folded_gh_ppm_out_res_hist_9_folded_hist; // @[BPU.scala 266:26 668:17]
  wire [7:0] s0_folded_gh_hist_8_folded_hist = s0_folded_gh_ppm_out_res_hist_8_folded_hist; // @[BPU.scala 266:26 668:17]
  wire [8:0] s0_folded_gh_hist_7_folded_hist = s0_folded_gh_ppm_out_res_hist_7_folded_hist; // @[BPU.scala 266:26 668:17]
  wire [8:0] s0_folded_gh_hist_6_folded_hist = s0_folded_gh_ppm_out_res_hist_6_folded_hist; // @[BPU.scala 266:26 668:17]
  wire [10:0] s0_folded_gh_hist_5_folded_hist = s0_folded_gh_ppm_out_res_hist_5_folded_hist; // @[BPU.scala 266:26 668:17]
  wire [3:0] s0_folded_gh_hist_4_folded_hist = s0_folded_gh_ppm_out_res_hist_4_folded_hist; // @[BPU.scala 266:26 668:17]
  wire [10:0] s0_folded_gh_hist_3_folded_hist = s0_folded_gh_ppm_out_res_hist_3_folded_hist; // @[BPU.scala 266:26 668:17]
  wire [7:0] s0_folded_gh_hist_2_folded_hist = s0_folded_gh_ppm_out_res_hist_2_folded_hist; // @[BPU.scala 266:26 668:17]
  wire [7:0] s0_folded_gh_hist_1_folded_hist = s0_folded_gh_ppm_out_res_hist_1_folded_hist; // @[BPU.scala 266:26 668:17]
  wire [7:0] s0_folded_gh_hist_0_folded_hist = s0_folded_gh_ppm_out_res_hist_0_folded_hist; // @[BPU.scala 266:26 668:17]
  reg [7:0] s2_folded_gh_hist_17_folded_hist; // @[Reg.scala 28:20]
  reg [7:0] s2_folded_gh_hist_16_folded_hist; // @[Reg.scala 28:20]
  reg [10:0] s2_folded_gh_hist_15_folded_hist; // @[Reg.scala 28:20]
  reg [6:0] s2_folded_gh_hist_14_folded_hist; // @[Reg.scala 28:20]
  reg [6:0] s2_folded_gh_hist_13_folded_hist; // @[Reg.scala 28:20]
  reg [6:0] s2_folded_gh_hist_12_folded_hist; // @[Reg.scala 28:20]
  reg [7:0] s2_folded_gh_hist_11_folded_hist; // @[Reg.scala 28:20]
  reg [8:0] s2_folded_gh_hist_10_folded_hist; // @[Reg.scala 28:20]
  reg [6:0] s2_folded_gh_hist_9_folded_hist; // @[Reg.scala 28:20]
  reg [7:0] s2_folded_gh_hist_8_folded_hist; // @[Reg.scala 28:20]
  reg [8:0] s2_folded_gh_hist_7_folded_hist; // @[Reg.scala 28:20]
  reg [8:0] s2_folded_gh_hist_6_folded_hist; // @[Reg.scala 28:20]
  reg [10:0] s2_folded_gh_hist_5_folded_hist; // @[Reg.scala 28:20]
  reg [3:0] s2_folded_gh_hist_4_folded_hist; // @[Reg.scala 28:20]
  reg [10:0] s2_folded_gh_hist_3_folded_hist; // @[Reg.scala 28:20]
  reg [7:0] s2_folded_gh_hist_2_folded_hist; // @[Reg.scala 28:20]
  reg [7:0] s2_folded_gh_hist_1_folded_hist; // @[Reg.scala 28:20]
  reg [7:0] s2_folded_gh_hist_0_folded_hist; // @[Reg.scala 28:20]
  reg [7:0] s3_folded_gh_hist_17_folded_hist; // @[Reg.scala 28:20]
  reg [7:0] s3_folded_gh_hist_16_folded_hist; // @[Reg.scala 28:20]
  reg [10:0] s3_folded_gh_hist_15_folded_hist; // @[Reg.scala 28:20]
  reg [6:0] s3_folded_gh_hist_14_folded_hist; // @[Reg.scala 28:20]
  reg [6:0] s3_folded_gh_hist_13_folded_hist; // @[Reg.scala 28:20]
  reg [6:0] s3_folded_gh_hist_12_folded_hist; // @[Reg.scala 28:20]
  reg [7:0] s3_folded_gh_hist_11_folded_hist; // @[Reg.scala 28:20]
  reg [8:0] s3_folded_gh_hist_10_folded_hist; // @[Reg.scala 28:20]
  reg [6:0] s3_folded_gh_hist_9_folded_hist; // @[Reg.scala 28:20]
  reg [7:0] s3_folded_gh_hist_8_folded_hist; // @[Reg.scala 28:20]
  reg [8:0] s3_folded_gh_hist_7_folded_hist; // @[Reg.scala 28:20]
  reg [8:0] s3_folded_gh_hist_6_folded_hist; // @[Reg.scala 28:20]
  reg [10:0] s3_folded_gh_hist_5_folded_hist; // @[Reg.scala 28:20]
  reg [3:0] s3_folded_gh_hist_4_folded_hist; // @[Reg.scala 28:20]
  reg [10:0] s3_folded_gh_hist_3_folded_hist; // @[Reg.scala 28:20]
  reg [7:0] s3_folded_gh_hist_2_folded_hist; // @[Reg.scala 28:20]
  reg [7:0] s3_folded_gh_hist_1_folded_hist; // @[Reg.scala 28:20]
  reg [7:0] s3_folded_gh_hist_0_folded_hist; // @[Reg.scala 28:20]
  reg [2:0] s0_last_br_num_oh_reg; // @[BPU.scala 273:38]
  reg [2:0] s1_last_br_num_oh; // @[Reg.scala 28:20]
  wire [2:0] s0_last_br_num_oh = s0_last_br_num_oh_ppm_out_res; // @[BPU.scala 272:31 671:21]
  reg [2:0] s2_last_br_num_oh; // @[Reg.scala 28:20]
  reg [2:0] s3_last_br_num_oh; // @[Reg.scala 28:20]
  reg  s0_ahead_fh_oldest_bits_reg_afhob_5_bits_0; // @[BPU.scala 279:44]
  reg  s0_ahead_fh_oldest_bits_reg_afhob_5_bits_1; // @[BPU.scala 279:44]
  reg  s0_ahead_fh_oldest_bits_reg_afhob_5_bits_2; // @[BPU.scala 279:44]
  reg  s0_ahead_fh_oldest_bits_reg_afhob_5_bits_3; // @[BPU.scala 279:44]
  reg  s0_ahead_fh_oldest_bits_reg_afhob_4_bits_0; // @[BPU.scala 279:44]
  reg  s0_ahead_fh_oldest_bits_reg_afhob_4_bits_1; // @[BPU.scala 279:44]
  reg  s0_ahead_fh_oldest_bits_reg_afhob_4_bits_2; // @[BPU.scala 279:44]
  reg  s0_ahead_fh_oldest_bits_reg_afhob_4_bits_3; // @[BPU.scala 279:44]
  reg  s0_ahead_fh_oldest_bits_reg_afhob_3_bits_0; // @[BPU.scala 279:44]
  reg  s0_ahead_fh_oldest_bits_reg_afhob_3_bits_1; // @[BPU.scala 279:44]
  reg  s0_ahead_fh_oldest_bits_reg_afhob_3_bits_2; // @[BPU.scala 279:44]
  reg  s0_ahead_fh_oldest_bits_reg_afhob_3_bits_3; // @[BPU.scala 279:44]
  reg  s0_ahead_fh_oldest_bits_reg_afhob_2_bits_0; // @[BPU.scala 279:44]
  reg  s0_ahead_fh_oldest_bits_reg_afhob_2_bits_1; // @[BPU.scala 279:44]
  reg  s0_ahead_fh_oldest_bits_reg_afhob_2_bits_2; // @[BPU.scala 279:44]
  reg  s0_ahead_fh_oldest_bits_reg_afhob_2_bits_3; // @[BPU.scala 279:44]
  reg  s0_ahead_fh_oldest_bits_reg_afhob_1_bits_0; // @[BPU.scala 279:44]
  reg  s0_ahead_fh_oldest_bits_reg_afhob_1_bits_1; // @[BPU.scala 279:44]
  reg  s0_ahead_fh_oldest_bits_reg_afhob_1_bits_2; // @[BPU.scala 279:44]
  reg  s0_ahead_fh_oldest_bits_reg_afhob_1_bits_3; // @[BPU.scala 279:44]
  reg  s0_ahead_fh_oldest_bits_reg_afhob_0_bits_0; // @[BPU.scala 279:44]
  reg  s0_ahead_fh_oldest_bits_reg_afhob_0_bits_1; // @[BPU.scala 279:44]
  reg  s0_ahead_fh_oldest_bits_reg_afhob_0_bits_2; // @[BPU.scala 279:44]
  reg  s0_ahead_fh_oldest_bits_reg_afhob_0_bits_3; // @[BPU.scala 279:44]
  reg  s1_ahead_fh_oldest_bits_afhob_5_bits_0; // @[Reg.scala 28:20]
  reg  s1_ahead_fh_oldest_bits_afhob_5_bits_1; // @[Reg.scala 28:20]
  reg  s1_ahead_fh_oldest_bits_afhob_5_bits_2; // @[Reg.scala 28:20]
  reg  s1_ahead_fh_oldest_bits_afhob_5_bits_3; // @[Reg.scala 28:20]
  reg  s1_ahead_fh_oldest_bits_afhob_4_bits_0; // @[Reg.scala 28:20]
  reg  s1_ahead_fh_oldest_bits_afhob_4_bits_1; // @[Reg.scala 28:20]
  reg  s1_ahead_fh_oldest_bits_afhob_4_bits_2; // @[Reg.scala 28:20]
  reg  s1_ahead_fh_oldest_bits_afhob_4_bits_3; // @[Reg.scala 28:20]
  reg  s1_ahead_fh_oldest_bits_afhob_3_bits_0; // @[Reg.scala 28:20]
  reg  s1_ahead_fh_oldest_bits_afhob_3_bits_1; // @[Reg.scala 28:20]
  reg  s1_ahead_fh_oldest_bits_afhob_3_bits_2; // @[Reg.scala 28:20]
  reg  s1_ahead_fh_oldest_bits_afhob_3_bits_3; // @[Reg.scala 28:20]
  reg  s1_ahead_fh_oldest_bits_afhob_2_bits_0; // @[Reg.scala 28:20]
  reg  s1_ahead_fh_oldest_bits_afhob_2_bits_1; // @[Reg.scala 28:20]
  reg  s1_ahead_fh_oldest_bits_afhob_2_bits_2; // @[Reg.scala 28:20]
  reg  s1_ahead_fh_oldest_bits_afhob_2_bits_3; // @[Reg.scala 28:20]
  reg  s1_ahead_fh_oldest_bits_afhob_1_bits_0; // @[Reg.scala 28:20]
  reg  s1_ahead_fh_oldest_bits_afhob_1_bits_1; // @[Reg.scala 28:20]
  reg  s1_ahead_fh_oldest_bits_afhob_1_bits_2; // @[Reg.scala 28:20]
  reg  s1_ahead_fh_oldest_bits_afhob_1_bits_3; // @[Reg.scala 28:20]
  reg  s1_ahead_fh_oldest_bits_afhob_0_bits_0; // @[Reg.scala 28:20]
  reg  s1_ahead_fh_oldest_bits_afhob_0_bits_1; // @[Reg.scala 28:20]
  reg  s1_ahead_fh_oldest_bits_afhob_0_bits_2; // @[Reg.scala 28:20]
  reg  s1_ahead_fh_oldest_bits_afhob_0_bits_3; // @[Reg.scala 28:20]
  wire  s0_ahead_fh_oldest_bits_afhob_5_bits_0 = s0_ahead_fh_oldest_bits_ppm_out_res_afhob_5_bits_0; // @[BPU.scala 278:37 670:27]
  wire  s0_ahead_fh_oldest_bits_afhob_5_bits_1 = s0_ahead_fh_oldest_bits_ppm_out_res_afhob_5_bits_1; // @[BPU.scala 278:37 670:27]
  wire  s0_ahead_fh_oldest_bits_afhob_5_bits_2 = s0_ahead_fh_oldest_bits_ppm_out_res_afhob_5_bits_2; // @[BPU.scala 278:37 670:27]
  wire  s0_ahead_fh_oldest_bits_afhob_5_bits_3 = s0_ahead_fh_oldest_bits_ppm_out_res_afhob_5_bits_3; // @[BPU.scala 278:37 670:27]
  wire  s0_ahead_fh_oldest_bits_afhob_4_bits_0 = s0_ahead_fh_oldest_bits_ppm_out_res_afhob_4_bits_0; // @[BPU.scala 278:37 670:27]
  wire  s0_ahead_fh_oldest_bits_afhob_4_bits_1 = s0_ahead_fh_oldest_bits_ppm_out_res_afhob_4_bits_1; // @[BPU.scala 278:37 670:27]
  wire  s0_ahead_fh_oldest_bits_afhob_4_bits_2 = s0_ahead_fh_oldest_bits_ppm_out_res_afhob_4_bits_2; // @[BPU.scala 278:37 670:27]
  wire  s0_ahead_fh_oldest_bits_afhob_4_bits_3 = s0_ahead_fh_oldest_bits_ppm_out_res_afhob_4_bits_3; // @[BPU.scala 278:37 670:27]
  wire  s0_ahead_fh_oldest_bits_afhob_3_bits_0 = s0_ahead_fh_oldest_bits_ppm_out_res_afhob_3_bits_0; // @[BPU.scala 278:37 670:27]
  wire  s0_ahead_fh_oldest_bits_afhob_3_bits_1 = s0_ahead_fh_oldest_bits_ppm_out_res_afhob_3_bits_1; // @[BPU.scala 278:37 670:27]
  wire  s0_ahead_fh_oldest_bits_afhob_3_bits_2 = s0_ahead_fh_oldest_bits_ppm_out_res_afhob_3_bits_2; // @[BPU.scala 278:37 670:27]
  wire  s0_ahead_fh_oldest_bits_afhob_3_bits_3 = s0_ahead_fh_oldest_bits_ppm_out_res_afhob_3_bits_3; // @[BPU.scala 278:37 670:27]
  wire  s0_ahead_fh_oldest_bits_afhob_2_bits_0 = s0_ahead_fh_oldest_bits_ppm_out_res_afhob_2_bits_0; // @[BPU.scala 278:37 670:27]
  wire  s0_ahead_fh_oldest_bits_afhob_2_bits_1 = s0_ahead_fh_oldest_bits_ppm_out_res_afhob_2_bits_1; // @[BPU.scala 278:37 670:27]
  wire  s0_ahead_fh_oldest_bits_afhob_2_bits_2 = s0_ahead_fh_oldest_bits_ppm_out_res_afhob_2_bits_2; // @[BPU.scala 278:37 670:27]
  wire  s0_ahead_fh_oldest_bits_afhob_2_bits_3 = s0_ahead_fh_oldest_bits_ppm_out_res_afhob_2_bits_3; // @[BPU.scala 278:37 670:27]
  wire  s0_ahead_fh_oldest_bits_afhob_1_bits_0 = s0_ahead_fh_oldest_bits_ppm_out_res_afhob_1_bits_0; // @[BPU.scala 278:37 670:27]
  wire  s0_ahead_fh_oldest_bits_afhob_1_bits_1 = s0_ahead_fh_oldest_bits_ppm_out_res_afhob_1_bits_1; // @[BPU.scala 278:37 670:27]
  wire  s0_ahead_fh_oldest_bits_afhob_1_bits_2 = s0_ahead_fh_oldest_bits_ppm_out_res_afhob_1_bits_2; // @[BPU.scala 278:37 670:27]
  wire  s0_ahead_fh_oldest_bits_afhob_1_bits_3 = s0_ahead_fh_oldest_bits_ppm_out_res_afhob_1_bits_3; // @[BPU.scala 278:37 670:27]
  wire  s0_ahead_fh_oldest_bits_afhob_0_bits_0 = s0_ahead_fh_oldest_bits_ppm_out_res_afhob_0_bits_0; // @[BPU.scala 278:37 670:27]
  wire  s0_ahead_fh_oldest_bits_afhob_0_bits_1 = s0_ahead_fh_oldest_bits_ppm_out_res_afhob_0_bits_1; // @[BPU.scala 278:37 670:27]
  wire  s0_ahead_fh_oldest_bits_afhob_0_bits_2 = s0_ahead_fh_oldest_bits_ppm_out_res_afhob_0_bits_2; // @[BPU.scala 278:37 670:27]
  wire  s0_ahead_fh_oldest_bits_afhob_0_bits_3 = s0_ahead_fh_oldest_bits_ppm_out_res_afhob_0_bits_3; // @[BPU.scala 278:37 670:27]
  reg  s2_ahead_fh_oldest_bits_afhob_5_bits_0; // @[Reg.scala 28:20]
  reg  s2_ahead_fh_oldest_bits_afhob_5_bits_1; // @[Reg.scala 28:20]
  reg  s2_ahead_fh_oldest_bits_afhob_5_bits_2; // @[Reg.scala 28:20]
  reg  s2_ahead_fh_oldest_bits_afhob_5_bits_3; // @[Reg.scala 28:20]
  reg  s2_ahead_fh_oldest_bits_afhob_4_bits_0; // @[Reg.scala 28:20]
  reg  s2_ahead_fh_oldest_bits_afhob_4_bits_1; // @[Reg.scala 28:20]
  reg  s2_ahead_fh_oldest_bits_afhob_4_bits_2; // @[Reg.scala 28:20]
  reg  s2_ahead_fh_oldest_bits_afhob_4_bits_3; // @[Reg.scala 28:20]
  reg  s2_ahead_fh_oldest_bits_afhob_3_bits_0; // @[Reg.scala 28:20]
  reg  s2_ahead_fh_oldest_bits_afhob_3_bits_1; // @[Reg.scala 28:20]
  reg  s2_ahead_fh_oldest_bits_afhob_3_bits_2; // @[Reg.scala 28:20]
  reg  s2_ahead_fh_oldest_bits_afhob_3_bits_3; // @[Reg.scala 28:20]
  reg  s2_ahead_fh_oldest_bits_afhob_2_bits_0; // @[Reg.scala 28:20]
  reg  s2_ahead_fh_oldest_bits_afhob_2_bits_1; // @[Reg.scala 28:20]
  reg  s2_ahead_fh_oldest_bits_afhob_2_bits_2; // @[Reg.scala 28:20]
  reg  s2_ahead_fh_oldest_bits_afhob_2_bits_3; // @[Reg.scala 28:20]
  reg  s2_ahead_fh_oldest_bits_afhob_1_bits_0; // @[Reg.scala 28:20]
  reg  s2_ahead_fh_oldest_bits_afhob_1_bits_1; // @[Reg.scala 28:20]
  reg  s2_ahead_fh_oldest_bits_afhob_1_bits_2; // @[Reg.scala 28:20]
  reg  s2_ahead_fh_oldest_bits_afhob_1_bits_3; // @[Reg.scala 28:20]
  reg  s2_ahead_fh_oldest_bits_afhob_0_bits_0; // @[Reg.scala 28:20]
  reg  s2_ahead_fh_oldest_bits_afhob_0_bits_1; // @[Reg.scala 28:20]
  reg  s2_ahead_fh_oldest_bits_afhob_0_bits_2; // @[Reg.scala 28:20]
  reg  s2_ahead_fh_oldest_bits_afhob_0_bits_3; // @[Reg.scala 28:20]
  reg  s3_ahead_fh_oldest_bits_afhob_5_bits_0; // @[Reg.scala 28:20]
  reg  s3_ahead_fh_oldest_bits_afhob_5_bits_1; // @[Reg.scala 28:20]
  reg  s3_ahead_fh_oldest_bits_afhob_5_bits_2; // @[Reg.scala 28:20]
  reg  s3_ahead_fh_oldest_bits_afhob_5_bits_3; // @[Reg.scala 28:20]
  reg  s3_ahead_fh_oldest_bits_afhob_4_bits_0; // @[Reg.scala 28:20]
  reg  s3_ahead_fh_oldest_bits_afhob_4_bits_1; // @[Reg.scala 28:20]
  reg  s3_ahead_fh_oldest_bits_afhob_4_bits_2; // @[Reg.scala 28:20]
  reg  s3_ahead_fh_oldest_bits_afhob_4_bits_3; // @[Reg.scala 28:20]
  reg  s3_ahead_fh_oldest_bits_afhob_3_bits_0; // @[Reg.scala 28:20]
  reg  s3_ahead_fh_oldest_bits_afhob_3_bits_1; // @[Reg.scala 28:20]
  reg  s3_ahead_fh_oldest_bits_afhob_3_bits_2; // @[Reg.scala 28:20]
  reg  s3_ahead_fh_oldest_bits_afhob_3_bits_3; // @[Reg.scala 28:20]
  reg  s3_ahead_fh_oldest_bits_afhob_2_bits_0; // @[Reg.scala 28:20]
  reg  s3_ahead_fh_oldest_bits_afhob_2_bits_1; // @[Reg.scala 28:20]
  reg  s3_ahead_fh_oldest_bits_afhob_2_bits_2; // @[Reg.scala 28:20]
  reg  s3_ahead_fh_oldest_bits_afhob_2_bits_3; // @[Reg.scala 28:20]
  reg  s3_ahead_fh_oldest_bits_afhob_1_bits_0; // @[Reg.scala 28:20]
  reg  s3_ahead_fh_oldest_bits_afhob_1_bits_1; // @[Reg.scala 28:20]
  reg  s3_ahead_fh_oldest_bits_afhob_1_bits_2; // @[Reg.scala 28:20]
  reg  s3_ahead_fh_oldest_bits_afhob_1_bits_3; // @[Reg.scala 28:20]
  reg  s3_ahead_fh_oldest_bits_afhob_0_bits_0; // @[Reg.scala 28:20]
  reg  s3_ahead_fh_oldest_bits_afhob_0_bits_1; // @[Reg.scala 28:20]
  reg  s3_ahead_fh_oldest_bits_afhob_0_bits_2; // @[Reg.scala 28:20]
  reg  s3_ahead_fh_oldest_bits_afhob_0_bits_3; // @[Reg.scala 28:20]
  reg  ghv_0; // @[BPU.scala 293:20]
  reg  ghv_1; // @[BPU.scala 293:20]
  reg  ghv_2; // @[BPU.scala 293:20]
  reg  ghv_3; // @[BPU.scala 293:20]
  reg  ghv_4; // @[BPU.scala 293:20]
  reg  ghv_5; // @[BPU.scala 293:20]
  reg  ghv_6; // @[BPU.scala 293:20]
  reg  ghv_7; // @[BPU.scala 293:20]
  reg  ghv_8; // @[BPU.scala 293:20]
  reg  ghv_9; // @[BPU.scala 293:20]
  reg  ghv_10; // @[BPU.scala 293:20]
  reg  ghv_11; // @[BPU.scala 293:20]
  reg  ghv_12; // @[BPU.scala 293:20]
  reg  ghv_13; // @[BPU.scala 293:20]
  reg  ghv_14; // @[BPU.scala 293:20]
  reg  ghv_15; // @[BPU.scala 293:20]
  reg  ghv_16; // @[BPU.scala 293:20]
  reg  ghv_17; // @[BPU.scala 293:20]
  reg  ghv_18; // @[BPU.scala 293:20]
  reg  ghv_19; // @[BPU.scala 293:20]
  reg  ghv_20; // @[BPU.scala 293:20]
  reg  ghv_21; // @[BPU.scala 293:20]
  reg  ghv_22; // @[BPU.scala 293:20]
  reg  ghv_23; // @[BPU.scala 293:20]
  reg  ghv_24; // @[BPU.scala 293:20]
  reg  ghv_25; // @[BPU.scala 293:20]
  reg  ghv_26; // @[BPU.scala 293:20]
  reg  ghv_27; // @[BPU.scala 293:20]
  reg  ghv_28; // @[BPU.scala 293:20]
  reg  ghv_29; // @[BPU.scala 293:20]
  reg  ghv_30; // @[BPU.scala 293:20]
  reg  ghv_31; // @[BPU.scala 293:20]
  reg  ghv_32; // @[BPU.scala 293:20]
  reg  ghv_33; // @[BPU.scala 293:20]
  reg  ghv_34; // @[BPU.scala 293:20]
  reg  ghv_35; // @[BPU.scala 293:20]
  reg  ghv_36; // @[BPU.scala 293:20]
  reg  ghv_37; // @[BPU.scala 293:20]
  reg  ghv_38; // @[BPU.scala 293:20]
  reg  ghv_39; // @[BPU.scala 293:20]
  reg  ghv_40; // @[BPU.scala 293:20]
  reg  ghv_41; // @[BPU.scala 293:20]
  reg  ghv_42; // @[BPU.scala 293:20]
  reg  ghv_43; // @[BPU.scala 293:20]
  reg  ghv_44; // @[BPU.scala 293:20]
  reg  ghv_45; // @[BPU.scala 293:20]
  reg  ghv_46; // @[BPU.scala 293:20]
  reg  ghv_47; // @[BPU.scala 293:20]
  reg  ghv_48; // @[BPU.scala 293:20]
  reg  ghv_49; // @[BPU.scala 293:20]
  reg  ghv_50; // @[BPU.scala 293:20]
  reg  ghv_51; // @[BPU.scala 293:20]
  reg  ghv_52; // @[BPU.scala 293:20]
  reg  ghv_53; // @[BPU.scala 293:20]
  reg  ghv_54; // @[BPU.scala 293:20]
  reg  ghv_55; // @[BPU.scala 293:20]
  reg  ghv_56; // @[BPU.scala 293:20]
  reg  ghv_57; // @[BPU.scala 293:20]
  reg  ghv_58; // @[BPU.scala 293:20]
  reg  ghv_59; // @[BPU.scala 293:20]
  reg  ghv_60; // @[BPU.scala 293:20]
  reg  ghv_61; // @[BPU.scala 293:20]
  reg  ghv_62; // @[BPU.scala 293:20]
  reg  ghv_63; // @[BPU.scala 293:20]
  reg  ghv_64; // @[BPU.scala 293:20]
  reg  ghv_65; // @[BPU.scala 293:20]
  reg  ghv_66; // @[BPU.scala 293:20]
  reg  ghv_67; // @[BPU.scala 293:20]
  reg  ghv_68; // @[BPU.scala 293:20]
  reg  ghv_69; // @[BPU.scala 293:20]
  reg  ghv_70; // @[BPU.scala 293:20]
  reg  ghv_71; // @[BPU.scala 293:20]
  reg  ghv_72; // @[BPU.scala 293:20]
  reg  ghv_73; // @[BPU.scala 293:20]
  reg  ghv_74; // @[BPU.scala 293:20]
  reg  ghv_75; // @[BPU.scala 293:20]
  reg  ghv_76; // @[BPU.scala 293:20]
  reg  ghv_77; // @[BPU.scala 293:20]
  reg  ghv_78; // @[BPU.scala 293:20]
  reg  ghv_79; // @[BPU.scala 293:20]
  reg  ghv_80; // @[BPU.scala 293:20]
  reg  ghv_81; // @[BPU.scala 293:20]
  reg  ghv_82; // @[BPU.scala 293:20]
  reg  ghv_83; // @[BPU.scala 293:20]
  reg  ghv_84; // @[BPU.scala 293:20]
  reg  ghv_85; // @[BPU.scala 293:20]
  reg  ghv_86; // @[BPU.scala 293:20]
  reg  ghv_87; // @[BPU.scala 293:20]
  reg  ghv_88; // @[BPU.scala 293:20]
  reg  ghv_89; // @[BPU.scala 293:20]
  reg  ghv_90; // @[BPU.scala 293:20]
  reg  ghv_91; // @[BPU.scala 293:20]
  reg  ghv_92; // @[BPU.scala 293:20]
  reg  ghv_93; // @[BPU.scala 293:20]
  reg  ghv_94; // @[BPU.scala 293:20]
  reg  ghv_95; // @[BPU.scala 293:20]
  reg  ghv_96; // @[BPU.scala 293:20]
  reg  ghv_97; // @[BPU.scala 293:20]
  reg  ghv_98; // @[BPU.scala 293:20]
  reg  ghv_99; // @[BPU.scala 293:20]
  reg  ghv_100; // @[BPU.scala 293:20]
  reg  ghv_101; // @[BPU.scala 293:20]
  reg  ghv_102; // @[BPU.scala 293:20]
  reg  ghv_103; // @[BPU.scala 293:20]
  reg  ghv_104; // @[BPU.scala 293:20]
  reg  ghv_105; // @[BPU.scala 293:20]
  reg  ghv_106; // @[BPU.scala 293:20]
  reg  ghv_107; // @[BPU.scala 293:20]
  reg  ghv_108; // @[BPU.scala 293:20]
  reg  ghv_109; // @[BPU.scala 293:20]
  reg  ghv_110; // @[BPU.scala 293:20]
  reg  ghv_111; // @[BPU.scala 293:20]
  reg  ghv_112; // @[BPU.scala 293:20]
  reg  ghv_113; // @[BPU.scala 293:20]
  reg  ghv_114; // @[BPU.scala 293:20]
  reg  ghv_115; // @[BPU.scala 293:20]
  reg  ghv_116; // @[BPU.scala 293:20]
  reg  ghv_117; // @[BPU.scala 293:20]
  reg  ghv_118; // @[BPU.scala 293:20]
  reg  ghv_119; // @[BPU.scala 293:20]
  reg  ghv_120; // @[BPU.scala 293:20]
  reg  ghv_121; // @[BPU.scala 293:20]
  reg  ghv_122; // @[BPU.scala 293:20]
  reg  ghv_123; // @[BPU.scala 293:20]
  reg  ghv_124; // @[BPU.scala 293:20]
  reg  ghv_125; // @[BPU.scala 293:20]
  reg  ghv_126; // @[BPU.scala 293:20]
  reg  ghv_127; // @[BPU.scala 293:20]
  reg  ghv_128; // @[BPU.scala 293:20]
  reg  ghv_129; // @[BPU.scala 293:20]
  reg  ghv_130; // @[BPU.scala 293:20]
  reg  ghv_131; // @[BPU.scala 293:20]
  reg  ghv_132; // @[BPU.scala 293:20]
  reg  ghv_133; // @[BPU.scala 293:20]
  reg  ghv_134; // @[BPU.scala 293:20]
  reg  ghv_135; // @[BPU.scala 293:20]
  reg  ghv_136; // @[BPU.scala 293:20]
  reg  ghv_137; // @[BPU.scala 293:20]
  reg  ghv_138; // @[BPU.scala 293:20]
  reg  ghv_139; // @[BPU.scala 293:20]
  reg  ghv_140; // @[BPU.scala 293:20]
  reg  ghv_141; // @[BPU.scala 293:20]
  reg  ghv_142; // @[BPU.scala 293:20]
  reg  ghv_143; // @[BPU.scala 293:20]
  reg  s0_ghist_ptr_reg_flag; // @[BPU.scala 304:33]
  reg [7:0] s0_ghist_ptr_reg_value; // @[BPU.scala 304:33]
  reg  s1_ghist_ptr_flag; // @[Reg.scala 28:20]
  reg [7:0] s1_ghist_ptr_value; // @[Reg.scala 28:20]
  wire  s0_ghist_ptr_flag = s0_ghist_ptr_ppm_out_res_flag; // @[BPU.scala 303:26 669:17]
  wire [7:0] s0_ghist_ptr_value = s0_ghist_ptr_ppm_out_res_value; // @[BPU.scala 303:26 669:17]
  reg  s2_ghist_ptr_flag; // @[Reg.scala 28:20]
  reg [7:0] s2_ghist_ptr_value; // @[Reg.scala 28:20]
  reg  s3_ghist_ptr_flag; // @[Reg.scala 28:20]
  reg [7:0] s3_ghist_ptr_value; // @[Reg.scala 28:20]
  reg  do_redirect_valid; // @[BPU.scala 332:28]
  reg  do_redirect_bits_level; // @[BPU.scala 332:28]
  reg [38:0] do_redirect_bits_cfiUpdate_pc; // @[BPU.scala 332:28]
  reg  do_redirect_bits_cfiUpdate_pd_isRVC; // @[BPU.scala 332:28]
  reg  do_redirect_bits_cfiUpdate_pd_isCall; // @[BPU.scala 332:28]
  reg  do_redirect_bits_cfiUpdate_pd_isRet; // @[BPU.scala 332:28]
  reg [4:0] do_redirect_bits_cfiUpdate_rasSp; // @[BPU.scala 332:28]
  reg [38:0] do_redirect_bits_cfiUpdate_rasEntry_retAddr; // @[BPU.scala 332:28]
  reg [7:0] do_redirect_bits_cfiUpdate_rasEntry_ctr; // @[BPU.scala 332:28]
  reg [7:0] do_redirect_bits_cfiUpdate_folded_hist_hist_17_folded_hist; // @[BPU.scala 332:28]
  reg [7:0] do_redirect_bits_cfiUpdate_folded_hist_hist_16_folded_hist; // @[BPU.scala 332:28]
  reg [10:0] do_redirect_bits_cfiUpdate_folded_hist_hist_15_folded_hist; // @[BPU.scala 332:28]
  reg [6:0] do_redirect_bits_cfiUpdate_folded_hist_hist_14_folded_hist; // @[BPU.scala 332:28]
  reg [6:0] do_redirect_bits_cfiUpdate_folded_hist_hist_13_folded_hist; // @[BPU.scala 332:28]
  reg [6:0] do_redirect_bits_cfiUpdate_folded_hist_hist_12_folded_hist; // @[BPU.scala 332:28]
  reg [7:0] do_redirect_bits_cfiUpdate_folded_hist_hist_11_folded_hist; // @[BPU.scala 332:28]
  reg [8:0] do_redirect_bits_cfiUpdate_folded_hist_hist_10_folded_hist; // @[BPU.scala 332:28]
  reg [6:0] do_redirect_bits_cfiUpdate_folded_hist_hist_9_folded_hist; // @[BPU.scala 332:28]
  reg [7:0] do_redirect_bits_cfiUpdate_folded_hist_hist_8_folded_hist; // @[BPU.scala 332:28]
  reg [8:0] do_redirect_bits_cfiUpdate_folded_hist_hist_7_folded_hist; // @[BPU.scala 332:28]
  reg [8:0] do_redirect_bits_cfiUpdate_folded_hist_hist_6_folded_hist; // @[BPU.scala 332:28]
  reg [10:0] do_redirect_bits_cfiUpdate_folded_hist_hist_5_folded_hist; // @[BPU.scala 332:28]
  reg [3:0] do_redirect_bits_cfiUpdate_folded_hist_hist_4_folded_hist; // @[BPU.scala 332:28]
  reg [10:0] do_redirect_bits_cfiUpdate_folded_hist_hist_3_folded_hist; // @[BPU.scala 332:28]
  reg [7:0] do_redirect_bits_cfiUpdate_folded_hist_hist_2_folded_hist; // @[BPU.scala 332:28]
  reg [7:0] do_redirect_bits_cfiUpdate_folded_hist_hist_1_folded_hist; // @[BPU.scala 332:28]
  reg [7:0] do_redirect_bits_cfiUpdate_folded_hist_hist_0_folded_hist; // @[BPU.scala 332:28]
  reg  do_redirect_bits_cfiUpdate_afhob_afhob_5_bits_0; // @[BPU.scala 332:28]
  reg  do_redirect_bits_cfiUpdate_afhob_afhob_5_bits_1; // @[BPU.scala 332:28]
  reg  do_redirect_bits_cfiUpdate_afhob_afhob_5_bits_2; // @[BPU.scala 332:28]
  reg  do_redirect_bits_cfiUpdate_afhob_afhob_5_bits_3; // @[BPU.scala 332:28]
  reg  do_redirect_bits_cfiUpdate_afhob_afhob_4_bits_0; // @[BPU.scala 332:28]
  reg  do_redirect_bits_cfiUpdate_afhob_afhob_4_bits_1; // @[BPU.scala 332:28]
  reg  do_redirect_bits_cfiUpdate_afhob_afhob_4_bits_2; // @[BPU.scala 332:28]
  reg  do_redirect_bits_cfiUpdate_afhob_afhob_3_bits_0; // @[BPU.scala 332:28]
  reg  do_redirect_bits_cfiUpdate_afhob_afhob_3_bits_1; // @[BPU.scala 332:28]
  reg  do_redirect_bits_cfiUpdate_afhob_afhob_3_bits_2; // @[BPU.scala 332:28]
  reg  do_redirect_bits_cfiUpdate_afhob_afhob_3_bits_3; // @[BPU.scala 332:28]
  reg  do_redirect_bits_cfiUpdate_afhob_afhob_2_bits_0; // @[BPU.scala 332:28]
  reg  do_redirect_bits_cfiUpdate_afhob_afhob_2_bits_1; // @[BPU.scala 332:28]
  reg  do_redirect_bits_cfiUpdate_afhob_afhob_2_bits_2; // @[BPU.scala 332:28]
  reg  do_redirect_bits_cfiUpdate_afhob_afhob_2_bits_3; // @[BPU.scala 332:28]
  reg  do_redirect_bits_cfiUpdate_afhob_afhob_1_bits_0; // @[BPU.scala 332:28]
  reg  do_redirect_bits_cfiUpdate_afhob_afhob_1_bits_1; // @[BPU.scala 332:28]
  reg  do_redirect_bits_cfiUpdate_afhob_afhob_1_bits_2; // @[BPU.scala 332:28]
  reg  do_redirect_bits_cfiUpdate_afhob_afhob_1_bits_3; // @[BPU.scala 332:28]
  reg  do_redirect_bits_cfiUpdate_afhob_afhob_0_bits_0; // @[BPU.scala 332:28]
  reg  do_redirect_bits_cfiUpdate_afhob_afhob_0_bits_1; // @[BPU.scala 332:28]
  reg  do_redirect_bits_cfiUpdate_afhob_afhob_0_bits_2; // @[BPU.scala 332:28]
  reg  do_redirect_bits_cfiUpdate_afhob_afhob_0_bits_3; // @[BPU.scala 332:28]
  reg [2:0] do_redirect_bits_cfiUpdate_lastBrNumOH; // @[BPU.scala 332:28]
  reg  do_redirect_bits_cfiUpdate_histPtr_flag; // @[BPU.scala 332:28]
  reg [7:0] do_redirect_bits_cfiUpdate_histPtr_value; // @[BPU.scala 332:28]
  reg [38:0] do_redirect_bits_cfiUpdate_target; // @[BPU.scala 332:28]
  reg  do_redirect_bits_cfiUpdate_taken; // @[BPU.scala 332:28]
  reg [1:0] do_redirect_bits_cfiUpdate_shift; // @[BPU.scala 332:28]
  reg  do_redirect_bits_cfiUpdate_addIntoHist; // @[BPU.scala 332:28]
  wire  _s3_redirect_on_br_taken_T_9 = predictors_io_out_s3_full_pred_br_taken_mask_1 &
    predictors_io_out_s3_full_pred_slot_valids_1 & predictors_io_out_s3_full_pred_is_br_sharing &
    predictors_io_out_s3_full_pred_hit; // @[FrontendBundle.scala 451:63]
  wire  _s3_redirect_on_br_taken_T = predictors_io_out_s3_full_pred_slot_valids_0 &
    predictors_io_out_s3_full_pred_br_taken_mask_0; // @[FrontendBundle.scala 435:69]
  wire  _s3_redirect_on_br_taken_T_5 = _s3_redirect_on_br_taken_T & predictors_io_out_s3_full_pred_hit; // @[FrontendBundle.scala 450:32]
  wire [1:0] _s3_redirect_on_br_taken_T_10 = {_s3_redirect_on_br_taken_T_9,_s3_redirect_on_br_taken_T_5}; // @[BPU.scala 563:72]
  reg  previous_s2_pred_full_pred_br_taken_mask_1; // @[Reg.scala 28:20]
  reg  previous_s2_pred_full_pred_slot_valids_1; // @[Reg.scala 28:20]
  reg  previous_s2_pred_full_pred_is_br_sharing; // @[Reg.scala 28:20]
  reg  previous_s2_pred_full_pred_hit; // @[Reg.scala 28:20]
  wire  _s3_redirect_on_br_taken_T_20 = previous_s2_pred_full_pred_br_taken_mask_1 &
    previous_s2_pred_full_pred_slot_valids_1 & previous_s2_pred_full_pred_is_br_sharing & previous_s2_pred_full_pred_hit
    ; // @[FrontendBundle.scala 451:63]
  reg  previous_s2_pred_full_pred_slot_valids_0; // @[Reg.scala 28:20]
  reg  previous_s2_pred_full_pred_br_taken_mask_0; // @[Reg.scala 28:20]
  wire  _s3_redirect_on_br_taken_T_11 = previous_s2_pred_full_pred_slot_valids_0 &
    previous_s2_pred_full_pred_br_taken_mask_0; // @[FrontendBundle.scala 435:69]
  wire  _s3_redirect_on_br_taken_T_16 = _s3_redirect_on_br_taken_T_11 & previous_s2_pred_full_pred_hit; // @[FrontendBundle.scala 450:32]
  wire [1:0] _s3_redirect_on_br_taken_T_21 = {_s3_redirect_on_br_taken_T_20,_s3_redirect_on_br_taken_T_16}; // @[BPU.scala 563:131]
  wire  s3_redirect_on_br_taken = _s3_redirect_on_br_taken_T_10 != _s3_redirect_on_br_taken_T_21; // @[BPU.scala 563:79]
  wire [38:0] _s3_redirect_on_target_T = _s3_redirect_on_br_taken_T_5 ? predictors_io_out_s3_full_pred_targets_0 : 39'h0
    ; // @[Mux.scala 27:73]
  wire  _s3_redirect_on_target_tm_T_3 = predictors_io_out_s3_full_pred_is_br_sharing &
    predictors_io_out_s3_full_pred_br_taken_mask_1 | ~predictors_io_out_s3_full_pred_is_br_sharing; // @[FrontendBundle.scala 437:47]
  wire  tm_3_1 = predictors_io_out_s3_full_pred_slot_valids_1 & _s3_redirect_on_target_tm_T_3; // @[FrontendBundle.scala 436:25]
  wire  selVecOH_1_3 = ~_s3_redirect_on_br_taken_T & tm_3_1 & predictors_io_out_s3_full_pred_hit; // @[FrontendBundle.scala 476:80]
  wire [38:0] _s3_redirect_on_target_T_1 = selVecOH_1_3 ? predictors_io_out_s3_full_pred_targets_1 : 39'h0; // @[Mux.scala 27:73]
  wire [38:0] _s3_redirect_on_target_T_4 = _s3_redirect_on_target_T | _s3_redirect_on_target_T_1; // @[Mux.scala 27:73]
  wire [1:0] _s3_redirect_on_target_selVecOH_T_5 = {tm_3_1,_s3_redirect_on_br_taken_T}; // @[FrontendBundle.scala 477:12]
  wire  selVecOH_2_3 = ~(|_s3_redirect_on_target_selVecOH_T_5) & predictors_io_out_s3_full_pred_hit; // @[FrontendBundle.scala 477:23]
  wire [38:0] _s3_redirect_on_target_T_2 = selVecOH_2_3 ? predictors_io_out_s3_full_pred_fallThroughAddr : 39'h0; // @[Mux.scala 27:73]
  wire [38:0] _s3_redirect_on_target_T_5 = _s3_redirect_on_target_T_4 | _s3_redirect_on_target_T_2; // @[Mux.scala 27:73]
  wire  selVecOH_3_3 = ~predictors_io_out_s3_full_pred_hit; // @[FrontendBundle.scala 477:34]
  wire [38:0] targetVec_3_3 = predictors_io_out_s3_pc + 39'h10; // @[FrontendBundle.scala 473:55]
  wire [38:0] _s3_redirect_on_target_T_3 = selVecOH_3_3 ? targetVec_3_3 : 39'h0; // @[Mux.scala 27:73]
  wire [38:0] _s3_redirect_on_target_T_6 = _s3_redirect_on_target_T_5 | _s3_redirect_on_target_T_3; // @[Mux.scala 27:73]
  reg [38:0] previous_s2_pred_full_pred_targets_0; // @[Reg.scala 28:20]
  wire [38:0] _s3_redirect_on_target_T_7 = _s3_redirect_on_br_taken_T_16 ? previous_s2_pred_full_pred_targets_0 : 39'h0; // @[Mux.scala 27:73]
  wire  _s3_redirect_on_target_tm_T_8 = previous_s2_pred_full_pred_is_br_sharing &
    previous_s2_pred_full_pred_br_taken_mask_1 | ~previous_s2_pred_full_pred_is_br_sharing; // @[FrontendBundle.scala 437:47]
  wire  tm_4_1 = previous_s2_pred_full_pred_slot_valids_1 & _s3_redirect_on_target_tm_T_8; // @[FrontendBundle.scala 436:25]
  wire  selVecOH_1_4 = ~_s3_redirect_on_br_taken_T_11 & tm_4_1 & previous_s2_pred_full_pred_hit; // @[FrontendBundle.scala 476:80]
  reg [38:0] previous_s2_pred_full_pred_targets_1; // @[Reg.scala 28:20]
  wire [38:0] _s3_redirect_on_target_T_8 = selVecOH_1_4 ? previous_s2_pred_full_pred_targets_1 : 39'h0; // @[Mux.scala 27:73]
  wire [38:0] _s3_redirect_on_target_T_11 = _s3_redirect_on_target_T_7 | _s3_redirect_on_target_T_8; // @[Mux.scala 27:73]
  wire [1:0] _s3_redirect_on_target_selVecOH_T_13 = {tm_4_1,_s3_redirect_on_br_taken_T_11}; // @[FrontendBundle.scala 477:12]
  wire  selVecOH_2_4 = ~(|_s3_redirect_on_target_selVecOH_T_13) & previous_s2_pred_full_pred_hit; // @[FrontendBundle.scala 477:23]
  reg [38:0] previous_s2_pred_full_pred_fallThroughAddr; // @[Reg.scala 28:20]
  wire [38:0] _s3_redirect_on_target_T_9 = selVecOH_2_4 ? previous_s2_pred_full_pred_fallThroughAddr : 39'h0; // @[Mux.scala 27:73]
  wire [38:0] _s3_redirect_on_target_T_12 = _s3_redirect_on_target_T_11 | _s3_redirect_on_target_T_9; // @[Mux.scala 27:73]
  wire  selVecOH_3_4 = ~previous_s2_pred_full_pred_hit; // @[FrontendBundle.scala 477:34]
  reg [38:0] previous_s2_pred_pc; // @[Reg.scala 28:20]
  wire [38:0] targetVec_3_4 = previous_s2_pred_pc + 39'h10; // @[FrontendBundle.scala 473:55]
  wire [38:0] _s3_redirect_on_target_T_10 = selVecOH_3_4 ? targetVec_3_4 : 39'h0; // @[Mux.scala 27:73]
  wire [38:0] _s3_redirect_on_target_T_13 = _s3_redirect_on_target_T_12 | _s3_redirect_on_target_T_10; // @[Mux.scala 27:73]
  wire  s3_redirect_on_target = _s3_redirect_on_target_T_6 != _s3_redirect_on_target_T_13; // @[BPU.scala 564:49]
  wire  s3_redirect_on_fall_thru_error = predictors_io_out_s3_full_pred_hit &
    predictors_io_out_s3_full_pred_fallThroughErr; // @[FrontendBundle.scala 481:33]
  wire  _s3_redirect_T_1 = s3_redirect_on_br_taken | s3_redirect_on_target | s3_redirect_on_fall_thru_error; // @[BPU.scala 569:54]
  wire  s3_redirect = s3_valid & _s3_redirect_T_1; // @[BPU.scala 568:26]
  wire  s2_flush = io_ftq_to_bpu_redirect_valid | s3_redirect; // @[BPU.scala 339:24]
  reg [38:0] previous_s1_pred_info_target; // @[Reg.scala 28:20]
  wire  s2_redirect_s1_last_pred_vec_tm_0 = predictors_io_out_s2_full_pred_slot_valids_0 &
    predictors_io_out_s2_full_pred_br_taken_mask_0; // @[FrontendBundle.scala 435:69]
  wire  s2_redirect_s1_last_pred_vec_selVecOH_0 = s2_redirect_s1_last_pred_vec_tm_0 & predictors_io_out_s2_full_pred_hit
    ; // @[FrontendBundle.scala 476:80]
  wire [38:0] _s2_redirect_s1_last_pred_vec_T = s2_redirect_s1_last_pred_vec_selVecOH_0 ?
    predictors_io_out_s2_full_pred_targets_0 : 39'h0; // @[Mux.scala 27:73]
  wire  _s2_redirect_s1_last_pred_vec_tm_T_3 = predictors_io_out_s2_full_pred_is_br_sharing &
    predictors_io_out_s2_full_pred_br_taken_mask_1 | ~predictors_io_out_s2_full_pred_is_br_sharing; // @[FrontendBundle.scala 437:47]
  wire  s2_redirect_s1_last_pred_vec_tm_1 = predictors_io_out_s2_full_pred_slot_valids_1 &
    _s2_redirect_s1_last_pred_vec_tm_T_3; // @[FrontendBundle.scala 436:25]
  wire  s2_redirect_s1_last_pred_vec_selVecOH_1 = ~s2_redirect_s1_last_pred_vec_tm_0 & s2_redirect_s1_last_pred_vec_tm_1
     & predictors_io_out_s2_full_pred_hit; // @[FrontendBundle.scala 476:80]
  wire [38:0] _s2_redirect_s1_last_pred_vec_T_1 = s2_redirect_s1_last_pred_vec_selVecOH_1 ?
    predictors_io_out_s2_full_pred_targets_1 : 39'h0; // @[Mux.scala 27:73]
  wire [38:0] _s2_redirect_s1_last_pred_vec_T_4 = _s2_redirect_s1_last_pred_vec_T | _s2_redirect_s1_last_pred_vec_T_1; // @[Mux.scala 27:73]
  wire [1:0] _s2_redirect_s1_last_pred_vec_selVecOH_T_5 = {s2_redirect_s1_last_pred_vec_tm_1,
    s2_redirect_s1_last_pred_vec_tm_0}; // @[FrontendBundle.scala 477:12]
  wire  s2_redirect_s1_last_pred_vec_selVecOH_2 = ~(|_s2_redirect_s1_last_pred_vec_selVecOH_T_5) &
    predictors_io_out_s2_full_pred_hit; // @[FrontendBundle.scala 477:23]
  wire [38:0] _s2_redirect_s1_last_pred_vec_T_2 = s2_redirect_s1_last_pred_vec_selVecOH_2 ?
    predictors_io_out_s2_full_pred_fallThroughAddr : 39'h0; // @[Mux.scala 27:73]
  wire [38:0] _s2_redirect_s1_last_pred_vec_T_5 = _s2_redirect_s1_last_pred_vec_T_4 | _s2_redirect_s1_last_pred_vec_T_2; // @[Mux.scala 27:73]
  wire  s2_redirect_s1_last_pred_vec_selVecOH_3 = ~predictors_io_out_s2_full_pred_hit; // @[FrontendBundle.scala 477:34]
  wire [38:0] s2_redirect_s1_last_pred_vec_targetVec_3 = predictors_io_out_s2_pc + 39'h10; // @[FrontendBundle.scala 473:55]
  wire [38:0] _s2_redirect_s1_last_pred_vec_T_3 = s2_redirect_s1_last_pred_vec_selVecOH_3 ?
    s2_redirect_s1_last_pred_vec_targetVec_3 : 39'h0; // @[Mux.scala 27:73]
  wire [38:0] _s2_redirect_s1_last_pred_vec_T_6 = _s2_redirect_s1_last_pred_vec_T_5 | _s2_redirect_s1_last_pred_vec_T_3; // @[Mux.scala 27:73]
  wire  s2_redirect_s1_last_pred_vec_0 = previous_s1_pred_info_target != _s2_redirect_s1_last_pred_vec_T_6; // @[BPU.scala 450:16]
  reg [2:0] previous_s1_pred_info_lastBrPosOH; // @[Reg.scala 28:20]
  wire  _s2_redirect_s1_last_pred_vec_T_41 = predictors_io_out_s2_full_pred_slot_valids_1 &
    predictors_io_out_s2_full_pred_is_br_sharing; // @[FrontendBundle.scala 430:48]
  wire  _s2_redirect_s1_last_pred_vec_T_52 = ~s2_redirect_s1_last_pred_vec_selVecOH_0; // @[FrontendBundle.scala 464:9]
  wire  _s2_redirect_s1_last_pred_vec_T_53 = _s2_redirect_s1_last_pred_vec_T_41 & _s2_redirect_s1_last_pred_vec_T_52; // @[FrontendBundle.scala 463:22]
  wire  _s2_redirect_s1_last_pred_vec_T_63 = predictors_io_out_s2_full_pred_br_taken_mask_1 &
    predictors_io_out_s2_full_pred_slot_valids_1 & predictors_io_out_s2_full_pred_is_br_sharing &
    predictors_io_out_s2_full_pred_hit; // @[FrontendBundle.scala 451:63]
  wire  _s2_redirect_s1_last_pred_vec_T_68 = _s2_redirect_s1_last_pred_vec_T_53 & predictors_io_out_s2_full_pred_hit; // @[FrontendBundle.scala 465:97]
  wire  _s2_redirect_s1_last_pred_vec_WIRE_2_0 = predictors_io_out_s2_full_pred_slot_valids_0; // @[FrontendBundle.scala 430:{12,12}]
  wire  _s2_redirect_s1_last_pred_vec_T_38 = s2_redirect_s1_last_pred_vec_selVecOH_0 | ~
    _s2_redirect_s1_last_pred_vec_T_41; // @[FrontendBundle.scala 465:34]
  wire  _s2_redirect_s1_last_pred_vec_T_39 = _s2_redirect_s1_last_pred_vec_WIRE_2_0 & _s2_redirect_s1_last_pred_vec_T_38
    ; // @[FrontendBundle.scala 464:75]
  wire  _s2_redirect_s1_last_pred_vec_T_40 = _s2_redirect_s1_last_pred_vec_T_39 & predictors_io_out_s2_full_pred_hit; // @[FrontendBundle.scala 465:97]
  wire [1:0] s2_redirect_s1_last_pred_vec_hi = {_s2_redirect_s1_last_pred_vec_T_68,_s2_redirect_s1_last_pred_vec_T_40}; // @[BPU.scala 451:39]
  wire  _s2_redirect_s1_last_pred_vec_T_12 = s2_redirect_s1_last_pred_vec_selVecOH_3 | ~(
    _s2_redirect_s1_last_pred_vec_WIRE_2_0 | _s2_redirect_s1_last_pred_vec_T_41); // @[FrontendBundle.scala 461:19]
  wire [2:0] _s2_redirect_s1_last_pred_vec_T_69 = {_s2_redirect_s1_last_pred_vec_T_68,_s2_redirect_s1_last_pred_vec_T_40
    ,_s2_redirect_s1_last_pred_vec_T_12}; // @[BPU.scala 451:39]
  wire  s2_redirect_s1_last_pred_vec_1 = previous_s1_pred_info_lastBrPosOH != _s2_redirect_s1_last_pred_vec_T_69; // @[BPU.scala 451:21]
  reg  previous_s1_pred_info_taken; // @[Reg.scala 28:20]
  wire  _s2_redirect_s1_last_pred_vec_cfiIndex_valid_T_6 = s2_redirect_s1_last_pred_vec_tm_1 &
    predictors_io_out_s2_full_pred_hit; // @[FrontendBundle.scala 444:38]
  wire [1:0] _s2_redirect_s1_last_pred_vec_cfiIndex_valid_T_7 = {_s2_redirect_s1_last_pred_vec_cfiIndex_valid_T_6,
    s2_redirect_s1_last_pred_vec_selVecOH_0}; // @[FrontendBundle.scala 492:46]
  wire  s2_redirect_s1_last_pred_vec_cfiIndex_valid = |_s2_redirect_s1_last_pred_vec_cfiIndex_valid_T_7; // @[FrontendBundle.scala 492:53]
  wire  s2_redirect_s1_last_pred_vec_2 = previous_s1_pred_info_taken != s2_redirect_s1_last_pred_vec_cfiIndex_valid; // @[BPU.scala 452:15]
  reg [2:0] previous_s1_pred_info_cfiIndex; // @[Reg.scala 28:20]
  wire [2:0] _s2_redirect_s1_last_pred_vec_cfiIndex_bits_T_52 = s2_redirect_s1_last_pred_vec_selVecOH_0 ?
    predictors_io_out_s2_full_pred_offsets_0 : predictors_io_out_s2_full_pred_offsets_1; // @[ParallelMux.scala 90:77]
  wire  _s2_redirect_s1_last_pred_vec_cfiIndex_bits_T_62 = ~s2_redirect_s1_last_pred_vec_cfiIndex_valid; // @[FrontendBundle.scala 496:37]
  wire [2:0] _s2_redirect_s1_last_pred_vec_cfiIndex_bits_T_64 = _s2_redirect_s1_last_pred_vec_cfiIndex_bits_T_62 ? 3'h7
     : 3'h0; // @[Bitwise.scala 74:12]
  wire [2:0] s2_redirect_s1_last_pred_vec_cfiIndex_2_bits = _s2_redirect_s1_last_pred_vec_cfiIndex_bits_T_52 |
    _s2_redirect_s1_last_pred_vec_cfiIndex_bits_T_64; // @[FrontendBundle.scala 495:60]
  wire  s2_redirect_s1_last_pred_vec_3 = previous_s1_pred_info_taken & s2_redirect_s1_last_pred_vec_cfiIndex_valid &
    previous_s1_pred_info_cfiIndex != s2_redirect_s1_last_pred_vec_cfiIndex_2_bits; // @[BPU.scala 453:28]
  wire  s2_redirect = s2_valid & (s2_redirect_s1_last_pred_vec_0 | s2_redirect_s1_last_pred_vec_1 |
    s2_redirect_s1_last_pred_vec_2 | s2_redirect_s1_last_pred_vec_3); // @[BPU.scala 503:26]
  wire  s1_flush = s2_flush | s2_redirect; // @[BPU.scala 340:24]
  wire  _GEN_139 = s1_fire ? 1'h0 : s1_valid; // @[BPU.scala 358:{29,40} 252:45]
  wire  _GEN_140 = s1_flush ? 1'h0 : _GEN_139; // @[BPU.scala 357:{29,40}]
  wire  _GEN_141 = s0_fire | _GEN_140; // @[BPU.scala 356:{29,40}]
  wire  _s3_valid_T = ~s2_flush; // @[BPU.scala 374:38]
  wire  _io_bpu_to_ftq_resp_valid_T_2 = s2_valid & s2_redirect; // @[BPU.scala 383:13]
  wire  _io_bpu_to_ftq_resp_valid_T_3 = _s1_fire_T_1 | _io_bpu_to_ftq_resp_valid_T_2; // @[BPU.scala 382:49]
  wire  _io_bpu_to_ftq_resp_valid_T_4 = s3_valid & s3_redirect; // @[BPU.scala 384:13]
  wire [7:0] _s1_possible_predicted_ghist_ptrs_flipped_new_ptr_T_1 = 8'h90 - 8'h0; // @[CircularQueuePtr.scala 54:50]
  wire [8:0] s1_possible_predicted_ghist_ptrs_flipped_new_ptr_new_value = s1_ghist_ptr_value +
    _s1_possible_predicted_ghist_ptrs_flipped_new_ptr_T_1; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _s1_possible_predicted_ghist_ptrs_flipped_new_ptr_diff_T_1 = {1'h0,
    s1_possible_predicted_ghist_ptrs_flipped_new_ptr_new_value}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] s1_possible_predicted_ghist_ptrs_flipped_new_ptr_diff = $signed(
    _s1_possible_predicted_ghist_ptrs_flipped_new_ptr_diff_T_1) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_possible_predicted_ghist_ptrs_flipped_new_ptr_reverse_flag = $signed(
    s1_possible_predicted_ghist_ptrs_flipped_new_ptr_diff) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire  s1_possible_predicted_ghist_ptrs_flipped_new_ptr_flag =
    s1_possible_predicted_ghist_ptrs_flipped_new_ptr_reverse_flag ? ~s1_ghist_ptr_flag : s1_ghist_ptr_flag; // @[CircularQueuePtr.scala 44:26]
  wire [9:0] _s1_possible_predicted_ghist_ptrs_flipped_new_ptr_new_ptr_value_T = $signed(
    _s1_possible_predicted_ghist_ptrs_flipped_new_ptr_diff_T_1) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_possible_predicted_ghist_ptrs_flipped_new_ptr_new_ptr_value_T_1 =
    s1_possible_predicted_ghist_ptrs_flipped_new_ptr_reverse_flag ?
    _s1_possible_predicted_ghist_ptrs_flipped_new_ptr_new_ptr_value_T : {{1'd0},
    s1_possible_predicted_ghist_ptrs_flipped_new_ptr_new_value}; // @[CircularQueuePtr.scala 45:27]
  wire  s1_possible_predicted_ghist_ptrs_0_flag = ~s1_possible_predicted_ghist_ptrs_flipped_new_ptr_flag; // @[CircularQueuePtr.scala 56:21]
  wire [7:0] _s1_possible_predicted_ghist_ptrs_flipped_new_ptr_T_3 = 8'h90 - 8'h1; // @[CircularQueuePtr.scala 54:50]
  wire [8:0] s1_possible_predicted_ghist_ptrs_flipped_new_ptr_new_value_1 = s1_ghist_ptr_value +
    _s1_possible_predicted_ghist_ptrs_flipped_new_ptr_T_3; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _s1_possible_predicted_ghist_ptrs_flipped_new_ptr_diff_T_7 = {1'h0,
    s1_possible_predicted_ghist_ptrs_flipped_new_ptr_new_value_1}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] s1_possible_predicted_ghist_ptrs_flipped_new_ptr_diff_1 = $signed(
    _s1_possible_predicted_ghist_ptrs_flipped_new_ptr_diff_T_7) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_possible_predicted_ghist_ptrs_flipped_new_ptr_reverse_flag_1 = $signed(
    s1_possible_predicted_ghist_ptrs_flipped_new_ptr_diff_1) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire  s1_possible_predicted_ghist_ptrs_flipped_new_ptr_1_flag =
    s1_possible_predicted_ghist_ptrs_flipped_new_ptr_reverse_flag_1 ? ~s1_ghist_ptr_flag : s1_ghist_ptr_flag; // @[CircularQueuePtr.scala 44:26]
  wire [9:0] _s1_possible_predicted_ghist_ptrs_flipped_new_ptr_new_ptr_value_T_2 = $signed(
    _s1_possible_predicted_ghist_ptrs_flipped_new_ptr_diff_T_7) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_possible_predicted_ghist_ptrs_flipped_new_ptr_new_ptr_value_T_3 =
    s1_possible_predicted_ghist_ptrs_flipped_new_ptr_reverse_flag_1 ?
    _s1_possible_predicted_ghist_ptrs_flipped_new_ptr_new_ptr_value_T_2 : {{1'd0},
    s1_possible_predicted_ghist_ptrs_flipped_new_ptr_new_value_1}; // @[CircularQueuePtr.scala 45:27]
  wire  s1_possible_predicted_ghist_ptrs_1_flag = ~s1_possible_predicted_ghist_ptrs_flipped_new_ptr_1_flag; // @[CircularQueuePtr.scala 56:21]
  wire [7:0] _s1_possible_predicted_ghist_ptrs_flipped_new_ptr_T_5 = 8'h90 - 8'h2; // @[CircularQueuePtr.scala 54:50]
  wire [8:0] s1_possible_predicted_ghist_ptrs_flipped_new_ptr_new_value_2 = s1_ghist_ptr_value +
    _s1_possible_predicted_ghist_ptrs_flipped_new_ptr_T_5; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _s1_possible_predicted_ghist_ptrs_flipped_new_ptr_diff_T_13 = {1'h0,
    s1_possible_predicted_ghist_ptrs_flipped_new_ptr_new_value_2}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] s1_possible_predicted_ghist_ptrs_flipped_new_ptr_diff_2 = $signed(
    _s1_possible_predicted_ghist_ptrs_flipped_new_ptr_diff_T_13) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_possible_predicted_ghist_ptrs_flipped_new_ptr_reverse_flag_2 = $signed(
    s1_possible_predicted_ghist_ptrs_flipped_new_ptr_diff_2) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire  s1_possible_predicted_ghist_ptrs_flipped_new_ptr_2_flag =
    s1_possible_predicted_ghist_ptrs_flipped_new_ptr_reverse_flag_2 ? ~s1_ghist_ptr_flag : s1_ghist_ptr_flag; // @[CircularQueuePtr.scala 44:26]
  wire [9:0] _s1_possible_predicted_ghist_ptrs_flipped_new_ptr_new_ptr_value_T_4 = $signed(
    _s1_possible_predicted_ghist_ptrs_flipped_new_ptr_diff_T_13) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_possible_predicted_ghist_ptrs_flipped_new_ptr_new_ptr_value_T_5 =
    s1_possible_predicted_ghist_ptrs_flipped_new_ptr_reverse_flag_2 ?
    _s1_possible_predicted_ghist_ptrs_flipped_new_ptr_new_ptr_value_T_4 : {{1'd0},
    s1_possible_predicted_ghist_ptrs_flipped_new_ptr_new_value_2}; // @[CircularQueuePtr.scala 45:27]
  wire  s1_possible_predicted_ghist_ptrs_2_flag = ~s1_possible_predicted_ghist_ptrs_flipped_new_ptr_2_flag; // @[CircularQueuePtr.scala 56:21]
  wire  _s1_predicted_ghist_ptr_T = ~predictors_io_out_s1_full_pred_hit; // @[FrontendBundle.scala 461:14]
  wire  _s1_predicted_ghist_ptr_T_1 = predictors_io_out_s1_full_pred_slot_valids_1 &
    predictors_io_out_s1_full_pred_is_br_sharing; // @[FrontendBundle.scala 430:48]
  wire  _s1_predicted_ghist_ptr_WIRE__0 = predictors_io_out_s1_full_pred_slot_valids_0; // @[FrontendBundle.scala 430:{12,12}]
  wire  _s1_predicted_ghist_ptr_T_4 = ~predictors_io_out_s1_full_pred_hit | ~(_s1_predicted_ghist_ptr_WIRE__0 |
    _s1_predicted_ghist_ptr_T_1); // @[FrontendBundle.scala 461:19]
  wire  _s1_predicted_ghist_ptr_T_6 = predictors_io_out_s1_full_pred_slot_valids_0 &
    predictors_io_out_s1_full_pred_br_taken_mask_0; // @[FrontendBundle.scala 435:69]
  wire  _s1_predicted_ghist_ptr_T_9 = predictors_io_out_s1_full_pred_is_br_sharing &
    predictors_io_out_s1_full_pred_br_taken_mask_1 | ~predictors_io_out_s1_full_pred_is_br_sharing; // @[FrontendBundle.scala 437:47]
  wire  _s1_predicted_ghist_ptr_T_10 = predictors_io_out_s1_full_pred_slot_valids_1 & _s1_predicted_ghist_ptr_T_9; // @[FrontendBundle.scala 436:25]
  wire  _s1_predicted_ghist_ptr_T_11 = _s1_predicted_ghist_ptr_T_6 & predictors_io_out_s1_full_pred_hit; // @[FrontendBundle.scala 450:32]
  wire  _s1_predicted_ghist_ptr_T_12 = _s1_predicted_ghist_ptr_T_10 & predictors_io_out_s1_full_pred_hit; // @[FrontendBundle.scala 450:32]
  wire  _s1_predicted_ghist_ptr_T_30 = _s1_predicted_ghist_ptr_T_11 | ~_s1_predicted_ghist_ptr_T_1; // @[FrontendBundle.scala 465:34]
  wire  _s1_predicted_ghist_ptr_T_31 = _s1_predicted_ghist_ptr_WIRE__0 & _s1_predicted_ghist_ptr_T_30; // @[FrontendBundle.scala 464:75]
  wire  _s1_predicted_ghist_ptr_T_32 = _s1_predicted_ghist_ptr_T_31 & predictors_io_out_s1_full_pred_hit; // @[FrontendBundle.scala 465:97]
  wire  _s1_predicted_ghist_ptr_T_44 = ~_s1_predicted_ghist_ptr_T_11; // @[FrontendBundle.scala 464:9]
  wire  _s1_predicted_ghist_ptr_T_45 = _s1_predicted_ghist_ptr_T_1 & _s1_predicted_ghist_ptr_T_44; // @[FrontendBundle.scala 463:22]
  wire  _s1_predicted_ghist_ptr_T_60 = _s1_predicted_ghist_ptr_T_45 & predictors_io_out_s1_full_pred_hit; // @[FrontendBundle.scala 465:97]
  wire [7:0] s1_possible_predicted_ghist_ptrs_flipped_new_ptr_value =
    _s1_possible_predicted_ghist_ptrs_flipped_new_ptr_new_ptr_value_T_1[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire [7:0] _s1_predicted_ghist_ptr_T_61 = _s1_predicted_ghist_ptr_T_4 ?
    s1_possible_predicted_ghist_ptrs_flipped_new_ptr_value : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] s1_possible_predicted_ghist_ptrs_flipped_new_ptr_1_value =
    _s1_possible_predicted_ghist_ptrs_flipped_new_ptr_new_ptr_value_T_3[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire [7:0] _s1_predicted_ghist_ptr_T_62 = _s1_predicted_ghist_ptr_T_32 ?
    s1_possible_predicted_ghist_ptrs_flipped_new_ptr_1_value : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] s1_possible_predicted_ghist_ptrs_flipped_new_ptr_2_value =
    _s1_possible_predicted_ghist_ptrs_flipped_new_ptr_new_ptr_value_T_5[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire [7:0] _s1_predicted_ghist_ptr_T_63 = _s1_predicted_ghist_ptr_T_60 ?
    s1_possible_predicted_ghist_ptrs_flipped_new_ptr_2_value : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _s1_predicted_ghist_ptr_T_64 = _s1_predicted_ghist_ptr_T_61 | _s1_predicted_ghist_ptr_T_62; // @[Mux.scala 27:73]
  wire  _s1_possible_predicted_fhs_T_5 = _s1_predicted_ghist_ptr_WIRE__0 &
    predictors_io_out_s1_full_pred_br_taken_mask_0 & predictors_io_out_s1_full_pred_hit | _s1_predicted_ghist_ptr_T_1 &
    predictors_io_out_s1_full_pred_br_taken_mask_1 & predictors_io_out_s1_full_pred_hit; // @[FrontendBundle.scala 470:90]
  wire  _s1_possible_predicted_fhs_T_67 = _s1_possible_predicted_fhs_T_5 & _s1_predicted_ghist_ptr_T_4; // @[BPU.scala 403:88]
  wire  s1_possible_predicted_fhs_ob__0 = s1_last_br_num_oh[0] & s1_ahead_fh_oldest_bits_afhob_3_bits_0 |
    s1_last_br_num_oh[1] & s1_ahead_fh_oldest_bits_afhob_3_bits_1 | s1_last_br_num_oh[2] &
    s1_ahead_fh_oldest_bits_afhob_3_bits_2; // @[Mux.scala 27:73]
  wire  s1_possible_predicted_fhs_ob__1 = s1_last_br_num_oh[0] & s1_ahead_fh_oldest_bits_afhob_3_bits_1 |
    s1_last_br_num_oh[1] & s1_ahead_fh_oldest_bits_afhob_3_bits_2 | s1_last_br_num_oh[2] &
    s1_ahead_fh_oldest_bits_afhob_3_bits_3; // @[Mux.scala 27:73]
  wire  s1_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__0 = s1_folded_gh_hist_0_folded_hist[0
    ]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__1 = s1_folded_gh_hist_0_folded_hist[1
    ]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__2 = s1_folded_gh_hist_0_folded_hist[2
    ]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__3 = s1_folded_gh_hist_0_folded_hist[3
    ]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__4 = s1_folded_gh_hist_0_folded_hist[4
    ]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__5 = s1_folded_gh_hist_0_folded_hist[5
    ]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__6 = s1_folded_gh_hist_0_folded_hist[6
    ]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__7 = s1_folded_gh_hist_0_folded_hist[7
    ]; // @[FrontendBundle.scala 280:54]
  wire [7:0] s1_possible_predicted_fhs_res_hist_0_new_folded_hist_xored = {
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__7,
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__6,
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__5,
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__4,
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__3,
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__1,
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [15:0] s1_possible_predicted_fhs_res_hist_0_new_folded_hist_src_doubled = {
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__7,
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__6,
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__5,
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__4,
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__3,
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__1,
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__0,
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_xored}; // @[Cat.scala 31:58]
  wire [7:0] s1_possible_predicted_fhs_res_hist_0_new_folded_hist =
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_src_doubled[15:8]; // @[FrontendBundle.scala 221:30]
  wire  s1_possible_predicted_fhs_ob_1_0 = s1_last_br_num_oh[0] & s1_ahead_fh_oldest_bits_afhob_2_bits_0 |
    s1_last_br_num_oh[1] & s1_ahead_fh_oldest_bits_afhob_2_bits_1 | s1_last_br_num_oh[2] &
    s1_ahead_fh_oldest_bits_afhob_2_bits_2; // @[Mux.scala 27:73]
  wire  s1_possible_predicted_fhs_ob_1_1 = s1_last_br_num_oh[0] & s1_ahead_fh_oldest_bits_afhob_2_bits_1 |
    s1_last_br_num_oh[1] & s1_ahead_fh_oldest_bits_afhob_2_bits_2 | s1_last_br_num_oh[2] &
    s1_ahead_fh_oldest_bits_afhob_2_bits_3; // @[Mux.scala 27:73]
  wire  s1_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__0 = s1_folded_gh_hist_1_folded_hist[0
    ]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__1 = s1_folded_gh_hist_1_folded_hist[1
    ]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__2 = s1_folded_gh_hist_1_folded_hist[2
    ]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__3 = s1_folded_gh_hist_1_folded_hist[3
    ]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__4 = s1_folded_gh_hist_1_folded_hist[4
    ]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__5 = s1_folded_gh_hist_1_folded_hist[5
    ]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__6 = s1_folded_gh_hist_1_folded_hist[6
    ]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__7 = s1_folded_gh_hist_1_folded_hist[7
    ]; // @[FrontendBundle.scala 280:54]
  wire [7:0] s1_possible_predicted_fhs_res_hist_1_new_folded_hist_xored = {
    s1_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__7,
    s1_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__6,
    s1_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__5,
    s1_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__4,
    s1_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__3,
    s1_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__1,
    s1_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [15:0] s1_possible_predicted_fhs_res_hist_1_new_folded_hist_src_doubled = {
    s1_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__7,
    s1_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__6,
    s1_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__5,
    s1_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__4,
    s1_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__3,
    s1_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__1,
    s1_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__0,
    s1_possible_predicted_fhs_res_hist_1_new_folded_hist_xored}; // @[Cat.scala 31:58]
  wire [7:0] s1_possible_predicted_fhs_res_hist_1_new_folded_hist =
    s1_possible_predicted_fhs_res_hist_1_new_folded_hist_src_doubled[15:8]; // @[FrontendBundle.scala 221:30]
  wire  s1_possible_predicted_fhs_ob_2_0 = s1_last_br_num_oh[0] & s1_ahead_fh_oldest_bits_afhob_5_bits_0 |
    s1_last_br_num_oh[1] & s1_ahead_fh_oldest_bits_afhob_5_bits_1 | s1_last_br_num_oh[2] &
    s1_ahead_fh_oldest_bits_afhob_5_bits_2; // @[Mux.scala 27:73]
  wire  s1_possible_predicted_fhs_ob_2_1 = s1_last_br_num_oh[0] & s1_ahead_fh_oldest_bits_afhob_5_bits_1 |
    s1_last_br_num_oh[1] & s1_ahead_fh_oldest_bits_afhob_5_bits_2 | s1_last_br_num_oh[2] &
    s1_ahead_fh_oldest_bits_afhob_5_bits_3; // @[Mux.scala 27:73]
  wire  s1_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__0 = s1_folded_gh_hist_2_folded_hist[0
    ]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__1 = s1_folded_gh_hist_2_folded_hist[1
    ]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__2 = s1_folded_gh_hist_2_folded_hist[2
    ]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__3 = s1_folded_gh_hist_2_folded_hist[3
    ]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__4 = s1_folded_gh_hist_2_folded_hist[4
    ]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__5 = s1_folded_gh_hist_2_folded_hist[5
    ]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__6 = s1_folded_gh_hist_2_folded_hist[6
    ]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__7 = s1_folded_gh_hist_2_folded_hist[7
    ]; // @[FrontendBundle.scala 280:54]
  wire [7:0] s1_possible_predicted_fhs_res_hist_2_new_folded_hist_xored = {
    s1_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__7,
    s1_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__6,
    s1_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__5,
    s1_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__4,
    s1_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__3,
    s1_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__1,
    s1_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [15:0] s1_possible_predicted_fhs_res_hist_2_new_folded_hist_src_doubled = {
    s1_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__7,
    s1_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__6,
    s1_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__5,
    s1_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__4,
    s1_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__3,
    s1_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__1,
    s1_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__0,
    s1_possible_predicted_fhs_res_hist_2_new_folded_hist_xored}; // @[Cat.scala 31:58]
  wire [7:0] s1_possible_predicted_fhs_res_hist_2_new_folded_hist =
    s1_possible_predicted_fhs_res_hist_2_new_folded_hist_src_doubled[15:8]; // @[FrontendBundle.scala 221:30]
  wire  s1_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__0 = s1_folded_gh_hist_3_folded_hist[0
    ]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__1 = s1_folded_gh_hist_3_folded_hist[1
    ]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__2 = s1_folded_gh_hist_3_folded_hist[2
    ]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__3 = s1_folded_gh_hist_3_folded_hist[3
    ]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__4 = s1_folded_gh_hist_3_folded_hist[4
    ]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__5 = s1_folded_gh_hist_3_folded_hist[5
    ]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__6 = s1_folded_gh_hist_3_folded_hist[6
    ]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__7 = s1_folded_gh_hist_3_folded_hist[7
    ]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__8 = s1_folded_gh_hist_3_folded_hist[8
    ]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__9 = s1_folded_gh_hist_3_folded_hist[9
    ]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__10 = s1_folded_gh_hist_3_folded_hist[
    10]; // @[FrontendBundle.scala 280:54]
  wire [4:0] s1_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_lo = {
    s1_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__4,
    s1_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__3,
    s1_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__1,
    s1_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [10:0] s1_possible_predicted_fhs_res_hist_3_new_folded_hist_xored = {
    s1_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__10,
    s1_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__9,
    s1_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__8,
    s1_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__7,
    s1_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__6,
    s1_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__5,
    s1_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_lo}; // @[FrontendBundle.scala 258:11]
  wire [21:0] s1_possible_predicted_fhs_res_hist_3_new_folded_hist_src_doubled = {
    s1_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__10,
    s1_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__9,
    s1_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__8,
    s1_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__7,
    s1_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__6,
    s1_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__5,
    s1_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_lo,
    s1_possible_predicted_fhs_res_hist_3_new_folded_hist_xored}; // @[Cat.scala 31:58]
  wire [10:0] s1_possible_predicted_fhs_res_hist_3_new_folded_hist =
    s1_possible_predicted_fhs_res_hist_3_new_folded_hist_src_doubled[21:11]; // @[FrontendBundle.scala 221:30]
  wire [3:0] _GEN_11910 = {{3'd0}, _s1_possible_predicted_fhs_T_67}; // @[FrontendBundle.scala 290:29]
  wire [3:0] s1_possible_predicted_fhs_res_hist_4_new_folded_hist = s1_folded_gh_hist_4_folded_hist | _GEN_11910; // @[FrontendBundle.scala 290:29]
  wire  s1_possible_predicted_fhs_ob_4_0 = s1_last_br_num_oh[0] & s1_ahead_fh_oldest_bits_afhob_1_bits_0 |
    s1_last_br_num_oh[1] & s1_ahead_fh_oldest_bits_afhob_1_bits_1 | s1_last_br_num_oh[2] &
    s1_ahead_fh_oldest_bits_afhob_1_bits_2; // @[Mux.scala 27:73]
  wire  s1_possible_predicted_fhs_ob_4_1 = s1_last_br_num_oh[0] & s1_ahead_fh_oldest_bits_afhob_1_bits_1 |
    s1_last_br_num_oh[1] & s1_ahead_fh_oldest_bits_afhob_1_bits_2 | s1_last_br_num_oh[2] &
    s1_ahead_fh_oldest_bits_afhob_1_bits_3; // @[Mux.scala 27:73]
  wire  s1_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__0 = s1_folded_gh_hist_5_folded_hist[0
    ]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__1 = s1_folded_gh_hist_5_folded_hist[1
    ]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__2 = s1_folded_gh_hist_5_folded_hist[2
    ]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__3 = s1_folded_gh_hist_5_folded_hist[3
    ]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__4 = s1_folded_gh_hist_5_folded_hist[4
    ]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__5 = s1_folded_gh_hist_5_folded_hist[5
    ]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__6 = s1_folded_gh_hist_5_folded_hist[6
    ]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__7 = s1_folded_gh_hist_5_folded_hist[7
    ]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__8 = s1_folded_gh_hist_5_folded_hist[8
    ]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__9 = s1_folded_gh_hist_5_folded_hist[9
    ]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__10 = s1_folded_gh_hist_5_folded_hist[
    10]; // @[FrontendBundle.scala 280:54]
  wire [4:0] s1_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_lo = {
    s1_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__4,
    s1_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__3,
    s1_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__1,
    s1_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [10:0] s1_possible_predicted_fhs_res_hist_5_new_folded_hist_xored = {
    s1_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__10,
    s1_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__9,
    s1_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__8,
    s1_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__7,
    s1_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__6,
    s1_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__5,
    s1_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_lo}; // @[FrontendBundle.scala 258:11]
  wire [21:0] s1_possible_predicted_fhs_res_hist_5_new_folded_hist_src_doubled = {
    s1_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__10,
    s1_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__9,
    s1_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__8,
    s1_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__7,
    s1_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__6,
    s1_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__5,
    s1_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_lo,
    s1_possible_predicted_fhs_res_hist_5_new_folded_hist_xored}; // @[Cat.scala 31:58]
  wire [10:0] s1_possible_predicted_fhs_res_hist_5_new_folded_hist =
    s1_possible_predicted_fhs_res_hist_5_new_folded_hist_src_doubled[21:11]; // @[FrontendBundle.scala 221:30]
  wire  s1_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__0 = s1_folded_gh_hist_6_folded_hist[0
    ]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__1 = s1_folded_gh_hist_6_folded_hist[1
    ]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__2 = s1_folded_gh_hist_6_folded_hist[2
    ]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__3 = s1_folded_gh_hist_6_folded_hist[3
    ]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__4 = s1_folded_gh_hist_6_folded_hist[4
    ]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__5 = s1_folded_gh_hist_6_folded_hist[5
    ]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__6 = s1_folded_gh_hist_6_folded_hist[6
    ]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__7 = s1_folded_gh_hist_6_folded_hist[7
    ]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__8 = s1_folded_gh_hist_6_folded_hist[8
    ]; // @[FrontendBundle.scala 280:54]
  wire [8:0] s1_possible_predicted_fhs_res_hist_6_new_folded_hist_xored = {
    s1_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__8,
    s1_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__7,
    s1_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__6,
    s1_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__5,
    s1_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__4,
    s1_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__3,
    s1_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__1,
    s1_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [17:0] s1_possible_predicted_fhs_res_hist_6_new_folded_hist_src_doubled = {
    s1_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__8,
    s1_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__7,
    s1_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__6,
    s1_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__5,
    s1_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__4,
    s1_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__3,
    s1_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__1,
    s1_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__0,
    s1_possible_predicted_fhs_res_hist_6_new_folded_hist_xored}; // @[Cat.scala 31:58]
  wire [8:0] s1_possible_predicted_fhs_res_hist_6_new_folded_hist =
    s1_possible_predicted_fhs_res_hist_6_new_folded_hist_src_doubled[17:9]; // @[FrontendBundle.scala 221:30]
  wire  s1_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__0 = s1_folded_gh_hist_7_folded_hist[0
    ]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__1 = s1_folded_gh_hist_7_folded_hist[1
    ]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__2 = s1_folded_gh_hist_7_folded_hist[2
    ]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__3 = s1_folded_gh_hist_7_folded_hist[3
    ]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__4 = s1_folded_gh_hist_7_folded_hist[4
    ]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__5 = s1_folded_gh_hist_7_folded_hist[5
    ]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__6 = s1_folded_gh_hist_7_folded_hist[6
    ]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__7 = s1_folded_gh_hist_7_folded_hist[7
    ]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__8 = s1_folded_gh_hist_7_folded_hist[8
    ]; // @[FrontendBundle.scala 280:54]
  wire [8:0] s1_possible_predicted_fhs_res_hist_7_new_folded_hist_xored = {
    s1_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__8,
    s1_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__7,
    s1_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__6,
    s1_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__5,
    s1_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__4,
    s1_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__3,
    s1_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__1,
    s1_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [17:0] s1_possible_predicted_fhs_res_hist_7_new_folded_hist_src_doubled = {
    s1_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__8,
    s1_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__7,
    s1_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__6,
    s1_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__5,
    s1_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__4,
    s1_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__3,
    s1_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__1,
    s1_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__0,
    s1_possible_predicted_fhs_res_hist_7_new_folded_hist_xored}; // @[Cat.scala 31:58]
  wire [8:0] s1_possible_predicted_fhs_res_hist_7_new_folded_hist =
    s1_possible_predicted_fhs_res_hist_7_new_folded_hist_src_doubled[17:9]; // @[FrontendBundle.scala 221:30]
  wire [7:0] _GEN_11911 = {{7'd0}, _s1_possible_predicted_fhs_T_67}; // @[FrontendBundle.scala 290:29]
  wire [7:0] s1_possible_predicted_fhs_res_hist_8_new_folded_hist = s1_folded_gh_hist_8_folded_hist | _GEN_11911; // @[FrontendBundle.scala 290:29]
  wire  s1_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__0 = s1_folded_gh_hist_9_folded_hist[0
    ]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__1 = s1_folded_gh_hist_9_folded_hist[1
    ]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__2 = s1_folded_gh_hist_9_folded_hist[2
    ]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__3 = s1_folded_gh_hist_9_folded_hist[3
    ]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__4 = s1_folded_gh_hist_9_folded_hist[4
    ]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__5 = s1_folded_gh_hist_9_folded_hist[5
    ]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__6 = s1_folded_gh_hist_9_folded_hist[6
    ]; // @[FrontendBundle.scala 280:54]
  wire [6:0] s1_possible_predicted_fhs_res_hist_9_new_folded_hist_xored = {
    s1_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__6,
    s1_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__5,
    s1_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__4,
    s1_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__3,
    s1_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__1,
    s1_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [13:0] s1_possible_predicted_fhs_res_hist_9_new_folded_hist_src_doubled = {
    s1_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__6,
    s1_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__5,
    s1_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__4,
    s1_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__3,
    s1_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__1,
    s1_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__0,
    s1_possible_predicted_fhs_res_hist_9_new_folded_hist_xored}; // @[Cat.scala 31:58]
  wire [6:0] s1_possible_predicted_fhs_res_hist_9_new_folded_hist =
    s1_possible_predicted_fhs_res_hist_9_new_folded_hist_src_doubled[13:7]; // @[FrontendBundle.scala 221:30]
  wire  s1_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__0 = s1_folded_gh_hist_10_folded_hist
    [0]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__1 = s1_folded_gh_hist_10_folded_hist
    [1]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__2 = s1_folded_gh_hist_10_folded_hist
    [2]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__3 = s1_folded_gh_hist_10_folded_hist
    [3]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__4 = s1_folded_gh_hist_10_folded_hist
    [4]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__5 = s1_folded_gh_hist_10_folded_hist
    [5]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__6 = s1_folded_gh_hist_10_folded_hist
    [6]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__7 = s1_folded_gh_hist_10_folded_hist
    [7]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__8 = s1_folded_gh_hist_10_folded_hist
    [8]; // @[FrontendBundle.scala 280:54]
  wire [8:0] s1_possible_predicted_fhs_res_hist_10_new_folded_hist_xored = {
    s1_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__8,
    s1_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__7,
    s1_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__6,
    s1_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__5,
    s1_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__4,
    s1_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__3,
    s1_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__1,
    s1_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [17:0] s1_possible_predicted_fhs_res_hist_10_new_folded_hist_src_doubled = {
    s1_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__8,
    s1_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__7,
    s1_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__6,
    s1_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__5,
    s1_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__4,
    s1_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__3,
    s1_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__1,
    s1_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__0,
    s1_possible_predicted_fhs_res_hist_10_new_folded_hist_xored}; // @[Cat.scala 31:58]
  wire [8:0] s1_possible_predicted_fhs_res_hist_10_new_folded_hist =
    s1_possible_predicted_fhs_res_hist_10_new_folded_hist_src_doubled[17:9]; // @[FrontendBundle.scala 221:30]
  wire [7:0] s1_possible_predicted_fhs_res_hist_11_new_folded_hist = s1_folded_gh_hist_11_folded_hist | _GEN_11911; // @[FrontendBundle.scala 290:29]
  wire  s1_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__0 = s1_folded_gh_hist_12_folded_hist
    [0]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__1 = s1_folded_gh_hist_12_folded_hist
    [1]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__2 = s1_folded_gh_hist_12_folded_hist
    [2]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__3 = s1_folded_gh_hist_12_folded_hist
    [3]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__4 = s1_folded_gh_hist_12_folded_hist
    [4]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__5 = s1_folded_gh_hist_12_folded_hist
    [5]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__6 = s1_folded_gh_hist_12_folded_hist
    [6]; // @[FrontendBundle.scala 280:54]
  wire [6:0] s1_possible_predicted_fhs_res_hist_12_new_folded_hist_xored = {
    s1_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__6,
    s1_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__5,
    s1_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__4,
    s1_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__3,
    s1_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__1,
    s1_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [13:0] s1_possible_predicted_fhs_res_hist_12_new_folded_hist_src_doubled = {
    s1_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__6,
    s1_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__5,
    s1_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__4,
    s1_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__3,
    s1_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__1,
    s1_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__0,
    s1_possible_predicted_fhs_res_hist_12_new_folded_hist_xored}; // @[Cat.scala 31:58]
  wire [6:0] s1_possible_predicted_fhs_res_hist_12_new_folded_hist =
    s1_possible_predicted_fhs_res_hist_12_new_folded_hist_src_doubled[13:7]; // @[FrontendBundle.scala 221:30]
  wire  s1_possible_predicted_fhs_ob_10_0 = s1_last_br_num_oh[0] & s1_ahead_fh_oldest_bits_afhob_4_bits_0 |
    s1_last_br_num_oh[1] & s1_ahead_fh_oldest_bits_afhob_4_bits_1 | s1_last_br_num_oh[2] &
    s1_ahead_fh_oldest_bits_afhob_4_bits_2; // @[Mux.scala 27:73]
  wire  s1_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__0 = s1_folded_gh_hist_13_folded_hist
    [0]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__1 = s1_folded_gh_hist_13_folded_hist
    [1]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__2 = s1_folded_gh_hist_13_folded_hist
    [2]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__3 = s1_folded_gh_hist_13_folded_hist
    [3]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__4 = s1_folded_gh_hist_13_folded_hist
    [4]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__5 = s1_folded_gh_hist_13_folded_hist
    [5]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__6 = s1_folded_gh_hist_13_folded_hist
    [6]; // @[FrontendBundle.scala 280:54]
  wire [6:0] s1_possible_predicted_fhs_res_hist_13_new_folded_hist_xored = {
    s1_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__6,
    s1_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__5,
    s1_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__4,
    s1_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__3,
    s1_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__1,
    s1_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [13:0] s1_possible_predicted_fhs_res_hist_13_new_folded_hist_src_doubled = {
    s1_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__6,
    s1_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__5,
    s1_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__4,
    s1_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__3,
    s1_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__1,
    s1_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__0,
    s1_possible_predicted_fhs_res_hist_13_new_folded_hist_xored}; // @[Cat.scala 31:58]
  wire [6:0] s1_possible_predicted_fhs_res_hist_13_new_folded_hist =
    s1_possible_predicted_fhs_res_hist_13_new_folded_hist_src_doubled[13:7]; // @[FrontendBundle.scala 221:30]
  wire  s1_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__0 = s1_folded_gh_hist_14_folded_hist
    [0]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__1 = s1_folded_gh_hist_14_folded_hist
    [1]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__2 = s1_folded_gh_hist_14_folded_hist
    [2]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__3 = s1_folded_gh_hist_14_folded_hist
    [3]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__4 = s1_folded_gh_hist_14_folded_hist
    [4]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__5 = s1_folded_gh_hist_14_folded_hist
    [5]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__6 = s1_folded_gh_hist_14_folded_hist
    [6]; // @[FrontendBundle.scala 280:54]
  wire [6:0] s1_possible_predicted_fhs_res_hist_14_new_folded_hist_xored = {
    s1_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__6,
    s1_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__5,
    s1_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__4,
    s1_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__3,
    s1_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__1,
    s1_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [13:0] s1_possible_predicted_fhs_res_hist_14_new_folded_hist_src_doubled = {
    s1_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__6,
    s1_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__5,
    s1_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__4,
    s1_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__3,
    s1_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__1,
    s1_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__0,
    s1_possible_predicted_fhs_res_hist_14_new_folded_hist_xored}; // @[Cat.scala 31:58]
  wire [6:0] s1_possible_predicted_fhs_res_hist_14_new_folded_hist =
    s1_possible_predicted_fhs_res_hist_14_new_folded_hist_src_doubled[13:7]; // @[FrontendBundle.scala 221:30]
  wire  s1_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__0 = s1_folded_gh_hist_15_folded_hist
    [0]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__1 = s1_folded_gh_hist_15_folded_hist
    [1]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__2 = s1_folded_gh_hist_15_folded_hist
    [2]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__3 = s1_folded_gh_hist_15_folded_hist
    [3]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__4 = s1_folded_gh_hist_15_folded_hist
    [4]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__5 = s1_folded_gh_hist_15_folded_hist
    [5]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__6 = s1_folded_gh_hist_15_folded_hist
    [6]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__7 = s1_folded_gh_hist_15_folded_hist
    [7]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__8 = s1_folded_gh_hist_15_folded_hist
    [8]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__9 = s1_folded_gh_hist_15_folded_hist
    [9]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__10 =
    s1_folded_gh_hist_15_folded_hist[10]; // @[FrontendBundle.scala 280:54]
  wire [4:0] s1_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_lo = {
    s1_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__4,
    s1_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__3,
    s1_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__1,
    s1_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [10:0] s1_possible_predicted_fhs_res_hist_15_new_folded_hist_xored = {
    s1_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__10,
    s1_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__9,
    s1_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__8,
    s1_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__7,
    s1_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__6,
    s1_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__5,
    s1_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_lo}; // @[FrontendBundle.scala 258:11]
  wire [21:0] s1_possible_predicted_fhs_res_hist_15_new_folded_hist_src_doubled = {
    s1_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__10,
    s1_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__9,
    s1_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__8,
    s1_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__7,
    s1_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__6,
    s1_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__5,
    s1_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_lo,
    s1_possible_predicted_fhs_res_hist_15_new_folded_hist_xored}; // @[Cat.scala 31:58]
  wire [10:0] s1_possible_predicted_fhs_res_hist_15_new_folded_hist =
    s1_possible_predicted_fhs_res_hist_15_new_folded_hist_src_doubled[21:11]; // @[FrontendBundle.scala 221:30]
  wire  s1_possible_predicted_fhs_ob_13_0 = s1_last_br_num_oh[0] & s1_ahead_fh_oldest_bits_afhob_0_bits_0 |
    s1_last_br_num_oh[1] & s1_ahead_fh_oldest_bits_afhob_0_bits_1 | s1_last_br_num_oh[2] &
    s1_ahead_fh_oldest_bits_afhob_0_bits_2; // @[Mux.scala 27:73]
  wire  s1_possible_predicted_fhs_ob_13_1 = s1_last_br_num_oh[0] & s1_ahead_fh_oldest_bits_afhob_0_bits_1 |
    s1_last_br_num_oh[1] & s1_ahead_fh_oldest_bits_afhob_0_bits_2 | s1_last_br_num_oh[2] &
    s1_ahead_fh_oldest_bits_afhob_0_bits_3; // @[Mux.scala 27:73]
  wire  s1_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__0 = s1_folded_gh_hist_16_folded_hist
    [0]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__1 = s1_folded_gh_hist_16_folded_hist
    [1]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__2 = s1_folded_gh_hist_16_folded_hist
    [2]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__3 = s1_folded_gh_hist_16_folded_hist
    [3]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__4 = s1_folded_gh_hist_16_folded_hist
    [4]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__5 = s1_folded_gh_hist_16_folded_hist
    [5]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__6 = s1_folded_gh_hist_16_folded_hist
    [6]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__7 = s1_folded_gh_hist_16_folded_hist
    [7]; // @[FrontendBundle.scala 280:54]
  wire [7:0] s1_possible_predicted_fhs_res_hist_16_new_folded_hist_xored = {
    s1_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__7,
    s1_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__6,
    s1_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__5,
    s1_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__4,
    s1_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__3,
    s1_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__1,
    s1_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [15:0] s1_possible_predicted_fhs_res_hist_16_new_folded_hist_src_doubled = {
    s1_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__7,
    s1_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__6,
    s1_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__5,
    s1_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__4,
    s1_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__3,
    s1_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__1,
    s1_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__0,
    s1_possible_predicted_fhs_res_hist_16_new_folded_hist_xored}; // @[Cat.scala 31:58]
  wire [7:0] s1_possible_predicted_fhs_res_hist_16_new_folded_hist =
    s1_possible_predicted_fhs_res_hist_16_new_folded_hist_src_doubled[15:8]; // @[FrontendBundle.scala 221:30]
  wire  s1_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__0 = s1_folded_gh_hist_17_folded_hist
    [0]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__1 = s1_folded_gh_hist_17_folded_hist
    [1]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__2 = s1_folded_gh_hist_17_folded_hist
    [2]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__3 = s1_folded_gh_hist_17_folded_hist
    [3]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__4 = s1_folded_gh_hist_17_folded_hist
    [4]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__5 = s1_folded_gh_hist_17_folded_hist
    [5]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__6 = s1_folded_gh_hist_17_folded_hist
    [6]; // @[FrontendBundle.scala 280:54]
  wire  s1_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__7 = s1_folded_gh_hist_17_folded_hist
    [7]; // @[FrontendBundle.scala 280:54]
  wire [7:0] s1_possible_predicted_fhs_res_hist_17_new_folded_hist_xored = {
    s1_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__7,
    s1_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__6,
    s1_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__5,
    s1_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__4,
    s1_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__3,
    s1_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__1,
    s1_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [15:0] s1_possible_predicted_fhs_res_hist_17_new_folded_hist_src_doubled = {
    s1_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__7,
    s1_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__6,
    s1_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__5,
    s1_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__4,
    s1_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__3,
    s1_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__1,
    s1_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__0,
    s1_possible_predicted_fhs_res_hist_17_new_folded_hist_xored}; // @[Cat.scala 31:58]
  wire [7:0] s1_possible_predicted_fhs_res_hist_17_new_folded_hist =
    s1_possible_predicted_fhs_res_hist_17_new_folded_hist_src_doubled[15:8]; // @[FrontendBundle.scala 221:30]
  wire  _s1_possible_predicted_fhs_T_135 = _s1_possible_predicted_fhs_T_5 & _s1_predicted_ghist_ptr_T_32; // @[BPU.scala 403:88]
  wire [1:0] s1_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1 = {1'h0,
    _s1_possible_predicted_fhs_T_135}; // @[FrontendBundle.scala 274:102]
  wire  s1_possible_predicted_fhs_res_hist_0_new_folded_hist_xored_res_1_6 =
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[1] ^
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__6; // @[FrontendBundle.scala 256:48]
  wire  s1_possible_predicted_fhs_res_hist_0_new_folded_hist_xored_res_1_7 =
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[0] ^ s1_possible_predicted_fhs_ob__0 ^
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__7; // @[FrontendBundle.scala 256:48]
  wire [7:0] s1_possible_predicted_fhs_res_hist_0_new_folded_hist_xored_1 = {
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_xored_res_1_7,
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_xored_res_1_6,
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__5,
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__4,
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__3,
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__1,
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [15:0] s1_possible_predicted_fhs_res_hist_0_new_folded_hist_src_doubled_1 = {
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_xored_res_1_7,
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_xored_res_1_6,
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__5,
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__4,
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__3,
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__1,
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__0,
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_xored_1}; // @[Cat.scala 31:58]
  wire [7:0] s1_possible_predicted_fhs_res_hist_0_new_folded_hist_1 =
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_src_doubled_1[14:7]; // @[FrontendBundle.scala 221:30]
  wire  s1_possible_predicted_fhs_res_hist_1_new_folded_hist_xored_res_1_6 =
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[1] ^
    s1_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__6; // @[FrontendBundle.scala 256:48]
  wire  s1_possible_predicted_fhs_res_hist_1_new_folded_hist_xored_res_1_7 =
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[0] ^ s1_possible_predicted_fhs_ob_1_0 ^
    s1_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__7; // @[FrontendBundle.scala 256:48]
  wire [7:0] s1_possible_predicted_fhs_res_hist_1_new_folded_hist_xored_1 = {
    s1_possible_predicted_fhs_res_hist_1_new_folded_hist_xored_res_1_7,
    s1_possible_predicted_fhs_res_hist_1_new_folded_hist_xored_res_1_6,
    s1_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__5,
    s1_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__4,
    s1_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__3,
    s1_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__1,
    s1_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [15:0] s1_possible_predicted_fhs_res_hist_1_new_folded_hist_src_doubled_1 = {
    s1_possible_predicted_fhs_res_hist_1_new_folded_hist_xored_res_1_7,
    s1_possible_predicted_fhs_res_hist_1_new_folded_hist_xored_res_1_6,
    s1_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__5,
    s1_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__4,
    s1_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__3,
    s1_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__1,
    s1_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__0,
    s1_possible_predicted_fhs_res_hist_1_new_folded_hist_xored_1}; // @[Cat.scala 31:58]
  wire [7:0] s1_possible_predicted_fhs_res_hist_1_new_folded_hist_1 =
    s1_possible_predicted_fhs_res_hist_1_new_folded_hist_src_doubled_1[14:7]; // @[FrontendBundle.scala 221:30]
  wire  s1_possible_predicted_fhs_res_hist_2_new_folded_hist_xored_res_1_6 =
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[1] ^ s1_possible_predicted_fhs_ob_2_0 ^
    s1_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__6; // @[FrontendBundle.scala 256:48]
  wire  s1_possible_predicted_fhs_res_hist_2_new_folded_hist_xored_res_1_7 =
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[0] ^
    s1_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__7; // @[FrontendBundle.scala 256:48]
  wire [7:0] s1_possible_predicted_fhs_res_hist_2_new_folded_hist_xored_1 = {
    s1_possible_predicted_fhs_res_hist_2_new_folded_hist_xored_res_1_7,
    s1_possible_predicted_fhs_res_hist_2_new_folded_hist_xored_res_1_6,
    s1_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__5,
    s1_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__4,
    s1_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__3,
    s1_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__1,
    s1_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [15:0] s1_possible_predicted_fhs_res_hist_2_new_folded_hist_src_doubled_1 = {
    s1_possible_predicted_fhs_res_hist_2_new_folded_hist_xored_res_1_7,
    s1_possible_predicted_fhs_res_hist_2_new_folded_hist_xored_res_1_6,
    s1_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__5,
    s1_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__4,
    s1_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__3,
    s1_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__1,
    s1_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__0,
    s1_possible_predicted_fhs_res_hist_2_new_folded_hist_xored_1}; // @[Cat.scala 31:58]
  wire [7:0] s1_possible_predicted_fhs_res_hist_2_new_folded_hist_1 =
    s1_possible_predicted_fhs_res_hist_2_new_folded_hist_src_doubled_1[14:7]; // @[FrontendBundle.scala 221:30]
  wire  s1_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_res_1_9 =
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[1] ^ s1_possible_predicted_fhs_ob_1_0 ^
    s1_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__9; // @[FrontendBundle.scala 256:48]
  wire  s1_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_res_1_10 =
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[0] ^
    s1_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__10; // @[FrontendBundle.scala 256:48]
  wire [10:0] s1_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_1 = {
    s1_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_res_1_10,
    s1_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_res_1_9,
    s1_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__8,
    s1_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__7,
    s1_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__6,
    s1_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__5,
    s1_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_lo}; // @[FrontendBundle.scala 258:11]
  wire [21:0] s1_possible_predicted_fhs_res_hist_3_new_folded_hist_src_doubled_1 = {
    s1_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_res_1_10,
    s1_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_res_1_9,
    s1_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__8,
    s1_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__7,
    s1_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__6,
    s1_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__5,
    s1_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_lo,
    s1_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_1}; // @[Cat.scala 31:58]
  wire [10:0] s1_possible_predicted_fhs_res_hist_3_new_folded_hist_1 =
    s1_possible_predicted_fhs_res_hist_3_new_folded_hist_src_doubled_1[20:10]; // @[FrontendBundle.scala 221:30]
  wire [4:0] _s1_possible_predicted_fhs_res_hist_4_new_folded_hist_T_2 = {s1_folded_gh_hist_4_folded_hist, 1'h0}; // @[FrontendBundle.scala 290:21]
  wire [4:0] _GEN_11913 = {{4'd0}, _s1_possible_predicted_fhs_T_135}; // @[FrontendBundle.scala 290:29]
  wire [4:0] _s1_possible_predicted_fhs_res_hist_4_new_folded_hist_T_3 =
    _s1_possible_predicted_fhs_res_hist_4_new_folded_hist_T_2 | _GEN_11913; // @[FrontendBundle.scala 290:29]
  wire [3:0] s1_possible_predicted_fhs_res_hist_4_new_folded_hist_1 =
    _s1_possible_predicted_fhs_res_hist_4_new_folded_hist_T_3[3:0]; // @[FrontendBundle.scala 290:37]
  wire  s1_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_res_1_1 = s1_possible_predicted_fhs_ob_4_0 ^
    s1_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__1; // @[FrontendBundle.scala 256:48]
  wire  s1_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_res_1_9 =
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[1] ^
    s1_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__9; // @[FrontendBundle.scala 256:48]
  wire  s1_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_res_1_10 =
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[0] ^
    s1_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__10; // @[FrontendBundle.scala 256:48]
  wire [4:0] s1_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_lo_1 = {
    s1_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__4,
    s1_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__3,
    s1_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_res_1_1,
    s1_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [10:0] s1_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_1 = {
    s1_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_res_1_10,
    s1_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_res_1_9,
    s1_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__8,
    s1_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__7,
    s1_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__6,
    s1_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__5,
    s1_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_lo_1}; // @[FrontendBundle.scala 258:11]
  wire [21:0] s1_possible_predicted_fhs_res_hist_5_new_folded_hist_src_doubled_1 = {
    s1_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_res_1_10,
    s1_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_res_1_9,
    s1_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__8,
    s1_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__7,
    s1_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__6,
    s1_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__5,
    s1_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_lo_1,
    s1_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_1}; // @[Cat.scala 31:58]
  wire [10:0] s1_possible_predicted_fhs_res_hist_5_new_folded_hist_1 =
    s1_possible_predicted_fhs_res_hist_5_new_folded_hist_src_doubled_1[20:10]; // @[FrontendBundle.scala 221:30]
  wire  s1_possible_predicted_fhs_res_hist_6_new_folded_hist_xored_res_1_3 = s1_possible_predicted_fhs_ob_4_0 ^
    s1_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__3; // @[FrontendBundle.scala 256:48]
  wire  s1_possible_predicted_fhs_res_hist_6_new_folded_hist_xored_res_1_7 =
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[1] ^
    s1_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__7; // @[FrontendBundle.scala 256:48]
  wire  s1_possible_predicted_fhs_res_hist_6_new_folded_hist_xored_res_1_8 =
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[0] ^
    s1_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__8; // @[FrontendBundle.scala 256:48]
  wire [8:0] s1_possible_predicted_fhs_res_hist_6_new_folded_hist_xored_1 = {
    s1_possible_predicted_fhs_res_hist_6_new_folded_hist_xored_res_1_8,
    s1_possible_predicted_fhs_res_hist_6_new_folded_hist_xored_res_1_7,
    s1_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__6,
    s1_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__5,
    s1_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__4,
    s1_possible_predicted_fhs_res_hist_6_new_folded_hist_xored_res_1_3,
    s1_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__1,
    s1_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [17:0] s1_possible_predicted_fhs_res_hist_6_new_folded_hist_src_doubled_1 = {
    s1_possible_predicted_fhs_res_hist_6_new_folded_hist_xored_res_1_8,
    s1_possible_predicted_fhs_res_hist_6_new_folded_hist_xored_res_1_7,
    s1_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__6,
    s1_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__5,
    s1_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__4,
    s1_possible_predicted_fhs_res_hist_6_new_folded_hist_xored_res_1_3,
    s1_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__1,
    s1_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__0,
    s1_possible_predicted_fhs_res_hist_6_new_folded_hist_xored_1}; // @[Cat.scala 31:58]
  wire [8:0] s1_possible_predicted_fhs_res_hist_6_new_folded_hist_1 =
    s1_possible_predicted_fhs_res_hist_6_new_folded_hist_src_doubled_1[16:8]; // @[FrontendBundle.scala 221:30]
  wire  s1_possible_predicted_fhs_res_hist_7_new_folded_hist_xored_res_1_6 = s1_possible_predicted_fhs_ob__0 ^
    s1_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__6; // @[FrontendBundle.scala 256:48]
  wire  s1_possible_predicted_fhs_res_hist_7_new_folded_hist_xored_res_1_7 =
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[1] ^
    s1_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__7; // @[FrontendBundle.scala 256:48]
  wire  s1_possible_predicted_fhs_res_hist_7_new_folded_hist_xored_res_1_8 =
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[0] ^
    s1_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__8; // @[FrontendBundle.scala 256:48]
  wire [8:0] s1_possible_predicted_fhs_res_hist_7_new_folded_hist_xored_1 = {
    s1_possible_predicted_fhs_res_hist_7_new_folded_hist_xored_res_1_8,
    s1_possible_predicted_fhs_res_hist_7_new_folded_hist_xored_res_1_7,
    s1_possible_predicted_fhs_res_hist_7_new_folded_hist_xored_res_1_6,
    s1_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__5,
    s1_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__4,
    s1_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__3,
    s1_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__1,
    s1_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [17:0] s1_possible_predicted_fhs_res_hist_7_new_folded_hist_src_doubled_1 = {
    s1_possible_predicted_fhs_res_hist_7_new_folded_hist_xored_res_1_8,
    s1_possible_predicted_fhs_res_hist_7_new_folded_hist_xored_res_1_7,
    s1_possible_predicted_fhs_res_hist_7_new_folded_hist_xored_res_1_6,
    s1_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__5,
    s1_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__4,
    s1_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__3,
    s1_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__1,
    s1_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__0,
    s1_possible_predicted_fhs_res_hist_7_new_folded_hist_xored_1}; // @[Cat.scala 31:58]
  wire [8:0] s1_possible_predicted_fhs_res_hist_7_new_folded_hist_1 =
    s1_possible_predicted_fhs_res_hist_7_new_folded_hist_src_doubled_1[16:8]; // @[FrontendBundle.scala 221:30]
  wire [8:0] _s1_possible_predicted_fhs_res_hist_8_new_folded_hist_T_2 = {s1_folded_gh_hist_8_folded_hist, 1'h0}; // @[FrontendBundle.scala 290:21]
  wire [8:0] _GEN_11914 = {{8'd0}, _s1_possible_predicted_fhs_T_135}; // @[FrontendBundle.scala 290:29]
  wire [8:0] _s1_possible_predicted_fhs_res_hist_8_new_folded_hist_T_3 =
    _s1_possible_predicted_fhs_res_hist_8_new_folded_hist_T_2 | _GEN_11914; // @[FrontendBundle.scala 290:29]
  wire [7:0] s1_possible_predicted_fhs_res_hist_8_new_folded_hist_1 =
    _s1_possible_predicted_fhs_res_hist_8_new_folded_hist_T_3[7:0]; // @[FrontendBundle.scala 290:37]
  wire  s1_possible_predicted_fhs_res_hist_9_new_folded_hist_xored_res_1_3 = s1_possible_predicted_fhs_ob_1_0 ^
    s1_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__3; // @[FrontendBundle.scala 256:48]
  wire  s1_possible_predicted_fhs_res_hist_9_new_folded_hist_xored_res_1_5 =
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[1] ^
    s1_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__5; // @[FrontendBundle.scala 256:48]
  wire  s1_possible_predicted_fhs_res_hist_9_new_folded_hist_xored_res_1_6 =
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[0] ^
    s1_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__6; // @[FrontendBundle.scala 256:48]
  wire [6:0] s1_possible_predicted_fhs_res_hist_9_new_folded_hist_xored_1 = {
    s1_possible_predicted_fhs_res_hist_9_new_folded_hist_xored_res_1_6,
    s1_possible_predicted_fhs_res_hist_9_new_folded_hist_xored_res_1_5,
    s1_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__4,
    s1_possible_predicted_fhs_res_hist_9_new_folded_hist_xored_res_1_3,
    s1_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__1,
    s1_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [13:0] s1_possible_predicted_fhs_res_hist_9_new_folded_hist_src_doubled_1 = {
    s1_possible_predicted_fhs_res_hist_9_new_folded_hist_xored_res_1_6,
    s1_possible_predicted_fhs_res_hist_9_new_folded_hist_xored_res_1_5,
    s1_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__4,
    s1_possible_predicted_fhs_res_hist_9_new_folded_hist_xored_res_1_3,
    s1_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__1,
    s1_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__0,
    s1_possible_predicted_fhs_res_hist_9_new_folded_hist_xored_1}; // @[Cat.scala 31:58]
  wire [6:0] s1_possible_predicted_fhs_res_hist_9_new_folded_hist_1 =
    s1_possible_predicted_fhs_res_hist_9_new_folded_hist_src_doubled_1[12:6]; // @[FrontendBundle.scala 221:30]
  wire  s1_possible_predicted_fhs_res_hist_10_new_folded_hist_xored_res_1_4 = s1_possible_predicted_fhs_ob_1_0 ^
    s1_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__4; // @[FrontendBundle.scala 256:48]
  wire  s1_possible_predicted_fhs_res_hist_10_new_folded_hist_xored_res_1_7 =
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[1] ^
    s1_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__7; // @[FrontendBundle.scala 256:48]
  wire  s1_possible_predicted_fhs_res_hist_10_new_folded_hist_xored_res_1_8 =
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[0] ^
    s1_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__8; // @[FrontendBundle.scala 256:48]
  wire [8:0] s1_possible_predicted_fhs_res_hist_10_new_folded_hist_xored_1 = {
    s1_possible_predicted_fhs_res_hist_10_new_folded_hist_xored_res_1_8,
    s1_possible_predicted_fhs_res_hist_10_new_folded_hist_xored_res_1_7,
    s1_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__6,
    s1_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__5,
    s1_possible_predicted_fhs_res_hist_10_new_folded_hist_xored_res_1_4,
    s1_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__3,
    s1_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__1,
    s1_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [17:0] s1_possible_predicted_fhs_res_hist_10_new_folded_hist_src_doubled_1 = {
    s1_possible_predicted_fhs_res_hist_10_new_folded_hist_xored_res_1_8,
    s1_possible_predicted_fhs_res_hist_10_new_folded_hist_xored_res_1_7,
    s1_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__6,
    s1_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__5,
    s1_possible_predicted_fhs_res_hist_10_new_folded_hist_xored_res_1_4,
    s1_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__3,
    s1_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__1,
    s1_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__0,
    s1_possible_predicted_fhs_res_hist_10_new_folded_hist_xored_1}; // @[Cat.scala 31:58]
  wire [8:0] s1_possible_predicted_fhs_res_hist_10_new_folded_hist_1 =
    s1_possible_predicted_fhs_res_hist_10_new_folded_hist_src_doubled_1[16:8]; // @[FrontendBundle.scala 221:30]
  wire [8:0] _s1_possible_predicted_fhs_res_hist_11_new_folded_hist_T_2 = {s1_folded_gh_hist_11_folded_hist, 1'h0}; // @[FrontendBundle.scala 290:21]
  wire [8:0] _s1_possible_predicted_fhs_res_hist_11_new_folded_hist_T_3 =
    _s1_possible_predicted_fhs_res_hist_11_new_folded_hist_T_2 | _GEN_11914; // @[FrontendBundle.scala 290:29]
  wire [7:0] s1_possible_predicted_fhs_res_hist_11_new_folded_hist_1 =
    _s1_possible_predicted_fhs_res_hist_11_new_folded_hist_T_3[7:0]; // @[FrontendBundle.scala 290:37]
  wire  s1_possible_predicted_fhs_res_hist_12_new_folded_hist_xored_res_1_5 =
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[1] ^ s1_possible_predicted_fhs_ob_4_0 ^
    s1_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__5; // @[FrontendBundle.scala 256:48]
  wire  s1_possible_predicted_fhs_res_hist_12_new_folded_hist_xored_res_1_6 =
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[0] ^
    s1_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__6; // @[FrontendBundle.scala 256:48]
  wire [6:0] s1_possible_predicted_fhs_res_hist_12_new_folded_hist_xored_1 = {
    s1_possible_predicted_fhs_res_hist_12_new_folded_hist_xored_res_1_6,
    s1_possible_predicted_fhs_res_hist_12_new_folded_hist_xored_res_1_5,
    s1_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__4,
    s1_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__3,
    s1_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__1,
    s1_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [13:0] s1_possible_predicted_fhs_res_hist_12_new_folded_hist_src_doubled_1 = {
    s1_possible_predicted_fhs_res_hist_12_new_folded_hist_xored_res_1_6,
    s1_possible_predicted_fhs_res_hist_12_new_folded_hist_xored_res_1_5,
    s1_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__4,
    s1_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__3,
    s1_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__1,
    s1_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__0,
    s1_possible_predicted_fhs_res_hist_12_new_folded_hist_xored_1}; // @[Cat.scala 31:58]
  wire [6:0] s1_possible_predicted_fhs_res_hist_12_new_folded_hist_1 =
    s1_possible_predicted_fhs_res_hist_12_new_folded_hist_src_doubled_1[12:6]; // @[FrontendBundle.scala 221:30]
  wire  s1_possible_predicted_fhs_res_hist_13_new_folded_hist_xored_res_1_0 = s1_possible_predicted_fhs_ob_10_0 ^
    s1_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__0; // @[FrontendBundle.scala 256:48]
  wire  s1_possible_predicted_fhs_res_hist_13_new_folded_hist_xored_res_1_5 =
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[1] ^
    s1_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__5; // @[FrontendBundle.scala 256:48]
  wire  s1_possible_predicted_fhs_res_hist_13_new_folded_hist_xored_res_1_6 =
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[0] ^
    s1_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__6; // @[FrontendBundle.scala 256:48]
  wire [6:0] s1_possible_predicted_fhs_res_hist_13_new_folded_hist_xored_1 = {
    s1_possible_predicted_fhs_res_hist_13_new_folded_hist_xored_res_1_6,
    s1_possible_predicted_fhs_res_hist_13_new_folded_hist_xored_res_1_5,
    s1_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__4,
    s1_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__3,
    s1_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__1,
    s1_possible_predicted_fhs_res_hist_13_new_folded_hist_xored_res_1_0}; // @[FrontendBundle.scala 258:11]
  wire [13:0] s1_possible_predicted_fhs_res_hist_13_new_folded_hist_src_doubled_1 = {
    s1_possible_predicted_fhs_res_hist_13_new_folded_hist_xored_res_1_6,
    s1_possible_predicted_fhs_res_hist_13_new_folded_hist_xored_res_1_5,
    s1_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__4,
    s1_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__3,
    s1_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__1,
    s1_possible_predicted_fhs_res_hist_13_new_folded_hist_xored_res_1_0,
    s1_possible_predicted_fhs_res_hist_13_new_folded_hist_xored_1}; // @[Cat.scala 31:58]
  wire [6:0] s1_possible_predicted_fhs_res_hist_13_new_folded_hist_1 =
    s1_possible_predicted_fhs_res_hist_13_new_folded_hist_src_doubled_1[12:6]; // @[FrontendBundle.scala 221:30]
  wire  s1_possible_predicted_fhs_res_hist_14_new_folded_hist_xored_res_1_5 =
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[1] ^
    s1_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__5; // @[FrontendBundle.scala 256:48]
  wire  s1_possible_predicted_fhs_res_hist_14_new_folded_hist_xored_res_1_6 =
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[0] ^ s1_possible_predicted_fhs_ob_2_0 ^
    s1_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__6; // @[FrontendBundle.scala 256:48]
  wire [6:0] s1_possible_predicted_fhs_res_hist_14_new_folded_hist_xored_1 = {
    s1_possible_predicted_fhs_res_hist_14_new_folded_hist_xored_res_1_6,
    s1_possible_predicted_fhs_res_hist_14_new_folded_hist_xored_res_1_5,
    s1_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__4,
    s1_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__3,
    s1_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__1,
    s1_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [13:0] s1_possible_predicted_fhs_res_hist_14_new_folded_hist_src_doubled_1 = {
    s1_possible_predicted_fhs_res_hist_14_new_folded_hist_xored_res_1_6,
    s1_possible_predicted_fhs_res_hist_14_new_folded_hist_xored_res_1_5,
    s1_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__4,
    s1_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__3,
    s1_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__1,
    s1_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__0,
    s1_possible_predicted_fhs_res_hist_14_new_folded_hist_xored_1}; // @[Cat.scala 31:58]
  wire [6:0] s1_possible_predicted_fhs_res_hist_14_new_folded_hist_1 =
    s1_possible_predicted_fhs_res_hist_14_new_folded_hist_src_doubled_1[12:6]; // @[FrontendBundle.scala 221:30]
  wire  s1_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_res_1_8 = s1_possible_predicted_fhs_ob_2_0 ^
    s1_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__8; // @[FrontendBundle.scala 256:48]
  wire  s1_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_res_1_9 =
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[1] ^
    s1_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__9; // @[FrontendBundle.scala 256:48]
  wire  s1_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_res_1_10 =
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[0] ^
    s1_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__10; // @[FrontendBundle.scala 256:48]
  wire [10:0] s1_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_1 = {
    s1_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_res_1_10,
    s1_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_res_1_9,
    s1_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_res_1_8,
    s1_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__7,
    s1_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__6,
    s1_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__5,
    s1_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_lo}; // @[FrontendBundle.scala 258:11]
  wire [21:0] s1_possible_predicted_fhs_res_hist_15_new_folded_hist_src_doubled_1 = {
    s1_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_res_1_10,
    s1_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_res_1_9,
    s1_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_res_1_8,
    s1_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__7,
    s1_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__6,
    s1_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__5,
    s1_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_lo,
    s1_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_1}; // @[Cat.scala 31:58]
  wire [10:0] s1_possible_predicted_fhs_res_hist_15_new_folded_hist_1 =
    s1_possible_predicted_fhs_res_hist_15_new_folded_hist_src_doubled_1[20:10]; // @[FrontendBundle.scala 221:30]
  wire  s1_possible_predicted_fhs_res_hist_16_new_folded_hist_xored_res_1_1 = s1_possible_predicted_fhs_ob_13_0 ^
    s1_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__1; // @[FrontendBundle.scala 256:48]
  wire  s1_possible_predicted_fhs_res_hist_16_new_folded_hist_xored_res_1_6 =
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[1] ^
    s1_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__6; // @[FrontendBundle.scala 256:48]
  wire  s1_possible_predicted_fhs_res_hist_16_new_folded_hist_xored_res_1_7 =
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[0] ^
    s1_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__7; // @[FrontendBundle.scala 256:48]
  wire [7:0] s1_possible_predicted_fhs_res_hist_16_new_folded_hist_xored_1 = {
    s1_possible_predicted_fhs_res_hist_16_new_folded_hist_xored_res_1_7,
    s1_possible_predicted_fhs_res_hist_16_new_folded_hist_xored_res_1_6,
    s1_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__5,
    s1_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__4,
    s1_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__3,
    s1_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_16_new_folded_hist_xored_res_1_1,
    s1_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [15:0] s1_possible_predicted_fhs_res_hist_16_new_folded_hist_src_doubled_1 = {
    s1_possible_predicted_fhs_res_hist_16_new_folded_hist_xored_res_1_7,
    s1_possible_predicted_fhs_res_hist_16_new_folded_hist_xored_res_1_6,
    s1_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__5,
    s1_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__4,
    s1_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__3,
    s1_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_16_new_folded_hist_xored_res_1_1,
    s1_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__0,
    s1_possible_predicted_fhs_res_hist_16_new_folded_hist_xored_1}; // @[Cat.scala 31:58]
  wire [7:0] s1_possible_predicted_fhs_res_hist_16_new_folded_hist_1 =
    s1_possible_predicted_fhs_res_hist_16_new_folded_hist_src_doubled_1[14:7]; // @[FrontendBundle.scala 221:30]
  wire  s1_possible_predicted_fhs_res_hist_17_new_folded_hist_xored_res_1_4 = s1_possible_predicted_fhs_ob_4_0 ^
    s1_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__4; // @[FrontendBundle.scala 256:48]
  wire  s1_possible_predicted_fhs_res_hist_17_new_folded_hist_xored_res_1_6 =
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[1] ^
    s1_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__6; // @[FrontendBundle.scala 256:48]
  wire  s1_possible_predicted_fhs_res_hist_17_new_folded_hist_xored_res_1_7 =
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[0] ^
    s1_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__7; // @[FrontendBundle.scala 256:48]
  wire [7:0] s1_possible_predicted_fhs_res_hist_17_new_folded_hist_xored_1 = {
    s1_possible_predicted_fhs_res_hist_17_new_folded_hist_xored_res_1_7,
    s1_possible_predicted_fhs_res_hist_17_new_folded_hist_xored_res_1_6,
    s1_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__5,
    s1_possible_predicted_fhs_res_hist_17_new_folded_hist_xored_res_1_4,
    s1_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__3,
    s1_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__1,
    s1_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [15:0] s1_possible_predicted_fhs_res_hist_17_new_folded_hist_src_doubled_1 = {
    s1_possible_predicted_fhs_res_hist_17_new_folded_hist_xored_res_1_7,
    s1_possible_predicted_fhs_res_hist_17_new_folded_hist_xored_res_1_6,
    s1_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__5,
    s1_possible_predicted_fhs_res_hist_17_new_folded_hist_xored_res_1_4,
    s1_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__3,
    s1_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__1,
    s1_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__0,
    s1_possible_predicted_fhs_res_hist_17_new_folded_hist_xored_1}; // @[Cat.scala 31:58]
  wire [7:0] s1_possible_predicted_fhs_res_hist_17_new_folded_hist_1 =
    s1_possible_predicted_fhs_res_hist_17_new_folded_hist_src_doubled_1[14:7]; // @[FrontendBundle.scala 221:30]
  wire  _s1_possible_predicted_fhs_T_203 = _s1_possible_predicted_fhs_T_5 & _s1_predicted_ghist_ptr_T_60; // @[BPU.scala 403:88]
  wire [1:0] s1_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2 = {
    _s1_possible_predicted_fhs_T_203,1'h0}; // @[FrontendBundle.scala 274:102]
  wire  s1_possible_predicted_fhs_res_hist_0_new_folded_hist_xored_res_2_6 =
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[1] ^ s1_possible_predicted_fhs_ob__1 ^
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__6; // @[FrontendBundle.scala 256:48]
  wire  s1_possible_predicted_fhs_res_hist_0_new_folded_hist_xored_res_2_7 =
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[0] ^ s1_possible_predicted_fhs_ob__0 ^
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__7; // @[FrontendBundle.scala 256:48]
  wire [7:0] s1_possible_predicted_fhs_res_hist_0_new_folded_hist_xored_2 = {
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_xored_res_2_7,
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_xored_res_2_6,
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__5,
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__4,
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__3,
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__1,
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [15:0] s1_possible_predicted_fhs_res_hist_0_new_folded_hist_src_doubled_2 = {
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_xored_res_2_7,
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_xored_res_2_6,
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__5,
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__4,
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__3,
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__1,
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__0,
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_xored_2}; // @[Cat.scala 31:58]
  wire [7:0] s1_possible_predicted_fhs_res_hist_0_new_folded_hist_2 =
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_src_doubled_2[13:6]; // @[FrontendBundle.scala 221:30]
  wire  s1_possible_predicted_fhs_res_hist_1_new_folded_hist_xored_res_2_6 =
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[1] ^ s1_possible_predicted_fhs_ob_1_1 ^
    s1_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__6; // @[FrontendBundle.scala 256:48]
  wire  s1_possible_predicted_fhs_res_hist_1_new_folded_hist_xored_res_2_7 =
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[0] ^ s1_possible_predicted_fhs_ob_1_0 ^
    s1_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__7; // @[FrontendBundle.scala 256:48]
  wire [7:0] s1_possible_predicted_fhs_res_hist_1_new_folded_hist_xored_2 = {
    s1_possible_predicted_fhs_res_hist_1_new_folded_hist_xored_res_2_7,
    s1_possible_predicted_fhs_res_hist_1_new_folded_hist_xored_res_2_6,
    s1_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__5,
    s1_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__4,
    s1_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__3,
    s1_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__1,
    s1_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [15:0] s1_possible_predicted_fhs_res_hist_1_new_folded_hist_src_doubled_2 = {
    s1_possible_predicted_fhs_res_hist_1_new_folded_hist_xored_res_2_7,
    s1_possible_predicted_fhs_res_hist_1_new_folded_hist_xored_res_2_6,
    s1_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__5,
    s1_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__4,
    s1_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__3,
    s1_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__1,
    s1_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__0,
    s1_possible_predicted_fhs_res_hist_1_new_folded_hist_xored_2}; // @[Cat.scala 31:58]
  wire [7:0] s1_possible_predicted_fhs_res_hist_1_new_folded_hist_2 =
    s1_possible_predicted_fhs_res_hist_1_new_folded_hist_src_doubled_2[13:6]; // @[FrontendBundle.scala 221:30]
  wire  s1_possible_predicted_fhs_res_hist_2_new_folded_hist_xored_res_2_5 = s1_possible_predicted_fhs_ob_2_1 ^
    s1_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__5; // @[FrontendBundle.scala 256:48]
  wire  s1_possible_predicted_fhs_res_hist_2_new_folded_hist_xored_res_2_6 =
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[1] ^ s1_possible_predicted_fhs_ob_2_0 ^
    s1_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__6; // @[FrontendBundle.scala 256:48]
  wire  s1_possible_predicted_fhs_res_hist_2_new_folded_hist_xored_res_2_7 =
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[0] ^
    s1_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__7; // @[FrontendBundle.scala 256:48]
  wire [7:0] s1_possible_predicted_fhs_res_hist_2_new_folded_hist_xored_2 = {
    s1_possible_predicted_fhs_res_hist_2_new_folded_hist_xored_res_2_7,
    s1_possible_predicted_fhs_res_hist_2_new_folded_hist_xored_res_2_6,
    s1_possible_predicted_fhs_res_hist_2_new_folded_hist_xored_res_2_5,
    s1_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__4,
    s1_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__3,
    s1_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__1,
    s1_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [15:0] s1_possible_predicted_fhs_res_hist_2_new_folded_hist_src_doubled_2 = {
    s1_possible_predicted_fhs_res_hist_2_new_folded_hist_xored_res_2_7,
    s1_possible_predicted_fhs_res_hist_2_new_folded_hist_xored_res_2_6,
    s1_possible_predicted_fhs_res_hist_2_new_folded_hist_xored_res_2_5,
    s1_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__4,
    s1_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__3,
    s1_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__1,
    s1_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__0,
    s1_possible_predicted_fhs_res_hist_2_new_folded_hist_xored_2}; // @[Cat.scala 31:58]
  wire [7:0] s1_possible_predicted_fhs_res_hist_2_new_folded_hist_2 =
    s1_possible_predicted_fhs_res_hist_2_new_folded_hist_src_doubled_2[13:6]; // @[FrontendBundle.scala 221:30]
  wire  s1_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_res_2_8 = s1_possible_predicted_fhs_ob_1_1 ^
    s1_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__8; // @[FrontendBundle.scala 256:48]
  wire  s1_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_res_2_9 =
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[1] ^ s1_possible_predicted_fhs_ob_1_0 ^
    s1_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__9; // @[FrontendBundle.scala 256:48]
  wire  s1_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_res_2_10 =
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[0] ^
    s1_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__10; // @[FrontendBundle.scala 256:48]
  wire [10:0] s1_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_2 = {
    s1_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_res_2_10,
    s1_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_res_2_9,
    s1_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_res_2_8,
    s1_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__7,
    s1_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__6,
    s1_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__5,
    s1_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_lo}; // @[FrontendBundle.scala 258:11]
  wire [21:0] s1_possible_predicted_fhs_res_hist_3_new_folded_hist_src_doubled_2 = {
    s1_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_res_2_10,
    s1_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_res_2_9,
    s1_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_res_2_8,
    s1_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__7,
    s1_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__6,
    s1_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__5,
    s1_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_lo,
    s1_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_2}; // @[Cat.scala 31:58]
  wire [10:0] s1_possible_predicted_fhs_res_hist_3_new_folded_hist_2 =
    s1_possible_predicted_fhs_res_hist_3_new_folded_hist_src_doubled_2[19:9]; // @[FrontendBundle.scala 221:30]
  wire [5:0] _s1_possible_predicted_fhs_res_hist_4_new_folded_hist_T_4 = {s1_folded_gh_hist_4_folded_hist, 2'h0}; // @[FrontendBundle.scala 290:21]
  wire [5:0] _GEN_11916 = {{5'd0}, _s1_possible_predicted_fhs_T_203}; // @[FrontendBundle.scala 290:29]
  wire [5:0] _s1_possible_predicted_fhs_res_hist_4_new_folded_hist_T_5 =
    _s1_possible_predicted_fhs_res_hist_4_new_folded_hist_T_4 | _GEN_11916; // @[FrontendBundle.scala 290:29]
  wire [3:0] s1_possible_predicted_fhs_res_hist_4_new_folded_hist_2 =
    _s1_possible_predicted_fhs_res_hist_4_new_folded_hist_T_5[3:0]; // @[FrontendBundle.scala 290:37]
  wire  s1_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_res_2_0 = s1_possible_predicted_fhs_ob_4_1 ^
    s1_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__0; // @[FrontendBundle.scala 256:48]
  wire  s1_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_res_2_9 =
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[1] ^
    s1_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__9; // @[FrontendBundle.scala 256:48]
  wire  s1_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_res_2_10 =
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[0] ^
    s1_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__10; // @[FrontendBundle.scala 256:48]
  wire [4:0] s1_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_lo_2 = {
    s1_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__4,
    s1_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__3,
    s1_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_res_1_1,
    s1_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_res_2_0}; // @[FrontendBundle.scala 258:11]
  wire [10:0] s1_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_2 = {
    s1_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_res_2_10,
    s1_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_res_2_9,
    s1_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__8,
    s1_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__7,
    s1_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__6,
    s1_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__5,
    s1_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_lo_2}; // @[FrontendBundle.scala 258:11]
  wire [21:0] s1_possible_predicted_fhs_res_hist_5_new_folded_hist_src_doubled_2 = {
    s1_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_res_2_10,
    s1_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_res_2_9,
    s1_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__8,
    s1_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__7,
    s1_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__6,
    s1_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__5,
    s1_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_lo_2,
    s1_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_2}; // @[Cat.scala 31:58]
  wire [10:0] s1_possible_predicted_fhs_res_hist_5_new_folded_hist_2 =
    s1_possible_predicted_fhs_res_hist_5_new_folded_hist_src_doubled_2[19:9]; // @[FrontendBundle.scala 221:30]
  wire  s1_possible_predicted_fhs_res_hist_6_new_folded_hist_xored_res_2_2 = s1_possible_predicted_fhs_ob_4_1 ^
    s1_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__2; // @[FrontendBundle.scala 256:48]
  wire  s1_possible_predicted_fhs_res_hist_6_new_folded_hist_xored_res_2_7 =
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[1] ^
    s1_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__7; // @[FrontendBundle.scala 256:48]
  wire  s1_possible_predicted_fhs_res_hist_6_new_folded_hist_xored_res_2_8 =
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[0] ^
    s1_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__8; // @[FrontendBundle.scala 256:48]
  wire [8:0] s1_possible_predicted_fhs_res_hist_6_new_folded_hist_xored_2 = {
    s1_possible_predicted_fhs_res_hist_6_new_folded_hist_xored_res_2_8,
    s1_possible_predicted_fhs_res_hist_6_new_folded_hist_xored_res_2_7,
    s1_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__6,
    s1_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__5,
    s1_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__4,
    s1_possible_predicted_fhs_res_hist_6_new_folded_hist_xored_res_1_3,
    s1_possible_predicted_fhs_res_hist_6_new_folded_hist_xored_res_2_2,
    s1_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__1,
    s1_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [17:0] s1_possible_predicted_fhs_res_hist_6_new_folded_hist_src_doubled_2 = {
    s1_possible_predicted_fhs_res_hist_6_new_folded_hist_xored_res_2_8,
    s1_possible_predicted_fhs_res_hist_6_new_folded_hist_xored_res_2_7,
    s1_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__6,
    s1_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__5,
    s1_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__4,
    s1_possible_predicted_fhs_res_hist_6_new_folded_hist_xored_res_1_3,
    s1_possible_predicted_fhs_res_hist_6_new_folded_hist_xored_res_2_2,
    s1_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__1,
    s1_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__0,
    s1_possible_predicted_fhs_res_hist_6_new_folded_hist_xored_2}; // @[Cat.scala 31:58]
  wire [8:0] s1_possible_predicted_fhs_res_hist_6_new_folded_hist_2 =
    s1_possible_predicted_fhs_res_hist_6_new_folded_hist_src_doubled_2[15:7]; // @[FrontendBundle.scala 221:30]
  wire  s1_possible_predicted_fhs_res_hist_7_new_folded_hist_xored_res_2_5 = s1_possible_predicted_fhs_ob__1 ^
    s1_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__5; // @[FrontendBundle.scala 256:48]
  wire  s1_possible_predicted_fhs_res_hist_7_new_folded_hist_xored_res_2_7 =
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[1] ^
    s1_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__7; // @[FrontendBundle.scala 256:48]
  wire  s1_possible_predicted_fhs_res_hist_7_new_folded_hist_xored_res_2_8 =
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[0] ^
    s1_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__8; // @[FrontendBundle.scala 256:48]
  wire [8:0] s1_possible_predicted_fhs_res_hist_7_new_folded_hist_xored_2 = {
    s1_possible_predicted_fhs_res_hist_7_new_folded_hist_xored_res_2_8,
    s1_possible_predicted_fhs_res_hist_7_new_folded_hist_xored_res_2_7,
    s1_possible_predicted_fhs_res_hist_7_new_folded_hist_xored_res_1_6,
    s1_possible_predicted_fhs_res_hist_7_new_folded_hist_xored_res_2_5,
    s1_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__4,
    s1_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__3,
    s1_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__1,
    s1_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [17:0] s1_possible_predicted_fhs_res_hist_7_new_folded_hist_src_doubled_2 = {
    s1_possible_predicted_fhs_res_hist_7_new_folded_hist_xored_res_2_8,
    s1_possible_predicted_fhs_res_hist_7_new_folded_hist_xored_res_2_7,
    s1_possible_predicted_fhs_res_hist_7_new_folded_hist_xored_res_1_6,
    s1_possible_predicted_fhs_res_hist_7_new_folded_hist_xored_res_2_5,
    s1_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__4,
    s1_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__3,
    s1_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__1,
    s1_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__0,
    s1_possible_predicted_fhs_res_hist_7_new_folded_hist_xored_2}; // @[Cat.scala 31:58]
  wire [8:0] s1_possible_predicted_fhs_res_hist_7_new_folded_hist_2 =
    s1_possible_predicted_fhs_res_hist_7_new_folded_hist_src_doubled_2[15:7]; // @[FrontendBundle.scala 221:30]
  wire [9:0] _s1_possible_predicted_fhs_res_hist_8_new_folded_hist_T_4 = {s1_folded_gh_hist_8_folded_hist, 2'h0}; // @[FrontendBundle.scala 290:21]
  wire [9:0] _GEN_11917 = {{9'd0}, _s1_possible_predicted_fhs_T_203}; // @[FrontendBundle.scala 290:29]
  wire [9:0] _s1_possible_predicted_fhs_res_hist_8_new_folded_hist_T_5 =
    _s1_possible_predicted_fhs_res_hist_8_new_folded_hist_T_4 | _GEN_11917; // @[FrontendBundle.scala 290:29]
  wire [7:0] s1_possible_predicted_fhs_res_hist_8_new_folded_hist_2 =
    _s1_possible_predicted_fhs_res_hist_8_new_folded_hist_T_5[7:0]; // @[FrontendBundle.scala 290:37]
  wire  s1_possible_predicted_fhs_res_hist_9_new_folded_hist_xored_res_2_2 = s1_possible_predicted_fhs_ob_1_1 ^
    s1_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__2; // @[FrontendBundle.scala 256:48]
  wire  s1_possible_predicted_fhs_res_hist_9_new_folded_hist_xored_res_2_5 =
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[1] ^
    s1_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__5; // @[FrontendBundle.scala 256:48]
  wire  s1_possible_predicted_fhs_res_hist_9_new_folded_hist_xored_res_2_6 =
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[0] ^
    s1_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__6; // @[FrontendBundle.scala 256:48]
  wire [6:0] s1_possible_predicted_fhs_res_hist_9_new_folded_hist_xored_2 = {
    s1_possible_predicted_fhs_res_hist_9_new_folded_hist_xored_res_2_6,
    s1_possible_predicted_fhs_res_hist_9_new_folded_hist_xored_res_2_5,
    s1_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__4,
    s1_possible_predicted_fhs_res_hist_9_new_folded_hist_xored_res_1_3,
    s1_possible_predicted_fhs_res_hist_9_new_folded_hist_xored_res_2_2,
    s1_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__1,
    s1_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [13:0] s1_possible_predicted_fhs_res_hist_9_new_folded_hist_src_doubled_2 = {
    s1_possible_predicted_fhs_res_hist_9_new_folded_hist_xored_res_2_6,
    s1_possible_predicted_fhs_res_hist_9_new_folded_hist_xored_res_2_5,
    s1_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__4,
    s1_possible_predicted_fhs_res_hist_9_new_folded_hist_xored_res_1_3,
    s1_possible_predicted_fhs_res_hist_9_new_folded_hist_xored_res_2_2,
    s1_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__1,
    s1_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__0,
    s1_possible_predicted_fhs_res_hist_9_new_folded_hist_xored_2}; // @[Cat.scala 31:58]
  wire [6:0] s1_possible_predicted_fhs_res_hist_9_new_folded_hist_2 =
    s1_possible_predicted_fhs_res_hist_9_new_folded_hist_src_doubled_2[11:5]; // @[FrontendBundle.scala 221:30]
  wire  s1_possible_predicted_fhs_res_hist_10_new_folded_hist_xored_res_2_3 = s1_possible_predicted_fhs_ob_1_1 ^
    s1_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__3; // @[FrontendBundle.scala 256:48]
  wire  s1_possible_predicted_fhs_res_hist_10_new_folded_hist_xored_res_2_7 =
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[1] ^
    s1_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__7; // @[FrontendBundle.scala 256:48]
  wire  s1_possible_predicted_fhs_res_hist_10_new_folded_hist_xored_res_2_8 =
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[0] ^
    s1_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__8; // @[FrontendBundle.scala 256:48]
  wire [8:0] s1_possible_predicted_fhs_res_hist_10_new_folded_hist_xored_2 = {
    s1_possible_predicted_fhs_res_hist_10_new_folded_hist_xored_res_2_8,
    s1_possible_predicted_fhs_res_hist_10_new_folded_hist_xored_res_2_7,
    s1_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__6,
    s1_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__5,
    s1_possible_predicted_fhs_res_hist_10_new_folded_hist_xored_res_1_4,
    s1_possible_predicted_fhs_res_hist_10_new_folded_hist_xored_res_2_3,
    s1_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__1,
    s1_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [17:0] s1_possible_predicted_fhs_res_hist_10_new_folded_hist_src_doubled_2 = {
    s1_possible_predicted_fhs_res_hist_10_new_folded_hist_xored_res_2_8,
    s1_possible_predicted_fhs_res_hist_10_new_folded_hist_xored_res_2_7,
    s1_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__6,
    s1_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__5,
    s1_possible_predicted_fhs_res_hist_10_new_folded_hist_xored_res_1_4,
    s1_possible_predicted_fhs_res_hist_10_new_folded_hist_xored_res_2_3,
    s1_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__1,
    s1_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__0,
    s1_possible_predicted_fhs_res_hist_10_new_folded_hist_xored_2}; // @[Cat.scala 31:58]
  wire [8:0] s1_possible_predicted_fhs_res_hist_10_new_folded_hist_2 =
    s1_possible_predicted_fhs_res_hist_10_new_folded_hist_src_doubled_2[15:7]; // @[FrontendBundle.scala 221:30]
  wire [9:0] _s1_possible_predicted_fhs_res_hist_11_new_folded_hist_T_4 = {s1_folded_gh_hist_11_folded_hist, 2'h0}; // @[FrontendBundle.scala 290:21]
  wire [9:0] _s1_possible_predicted_fhs_res_hist_11_new_folded_hist_T_5 =
    _s1_possible_predicted_fhs_res_hist_11_new_folded_hist_T_4 | _GEN_11917; // @[FrontendBundle.scala 290:29]
  wire [7:0] s1_possible_predicted_fhs_res_hist_11_new_folded_hist_2 =
    _s1_possible_predicted_fhs_res_hist_11_new_folded_hist_T_5[7:0]; // @[FrontendBundle.scala 290:37]
  wire  s1_possible_predicted_fhs_res_hist_12_new_folded_hist_xored_res_2_4 = s1_possible_predicted_fhs_ob_4_1 ^
    s1_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__4; // @[FrontendBundle.scala 256:48]
  wire  s1_possible_predicted_fhs_res_hist_12_new_folded_hist_xored_res_2_5 =
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[1] ^ s1_possible_predicted_fhs_ob_4_0 ^
    s1_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__5; // @[FrontendBundle.scala 256:48]
  wire  s1_possible_predicted_fhs_res_hist_12_new_folded_hist_xored_res_2_6 =
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[0] ^
    s1_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__6; // @[FrontendBundle.scala 256:48]
  wire [6:0] s1_possible_predicted_fhs_res_hist_12_new_folded_hist_xored_2 = {
    s1_possible_predicted_fhs_res_hist_12_new_folded_hist_xored_res_2_6,
    s1_possible_predicted_fhs_res_hist_12_new_folded_hist_xored_res_2_5,
    s1_possible_predicted_fhs_res_hist_12_new_folded_hist_xored_res_2_4,
    s1_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__3,
    s1_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__1,
    s1_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [13:0] s1_possible_predicted_fhs_res_hist_12_new_folded_hist_src_doubled_2 = {
    s1_possible_predicted_fhs_res_hist_12_new_folded_hist_xored_res_2_6,
    s1_possible_predicted_fhs_res_hist_12_new_folded_hist_xored_res_2_5,
    s1_possible_predicted_fhs_res_hist_12_new_folded_hist_xored_res_2_4,
    s1_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__3,
    s1_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__1,
    s1_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__0,
    s1_possible_predicted_fhs_res_hist_12_new_folded_hist_xored_2}; // @[Cat.scala 31:58]
  wire [6:0] s1_possible_predicted_fhs_res_hist_12_new_folded_hist_2 =
    s1_possible_predicted_fhs_res_hist_12_new_folded_hist_src_doubled_2[11:5]; // @[FrontendBundle.scala 221:30]
  wire  s1_possible_predicted_fhs_res_hist_13_new_folded_hist_xored_res_2_5 =
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[1] ^
    s1_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__5; // @[FrontendBundle.scala 256:48]
  wire [6:0] s1_possible_predicted_fhs_res_hist_13_new_folded_hist_xored_2 = {
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[0],
    s1_possible_predicted_fhs_res_hist_13_new_folded_hist_xored_res_2_5,
    s1_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__4,
    s1_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__3,
    s1_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__1,
    s1_possible_predicted_fhs_res_hist_13_new_folded_hist_xored_res_1_0}; // @[FrontendBundle.scala 258:11]
  wire [13:0] s1_possible_predicted_fhs_res_hist_13_new_folded_hist_src_doubled_2 = {
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[0],
    s1_possible_predicted_fhs_res_hist_13_new_folded_hist_xored_res_2_5,
    s1_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__4,
    s1_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__3,
    s1_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__1,
    s1_possible_predicted_fhs_res_hist_13_new_folded_hist_xored_res_1_0,
    s1_possible_predicted_fhs_res_hist_13_new_folded_hist_xored_2}; // @[Cat.scala 31:58]
  wire [6:0] s1_possible_predicted_fhs_res_hist_13_new_folded_hist_2 =
    s1_possible_predicted_fhs_res_hist_13_new_folded_hist_src_doubled_2[11:5]; // @[FrontendBundle.scala 221:30]
  wire  s1_possible_predicted_fhs_res_hist_14_new_folded_hist_xored_res_2_5 =
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[1] ^ s1_possible_predicted_fhs_ob_2_1 ^
    s1_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__5; // @[FrontendBundle.scala 256:48]
  wire  s1_possible_predicted_fhs_res_hist_14_new_folded_hist_xored_res_2_6 =
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[0] ^ s1_possible_predicted_fhs_ob_2_0 ^
    s1_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__6; // @[FrontendBundle.scala 256:48]
  wire [6:0] s1_possible_predicted_fhs_res_hist_14_new_folded_hist_xored_2 = {
    s1_possible_predicted_fhs_res_hist_14_new_folded_hist_xored_res_2_6,
    s1_possible_predicted_fhs_res_hist_14_new_folded_hist_xored_res_2_5,
    s1_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__4,
    s1_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__3,
    s1_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__1,
    s1_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [13:0] s1_possible_predicted_fhs_res_hist_14_new_folded_hist_src_doubled_2 = {
    s1_possible_predicted_fhs_res_hist_14_new_folded_hist_xored_res_2_6,
    s1_possible_predicted_fhs_res_hist_14_new_folded_hist_xored_res_2_5,
    s1_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__4,
    s1_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__3,
    s1_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__1,
    s1_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__0,
    s1_possible_predicted_fhs_res_hist_14_new_folded_hist_xored_2}; // @[Cat.scala 31:58]
  wire [6:0] s1_possible_predicted_fhs_res_hist_14_new_folded_hist_2 =
    s1_possible_predicted_fhs_res_hist_14_new_folded_hist_src_doubled_2[11:5]; // @[FrontendBundle.scala 221:30]
  wire  s1_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_res_2_7 = s1_possible_predicted_fhs_ob_2_1 ^
    s1_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__7; // @[FrontendBundle.scala 256:48]
  wire  s1_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_res_2_9 =
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[1] ^
    s1_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__9; // @[FrontendBundle.scala 256:48]
  wire  s1_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_res_2_10 =
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[0] ^
    s1_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__10; // @[FrontendBundle.scala 256:48]
  wire [10:0] s1_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_2 = {
    s1_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_res_2_10,
    s1_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_res_2_9,
    s1_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_res_1_8,
    s1_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_res_2_7,
    s1_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__6,
    s1_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__5,
    s1_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_lo}; // @[FrontendBundle.scala 258:11]
  wire [21:0] s1_possible_predicted_fhs_res_hist_15_new_folded_hist_src_doubled_2 = {
    s1_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_res_2_10,
    s1_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_res_2_9,
    s1_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_res_1_8,
    s1_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_res_2_7,
    s1_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__6,
    s1_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__5,
    s1_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_lo,
    s1_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_2}; // @[Cat.scala 31:58]
  wire [10:0] s1_possible_predicted_fhs_res_hist_15_new_folded_hist_2 =
    s1_possible_predicted_fhs_res_hist_15_new_folded_hist_src_doubled_2[19:9]; // @[FrontendBundle.scala 221:30]
  wire  s1_possible_predicted_fhs_res_hist_16_new_folded_hist_xored_res_2_0 = s1_possible_predicted_fhs_ob_13_1 ^
    s1_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__0; // @[FrontendBundle.scala 256:48]
  wire  s1_possible_predicted_fhs_res_hist_16_new_folded_hist_xored_res_2_6 =
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[1] ^
    s1_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__6; // @[FrontendBundle.scala 256:48]
  wire  s1_possible_predicted_fhs_res_hist_16_new_folded_hist_xored_res_2_7 =
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[0] ^
    s1_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__7; // @[FrontendBundle.scala 256:48]
  wire [7:0] s1_possible_predicted_fhs_res_hist_16_new_folded_hist_xored_2 = {
    s1_possible_predicted_fhs_res_hist_16_new_folded_hist_xored_res_2_7,
    s1_possible_predicted_fhs_res_hist_16_new_folded_hist_xored_res_2_6,
    s1_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__5,
    s1_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__4,
    s1_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__3,
    s1_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_16_new_folded_hist_xored_res_1_1,
    s1_possible_predicted_fhs_res_hist_16_new_folded_hist_xored_res_2_0}; // @[FrontendBundle.scala 258:11]
  wire [15:0] s1_possible_predicted_fhs_res_hist_16_new_folded_hist_src_doubled_2 = {
    s1_possible_predicted_fhs_res_hist_16_new_folded_hist_xored_res_2_7,
    s1_possible_predicted_fhs_res_hist_16_new_folded_hist_xored_res_2_6,
    s1_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__5,
    s1_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__4,
    s1_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__3,
    s1_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_16_new_folded_hist_xored_res_1_1,
    s1_possible_predicted_fhs_res_hist_16_new_folded_hist_xored_res_2_0,
    s1_possible_predicted_fhs_res_hist_16_new_folded_hist_xored_2}; // @[Cat.scala 31:58]
  wire [7:0] s1_possible_predicted_fhs_res_hist_16_new_folded_hist_2 =
    s1_possible_predicted_fhs_res_hist_16_new_folded_hist_src_doubled_2[13:6]; // @[FrontendBundle.scala 221:30]
  wire  s1_possible_predicted_fhs_res_hist_17_new_folded_hist_xored_res_2_3 = s1_possible_predicted_fhs_ob_4_1 ^
    s1_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__3; // @[FrontendBundle.scala 256:48]
  wire  s1_possible_predicted_fhs_res_hist_17_new_folded_hist_xored_res_2_6 =
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[1] ^
    s1_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__6; // @[FrontendBundle.scala 256:48]
  wire  s1_possible_predicted_fhs_res_hist_17_new_folded_hist_xored_res_2_7 =
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[0] ^
    s1_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__7; // @[FrontendBundle.scala 256:48]
  wire [7:0] s1_possible_predicted_fhs_res_hist_17_new_folded_hist_xored_2 = {
    s1_possible_predicted_fhs_res_hist_17_new_folded_hist_xored_res_2_7,
    s1_possible_predicted_fhs_res_hist_17_new_folded_hist_xored_res_2_6,
    s1_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__5,
    s1_possible_predicted_fhs_res_hist_17_new_folded_hist_xored_res_1_4,
    s1_possible_predicted_fhs_res_hist_17_new_folded_hist_xored_res_2_3,
    s1_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__1,
    s1_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [15:0] s1_possible_predicted_fhs_res_hist_17_new_folded_hist_src_doubled_2 = {
    s1_possible_predicted_fhs_res_hist_17_new_folded_hist_xored_res_2_7,
    s1_possible_predicted_fhs_res_hist_17_new_folded_hist_xored_res_2_6,
    s1_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__5,
    s1_possible_predicted_fhs_res_hist_17_new_folded_hist_xored_res_1_4,
    s1_possible_predicted_fhs_res_hist_17_new_folded_hist_xored_res_2_3,
    s1_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__2,
    s1_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__1,
    s1_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__0,
    s1_possible_predicted_fhs_res_hist_17_new_folded_hist_xored_2}; // @[Cat.scala 31:58]
  wire [7:0] s1_possible_predicted_fhs_res_hist_17_new_folded_hist_2 =
    s1_possible_predicted_fhs_res_hist_17_new_folded_hist_src_doubled_2[13:6]; // @[FrontendBundle.scala 221:30]
  wire [7:0] _s1_predicted_fh_T_61 = _s1_predicted_ghist_ptr_T_4 ? s1_possible_predicted_fhs_res_hist_0_new_folded_hist
     : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _s1_predicted_fh_T_62 = _s1_predicted_ghist_ptr_T_32 ?
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _s1_predicted_fh_T_63 = _s1_predicted_ghist_ptr_T_60 ?
    s1_possible_predicted_fhs_res_hist_0_new_folded_hist_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _s1_predicted_fh_T_64 = _s1_predicted_fh_T_61 | _s1_predicted_fh_T_62; // @[Mux.scala 27:73]
  wire [7:0] _s1_predicted_fh_T_66 = _s1_predicted_ghist_ptr_T_4 ? s1_possible_predicted_fhs_res_hist_1_new_folded_hist
     : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _s1_predicted_fh_T_67 = _s1_predicted_ghist_ptr_T_32 ?
    s1_possible_predicted_fhs_res_hist_1_new_folded_hist_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _s1_predicted_fh_T_68 = _s1_predicted_ghist_ptr_T_60 ?
    s1_possible_predicted_fhs_res_hist_1_new_folded_hist_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _s1_predicted_fh_T_69 = _s1_predicted_fh_T_66 | _s1_predicted_fh_T_67; // @[Mux.scala 27:73]
  wire [7:0] _s1_predicted_fh_T_71 = _s1_predicted_ghist_ptr_T_4 ? s1_possible_predicted_fhs_res_hist_2_new_folded_hist
     : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _s1_predicted_fh_T_72 = _s1_predicted_ghist_ptr_T_32 ?
    s1_possible_predicted_fhs_res_hist_2_new_folded_hist_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _s1_predicted_fh_T_73 = _s1_predicted_ghist_ptr_T_60 ?
    s1_possible_predicted_fhs_res_hist_2_new_folded_hist_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _s1_predicted_fh_T_74 = _s1_predicted_fh_T_71 | _s1_predicted_fh_T_72; // @[Mux.scala 27:73]
  wire [10:0] _s1_predicted_fh_T_76 = _s1_predicted_ghist_ptr_T_4 ? s1_possible_predicted_fhs_res_hist_3_new_folded_hist
     : 11'h0; // @[Mux.scala 27:73]
  wire [10:0] _s1_predicted_fh_T_77 = _s1_predicted_ghist_ptr_T_32 ?
    s1_possible_predicted_fhs_res_hist_3_new_folded_hist_1 : 11'h0; // @[Mux.scala 27:73]
  wire [10:0] _s1_predicted_fh_T_78 = _s1_predicted_ghist_ptr_T_60 ?
    s1_possible_predicted_fhs_res_hist_3_new_folded_hist_2 : 11'h0; // @[Mux.scala 27:73]
  wire [10:0] _s1_predicted_fh_T_79 = _s1_predicted_fh_T_76 | _s1_predicted_fh_T_77; // @[Mux.scala 27:73]
  wire [3:0] _s1_predicted_fh_T_81 = _s1_predicted_ghist_ptr_T_4 ? s1_possible_predicted_fhs_res_hist_4_new_folded_hist
     : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _s1_predicted_fh_T_82 = _s1_predicted_ghist_ptr_T_32 ?
    s1_possible_predicted_fhs_res_hist_4_new_folded_hist_1 : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _s1_predicted_fh_T_83 = _s1_predicted_ghist_ptr_T_60 ?
    s1_possible_predicted_fhs_res_hist_4_new_folded_hist_2 : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _s1_predicted_fh_T_84 = _s1_predicted_fh_T_81 | _s1_predicted_fh_T_82; // @[Mux.scala 27:73]
  wire [10:0] _s1_predicted_fh_T_86 = _s1_predicted_ghist_ptr_T_4 ? s1_possible_predicted_fhs_res_hist_5_new_folded_hist
     : 11'h0; // @[Mux.scala 27:73]
  wire [10:0] _s1_predicted_fh_T_87 = _s1_predicted_ghist_ptr_T_32 ?
    s1_possible_predicted_fhs_res_hist_5_new_folded_hist_1 : 11'h0; // @[Mux.scala 27:73]
  wire [10:0] _s1_predicted_fh_T_88 = _s1_predicted_ghist_ptr_T_60 ?
    s1_possible_predicted_fhs_res_hist_5_new_folded_hist_2 : 11'h0; // @[Mux.scala 27:73]
  wire [10:0] _s1_predicted_fh_T_89 = _s1_predicted_fh_T_86 | _s1_predicted_fh_T_87; // @[Mux.scala 27:73]
  wire [8:0] _s1_predicted_fh_T_91 = _s1_predicted_ghist_ptr_T_4 ? s1_possible_predicted_fhs_res_hist_6_new_folded_hist
     : 9'h0; // @[Mux.scala 27:73]
  wire [8:0] _s1_predicted_fh_T_92 = _s1_predicted_ghist_ptr_T_32 ?
    s1_possible_predicted_fhs_res_hist_6_new_folded_hist_1 : 9'h0; // @[Mux.scala 27:73]
  wire [8:0] _s1_predicted_fh_T_93 = _s1_predicted_ghist_ptr_T_60 ?
    s1_possible_predicted_fhs_res_hist_6_new_folded_hist_2 : 9'h0; // @[Mux.scala 27:73]
  wire [8:0] _s1_predicted_fh_T_94 = _s1_predicted_fh_T_91 | _s1_predicted_fh_T_92; // @[Mux.scala 27:73]
  wire [8:0] _s1_predicted_fh_T_96 = _s1_predicted_ghist_ptr_T_4 ? s1_possible_predicted_fhs_res_hist_7_new_folded_hist
     : 9'h0; // @[Mux.scala 27:73]
  wire [8:0] _s1_predicted_fh_T_97 = _s1_predicted_ghist_ptr_T_32 ?
    s1_possible_predicted_fhs_res_hist_7_new_folded_hist_1 : 9'h0; // @[Mux.scala 27:73]
  wire [8:0] _s1_predicted_fh_T_98 = _s1_predicted_ghist_ptr_T_60 ?
    s1_possible_predicted_fhs_res_hist_7_new_folded_hist_2 : 9'h0; // @[Mux.scala 27:73]
  wire [8:0] _s1_predicted_fh_T_99 = _s1_predicted_fh_T_96 | _s1_predicted_fh_T_97; // @[Mux.scala 27:73]
  wire [7:0] _s1_predicted_fh_T_101 = _s1_predicted_ghist_ptr_T_4 ? s1_possible_predicted_fhs_res_hist_8_new_folded_hist
     : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _s1_predicted_fh_T_102 = _s1_predicted_ghist_ptr_T_32 ?
    s1_possible_predicted_fhs_res_hist_8_new_folded_hist_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _s1_predicted_fh_T_103 = _s1_predicted_ghist_ptr_T_60 ?
    s1_possible_predicted_fhs_res_hist_8_new_folded_hist_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _s1_predicted_fh_T_104 = _s1_predicted_fh_T_101 | _s1_predicted_fh_T_102; // @[Mux.scala 27:73]
  wire [6:0] _s1_predicted_fh_T_106 = _s1_predicted_ghist_ptr_T_4 ? s1_possible_predicted_fhs_res_hist_9_new_folded_hist
     : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _s1_predicted_fh_T_107 = _s1_predicted_ghist_ptr_T_32 ?
    s1_possible_predicted_fhs_res_hist_9_new_folded_hist_1 : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _s1_predicted_fh_T_108 = _s1_predicted_ghist_ptr_T_60 ?
    s1_possible_predicted_fhs_res_hist_9_new_folded_hist_2 : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _s1_predicted_fh_T_109 = _s1_predicted_fh_T_106 | _s1_predicted_fh_T_107; // @[Mux.scala 27:73]
  wire [8:0] _s1_predicted_fh_T_111 = _s1_predicted_ghist_ptr_T_4 ?
    s1_possible_predicted_fhs_res_hist_10_new_folded_hist : 9'h0; // @[Mux.scala 27:73]
  wire [8:0] _s1_predicted_fh_T_112 = _s1_predicted_ghist_ptr_T_32 ?
    s1_possible_predicted_fhs_res_hist_10_new_folded_hist_1 : 9'h0; // @[Mux.scala 27:73]
  wire [8:0] _s1_predicted_fh_T_113 = _s1_predicted_ghist_ptr_T_60 ?
    s1_possible_predicted_fhs_res_hist_10_new_folded_hist_2 : 9'h0; // @[Mux.scala 27:73]
  wire [8:0] _s1_predicted_fh_T_114 = _s1_predicted_fh_T_111 | _s1_predicted_fh_T_112; // @[Mux.scala 27:73]
  wire [7:0] _s1_predicted_fh_T_116 = _s1_predicted_ghist_ptr_T_4 ?
    s1_possible_predicted_fhs_res_hist_11_new_folded_hist : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _s1_predicted_fh_T_117 = _s1_predicted_ghist_ptr_T_32 ?
    s1_possible_predicted_fhs_res_hist_11_new_folded_hist_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _s1_predicted_fh_T_118 = _s1_predicted_ghist_ptr_T_60 ?
    s1_possible_predicted_fhs_res_hist_11_new_folded_hist_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _s1_predicted_fh_T_119 = _s1_predicted_fh_T_116 | _s1_predicted_fh_T_117; // @[Mux.scala 27:73]
  wire [6:0] _s1_predicted_fh_T_121 = _s1_predicted_ghist_ptr_T_4 ?
    s1_possible_predicted_fhs_res_hist_12_new_folded_hist : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _s1_predicted_fh_T_122 = _s1_predicted_ghist_ptr_T_32 ?
    s1_possible_predicted_fhs_res_hist_12_new_folded_hist_1 : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _s1_predicted_fh_T_123 = _s1_predicted_ghist_ptr_T_60 ?
    s1_possible_predicted_fhs_res_hist_12_new_folded_hist_2 : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _s1_predicted_fh_T_124 = _s1_predicted_fh_T_121 | _s1_predicted_fh_T_122; // @[Mux.scala 27:73]
  wire [6:0] _s1_predicted_fh_T_126 = _s1_predicted_ghist_ptr_T_4 ?
    s1_possible_predicted_fhs_res_hist_13_new_folded_hist : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _s1_predicted_fh_T_127 = _s1_predicted_ghist_ptr_T_32 ?
    s1_possible_predicted_fhs_res_hist_13_new_folded_hist_1 : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _s1_predicted_fh_T_128 = _s1_predicted_ghist_ptr_T_60 ?
    s1_possible_predicted_fhs_res_hist_13_new_folded_hist_2 : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _s1_predicted_fh_T_129 = _s1_predicted_fh_T_126 | _s1_predicted_fh_T_127; // @[Mux.scala 27:73]
  wire [6:0] _s1_predicted_fh_T_131 = _s1_predicted_ghist_ptr_T_4 ?
    s1_possible_predicted_fhs_res_hist_14_new_folded_hist : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _s1_predicted_fh_T_132 = _s1_predicted_ghist_ptr_T_32 ?
    s1_possible_predicted_fhs_res_hist_14_new_folded_hist_1 : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _s1_predicted_fh_T_133 = _s1_predicted_ghist_ptr_T_60 ?
    s1_possible_predicted_fhs_res_hist_14_new_folded_hist_2 : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _s1_predicted_fh_T_134 = _s1_predicted_fh_T_131 | _s1_predicted_fh_T_132; // @[Mux.scala 27:73]
  wire [10:0] _s1_predicted_fh_T_136 = _s1_predicted_ghist_ptr_T_4 ?
    s1_possible_predicted_fhs_res_hist_15_new_folded_hist : 11'h0; // @[Mux.scala 27:73]
  wire [10:0] _s1_predicted_fh_T_137 = _s1_predicted_ghist_ptr_T_32 ?
    s1_possible_predicted_fhs_res_hist_15_new_folded_hist_1 : 11'h0; // @[Mux.scala 27:73]
  wire [10:0] _s1_predicted_fh_T_138 = _s1_predicted_ghist_ptr_T_60 ?
    s1_possible_predicted_fhs_res_hist_15_new_folded_hist_2 : 11'h0; // @[Mux.scala 27:73]
  wire [10:0] _s1_predicted_fh_T_139 = _s1_predicted_fh_T_136 | _s1_predicted_fh_T_137; // @[Mux.scala 27:73]
  wire [7:0] _s1_predicted_fh_T_141 = _s1_predicted_ghist_ptr_T_4 ?
    s1_possible_predicted_fhs_res_hist_16_new_folded_hist : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _s1_predicted_fh_T_142 = _s1_predicted_ghist_ptr_T_32 ?
    s1_possible_predicted_fhs_res_hist_16_new_folded_hist_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _s1_predicted_fh_T_143 = _s1_predicted_ghist_ptr_T_60 ?
    s1_possible_predicted_fhs_res_hist_16_new_folded_hist_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _s1_predicted_fh_T_144 = _s1_predicted_fh_T_141 | _s1_predicted_fh_T_142; // @[Mux.scala 27:73]
  wire [7:0] _s1_predicted_fh_T_146 = _s1_predicted_ghist_ptr_T_4 ?
    s1_possible_predicted_fhs_res_hist_17_new_folded_hist : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _s1_predicted_fh_T_147 = _s1_predicted_ghist_ptr_T_32 ?
    s1_possible_predicted_fhs_res_hist_17_new_folded_hist_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _s1_predicted_fh_T_148 = _s1_predicted_ghist_ptr_T_60 ?
    s1_possible_predicted_fhs_res_hist_17_new_folded_hist_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _s1_predicted_fh_T_149 = _s1_predicted_fh_T_146 | _s1_predicted_fh_T_147; // @[Mux.scala 27:73]
  wire [8:0] new_value = s1_ghist_ptr_value + 8'h74; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_1 = {1'h0,new_value}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff = $signed(_diff_T_1) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag = $signed(diff) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T = $signed(_diff_T_1) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_1 = reverse_flag ? _new_ptr_value_T : {{1'd0}, new_value}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_1 = s1_ghist_ptr_value + 8'h6; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_7 = {1'h0,new_value_1}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_1 = $signed(_diff_T_7) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_1 = $signed(diff_1) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_2 = $signed(_diff_T_7) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_3 = reverse_flag_1 ? _new_ptr_value_T_2 : {{1'd0}, new_value_1}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_2 = s1_ghist_ptr_value + 8'hb; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_13 = {1'h0,new_value_2}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_2 = $signed(_diff_T_13) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_2 = $signed(diff_2) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_4 = $signed(_diff_T_13) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_5 = reverse_flag_2 ? _new_ptr_value_T_4 : {{1'd0}, new_value_2}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_3 = s1_ghist_ptr_value + 8'hf; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_19 = {1'h0,new_value_3}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_3 = $signed(_diff_T_19) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_3 = $signed(diff_3) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_6 = $signed(_diff_T_19) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_7 = reverse_flag_3 ? _new_ptr_value_T_6 : {{1'd0}, new_value_3}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_4 = s1_ghist_ptr_value + 8'h1e; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_25 = {1'h0,new_value_4}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_4 = $signed(_diff_T_25) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_4 = $signed(diff_4) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_8 = $signed(_diff_T_25) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_9 = reverse_flag_4 ? _new_ptr_value_T_8 : {{1'd0}, new_value_4}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_5 = s1_ghist_ptr_value + 8'h75; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_31 = {1'h0,new_value_5}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_5 = $signed(_diff_T_31) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_5 = $signed(diff_5) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_10 = $signed(_diff_T_31) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_11 = reverse_flag_5 ? _new_ptr_value_T_10 : {{1'd0}, new_value_5}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_6 = s1_ghist_ptr_value + 8'h7; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_37 = {1'h0,new_value_6}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_6 = $signed(_diff_T_37) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_6 = $signed(diff_6) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_12 = $signed(_diff_T_37) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_13 = reverse_flag_6 ? _new_ptr_value_T_12 : {{1'd0}, new_value_6}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_7 = s1_ghist_ptr_value + 8'h76; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_43 = {1'h0,new_value_7}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_7 = $signed(_diff_T_43) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_7 = $signed(diff_7) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_14 = $signed(_diff_T_43) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_15 = reverse_flag_7 ? _new_ptr_value_T_14 : {{1'd0}, new_value_7}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_8 = s1_ghist_ptr_value + 8'h1d; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_49 = {1'h0,new_value_8}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_8 = $signed(_diff_T_49) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_8 = $signed(diff_8) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_16 = $signed(_diff_T_49) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_17 = reverse_flag_8 ? _new_ptr_value_T_16 : {{1'd0}, new_value_8}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_9 = s1_ghist_ptr_value + 8'ha; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_55 = {1'h0,new_value_9}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_9 = $signed(_diff_T_55) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_9 = $signed(diff_9) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_18 = $signed(_diff_T_55) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_19 = reverse_flag_9 ? _new_ptr_value_T_18 : {{1'd0}, new_value_9}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_10 = s1_ghist_ptr_value + 8'he; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_61 = {1'h0,new_value_10}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_10 = $signed(_diff_T_61) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_10 = $signed(diff_10) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_20 = $signed(_diff_T_61) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_21 = reverse_flag_10 ? _new_ptr_value_T_20 : {{1'd0}, new_value_10}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_11 = s1_ghist_ptr_value + 8'h77; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_67 = {1'h0,new_value_11}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_11 = $signed(_diff_T_67) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_11 = $signed(diff_11) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_22 = $signed(_diff_T_67) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_23 = reverse_flag_11 ? _new_ptr_value_T_22 : {{1'd0}, new_value_11}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_12 = s1_ghist_ptr_value + 8'hd; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_73 = {1'h0,new_value_12}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_12 = $signed(_diff_T_73) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_12 = $signed(diff_12) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_24 = $signed(_diff_T_73) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_25 = reverse_flag_12 ? _new_ptr_value_T_24 : {{1'd0}, new_value_12}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_13 = s1_ghist_ptr_value + 8'h8; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_79 = {1'h0,new_value_13}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_13 = $signed(_diff_T_79) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_13 = $signed(diff_13) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_26 = $signed(_diff_T_79) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_27 = reverse_flag_13 ? _new_ptr_value_T_26 : {{1'd0}, new_value_13}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_14 = s1_ghist_ptr_value + 8'h20; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_85 = {1'h0,new_value_14}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_14 = $signed(_diff_T_85) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_14 = $signed(diff_14) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_28 = $signed(_diff_T_85) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_29 = reverse_flag_14 ? _new_ptr_value_T_28 : {{1'd0}, new_value_14}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_15 = s1_ghist_ptr_value + 8'hc; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_91 = {1'h0,new_value_15}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_15 = $signed(_diff_T_91) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_15 = $signed(diff_15) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_30 = $signed(_diff_T_91) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_31 = reverse_flag_15 ? _new_ptr_value_T_30 : {{1'd0}, new_value_15}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_16 = s1_ghist_ptr_value + 8'h9; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_97 = {1'h0,new_value_16}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_16 = $signed(_diff_T_97) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_16 = $signed(diff_16) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_32 = $signed(_diff_T_97) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_33 = reverse_flag_16 ? _new_ptr_value_T_32 : {{1'd0}, new_value_16}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_17 = s1_ghist_ptr_value + 8'h1f; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_103 = {1'h0,new_value_17}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_17 = $signed(_diff_T_103) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_17 = $signed(diff_17) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_34 = $signed(_diff_T_103) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_35 = reverse_flag_17 ? _new_ptr_value_T_34 : {{1'd0}, new_value_17}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_18 = s1_ghist_ptr_value + 8'h5; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_109 = {1'h0,new_value_18}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_18 = $signed(_diff_T_109) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_18 = $signed(diff_18) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_36 = $signed(_diff_T_109) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_37 = reverse_flag_18 ? _new_ptr_value_T_36 : {{1'd0}, new_value_18}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_19 = s1_ghist_ptr_value + 8'h10; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_115 = {1'h0,new_value_19}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_19 = $signed(_diff_T_115) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_19 = $signed(diff_19) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_38 = $signed(_diff_T_115) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_39 = reverse_flag_19 ? _new_ptr_value_T_38 : {{1'd0}, new_value_19}; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] new_ptr_9_value = _new_ptr_value_T_19[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_150 = 8'h1 == new_ptr_9_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_151 = 8'h2 == new_ptr_9_value ? ghv_2 : _GEN_150; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_152 = 8'h3 == new_ptr_9_value ? ghv_3 : _GEN_151; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_153 = 8'h4 == new_ptr_9_value ? ghv_4 : _GEN_152; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_154 = 8'h5 == new_ptr_9_value ? ghv_5 : _GEN_153; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_155 = 8'h6 == new_ptr_9_value ? ghv_6 : _GEN_154; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_156 = 8'h7 == new_ptr_9_value ? ghv_7 : _GEN_155; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_157 = 8'h8 == new_ptr_9_value ? ghv_8 : _GEN_156; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_158 = 8'h9 == new_ptr_9_value ? ghv_9 : _GEN_157; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_159 = 8'ha == new_ptr_9_value ? ghv_10 : _GEN_158; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_160 = 8'hb == new_ptr_9_value ? ghv_11 : _GEN_159; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_161 = 8'hc == new_ptr_9_value ? ghv_12 : _GEN_160; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_162 = 8'hd == new_ptr_9_value ? ghv_13 : _GEN_161; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_163 = 8'he == new_ptr_9_value ? ghv_14 : _GEN_162; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_164 = 8'hf == new_ptr_9_value ? ghv_15 : _GEN_163; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_165 = 8'h10 == new_ptr_9_value ? ghv_16 : _GEN_164; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_166 = 8'h11 == new_ptr_9_value ? ghv_17 : _GEN_165; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_167 = 8'h12 == new_ptr_9_value ? ghv_18 : _GEN_166; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_168 = 8'h13 == new_ptr_9_value ? ghv_19 : _GEN_167; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_169 = 8'h14 == new_ptr_9_value ? ghv_20 : _GEN_168; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_170 = 8'h15 == new_ptr_9_value ? ghv_21 : _GEN_169; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_171 = 8'h16 == new_ptr_9_value ? ghv_22 : _GEN_170; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_172 = 8'h17 == new_ptr_9_value ? ghv_23 : _GEN_171; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_173 = 8'h18 == new_ptr_9_value ? ghv_24 : _GEN_172; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_174 = 8'h19 == new_ptr_9_value ? ghv_25 : _GEN_173; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_175 = 8'h1a == new_ptr_9_value ? ghv_26 : _GEN_174; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_176 = 8'h1b == new_ptr_9_value ? ghv_27 : _GEN_175; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_177 = 8'h1c == new_ptr_9_value ? ghv_28 : _GEN_176; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_178 = 8'h1d == new_ptr_9_value ? ghv_29 : _GEN_177; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_179 = 8'h1e == new_ptr_9_value ? ghv_30 : _GEN_178; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_180 = 8'h1f == new_ptr_9_value ? ghv_31 : _GEN_179; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_181 = 8'h20 == new_ptr_9_value ? ghv_32 : _GEN_180; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_182 = 8'h21 == new_ptr_9_value ? ghv_33 : _GEN_181; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_183 = 8'h22 == new_ptr_9_value ? ghv_34 : _GEN_182; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_184 = 8'h23 == new_ptr_9_value ? ghv_35 : _GEN_183; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_185 = 8'h24 == new_ptr_9_value ? ghv_36 : _GEN_184; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_186 = 8'h25 == new_ptr_9_value ? ghv_37 : _GEN_185; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_187 = 8'h26 == new_ptr_9_value ? ghv_38 : _GEN_186; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_188 = 8'h27 == new_ptr_9_value ? ghv_39 : _GEN_187; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_189 = 8'h28 == new_ptr_9_value ? ghv_40 : _GEN_188; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_190 = 8'h29 == new_ptr_9_value ? ghv_41 : _GEN_189; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_191 = 8'h2a == new_ptr_9_value ? ghv_42 : _GEN_190; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_192 = 8'h2b == new_ptr_9_value ? ghv_43 : _GEN_191; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_193 = 8'h2c == new_ptr_9_value ? ghv_44 : _GEN_192; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_194 = 8'h2d == new_ptr_9_value ? ghv_45 : _GEN_193; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_195 = 8'h2e == new_ptr_9_value ? ghv_46 : _GEN_194; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_196 = 8'h2f == new_ptr_9_value ? ghv_47 : _GEN_195; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_197 = 8'h30 == new_ptr_9_value ? ghv_48 : _GEN_196; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_198 = 8'h31 == new_ptr_9_value ? ghv_49 : _GEN_197; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_199 = 8'h32 == new_ptr_9_value ? ghv_50 : _GEN_198; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_200 = 8'h33 == new_ptr_9_value ? ghv_51 : _GEN_199; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_201 = 8'h34 == new_ptr_9_value ? ghv_52 : _GEN_200; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_202 = 8'h35 == new_ptr_9_value ? ghv_53 : _GEN_201; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_203 = 8'h36 == new_ptr_9_value ? ghv_54 : _GEN_202; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_204 = 8'h37 == new_ptr_9_value ? ghv_55 : _GEN_203; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_205 = 8'h38 == new_ptr_9_value ? ghv_56 : _GEN_204; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_206 = 8'h39 == new_ptr_9_value ? ghv_57 : _GEN_205; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_207 = 8'h3a == new_ptr_9_value ? ghv_58 : _GEN_206; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_208 = 8'h3b == new_ptr_9_value ? ghv_59 : _GEN_207; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_209 = 8'h3c == new_ptr_9_value ? ghv_60 : _GEN_208; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_210 = 8'h3d == new_ptr_9_value ? ghv_61 : _GEN_209; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_211 = 8'h3e == new_ptr_9_value ? ghv_62 : _GEN_210; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_212 = 8'h3f == new_ptr_9_value ? ghv_63 : _GEN_211; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_213 = 8'h40 == new_ptr_9_value ? ghv_64 : _GEN_212; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_214 = 8'h41 == new_ptr_9_value ? ghv_65 : _GEN_213; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_215 = 8'h42 == new_ptr_9_value ? ghv_66 : _GEN_214; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_216 = 8'h43 == new_ptr_9_value ? ghv_67 : _GEN_215; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_217 = 8'h44 == new_ptr_9_value ? ghv_68 : _GEN_216; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_218 = 8'h45 == new_ptr_9_value ? ghv_69 : _GEN_217; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_219 = 8'h46 == new_ptr_9_value ? ghv_70 : _GEN_218; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_220 = 8'h47 == new_ptr_9_value ? ghv_71 : _GEN_219; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_221 = 8'h48 == new_ptr_9_value ? ghv_72 : _GEN_220; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_222 = 8'h49 == new_ptr_9_value ? ghv_73 : _GEN_221; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_223 = 8'h4a == new_ptr_9_value ? ghv_74 : _GEN_222; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_224 = 8'h4b == new_ptr_9_value ? ghv_75 : _GEN_223; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_225 = 8'h4c == new_ptr_9_value ? ghv_76 : _GEN_224; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_226 = 8'h4d == new_ptr_9_value ? ghv_77 : _GEN_225; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_227 = 8'h4e == new_ptr_9_value ? ghv_78 : _GEN_226; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_228 = 8'h4f == new_ptr_9_value ? ghv_79 : _GEN_227; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_229 = 8'h50 == new_ptr_9_value ? ghv_80 : _GEN_228; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_230 = 8'h51 == new_ptr_9_value ? ghv_81 : _GEN_229; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_231 = 8'h52 == new_ptr_9_value ? ghv_82 : _GEN_230; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_232 = 8'h53 == new_ptr_9_value ? ghv_83 : _GEN_231; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_233 = 8'h54 == new_ptr_9_value ? ghv_84 : _GEN_232; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_234 = 8'h55 == new_ptr_9_value ? ghv_85 : _GEN_233; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_235 = 8'h56 == new_ptr_9_value ? ghv_86 : _GEN_234; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_236 = 8'h57 == new_ptr_9_value ? ghv_87 : _GEN_235; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_237 = 8'h58 == new_ptr_9_value ? ghv_88 : _GEN_236; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_238 = 8'h59 == new_ptr_9_value ? ghv_89 : _GEN_237; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_239 = 8'h5a == new_ptr_9_value ? ghv_90 : _GEN_238; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_240 = 8'h5b == new_ptr_9_value ? ghv_91 : _GEN_239; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_241 = 8'h5c == new_ptr_9_value ? ghv_92 : _GEN_240; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_242 = 8'h5d == new_ptr_9_value ? ghv_93 : _GEN_241; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_243 = 8'h5e == new_ptr_9_value ? ghv_94 : _GEN_242; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_244 = 8'h5f == new_ptr_9_value ? ghv_95 : _GEN_243; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_245 = 8'h60 == new_ptr_9_value ? ghv_96 : _GEN_244; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_246 = 8'h61 == new_ptr_9_value ? ghv_97 : _GEN_245; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_247 = 8'h62 == new_ptr_9_value ? ghv_98 : _GEN_246; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_248 = 8'h63 == new_ptr_9_value ? ghv_99 : _GEN_247; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_249 = 8'h64 == new_ptr_9_value ? ghv_100 : _GEN_248; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_250 = 8'h65 == new_ptr_9_value ? ghv_101 : _GEN_249; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_251 = 8'h66 == new_ptr_9_value ? ghv_102 : _GEN_250; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_252 = 8'h67 == new_ptr_9_value ? ghv_103 : _GEN_251; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_253 = 8'h68 == new_ptr_9_value ? ghv_104 : _GEN_252; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_254 = 8'h69 == new_ptr_9_value ? ghv_105 : _GEN_253; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_255 = 8'h6a == new_ptr_9_value ? ghv_106 : _GEN_254; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_256 = 8'h6b == new_ptr_9_value ? ghv_107 : _GEN_255; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_257 = 8'h6c == new_ptr_9_value ? ghv_108 : _GEN_256; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_258 = 8'h6d == new_ptr_9_value ? ghv_109 : _GEN_257; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_259 = 8'h6e == new_ptr_9_value ? ghv_110 : _GEN_258; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_260 = 8'h6f == new_ptr_9_value ? ghv_111 : _GEN_259; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_261 = 8'h70 == new_ptr_9_value ? ghv_112 : _GEN_260; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_262 = 8'h71 == new_ptr_9_value ? ghv_113 : _GEN_261; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_263 = 8'h72 == new_ptr_9_value ? ghv_114 : _GEN_262; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_264 = 8'h73 == new_ptr_9_value ? ghv_115 : _GEN_263; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_265 = 8'h74 == new_ptr_9_value ? ghv_116 : _GEN_264; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_266 = 8'h75 == new_ptr_9_value ? ghv_117 : _GEN_265; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_267 = 8'h76 == new_ptr_9_value ? ghv_118 : _GEN_266; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_268 = 8'h77 == new_ptr_9_value ? ghv_119 : _GEN_267; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_269 = 8'h78 == new_ptr_9_value ? ghv_120 : _GEN_268; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_270 = 8'h79 == new_ptr_9_value ? ghv_121 : _GEN_269; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_271 = 8'h7a == new_ptr_9_value ? ghv_122 : _GEN_270; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_272 = 8'h7b == new_ptr_9_value ? ghv_123 : _GEN_271; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_273 = 8'h7c == new_ptr_9_value ? ghv_124 : _GEN_272; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_274 = 8'h7d == new_ptr_9_value ? ghv_125 : _GEN_273; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_275 = 8'h7e == new_ptr_9_value ? ghv_126 : _GEN_274; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_276 = 8'h7f == new_ptr_9_value ? ghv_127 : _GEN_275; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_277 = 8'h80 == new_ptr_9_value ? ghv_128 : _GEN_276; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_278 = 8'h81 == new_ptr_9_value ? ghv_129 : _GEN_277; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_279 = 8'h82 == new_ptr_9_value ? ghv_130 : _GEN_278; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_280 = 8'h83 == new_ptr_9_value ? ghv_131 : _GEN_279; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_281 = 8'h84 == new_ptr_9_value ? ghv_132 : _GEN_280; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_282 = 8'h85 == new_ptr_9_value ? ghv_133 : _GEN_281; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_283 = 8'h86 == new_ptr_9_value ? ghv_134 : _GEN_282; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_284 = 8'h87 == new_ptr_9_value ? ghv_135 : _GEN_283; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_285 = 8'h88 == new_ptr_9_value ? ghv_136 : _GEN_284; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_286 = 8'h89 == new_ptr_9_value ? ghv_137 : _GEN_285; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_287 = 8'h8a == new_ptr_9_value ? ghv_138 : _GEN_286; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_288 = 8'h8b == new_ptr_9_value ? ghv_139 : _GEN_287; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_289 = 8'h8c == new_ptr_9_value ? ghv_140 : _GEN_288; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_290 = 8'h8d == new_ptr_9_value ? ghv_141 : _GEN_289; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_291 = 8'h8e == new_ptr_9_value ? ghv_142 : _GEN_290; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_16_value = _new_ptr_value_T_33[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_294 = 8'h1 == new_ptr_16_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_295 = 8'h2 == new_ptr_16_value ? ghv_2 : _GEN_294; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_296 = 8'h3 == new_ptr_16_value ? ghv_3 : _GEN_295; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_297 = 8'h4 == new_ptr_16_value ? ghv_4 : _GEN_296; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_298 = 8'h5 == new_ptr_16_value ? ghv_5 : _GEN_297; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_299 = 8'h6 == new_ptr_16_value ? ghv_6 : _GEN_298; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_300 = 8'h7 == new_ptr_16_value ? ghv_7 : _GEN_299; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_301 = 8'h8 == new_ptr_16_value ? ghv_8 : _GEN_300; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_302 = 8'h9 == new_ptr_16_value ? ghv_9 : _GEN_301; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_303 = 8'ha == new_ptr_16_value ? ghv_10 : _GEN_302; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_304 = 8'hb == new_ptr_16_value ? ghv_11 : _GEN_303; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_305 = 8'hc == new_ptr_16_value ? ghv_12 : _GEN_304; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_306 = 8'hd == new_ptr_16_value ? ghv_13 : _GEN_305; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_307 = 8'he == new_ptr_16_value ? ghv_14 : _GEN_306; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_308 = 8'hf == new_ptr_16_value ? ghv_15 : _GEN_307; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_309 = 8'h10 == new_ptr_16_value ? ghv_16 : _GEN_308; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_310 = 8'h11 == new_ptr_16_value ? ghv_17 : _GEN_309; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_311 = 8'h12 == new_ptr_16_value ? ghv_18 : _GEN_310; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_312 = 8'h13 == new_ptr_16_value ? ghv_19 : _GEN_311; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_313 = 8'h14 == new_ptr_16_value ? ghv_20 : _GEN_312; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_314 = 8'h15 == new_ptr_16_value ? ghv_21 : _GEN_313; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_315 = 8'h16 == new_ptr_16_value ? ghv_22 : _GEN_314; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_316 = 8'h17 == new_ptr_16_value ? ghv_23 : _GEN_315; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_317 = 8'h18 == new_ptr_16_value ? ghv_24 : _GEN_316; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_318 = 8'h19 == new_ptr_16_value ? ghv_25 : _GEN_317; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_319 = 8'h1a == new_ptr_16_value ? ghv_26 : _GEN_318; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_320 = 8'h1b == new_ptr_16_value ? ghv_27 : _GEN_319; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_321 = 8'h1c == new_ptr_16_value ? ghv_28 : _GEN_320; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_322 = 8'h1d == new_ptr_16_value ? ghv_29 : _GEN_321; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_323 = 8'h1e == new_ptr_16_value ? ghv_30 : _GEN_322; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_324 = 8'h1f == new_ptr_16_value ? ghv_31 : _GEN_323; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_325 = 8'h20 == new_ptr_16_value ? ghv_32 : _GEN_324; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_326 = 8'h21 == new_ptr_16_value ? ghv_33 : _GEN_325; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_327 = 8'h22 == new_ptr_16_value ? ghv_34 : _GEN_326; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_328 = 8'h23 == new_ptr_16_value ? ghv_35 : _GEN_327; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_329 = 8'h24 == new_ptr_16_value ? ghv_36 : _GEN_328; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_330 = 8'h25 == new_ptr_16_value ? ghv_37 : _GEN_329; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_331 = 8'h26 == new_ptr_16_value ? ghv_38 : _GEN_330; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_332 = 8'h27 == new_ptr_16_value ? ghv_39 : _GEN_331; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_333 = 8'h28 == new_ptr_16_value ? ghv_40 : _GEN_332; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_334 = 8'h29 == new_ptr_16_value ? ghv_41 : _GEN_333; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_335 = 8'h2a == new_ptr_16_value ? ghv_42 : _GEN_334; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_336 = 8'h2b == new_ptr_16_value ? ghv_43 : _GEN_335; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_337 = 8'h2c == new_ptr_16_value ? ghv_44 : _GEN_336; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_338 = 8'h2d == new_ptr_16_value ? ghv_45 : _GEN_337; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_339 = 8'h2e == new_ptr_16_value ? ghv_46 : _GEN_338; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_340 = 8'h2f == new_ptr_16_value ? ghv_47 : _GEN_339; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_341 = 8'h30 == new_ptr_16_value ? ghv_48 : _GEN_340; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_342 = 8'h31 == new_ptr_16_value ? ghv_49 : _GEN_341; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_343 = 8'h32 == new_ptr_16_value ? ghv_50 : _GEN_342; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_344 = 8'h33 == new_ptr_16_value ? ghv_51 : _GEN_343; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_345 = 8'h34 == new_ptr_16_value ? ghv_52 : _GEN_344; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_346 = 8'h35 == new_ptr_16_value ? ghv_53 : _GEN_345; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_347 = 8'h36 == new_ptr_16_value ? ghv_54 : _GEN_346; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_348 = 8'h37 == new_ptr_16_value ? ghv_55 : _GEN_347; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_349 = 8'h38 == new_ptr_16_value ? ghv_56 : _GEN_348; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_350 = 8'h39 == new_ptr_16_value ? ghv_57 : _GEN_349; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_351 = 8'h3a == new_ptr_16_value ? ghv_58 : _GEN_350; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_352 = 8'h3b == new_ptr_16_value ? ghv_59 : _GEN_351; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_353 = 8'h3c == new_ptr_16_value ? ghv_60 : _GEN_352; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_354 = 8'h3d == new_ptr_16_value ? ghv_61 : _GEN_353; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_355 = 8'h3e == new_ptr_16_value ? ghv_62 : _GEN_354; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_356 = 8'h3f == new_ptr_16_value ? ghv_63 : _GEN_355; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_357 = 8'h40 == new_ptr_16_value ? ghv_64 : _GEN_356; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_358 = 8'h41 == new_ptr_16_value ? ghv_65 : _GEN_357; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_359 = 8'h42 == new_ptr_16_value ? ghv_66 : _GEN_358; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_360 = 8'h43 == new_ptr_16_value ? ghv_67 : _GEN_359; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_361 = 8'h44 == new_ptr_16_value ? ghv_68 : _GEN_360; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_362 = 8'h45 == new_ptr_16_value ? ghv_69 : _GEN_361; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_363 = 8'h46 == new_ptr_16_value ? ghv_70 : _GEN_362; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_364 = 8'h47 == new_ptr_16_value ? ghv_71 : _GEN_363; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_365 = 8'h48 == new_ptr_16_value ? ghv_72 : _GEN_364; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_366 = 8'h49 == new_ptr_16_value ? ghv_73 : _GEN_365; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_367 = 8'h4a == new_ptr_16_value ? ghv_74 : _GEN_366; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_368 = 8'h4b == new_ptr_16_value ? ghv_75 : _GEN_367; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_369 = 8'h4c == new_ptr_16_value ? ghv_76 : _GEN_368; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_370 = 8'h4d == new_ptr_16_value ? ghv_77 : _GEN_369; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_371 = 8'h4e == new_ptr_16_value ? ghv_78 : _GEN_370; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_372 = 8'h4f == new_ptr_16_value ? ghv_79 : _GEN_371; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_373 = 8'h50 == new_ptr_16_value ? ghv_80 : _GEN_372; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_374 = 8'h51 == new_ptr_16_value ? ghv_81 : _GEN_373; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_375 = 8'h52 == new_ptr_16_value ? ghv_82 : _GEN_374; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_376 = 8'h53 == new_ptr_16_value ? ghv_83 : _GEN_375; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_377 = 8'h54 == new_ptr_16_value ? ghv_84 : _GEN_376; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_378 = 8'h55 == new_ptr_16_value ? ghv_85 : _GEN_377; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_379 = 8'h56 == new_ptr_16_value ? ghv_86 : _GEN_378; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_380 = 8'h57 == new_ptr_16_value ? ghv_87 : _GEN_379; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_381 = 8'h58 == new_ptr_16_value ? ghv_88 : _GEN_380; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_382 = 8'h59 == new_ptr_16_value ? ghv_89 : _GEN_381; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_383 = 8'h5a == new_ptr_16_value ? ghv_90 : _GEN_382; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_384 = 8'h5b == new_ptr_16_value ? ghv_91 : _GEN_383; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_385 = 8'h5c == new_ptr_16_value ? ghv_92 : _GEN_384; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_386 = 8'h5d == new_ptr_16_value ? ghv_93 : _GEN_385; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_387 = 8'h5e == new_ptr_16_value ? ghv_94 : _GEN_386; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_388 = 8'h5f == new_ptr_16_value ? ghv_95 : _GEN_387; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_389 = 8'h60 == new_ptr_16_value ? ghv_96 : _GEN_388; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_390 = 8'h61 == new_ptr_16_value ? ghv_97 : _GEN_389; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_391 = 8'h62 == new_ptr_16_value ? ghv_98 : _GEN_390; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_392 = 8'h63 == new_ptr_16_value ? ghv_99 : _GEN_391; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_393 = 8'h64 == new_ptr_16_value ? ghv_100 : _GEN_392; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_394 = 8'h65 == new_ptr_16_value ? ghv_101 : _GEN_393; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_395 = 8'h66 == new_ptr_16_value ? ghv_102 : _GEN_394; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_396 = 8'h67 == new_ptr_16_value ? ghv_103 : _GEN_395; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_397 = 8'h68 == new_ptr_16_value ? ghv_104 : _GEN_396; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_398 = 8'h69 == new_ptr_16_value ? ghv_105 : _GEN_397; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_399 = 8'h6a == new_ptr_16_value ? ghv_106 : _GEN_398; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_400 = 8'h6b == new_ptr_16_value ? ghv_107 : _GEN_399; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_401 = 8'h6c == new_ptr_16_value ? ghv_108 : _GEN_400; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_402 = 8'h6d == new_ptr_16_value ? ghv_109 : _GEN_401; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_403 = 8'h6e == new_ptr_16_value ? ghv_110 : _GEN_402; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_404 = 8'h6f == new_ptr_16_value ? ghv_111 : _GEN_403; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_405 = 8'h70 == new_ptr_16_value ? ghv_112 : _GEN_404; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_406 = 8'h71 == new_ptr_16_value ? ghv_113 : _GEN_405; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_407 = 8'h72 == new_ptr_16_value ? ghv_114 : _GEN_406; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_408 = 8'h73 == new_ptr_16_value ? ghv_115 : _GEN_407; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_409 = 8'h74 == new_ptr_16_value ? ghv_116 : _GEN_408; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_410 = 8'h75 == new_ptr_16_value ? ghv_117 : _GEN_409; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_411 = 8'h76 == new_ptr_16_value ? ghv_118 : _GEN_410; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_412 = 8'h77 == new_ptr_16_value ? ghv_119 : _GEN_411; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_413 = 8'h78 == new_ptr_16_value ? ghv_120 : _GEN_412; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_414 = 8'h79 == new_ptr_16_value ? ghv_121 : _GEN_413; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_415 = 8'h7a == new_ptr_16_value ? ghv_122 : _GEN_414; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_416 = 8'h7b == new_ptr_16_value ? ghv_123 : _GEN_415; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_417 = 8'h7c == new_ptr_16_value ? ghv_124 : _GEN_416; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_418 = 8'h7d == new_ptr_16_value ? ghv_125 : _GEN_417; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_419 = 8'h7e == new_ptr_16_value ? ghv_126 : _GEN_418; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_420 = 8'h7f == new_ptr_16_value ? ghv_127 : _GEN_419; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_421 = 8'h80 == new_ptr_16_value ? ghv_128 : _GEN_420; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_422 = 8'h81 == new_ptr_16_value ? ghv_129 : _GEN_421; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_423 = 8'h82 == new_ptr_16_value ? ghv_130 : _GEN_422; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_424 = 8'h83 == new_ptr_16_value ? ghv_131 : _GEN_423; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_425 = 8'h84 == new_ptr_16_value ? ghv_132 : _GEN_424; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_426 = 8'h85 == new_ptr_16_value ? ghv_133 : _GEN_425; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_427 = 8'h86 == new_ptr_16_value ? ghv_134 : _GEN_426; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_428 = 8'h87 == new_ptr_16_value ? ghv_135 : _GEN_427; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_429 = 8'h88 == new_ptr_16_value ? ghv_136 : _GEN_428; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_430 = 8'h89 == new_ptr_16_value ? ghv_137 : _GEN_429; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_431 = 8'h8a == new_ptr_16_value ? ghv_138 : _GEN_430; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_432 = 8'h8b == new_ptr_16_value ? ghv_139 : _GEN_431; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_433 = 8'h8c == new_ptr_16_value ? ghv_140 : _GEN_432; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_434 = 8'h8d == new_ptr_16_value ? ghv_141 : _GEN_433; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_435 = 8'h8e == new_ptr_16_value ? ghv_142 : _GEN_434; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_13_value = _new_ptr_value_T_27[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_438 = 8'h1 == new_ptr_13_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_439 = 8'h2 == new_ptr_13_value ? ghv_2 : _GEN_438; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_440 = 8'h3 == new_ptr_13_value ? ghv_3 : _GEN_439; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_441 = 8'h4 == new_ptr_13_value ? ghv_4 : _GEN_440; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_442 = 8'h5 == new_ptr_13_value ? ghv_5 : _GEN_441; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_443 = 8'h6 == new_ptr_13_value ? ghv_6 : _GEN_442; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_444 = 8'h7 == new_ptr_13_value ? ghv_7 : _GEN_443; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_445 = 8'h8 == new_ptr_13_value ? ghv_8 : _GEN_444; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_446 = 8'h9 == new_ptr_13_value ? ghv_9 : _GEN_445; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_447 = 8'ha == new_ptr_13_value ? ghv_10 : _GEN_446; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_448 = 8'hb == new_ptr_13_value ? ghv_11 : _GEN_447; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_449 = 8'hc == new_ptr_13_value ? ghv_12 : _GEN_448; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_450 = 8'hd == new_ptr_13_value ? ghv_13 : _GEN_449; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_451 = 8'he == new_ptr_13_value ? ghv_14 : _GEN_450; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_452 = 8'hf == new_ptr_13_value ? ghv_15 : _GEN_451; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_453 = 8'h10 == new_ptr_13_value ? ghv_16 : _GEN_452; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_454 = 8'h11 == new_ptr_13_value ? ghv_17 : _GEN_453; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_455 = 8'h12 == new_ptr_13_value ? ghv_18 : _GEN_454; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_456 = 8'h13 == new_ptr_13_value ? ghv_19 : _GEN_455; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_457 = 8'h14 == new_ptr_13_value ? ghv_20 : _GEN_456; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_458 = 8'h15 == new_ptr_13_value ? ghv_21 : _GEN_457; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_459 = 8'h16 == new_ptr_13_value ? ghv_22 : _GEN_458; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_460 = 8'h17 == new_ptr_13_value ? ghv_23 : _GEN_459; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_461 = 8'h18 == new_ptr_13_value ? ghv_24 : _GEN_460; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_462 = 8'h19 == new_ptr_13_value ? ghv_25 : _GEN_461; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_463 = 8'h1a == new_ptr_13_value ? ghv_26 : _GEN_462; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_464 = 8'h1b == new_ptr_13_value ? ghv_27 : _GEN_463; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_465 = 8'h1c == new_ptr_13_value ? ghv_28 : _GEN_464; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_466 = 8'h1d == new_ptr_13_value ? ghv_29 : _GEN_465; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_467 = 8'h1e == new_ptr_13_value ? ghv_30 : _GEN_466; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_468 = 8'h1f == new_ptr_13_value ? ghv_31 : _GEN_467; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_469 = 8'h20 == new_ptr_13_value ? ghv_32 : _GEN_468; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_470 = 8'h21 == new_ptr_13_value ? ghv_33 : _GEN_469; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_471 = 8'h22 == new_ptr_13_value ? ghv_34 : _GEN_470; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_472 = 8'h23 == new_ptr_13_value ? ghv_35 : _GEN_471; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_473 = 8'h24 == new_ptr_13_value ? ghv_36 : _GEN_472; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_474 = 8'h25 == new_ptr_13_value ? ghv_37 : _GEN_473; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_475 = 8'h26 == new_ptr_13_value ? ghv_38 : _GEN_474; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_476 = 8'h27 == new_ptr_13_value ? ghv_39 : _GEN_475; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_477 = 8'h28 == new_ptr_13_value ? ghv_40 : _GEN_476; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_478 = 8'h29 == new_ptr_13_value ? ghv_41 : _GEN_477; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_479 = 8'h2a == new_ptr_13_value ? ghv_42 : _GEN_478; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_480 = 8'h2b == new_ptr_13_value ? ghv_43 : _GEN_479; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_481 = 8'h2c == new_ptr_13_value ? ghv_44 : _GEN_480; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_482 = 8'h2d == new_ptr_13_value ? ghv_45 : _GEN_481; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_483 = 8'h2e == new_ptr_13_value ? ghv_46 : _GEN_482; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_484 = 8'h2f == new_ptr_13_value ? ghv_47 : _GEN_483; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_485 = 8'h30 == new_ptr_13_value ? ghv_48 : _GEN_484; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_486 = 8'h31 == new_ptr_13_value ? ghv_49 : _GEN_485; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_487 = 8'h32 == new_ptr_13_value ? ghv_50 : _GEN_486; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_488 = 8'h33 == new_ptr_13_value ? ghv_51 : _GEN_487; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_489 = 8'h34 == new_ptr_13_value ? ghv_52 : _GEN_488; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_490 = 8'h35 == new_ptr_13_value ? ghv_53 : _GEN_489; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_491 = 8'h36 == new_ptr_13_value ? ghv_54 : _GEN_490; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_492 = 8'h37 == new_ptr_13_value ? ghv_55 : _GEN_491; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_493 = 8'h38 == new_ptr_13_value ? ghv_56 : _GEN_492; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_494 = 8'h39 == new_ptr_13_value ? ghv_57 : _GEN_493; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_495 = 8'h3a == new_ptr_13_value ? ghv_58 : _GEN_494; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_496 = 8'h3b == new_ptr_13_value ? ghv_59 : _GEN_495; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_497 = 8'h3c == new_ptr_13_value ? ghv_60 : _GEN_496; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_498 = 8'h3d == new_ptr_13_value ? ghv_61 : _GEN_497; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_499 = 8'h3e == new_ptr_13_value ? ghv_62 : _GEN_498; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_500 = 8'h3f == new_ptr_13_value ? ghv_63 : _GEN_499; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_501 = 8'h40 == new_ptr_13_value ? ghv_64 : _GEN_500; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_502 = 8'h41 == new_ptr_13_value ? ghv_65 : _GEN_501; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_503 = 8'h42 == new_ptr_13_value ? ghv_66 : _GEN_502; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_504 = 8'h43 == new_ptr_13_value ? ghv_67 : _GEN_503; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_505 = 8'h44 == new_ptr_13_value ? ghv_68 : _GEN_504; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_506 = 8'h45 == new_ptr_13_value ? ghv_69 : _GEN_505; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_507 = 8'h46 == new_ptr_13_value ? ghv_70 : _GEN_506; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_508 = 8'h47 == new_ptr_13_value ? ghv_71 : _GEN_507; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_509 = 8'h48 == new_ptr_13_value ? ghv_72 : _GEN_508; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_510 = 8'h49 == new_ptr_13_value ? ghv_73 : _GEN_509; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_511 = 8'h4a == new_ptr_13_value ? ghv_74 : _GEN_510; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_512 = 8'h4b == new_ptr_13_value ? ghv_75 : _GEN_511; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_513 = 8'h4c == new_ptr_13_value ? ghv_76 : _GEN_512; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_514 = 8'h4d == new_ptr_13_value ? ghv_77 : _GEN_513; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_515 = 8'h4e == new_ptr_13_value ? ghv_78 : _GEN_514; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_516 = 8'h4f == new_ptr_13_value ? ghv_79 : _GEN_515; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_517 = 8'h50 == new_ptr_13_value ? ghv_80 : _GEN_516; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_518 = 8'h51 == new_ptr_13_value ? ghv_81 : _GEN_517; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_519 = 8'h52 == new_ptr_13_value ? ghv_82 : _GEN_518; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_520 = 8'h53 == new_ptr_13_value ? ghv_83 : _GEN_519; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_521 = 8'h54 == new_ptr_13_value ? ghv_84 : _GEN_520; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_522 = 8'h55 == new_ptr_13_value ? ghv_85 : _GEN_521; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_523 = 8'h56 == new_ptr_13_value ? ghv_86 : _GEN_522; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_524 = 8'h57 == new_ptr_13_value ? ghv_87 : _GEN_523; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_525 = 8'h58 == new_ptr_13_value ? ghv_88 : _GEN_524; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_526 = 8'h59 == new_ptr_13_value ? ghv_89 : _GEN_525; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_527 = 8'h5a == new_ptr_13_value ? ghv_90 : _GEN_526; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_528 = 8'h5b == new_ptr_13_value ? ghv_91 : _GEN_527; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_529 = 8'h5c == new_ptr_13_value ? ghv_92 : _GEN_528; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_530 = 8'h5d == new_ptr_13_value ? ghv_93 : _GEN_529; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_531 = 8'h5e == new_ptr_13_value ? ghv_94 : _GEN_530; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_532 = 8'h5f == new_ptr_13_value ? ghv_95 : _GEN_531; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_533 = 8'h60 == new_ptr_13_value ? ghv_96 : _GEN_532; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_534 = 8'h61 == new_ptr_13_value ? ghv_97 : _GEN_533; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_535 = 8'h62 == new_ptr_13_value ? ghv_98 : _GEN_534; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_536 = 8'h63 == new_ptr_13_value ? ghv_99 : _GEN_535; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_537 = 8'h64 == new_ptr_13_value ? ghv_100 : _GEN_536; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_538 = 8'h65 == new_ptr_13_value ? ghv_101 : _GEN_537; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_539 = 8'h66 == new_ptr_13_value ? ghv_102 : _GEN_538; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_540 = 8'h67 == new_ptr_13_value ? ghv_103 : _GEN_539; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_541 = 8'h68 == new_ptr_13_value ? ghv_104 : _GEN_540; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_542 = 8'h69 == new_ptr_13_value ? ghv_105 : _GEN_541; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_543 = 8'h6a == new_ptr_13_value ? ghv_106 : _GEN_542; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_544 = 8'h6b == new_ptr_13_value ? ghv_107 : _GEN_543; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_545 = 8'h6c == new_ptr_13_value ? ghv_108 : _GEN_544; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_546 = 8'h6d == new_ptr_13_value ? ghv_109 : _GEN_545; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_547 = 8'h6e == new_ptr_13_value ? ghv_110 : _GEN_546; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_548 = 8'h6f == new_ptr_13_value ? ghv_111 : _GEN_547; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_549 = 8'h70 == new_ptr_13_value ? ghv_112 : _GEN_548; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_550 = 8'h71 == new_ptr_13_value ? ghv_113 : _GEN_549; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_551 = 8'h72 == new_ptr_13_value ? ghv_114 : _GEN_550; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_552 = 8'h73 == new_ptr_13_value ? ghv_115 : _GEN_551; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_553 = 8'h74 == new_ptr_13_value ? ghv_116 : _GEN_552; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_554 = 8'h75 == new_ptr_13_value ? ghv_117 : _GEN_553; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_555 = 8'h76 == new_ptr_13_value ? ghv_118 : _GEN_554; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_556 = 8'h77 == new_ptr_13_value ? ghv_119 : _GEN_555; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_557 = 8'h78 == new_ptr_13_value ? ghv_120 : _GEN_556; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_558 = 8'h79 == new_ptr_13_value ? ghv_121 : _GEN_557; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_559 = 8'h7a == new_ptr_13_value ? ghv_122 : _GEN_558; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_560 = 8'h7b == new_ptr_13_value ? ghv_123 : _GEN_559; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_561 = 8'h7c == new_ptr_13_value ? ghv_124 : _GEN_560; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_562 = 8'h7d == new_ptr_13_value ? ghv_125 : _GEN_561; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_563 = 8'h7e == new_ptr_13_value ? ghv_126 : _GEN_562; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_564 = 8'h7f == new_ptr_13_value ? ghv_127 : _GEN_563; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_565 = 8'h80 == new_ptr_13_value ? ghv_128 : _GEN_564; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_566 = 8'h81 == new_ptr_13_value ? ghv_129 : _GEN_565; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_567 = 8'h82 == new_ptr_13_value ? ghv_130 : _GEN_566; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_568 = 8'h83 == new_ptr_13_value ? ghv_131 : _GEN_567; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_569 = 8'h84 == new_ptr_13_value ? ghv_132 : _GEN_568; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_570 = 8'h85 == new_ptr_13_value ? ghv_133 : _GEN_569; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_571 = 8'h86 == new_ptr_13_value ? ghv_134 : _GEN_570; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_572 = 8'h87 == new_ptr_13_value ? ghv_135 : _GEN_571; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_573 = 8'h88 == new_ptr_13_value ? ghv_136 : _GEN_572; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_574 = 8'h89 == new_ptr_13_value ? ghv_137 : _GEN_573; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_575 = 8'h8a == new_ptr_13_value ? ghv_138 : _GEN_574; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_576 = 8'h8b == new_ptr_13_value ? ghv_139 : _GEN_575; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_577 = 8'h8c == new_ptr_13_value ? ghv_140 : _GEN_576; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_578 = 8'h8d == new_ptr_13_value ? ghv_141 : _GEN_577; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_579 = 8'h8e == new_ptr_13_value ? ghv_142 : _GEN_578; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_6_value = _new_ptr_value_T_13[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_582 = 8'h1 == new_ptr_6_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_583 = 8'h2 == new_ptr_6_value ? ghv_2 : _GEN_582; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_584 = 8'h3 == new_ptr_6_value ? ghv_3 : _GEN_583; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_585 = 8'h4 == new_ptr_6_value ? ghv_4 : _GEN_584; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_586 = 8'h5 == new_ptr_6_value ? ghv_5 : _GEN_585; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_587 = 8'h6 == new_ptr_6_value ? ghv_6 : _GEN_586; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_588 = 8'h7 == new_ptr_6_value ? ghv_7 : _GEN_587; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_589 = 8'h8 == new_ptr_6_value ? ghv_8 : _GEN_588; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_590 = 8'h9 == new_ptr_6_value ? ghv_9 : _GEN_589; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_591 = 8'ha == new_ptr_6_value ? ghv_10 : _GEN_590; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_592 = 8'hb == new_ptr_6_value ? ghv_11 : _GEN_591; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_593 = 8'hc == new_ptr_6_value ? ghv_12 : _GEN_592; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_594 = 8'hd == new_ptr_6_value ? ghv_13 : _GEN_593; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_595 = 8'he == new_ptr_6_value ? ghv_14 : _GEN_594; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_596 = 8'hf == new_ptr_6_value ? ghv_15 : _GEN_595; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_597 = 8'h10 == new_ptr_6_value ? ghv_16 : _GEN_596; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_598 = 8'h11 == new_ptr_6_value ? ghv_17 : _GEN_597; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_599 = 8'h12 == new_ptr_6_value ? ghv_18 : _GEN_598; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_600 = 8'h13 == new_ptr_6_value ? ghv_19 : _GEN_599; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_601 = 8'h14 == new_ptr_6_value ? ghv_20 : _GEN_600; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_602 = 8'h15 == new_ptr_6_value ? ghv_21 : _GEN_601; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_603 = 8'h16 == new_ptr_6_value ? ghv_22 : _GEN_602; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_604 = 8'h17 == new_ptr_6_value ? ghv_23 : _GEN_603; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_605 = 8'h18 == new_ptr_6_value ? ghv_24 : _GEN_604; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_606 = 8'h19 == new_ptr_6_value ? ghv_25 : _GEN_605; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_607 = 8'h1a == new_ptr_6_value ? ghv_26 : _GEN_606; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_608 = 8'h1b == new_ptr_6_value ? ghv_27 : _GEN_607; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_609 = 8'h1c == new_ptr_6_value ? ghv_28 : _GEN_608; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_610 = 8'h1d == new_ptr_6_value ? ghv_29 : _GEN_609; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_611 = 8'h1e == new_ptr_6_value ? ghv_30 : _GEN_610; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_612 = 8'h1f == new_ptr_6_value ? ghv_31 : _GEN_611; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_613 = 8'h20 == new_ptr_6_value ? ghv_32 : _GEN_612; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_614 = 8'h21 == new_ptr_6_value ? ghv_33 : _GEN_613; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_615 = 8'h22 == new_ptr_6_value ? ghv_34 : _GEN_614; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_616 = 8'h23 == new_ptr_6_value ? ghv_35 : _GEN_615; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_617 = 8'h24 == new_ptr_6_value ? ghv_36 : _GEN_616; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_618 = 8'h25 == new_ptr_6_value ? ghv_37 : _GEN_617; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_619 = 8'h26 == new_ptr_6_value ? ghv_38 : _GEN_618; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_620 = 8'h27 == new_ptr_6_value ? ghv_39 : _GEN_619; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_621 = 8'h28 == new_ptr_6_value ? ghv_40 : _GEN_620; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_622 = 8'h29 == new_ptr_6_value ? ghv_41 : _GEN_621; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_623 = 8'h2a == new_ptr_6_value ? ghv_42 : _GEN_622; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_624 = 8'h2b == new_ptr_6_value ? ghv_43 : _GEN_623; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_625 = 8'h2c == new_ptr_6_value ? ghv_44 : _GEN_624; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_626 = 8'h2d == new_ptr_6_value ? ghv_45 : _GEN_625; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_627 = 8'h2e == new_ptr_6_value ? ghv_46 : _GEN_626; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_628 = 8'h2f == new_ptr_6_value ? ghv_47 : _GEN_627; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_629 = 8'h30 == new_ptr_6_value ? ghv_48 : _GEN_628; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_630 = 8'h31 == new_ptr_6_value ? ghv_49 : _GEN_629; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_631 = 8'h32 == new_ptr_6_value ? ghv_50 : _GEN_630; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_632 = 8'h33 == new_ptr_6_value ? ghv_51 : _GEN_631; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_633 = 8'h34 == new_ptr_6_value ? ghv_52 : _GEN_632; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_634 = 8'h35 == new_ptr_6_value ? ghv_53 : _GEN_633; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_635 = 8'h36 == new_ptr_6_value ? ghv_54 : _GEN_634; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_636 = 8'h37 == new_ptr_6_value ? ghv_55 : _GEN_635; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_637 = 8'h38 == new_ptr_6_value ? ghv_56 : _GEN_636; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_638 = 8'h39 == new_ptr_6_value ? ghv_57 : _GEN_637; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_639 = 8'h3a == new_ptr_6_value ? ghv_58 : _GEN_638; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_640 = 8'h3b == new_ptr_6_value ? ghv_59 : _GEN_639; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_641 = 8'h3c == new_ptr_6_value ? ghv_60 : _GEN_640; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_642 = 8'h3d == new_ptr_6_value ? ghv_61 : _GEN_641; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_643 = 8'h3e == new_ptr_6_value ? ghv_62 : _GEN_642; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_644 = 8'h3f == new_ptr_6_value ? ghv_63 : _GEN_643; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_645 = 8'h40 == new_ptr_6_value ? ghv_64 : _GEN_644; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_646 = 8'h41 == new_ptr_6_value ? ghv_65 : _GEN_645; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_647 = 8'h42 == new_ptr_6_value ? ghv_66 : _GEN_646; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_648 = 8'h43 == new_ptr_6_value ? ghv_67 : _GEN_647; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_649 = 8'h44 == new_ptr_6_value ? ghv_68 : _GEN_648; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_650 = 8'h45 == new_ptr_6_value ? ghv_69 : _GEN_649; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_651 = 8'h46 == new_ptr_6_value ? ghv_70 : _GEN_650; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_652 = 8'h47 == new_ptr_6_value ? ghv_71 : _GEN_651; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_653 = 8'h48 == new_ptr_6_value ? ghv_72 : _GEN_652; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_654 = 8'h49 == new_ptr_6_value ? ghv_73 : _GEN_653; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_655 = 8'h4a == new_ptr_6_value ? ghv_74 : _GEN_654; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_656 = 8'h4b == new_ptr_6_value ? ghv_75 : _GEN_655; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_657 = 8'h4c == new_ptr_6_value ? ghv_76 : _GEN_656; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_658 = 8'h4d == new_ptr_6_value ? ghv_77 : _GEN_657; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_659 = 8'h4e == new_ptr_6_value ? ghv_78 : _GEN_658; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_660 = 8'h4f == new_ptr_6_value ? ghv_79 : _GEN_659; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_661 = 8'h50 == new_ptr_6_value ? ghv_80 : _GEN_660; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_662 = 8'h51 == new_ptr_6_value ? ghv_81 : _GEN_661; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_663 = 8'h52 == new_ptr_6_value ? ghv_82 : _GEN_662; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_664 = 8'h53 == new_ptr_6_value ? ghv_83 : _GEN_663; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_665 = 8'h54 == new_ptr_6_value ? ghv_84 : _GEN_664; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_666 = 8'h55 == new_ptr_6_value ? ghv_85 : _GEN_665; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_667 = 8'h56 == new_ptr_6_value ? ghv_86 : _GEN_666; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_668 = 8'h57 == new_ptr_6_value ? ghv_87 : _GEN_667; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_669 = 8'h58 == new_ptr_6_value ? ghv_88 : _GEN_668; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_670 = 8'h59 == new_ptr_6_value ? ghv_89 : _GEN_669; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_671 = 8'h5a == new_ptr_6_value ? ghv_90 : _GEN_670; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_672 = 8'h5b == new_ptr_6_value ? ghv_91 : _GEN_671; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_673 = 8'h5c == new_ptr_6_value ? ghv_92 : _GEN_672; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_674 = 8'h5d == new_ptr_6_value ? ghv_93 : _GEN_673; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_675 = 8'h5e == new_ptr_6_value ? ghv_94 : _GEN_674; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_676 = 8'h5f == new_ptr_6_value ? ghv_95 : _GEN_675; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_677 = 8'h60 == new_ptr_6_value ? ghv_96 : _GEN_676; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_678 = 8'h61 == new_ptr_6_value ? ghv_97 : _GEN_677; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_679 = 8'h62 == new_ptr_6_value ? ghv_98 : _GEN_678; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_680 = 8'h63 == new_ptr_6_value ? ghv_99 : _GEN_679; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_681 = 8'h64 == new_ptr_6_value ? ghv_100 : _GEN_680; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_682 = 8'h65 == new_ptr_6_value ? ghv_101 : _GEN_681; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_683 = 8'h66 == new_ptr_6_value ? ghv_102 : _GEN_682; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_684 = 8'h67 == new_ptr_6_value ? ghv_103 : _GEN_683; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_685 = 8'h68 == new_ptr_6_value ? ghv_104 : _GEN_684; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_686 = 8'h69 == new_ptr_6_value ? ghv_105 : _GEN_685; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_687 = 8'h6a == new_ptr_6_value ? ghv_106 : _GEN_686; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_688 = 8'h6b == new_ptr_6_value ? ghv_107 : _GEN_687; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_689 = 8'h6c == new_ptr_6_value ? ghv_108 : _GEN_688; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_690 = 8'h6d == new_ptr_6_value ? ghv_109 : _GEN_689; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_691 = 8'h6e == new_ptr_6_value ? ghv_110 : _GEN_690; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_692 = 8'h6f == new_ptr_6_value ? ghv_111 : _GEN_691; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_693 = 8'h70 == new_ptr_6_value ? ghv_112 : _GEN_692; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_694 = 8'h71 == new_ptr_6_value ? ghv_113 : _GEN_693; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_695 = 8'h72 == new_ptr_6_value ? ghv_114 : _GEN_694; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_696 = 8'h73 == new_ptr_6_value ? ghv_115 : _GEN_695; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_697 = 8'h74 == new_ptr_6_value ? ghv_116 : _GEN_696; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_698 = 8'h75 == new_ptr_6_value ? ghv_117 : _GEN_697; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_699 = 8'h76 == new_ptr_6_value ? ghv_118 : _GEN_698; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_700 = 8'h77 == new_ptr_6_value ? ghv_119 : _GEN_699; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_701 = 8'h78 == new_ptr_6_value ? ghv_120 : _GEN_700; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_702 = 8'h79 == new_ptr_6_value ? ghv_121 : _GEN_701; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_703 = 8'h7a == new_ptr_6_value ? ghv_122 : _GEN_702; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_704 = 8'h7b == new_ptr_6_value ? ghv_123 : _GEN_703; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_705 = 8'h7c == new_ptr_6_value ? ghv_124 : _GEN_704; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_706 = 8'h7d == new_ptr_6_value ? ghv_125 : _GEN_705; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_707 = 8'h7e == new_ptr_6_value ? ghv_126 : _GEN_706; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_708 = 8'h7f == new_ptr_6_value ? ghv_127 : _GEN_707; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_709 = 8'h80 == new_ptr_6_value ? ghv_128 : _GEN_708; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_710 = 8'h81 == new_ptr_6_value ? ghv_129 : _GEN_709; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_711 = 8'h82 == new_ptr_6_value ? ghv_130 : _GEN_710; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_712 = 8'h83 == new_ptr_6_value ? ghv_131 : _GEN_711; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_713 = 8'h84 == new_ptr_6_value ? ghv_132 : _GEN_712; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_714 = 8'h85 == new_ptr_6_value ? ghv_133 : _GEN_713; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_715 = 8'h86 == new_ptr_6_value ? ghv_134 : _GEN_714; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_716 = 8'h87 == new_ptr_6_value ? ghv_135 : _GEN_715; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_717 = 8'h88 == new_ptr_6_value ? ghv_136 : _GEN_716; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_718 = 8'h89 == new_ptr_6_value ? ghv_137 : _GEN_717; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_719 = 8'h8a == new_ptr_6_value ? ghv_138 : _GEN_718; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_720 = 8'h8b == new_ptr_6_value ? ghv_139 : _GEN_719; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_721 = 8'h8c == new_ptr_6_value ? ghv_140 : _GEN_720; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_722 = 8'h8d == new_ptr_6_value ? ghv_141 : _GEN_721; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_723 = 8'h8e == new_ptr_6_value ? ghv_142 : _GEN_722; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_12_value = _new_ptr_value_T_25[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_726 = 8'h1 == new_ptr_12_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_727 = 8'h2 == new_ptr_12_value ? ghv_2 : _GEN_726; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_728 = 8'h3 == new_ptr_12_value ? ghv_3 : _GEN_727; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_729 = 8'h4 == new_ptr_12_value ? ghv_4 : _GEN_728; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_730 = 8'h5 == new_ptr_12_value ? ghv_5 : _GEN_729; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_731 = 8'h6 == new_ptr_12_value ? ghv_6 : _GEN_730; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_732 = 8'h7 == new_ptr_12_value ? ghv_7 : _GEN_731; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_733 = 8'h8 == new_ptr_12_value ? ghv_8 : _GEN_732; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_734 = 8'h9 == new_ptr_12_value ? ghv_9 : _GEN_733; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_735 = 8'ha == new_ptr_12_value ? ghv_10 : _GEN_734; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_736 = 8'hb == new_ptr_12_value ? ghv_11 : _GEN_735; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_737 = 8'hc == new_ptr_12_value ? ghv_12 : _GEN_736; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_738 = 8'hd == new_ptr_12_value ? ghv_13 : _GEN_737; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_739 = 8'he == new_ptr_12_value ? ghv_14 : _GEN_738; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_740 = 8'hf == new_ptr_12_value ? ghv_15 : _GEN_739; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_741 = 8'h10 == new_ptr_12_value ? ghv_16 : _GEN_740; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_742 = 8'h11 == new_ptr_12_value ? ghv_17 : _GEN_741; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_743 = 8'h12 == new_ptr_12_value ? ghv_18 : _GEN_742; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_744 = 8'h13 == new_ptr_12_value ? ghv_19 : _GEN_743; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_745 = 8'h14 == new_ptr_12_value ? ghv_20 : _GEN_744; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_746 = 8'h15 == new_ptr_12_value ? ghv_21 : _GEN_745; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_747 = 8'h16 == new_ptr_12_value ? ghv_22 : _GEN_746; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_748 = 8'h17 == new_ptr_12_value ? ghv_23 : _GEN_747; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_749 = 8'h18 == new_ptr_12_value ? ghv_24 : _GEN_748; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_750 = 8'h19 == new_ptr_12_value ? ghv_25 : _GEN_749; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_751 = 8'h1a == new_ptr_12_value ? ghv_26 : _GEN_750; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_752 = 8'h1b == new_ptr_12_value ? ghv_27 : _GEN_751; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_753 = 8'h1c == new_ptr_12_value ? ghv_28 : _GEN_752; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_754 = 8'h1d == new_ptr_12_value ? ghv_29 : _GEN_753; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_755 = 8'h1e == new_ptr_12_value ? ghv_30 : _GEN_754; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_756 = 8'h1f == new_ptr_12_value ? ghv_31 : _GEN_755; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_757 = 8'h20 == new_ptr_12_value ? ghv_32 : _GEN_756; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_758 = 8'h21 == new_ptr_12_value ? ghv_33 : _GEN_757; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_759 = 8'h22 == new_ptr_12_value ? ghv_34 : _GEN_758; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_760 = 8'h23 == new_ptr_12_value ? ghv_35 : _GEN_759; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_761 = 8'h24 == new_ptr_12_value ? ghv_36 : _GEN_760; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_762 = 8'h25 == new_ptr_12_value ? ghv_37 : _GEN_761; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_763 = 8'h26 == new_ptr_12_value ? ghv_38 : _GEN_762; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_764 = 8'h27 == new_ptr_12_value ? ghv_39 : _GEN_763; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_765 = 8'h28 == new_ptr_12_value ? ghv_40 : _GEN_764; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_766 = 8'h29 == new_ptr_12_value ? ghv_41 : _GEN_765; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_767 = 8'h2a == new_ptr_12_value ? ghv_42 : _GEN_766; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_768 = 8'h2b == new_ptr_12_value ? ghv_43 : _GEN_767; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_769 = 8'h2c == new_ptr_12_value ? ghv_44 : _GEN_768; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_770 = 8'h2d == new_ptr_12_value ? ghv_45 : _GEN_769; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_771 = 8'h2e == new_ptr_12_value ? ghv_46 : _GEN_770; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_772 = 8'h2f == new_ptr_12_value ? ghv_47 : _GEN_771; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_773 = 8'h30 == new_ptr_12_value ? ghv_48 : _GEN_772; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_774 = 8'h31 == new_ptr_12_value ? ghv_49 : _GEN_773; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_775 = 8'h32 == new_ptr_12_value ? ghv_50 : _GEN_774; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_776 = 8'h33 == new_ptr_12_value ? ghv_51 : _GEN_775; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_777 = 8'h34 == new_ptr_12_value ? ghv_52 : _GEN_776; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_778 = 8'h35 == new_ptr_12_value ? ghv_53 : _GEN_777; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_779 = 8'h36 == new_ptr_12_value ? ghv_54 : _GEN_778; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_780 = 8'h37 == new_ptr_12_value ? ghv_55 : _GEN_779; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_781 = 8'h38 == new_ptr_12_value ? ghv_56 : _GEN_780; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_782 = 8'h39 == new_ptr_12_value ? ghv_57 : _GEN_781; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_783 = 8'h3a == new_ptr_12_value ? ghv_58 : _GEN_782; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_784 = 8'h3b == new_ptr_12_value ? ghv_59 : _GEN_783; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_785 = 8'h3c == new_ptr_12_value ? ghv_60 : _GEN_784; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_786 = 8'h3d == new_ptr_12_value ? ghv_61 : _GEN_785; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_787 = 8'h3e == new_ptr_12_value ? ghv_62 : _GEN_786; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_788 = 8'h3f == new_ptr_12_value ? ghv_63 : _GEN_787; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_789 = 8'h40 == new_ptr_12_value ? ghv_64 : _GEN_788; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_790 = 8'h41 == new_ptr_12_value ? ghv_65 : _GEN_789; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_791 = 8'h42 == new_ptr_12_value ? ghv_66 : _GEN_790; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_792 = 8'h43 == new_ptr_12_value ? ghv_67 : _GEN_791; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_793 = 8'h44 == new_ptr_12_value ? ghv_68 : _GEN_792; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_794 = 8'h45 == new_ptr_12_value ? ghv_69 : _GEN_793; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_795 = 8'h46 == new_ptr_12_value ? ghv_70 : _GEN_794; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_796 = 8'h47 == new_ptr_12_value ? ghv_71 : _GEN_795; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_797 = 8'h48 == new_ptr_12_value ? ghv_72 : _GEN_796; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_798 = 8'h49 == new_ptr_12_value ? ghv_73 : _GEN_797; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_799 = 8'h4a == new_ptr_12_value ? ghv_74 : _GEN_798; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_800 = 8'h4b == new_ptr_12_value ? ghv_75 : _GEN_799; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_801 = 8'h4c == new_ptr_12_value ? ghv_76 : _GEN_800; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_802 = 8'h4d == new_ptr_12_value ? ghv_77 : _GEN_801; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_803 = 8'h4e == new_ptr_12_value ? ghv_78 : _GEN_802; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_804 = 8'h4f == new_ptr_12_value ? ghv_79 : _GEN_803; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_805 = 8'h50 == new_ptr_12_value ? ghv_80 : _GEN_804; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_806 = 8'h51 == new_ptr_12_value ? ghv_81 : _GEN_805; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_807 = 8'h52 == new_ptr_12_value ? ghv_82 : _GEN_806; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_808 = 8'h53 == new_ptr_12_value ? ghv_83 : _GEN_807; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_809 = 8'h54 == new_ptr_12_value ? ghv_84 : _GEN_808; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_810 = 8'h55 == new_ptr_12_value ? ghv_85 : _GEN_809; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_811 = 8'h56 == new_ptr_12_value ? ghv_86 : _GEN_810; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_812 = 8'h57 == new_ptr_12_value ? ghv_87 : _GEN_811; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_813 = 8'h58 == new_ptr_12_value ? ghv_88 : _GEN_812; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_814 = 8'h59 == new_ptr_12_value ? ghv_89 : _GEN_813; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_815 = 8'h5a == new_ptr_12_value ? ghv_90 : _GEN_814; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_816 = 8'h5b == new_ptr_12_value ? ghv_91 : _GEN_815; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_817 = 8'h5c == new_ptr_12_value ? ghv_92 : _GEN_816; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_818 = 8'h5d == new_ptr_12_value ? ghv_93 : _GEN_817; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_819 = 8'h5e == new_ptr_12_value ? ghv_94 : _GEN_818; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_820 = 8'h5f == new_ptr_12_value ? ghv_95 : _GEN_819; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_821 = 8'h60 == new_ptr_12_value ? ghv_96 : _GEN_820; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_822 = 8'h61 == new_ptr_12_value ? ghv_97 : _GEN_821; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_823 = 8'h62 == new_ptr_12_value ? ghv_98 : _GEN_822; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_824 = 8'h63 == new_ptr_12_value ? ghv_99 : _GEN_823; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_825 = 8'h64 == new_ptr_12_value ? ghv_100 : _GEN_824; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_826 = 8'h65 == new_ptr_12_value ? ghv_101 : _GEN_825; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_827 = 8'h66 == new_ptr_12_value ? ghv_102 : _GEN_826; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_828 = 8'h67 == new_ptr_12_value ? ghv_103 : _GEN_827; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_829 = 8'h68 == new_ptr_12_value ? ghv_104 : _GEN_828; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_830 = 8'h69 == new_ptr_12_value ? ghv_105 : _GEN_829; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_831 = 8'h6a == new_ptr_12_value ? ghv_106 : _GEN_830; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_832 = 8'h6b == new_ptr_12_value ? ghv_107 : _GEN_831; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_833 = 8'h6c == new_ptr_12_value ? ghv_108 : _GEN_832; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_834 = 8'h6d == new_ptr_12_value ? ghv_109 : _GEN_833; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_835 = 8'h6e == new_ptr_12_value ? ghv_110 : _GEN_834; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_836 = 8'h6f == new_ptr_12_value ? ghv_111 : _GEN_835; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_837 = 8'h70 == new_ptr_12_value ? ghv_112 : _GEN_836; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_838 = 8'h71 == new_ptr_12_value ? ghv_113 : _GEN_837; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_839 = 8'h72 == new_ptr_12_value ? ghv_114 : _GEN_838; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_840 = 8'h73 == new_ptr_12_value ? ghv_115 : _GEN_839; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_841 = 8'h74 == new_ptr_12_value ? ghv_116 : _GEN_840; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_842 = 8'h75 == new_ptr_12_value ? ghv_117 : _GEN_841; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_843 = 8'h76 == new_ptr_12_value ? ghv_118 : _GEN_842; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_844 = 8'h77 == new_ptr_12_value ? ghv_119 : _GEN_843; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_845 = 8'h78 == new_ptr_12_value ? ghv_120 : _GEN_844; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_846 = 8'h79 == new_ptr_12_value ? ghv_121 : _GEN_845; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_847 = 8'h7a == new_ptr_12_value ? ghv_122 : _GEN_846; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_848 = 8'h7b == new_ptr_12_value ? ghv_123 : _GEN_847; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_849 = 8'h7c == new_ptr_12_value ? ghv_124 : _GEN_848; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_850 = 8'h7d == new_ptr_12_value ? ghv_125 : _GEN_849; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_851 = 8'h7e == new_ptr_12_value ? ghv_126 : _GEN_850; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_852 = 8'h7f == new_ptr_12_value ? ghv_127 : _GEN_851; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_853 = 8'h80 == new_ptr_12_value ? ghv_128 : _GEN_852; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_854 = 8'h81 == new_ptr_12_value ? ghv_129 : _GEN_853; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_855 = 8'h82 == new_ptr_12_value ? ghv_130 : _GEN_854; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_856 = 8'h83 == new_ptr_12_value ? ghv_131 : _GEN_855; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_857 = 8'h84 == new_ptr_12_value ? ghv_132 : _GEN_856; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_858 = 8'h85 == new_ptr_12_value ? ghv_133 : _GEN_857; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_859 = 8'h86 == new_ptr_12_value ? ghv_134 : _GEN_858; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_860 = 8'h87 == new_ptr_12_value ? ghv_135 : _GEN_859; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_861 = 8'h88 == new_ptr_12_value ? ghv_136 : _GEN_860; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_862 = 8'h89 == new_ptr_12_value ? ghv_137 : _GEN_861; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_863 = 8'h8a == new_ptr_12_value ? ghv_138 : _GEN_862; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_864 = 8'h8b == new_ptr_12_value ? ghv_139 : _GEN_863; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_865 = 8'h8c == new_ptr_12_value ? ghv_140 : _GEN_864; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_866 = 8'h8d == new_ptr_12_value ? ghv_141 : _GEN_865; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_867 = 8'h8e == new_ptr_12_value ? ghv_142 : _GEN_866; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_15_value = _new_ptr_value_T_31[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_870 = 8'h1 == new_ptr_15_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_871 = 8'h2 == new_ptr_15_value ? ghv_2 : _GEN_870; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_872 = 8'h3 == new_ptr_15_value ? ghv_3 : _GEN_871; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_873 = 8'h4 == new_ptr_15_value ? ghv_4 : _GEN_872; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_874 = 8'h5 == new_ptr_15_value ? ghv_5 : _GEN_873; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_875 = 8'h6 == new_ptr_15_value ? ghv_6 : _GEN_874; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_876 = 8'h7 == new_ptr_15_value ? ghv_7 : _GEN_875; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_877 = 8'h8 == new_ptr_15_value ? ghv_8 : _GEN_876; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_878 = 8'h9 == new_ptr_15_value ? ghv_9 : _GEN_877; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_879 = 8'ha == new_ptr_15_value ? ghv_10 : _GEN_878; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_880 = 8'hb == new_ptr_15_value ? ghv_11 : _GEN_879; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_881 = 8'hc == new_ptr_15_value ? ghv_12 : _GEN_880; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_882 = 8'hd == new_ptr_15_value ? ghv_13 : _GEN_881; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_883 = 8'he == new_ptr_15_value ? ghv_14 : _GEN_882; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_884 = 8'hf == new_ptr_15_value ? ghv_15 : _GEN_883; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_885 = 8'h10 == new_ptr_15_value ? ghv_16 : _GEN_884; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_886 = 8'h11 == new_ptr_15_value ? ghv_17 : _GEN_885; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_887 = 8'h12 == new_ptr_15_value ? ghv_18 : _GEN_886; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_888 = 8'h13 == new_ptr_15_value ? ghv_19 : _GEN_887; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_889 = 8'h14 == new_ptr_15_value ? ghv_20 : _GEN_888; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_890 = 8'h15 == new_ptr_15_value ? ghv_21 : _GEN_889; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_891 = 8'h16 == new_ptr_15_value ? ghv_22 : _GEN_890; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_892 = 8'h17 == new_ptr_15_value ? ghv_23 : _GEN_891; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_893 = 8'h18 == new_ptr_15_value ? ghv_24 : _GEN_892; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_894 = 8'h19 == new_ptr_15_value ? ghv_25 : _GEN_893; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_895 = 8'h1a == new_ptr_15_value ? ghv_26 : _GEN_894; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_896 = 8'h1b == new_ptr_15_value ? ghv_27 : _GEN_895; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_897 = 8'h1c == new_ptr_15_value ? ghv_28 : _GEN_896; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_898 = 8'h1d == new_ptr_15_value ? ghv_29 : _GEN_897; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_899 = 8'h1e == new_ptr_15_value ? ghv_30 : _GEN_898; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_900 = 8'h1f == new_ptr_15_value ? ghv_31 : _GEN_899; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_901 = 8'h20 == new_ptr_15_value ? ghv_32 : _GEN_900; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_902 = 8'h21 == new_ptr_15_value ? ghv_33 : _GEN_901; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_903 = 8'h22 == new_ptr_15_value ? ghv_34 : _GEN_902; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_904 = 8'h23 == new_ptr_15_value ? ghv_35 : _GEN_903; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_905 = 8'h24 == new_ptr_15_value ? ghv_36 : _GEN_904; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_906 = 8'h25 == new_ptr_15_value ? ghv_37 : _GEN_905; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_907 = 8'h26 == new_ptr_15_value ? ghv_38 : _GEN_906; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_908 = 8'h27 == new_ptr_15_value ? ghv_39 : _GEN_907; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_909 = 8'h28 == new_ptr_15_value ? ghv_40 : _GEN_908; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_910 = 8'h29 == new_ptr_15_value ? ghv_41 : _GEN_909; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_911 = 8'h2a == new_ptr_15_value ? ghv_42 : _GEN_910; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_912 = 8'h2b == new_ptr_15_value ? ghv_43 : _GEN_911; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_913 = 8'h2c == new_ptr_15_value ? ghv_44 : _GEN_912; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_914 = 8'h2d == new_ptr_15_value ? ghv_45 : _GEN_913; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_915 = 8'h2e == new_ptr_15_value ? ghv_46 : _GEN_914; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_916 = 8'h2f == new_ptr_15_value ? ghv_47 : _GEN_915; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_917 = 8'h30 == new_ptr_15_value ? ghv_48 : _GEN_916; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_918 = 8'h31 == new_ptr_15_value ? ghv_49 : _GEN_917; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_919 = 8'h32 == new_ptr_15_value ? ghv_50 : _GEN_918; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_920 = 8'h33 == new_ptr_15_value ? ghv_51 : _GEN_919; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_921 = 8'h34 == new_ptr_15_value ? ghv_52 : _GEN_920; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_922 = 8'h35 == new_ptr_15_value ? ghv_53 : _GEN_921; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_923 = 8'h36 == new_ptr_15_value ? ghv_54 : _GEN_922; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_924 = 8'h37 == new_ptr_15_value ? ghv_55 : _GEN_923; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_925 = 8'h38 == new_ptr_15_value ? ghv_56 : _GEN_924; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_926 = 8'h39 == new_ptr_15_value ? ghv_57 : _GEN_925; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_927 = 8'h3a == new_ptr_15_value ? ghv_58 : _GEN_926; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_928 = 8'h3b == new_ptr_15_value ? ghv_59 : _GEN_927; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_929 = 8'h3c == new_ptr_15_value ? ghv_60 : _GEN_928; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_930 = 8'h3d == new_ptr_15_value ? ghv_61 : _GEN_929; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_931 = 8'h3e == new_ptr_15_value ? ghv_62 : _GEN_930; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_932 = 8'h3f == new_ptr_15_value ? ghv_63 : _GEN_931; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_933 = 8'h40 == new_ptr_15_value ? ghv_64 : _GEN_932; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_934 = 8'h41 == new_ptr_15_value ? ghv_65 : _GEN_933; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_935 = 8'h42 == new_ptr_15_value ? ghv_66 : _GEN_934; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_936 = 8'h43 == new_ptr_15_value ? ghv_67 : _GEN_935; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_937 = 8'h44 == new_ptr_15_value ? ghv_68 : _GEN_936; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_938 = 8'h45 == new_ptr_15_value ? ghv_69 : _GEN_937; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_939 = 8'h46 == new_ptr_15_value ? ghv_70 : _GEN_938; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_940 = 8'h47 == new_ptr_15_value ? ghv_71 : _GEN_939; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_941 = 8'h48 == new_ptr_15_value ? ghv_72 : _GEN_940; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_942 = 8'h49 == new_ptr_15_value ? ghv_73 : _GEN_941; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_943 = 8'h4a == new_ptr_15_value ? ghv_74 : _GEN_942; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_944 = 8'h4b == new_ptr_15_value ? ghv_75 : _GEN_943; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_945 = 8'h4c == new_ptr_15_value ? ghv_76 : _GEN_944; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_946 = 8'h4d == new_ptr_15_value ? ghv_77 : _GEN_945; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_947 = 8'h4e == new_ptr_15_value ? ghv_78 : _GEN_946; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_948 = 8'h4f == new_ptr_15_value ? ghv_79 : _GEN_947; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_949 = 8'h50 == new_ptr_15_value ? ghv_80 : _GEN_948; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_950 = 8'h51 == new_ptr_15_value ? ghv_81 : _GEN_949; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_951 = 8'h52 == new_ptr_15_value ? ghv_82 : _GEN_950; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_952 = 8'h53 == new_ptr_15_value ? ghv_83 : _GEN_951; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_953 = 8'h54 == new_ptr_15_value ? ghv_84 : _GEN_952; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_954 = 8'h55 == new_ptr_15_value ? ghv_85 : _GEN_953; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_955 = 8'h56 == new_ptr_15_value ? ghv_86 : _GEN_954; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_956 = 8'h57 == new_ptr_15_value ? ghv_87 : _GEN_955; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_957 = 8'h58 == new_ptr_15_value ? ghv_88 : _GEN_956; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_958 = 8'h59 == new_ptr_15_value ? ghv_89 : _GEN_957; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_959 = 8'h5a == new_ptr_15_value ? ghv_90 : _GEN_958; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_960 = 8'h5b == new_ptr_15_value ? ghv_91 : _GEN_959; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_961 = 8'h5c == new_ptr_15_value ? ghv_92 : _GEN_960; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_962 = 8'h5d == new_ptr_15_value ? ghv_93 : _GEN_961; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_963 = 8'h5e == new_ptr_15_value ? ghv_94 : _GEN_962; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_964 = 8'h5f == new_ptr_15_value ? ghv_95 : _GEN_963; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_965 = 8'h60 == new_ptr_15_value ? ghv_96 : _GEN_964; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_966 = 8'h61 == new_ptr_15_value ? ghv_97 : _GEN_965; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_967 = 8'h62 == new_ptr_15_value ? ghv_98 : _GEN_966; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_968 = 8'h63 == new_ptr_15_value ? ghv_99 : _GEN_967; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_969 = 8'h64 == new_ptr_15_value ? ghv_100 : _GEN_968; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_970 = 8'h65 == new_ptr_15_value ? ghv_101 : _GEN_969; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_971 = 8'h66 == new_ptr_15_value ? ghv_102 : _GEN_970; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_972 = 8'h67 == new_ptr_15_value ? ghv_103 : _GEN_971; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_973 = 8'h68 == new_ptr_15_value ? ghv_104 : _GEN_972; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_974 = 8'h69 == new_ptr_15_value ? ghv_105 : _GEN_973; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_975 = 8'h6a == new_ptr_15_value ? ghv_106 : _GEN_974; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_976 = 8'h6b == new_ptr_15_value ? ghv_107 : _GEN_975; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_977 = 8'h6c == new_ptr_15_value ? ghv_108 : _GEN_976; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_978 = 8'h6d == new_ptr_15_value ? ghv_109 : _GEN_977; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_979 = 8'h6e == new_ptr_15_value ? ghv_110 : _GEN_978; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_980 = 8'h6f == new_ptr_15_value ? ghv_111 : _GEN_979; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_981 = 8'h70 == new_ptr_15_value ? ghv_112 : _GEN_980; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_982 = 8'h71 == new_ptr_15_value ? ghv_113 : _GEN_981; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_983 = 8'h72 == new_ptr_15_value ? ghv_114 : _GEN_982; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_984 = 8'h73 == new_ptr_15_value ? ghv_115 : _GEN_983; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_985 = 8'h74 == new_ptr_15_value ? ghv_116 : _GEN_984; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_986 = 8'h75 == new_ptr_15_value ? ghv_117 : _GEN_985; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_987 = 8'h76 == new_ptr_15_value ? ghv_118 : _GEN_986; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_988 = 8'h77 == new_ptr_15_value ? ghv_119 : _GEN_987; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_989 = 8'h78 == new_ptr_15_value ? ghv_120 : _GEN_988; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_990 = 8'h79 == new_ptr_15_value ? ghv_121 : _GEN_989; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_991 = 8'h7a == new_ptr_15_value ? ghv_122 : _GEN_990; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_992 = 8'h7b == new_ptr_15_value ? ghv_123 : _GEN_991; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_993 = 8'h7c == new_ptr_15_value ? ghv_124 : _GEN_992; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_994 = 8'h7d == new_ptr_15_value ? ghv_125 : _GEN_993; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_995 = 8'h7e == new_ptr_15_value ? ghv_126 : _GEN_994; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_996 = 8'h7f == new_ptr_15_value ? ghv_127 : _GEN_995; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_997 = 8'h80 == new_ptr_15_value ? ghv_128 : _GEN_996; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_998 = 8'h81 == new_ptr_15_value ? ghv_129 : _GEN_997; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_999 = 8'h82 == new_ptr_15_value ? ghv_130 : _GEN_998; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1000 = 8'h83 == new_ptr_15_value ? ghv_131 : _GEN_999; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1001 = 8'h84 == new_ptr_15_value ? ghv_132 : _GEN_1000; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1002 = 8'h85 == new_ptr_15_value ? ghv_133 : _GEN_1001; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1003 = 8'h86 == new_ptr_15_value ? ghv_134 : _GEN_1002; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1004 = 8'h87 == new_ptr_15_value ? ghv_135 : _GEN_1003; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1005 = 8'h88 == new_ptr_15_value ? ghv_136 : _GEN_1004; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1006 = 8'h89 == new_ptr_15_value ? ghv_137 : _GEN_1005; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1007 = 8'h8a == new_ptr_15_value ? ghv_138 : _GEN_1006; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1008 = 8'h8b == new_ptr_15_value ? ghv_139 : _GEN_1007; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1009 = 8'h8c == new_ptr_15_value ? ghv_140 : _GEN_1008; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1010 = 8'h8d == new_ptr_15_value ? ghv_141 : _GEN_1009; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1011 = 8'h8e == new_ptr_15_value ? ghv_142 : _GEN_1010; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_2_value = _new_ptr_value_T_5[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_1014 = 8'h1 == new_ptr_2_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1015 = 8'h2 == new_ptr_2_value ? ghv_2 : _GEN_1014; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1016 = 8'h3 == new_ptr_2_value ? ghv_3 : _GEN_1015; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1017 = 8'h4 == new_ptr_2_value ? ghv_4 : _GEN_1016; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1018 = 8'h5 == new_ptr_2_value ? ghv_5 : _GEN_1017; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1019 = 8'h6 == new_ptr_2_value ? ghv_6 : _GEN_1018; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1020 = 8'h7 == new_ptr_2_value ? ghv_7 : _GEN_1019; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1021 = 8'h8 == new_ptr_2_value ? ghv_8 : _GEN_1020; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1022 = 8'h9 == new_ptr_2_value ? ghv_9 : _GEN_1021; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1023 = 8'ha == new_ptr_2_value ? ghv_10 : _GEN_1022; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1024 = 8'hb == new_ptr_2_value ? ghv_11 : _GEN_1023; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1025 = 8'hc == new_ptr_2_value ? ghv_12 : _GEN_1024; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1026 = 8'hd == new_ptr_2_value ? ghv_13 : _GEN_1025; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1027 = 8'he == new_ptr_2_value ? ghv_14 : _GEN_1026; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1028 = 8'hf == new_ptr_2_value ? ghv_15 : _GEN_1027; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1029 = 8'h10 == new_ptr_2_value ? ghv_16 : _GEN_1028; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1030 = 8'h11 == new_ptr_2_value ? ghv_17 : _GEN_1029; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1031 = 8'h12 == new_ptr_2_value ? ghv_18 : _GEN_1030; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1032 = 8'h13 == new_ptr_2_value ? ghv_19 : _GEN_1031; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1033 = 8'h14 == new_ptr_2_value ? ghv_20 : _GEN_1032; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1034 = 8'h15 == new_ptr_2_value ? ghv_21 : _GEN_1033; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1035 = 8'h16 == new_ptr_2_value ? ghv_22 : _GEN_1034; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1036 = 8'h17 == new_ptr_2_value ? ghv_23 : _GEN_1035; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1037 = 8'h18 == new_ptr_2_value ? ghv_24 : _GEN_1036; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1038 = 8'h19 == new_ptr_2_value ? ghv_25 : _GEN_1037; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1039 = 8'h1a == new_ptr_2_value ? ghv_26 : _GEN_1038; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1040 = 8'h1b == new_ptr_2_value ? ghv_27 : _GEN_1039; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1041 = 8'h1c == new_ptr_2_value ? ghv_28 : _GEN_1040; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1042 = 8'h1d == new_ptr_2_value ? ghv_29 : _GEN_1041; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1043 = 8'h1e == new_ptr_2_value ? ghv_30 : _GEN_1042; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1044 = 8'h1f == new_ptr_2_value ? ghv_31 : _GEN_1043; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1045 = 8'h20 == new_ptr_2_value ? ghv_32 : _GEN_1044; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1046 = 8'h21 == new_ptr_2_value ? ghv_33 : _GEN_1045; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1047 = 8'h22 == new_ptr_2_value ? ghv_34 : _GEN_1046; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1048 = 8'h23 == new_ptr_2_value ? ghv_35 : _GEN_1047; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1049 = 8'h24 == new_ptr_2_value ? ghv_36 : _GEN_1048; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1050 = 8'h25 == new_ptr_2_value ? ghv_37 : _GEN_1049; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1051 = 8'h26 == new_ptr_2_value ? ghv_38 : _GEN_1050; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1052 = 8'h27 == new_ptr_2_value ? ghv_39 : _GEN_1051; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1053 = 8'h28 == new_ptr_2_value ? ghv_40 : _GEN_1052; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1054 = 8'h29 == new_ptr_2_value ? ghv_41 : _GEN_1053; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1055 = 8'h2a == new_ptr_2_value ? ghv_42 : _GEN_1054; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1056 = 8'h2b == new_ptr_2_value ? ghv_43 : _GEN_1055; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1057 = 8'h2c == new_ptr_2_value ? ghv_44 : _GEN_1056; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1058 = 8'h2d == new_ptr_2_value ? ghv_45 : _GEN_1057; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1059 = 8'h2e == new_ptr_2_value ? ghv_46 : _GEN_1058; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1060 = 8'h2f == new_ptr_2_value ? ghv_47 : _GEN_1059; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1061 = 8'h30 == new_ptr_2_value ? ghv_48 : _GEN_1060; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1062 = 8'h31 == new_ptr_2_value ? ghv_49 : _GEN_1061; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1063 = 8'h32 == new_ptr_2_value ? ghv_50 : _GEN_1062; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1064 = 8'h33 == new_ptr_2_value ? ghv_51 : _GEN_1063; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1065 = 8'h34 == new_ptr_2_value ? ghv_52 : _GEN_1064; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1066 = 8'h35 == new_ptr_2_value ? ghv_53 : _GEN_1065; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1067 = 8'h36 == new_ptr_2_value ? ghv_54 : _GEN_1066; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1068 = 8'h37 == new_ptr_2_value ? ghv_55 : _GEN_1067; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1069 = 8'h38 == new_ptr_2_value ? ghv_56 : _GEN_1068; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1070 = 8'h39 == new_ptr_2_value ? ghv_57 : _GEN_1069; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1071 = 8'h3a == new_ptr_2_value ? ghv_58 : _GEN_1070; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1072 = 8'h3b == new_ptr_2_value ? ghv_59 : _GEN_1071; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1073 = 8'h3c == new_ptr_2_value ? ghv_60 : _GEN_1072; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1074 = 8'h3d == new_ptr_2_value ? ghv_61 : _GEN_1073; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1075 = 8'h3e == new_ptr_2_value ? ghv_62 : _GEN_1074; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1076 = 8'h3f == new_ptr_2_value ? ghv_63 : _GEN_1075; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1077 = 8'h40 == new_ptr_2_value ? ghv_64 : _GEN_1076; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1078 = 8'h41 == new_ptr_2_value ? ghv_65 : _GEN_1077; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1079 = 8'h42 == new_ptr_2_value ? ghv_66 : _GEN_1078; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1080 = 8'h43 == new_ptr_2_value ? ghv_67 : _GEN_1079; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1081 = 8'h44 == new_ptr_2_value ? ghv_68 : _GEN_1080; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1082 = 8'h45 == new_ptr_2_value ? ghv_69 : _GEN_1081; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1083 = 8'h46 == new_ptr_2_value ? ghv_70 : _GEN_1082; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1084 = 8'h47 == new_ptr_2_value ? ghv_71 : _GEN_1083; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1085 = 8'h48 == new_ptr_2_value ? ghv_72 : _GEN_1084; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1086 = 8'h49 == new_ptr_2_value ? ghv_73 : _GEN_1085; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1087 = 8'h4a == new_ptr_2_value ? ghv_74 : _GEN_1086; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1088 = 8'h4b == new_ptr_2_value ? ghv_75 : _GEN_1087; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1089 = 8'h4c == new_ptr_2_value ? ghv_76 : _GEN_1088; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1090 = 8'h4d == new_ptr_2_value ? ghv_77 : _GEN_1089; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1091 = 8'h4e == new_ptr_2_value ? ghv_78 : _GEN_1090; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1092 = 8'h4f == new_ptr_2_value ? ghv_79 : _GEN_1091; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1093 = 8'h50 == new_ptr_2_value ? ghv_80 : _GEN_1092; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1094 = 8'h51 == new_ptr_2_value ? ghv_81 : _GEN_1093; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1095 = 8'h52 == new_ptr_2_value ? ghv_82 : _GEN_1094; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1096 = 8'h53 == new_ptr_2_value ? ghv_83 : _GEN_1095; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1097 = 8'h54 == new_ptr_2_value ? ghv_84 : _GEN_1096; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1098 = 8'h55 == new_ptr_2_value ? ghv_85 : _GEN_1097; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1099 = 8'h56 == new_ptr_2_value ? ghv_86 : _GEN_1098; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1100 = 8'h57 == new_ptr_2_value ? ghv_87 : _GEN_1099; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1101 = 8'h58 == new_ptr_2_value ? ghv_88 : _GEN_1100; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1102 = 8'h59 == new_ptr_2_value ? ghv_89 : _GEN_1101; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1103 = 8'h5a == new_ptr_2_value ? ghv_90 : _GEN_1102; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1104 = 8'h5b == new_ptr_2_value ? ghv_91 : _GEN_1103; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1105 = 8'h5c == new_ptr_2_value ? ghv_92 : _GEN_1104; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1106 = 8'h5d == new_ptr_2_value ? ghv_93 : _GEN_1105; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1107 = 8'h5e == new_ptr_2_value ? ghv_94 : _GEN_1106; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1108 = 8'h5f == new_ptr_2_value ? ghv_95 : _GEN_1107; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1109 = 8'h60 == new_ptr_2_value ? ghv_96 : _GEN_1108; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1110 = 8'h61 == new_ptr_2_value ? ghv_97 : _GEN_1109; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1111 = 8'h62 == new_ptr_2_value ? ghv_98 : _GEN_1110; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1112 = 8'h63 == new_ptr_2_value ? ghv_99 : _GEN_1111; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1113 = 8'h64 == new_ptr_2_value ? ghv_100 : _GEN_1112; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1114 = 8'h65 == new_ptr_2_value ? ghv_101 : _GEN_1113; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1115 = 8'h66 == new_ptr_2_value ? ghv_102 : _GEN_1114; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1116 = 8'h67 == new_ptr_2_value ? ghv_103 : _GEN_1115; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1117 = 8'h68 == new_ptr_2_value ? ghv_104 : _GEN_1116; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1118 = 8'h69 == new_ptr_2_value ? ghv_105 : _GEN_1117; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1119 = 8'h6a == new_ptr_2_value ? ghv_106 : _GEN_1118; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1120 = 8'h6b == new_ptr_2_value ? ghv_107 : _GEN_1119; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1121 = 8'h6c == new_ptr_2_value ? ghv_108 : _GEN_1120; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1122 = 8'h6d == new_ptr_2_value ? ghv_109 : _GEN_1121; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1123 = 8'h6e == new_ptr_2_value ? ghv_110 : _GEN_1122; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1124 = 8'h6f == new_ptr_2_value ? ghv_111 : _GEN_1123; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1125 = 8'h70 == new_ptr_2_value ? ghv_112 : _GEN_1124; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1126 = 8'h71 == new_ptr_2_value ? ghv_113 : _GEN_1125; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1127 = 8'h72 == new_ptr_2_value ? ghv_114 : _GEN_1126; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1128 = 8'h73 == new_ptr_2_value ? ghv_115 : _GEN_1127; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1129 = 8'h74 == new_ptr_2_value ? ghv_116 : _GEN_1128; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1130 = 8'h75 == new_ptr_2_value ? ghv_117 : _GEN_1129; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1131 = 8'h76 == new_ptr_2_value ? ghv_118 : _GEN_1130; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1132 = 8'h77 == new_ptr_2_value ? ghv_119 : _GEN_1131; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1133 = 8'h78 == new_ptr_2_value ? ghv_120 : _GEN_1132; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1134 = 8'h79 == new_ptr_2_value ? ghv_121 : _GEN_1133; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1135 = 8'h7a == new_ptr_2_value ? ghv_122 : _GEN_1134; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1136 = 8'h7b == new_ptr_2_value ? ghv_123 : _GEN_1135; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1137 = 8'h7c == new_ptr_2_value ? ghv_124 : _GEN_1136; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1138 = 8'h7d == new_ptr_2_value ? ghv_125 : _GEN_1137; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1139 = 8'h7e == new_ptr_2_value ? ghv_126 : _GEN_1138; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1140 = 8'h7f == new_ptr_2_value ? ghv_127 : _GEN_1139; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1141 = 8'h80 == new_ptr_2_value ? ghv_128 : _GEN_1140; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1142 = 8'h81 == new_ptr_2_value ? ghv_129 : _GEN_1141; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1143 = 8'h82 == new_ptr_2_value ? ghv_130 : _GEN_1142; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1144 = 8'h83 == new_ptr_2_value ? ghv_131 : _GEN_1143; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1145 = 8'h84 == new_ptr_2_value ? ghv_132 : _GEN_1144; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1146 = 8'h85 == new_ptr_2_value ? ghv_133 : _GEN_1145; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1147 = 8'h86 == new_ptr_2_value ? ghv_134 : _GEN_1146; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1148 = 8'h87 == new_ptr_2_value ? ghv_135 : _GEN_1147; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1149 = 8'h88 == new_ptr_2_value ? ghv_136 : _GEN_1148; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1150 = 8'h89 == new_ptr_2_value ? ghv_137 : _GEN_1149; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1151 = 8'h8a == new_ptr_2_value ? ghv_138 : _GEN_1150; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1152 = 8'h8b == new_ptr_2_value ? ghv_139 : _GEN_1151; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1153 = 8'h8c == new_ptr_2_value ? ghv_140 : _GEN_1152; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1154 = 8'h8d == new_ptr_2_value ? ghv_141 : _GEN_1153; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1155 = 8'h8e == new_ptr_2_value ? ghv_142 : _GEN_1154; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_14_value = _new_ptr_value_T_29[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_1158 = 8'h1 == new_ptr_14_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1159 = 8'h2 == new_ptr_14_value ? ghv_2 : _GEN_1158; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1160 = 8'h3 == new_ptr_14_value ? ghv_3 : _GEN_1159; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1161 = 8'h4 == new_ptr_14_value ? ghv_4 : _GEN_1160; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1162 = 8'h5 == new_ptr_14_value ? ghv_5 : _GEN_1161; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1163 = 8'h6 == new_ptr_14_value ? ghv_6 : _GEN_1162; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1164 = 8'h7 == new_ptr_14_value ? ghv_7 : _GEN_1163; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1165 = 8'h8 == new_ptr_14_value ? ghv_8 : _GEN_1164; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1166 = 8'h9 == new_ptr_14_value ? ghv_9 : _GEN_1165; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1167 = 8'ha == new_ptr_14_value ? ghv_10 : _GEN_1166; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1168 = 8'hb == new_ptr_14_value ? ghv_11 : _GEN_1167; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1169 = 8'hc == new_ptr_14_value ? ghv_12 : _GEN_1168; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1170 = 8'hd == new_ptr_14_value ? ghv_13 : _GEN_1169; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1171 = 8'he == new_ptr_14_value ? ghv_14 : _GEN_1170; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1172 = 8'hf == new_ptr_14_value ? ghv_15 : _GEN_1171; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1173 = 8'h10 == new_ptr_14_value ? ghv_16 : _GEN_1172; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1174 = 8'h11 == new_ptr_14_value ? ghv_17 : _GEN_1173; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1175 = 8'h12 == new_ptr_14_value ? ghv_18 : _GEN_1174; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1176 = 8'h13 == new_ptr_14_value ? ghv_19 : _GEN_1175; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1177 = 8'h14 == new_ptr_14_value ? ghv_20 : _GEN_1176; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1178 = 8'h15 == new_ptr_14_value ? ghv_21 : _GEN_1177; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1179 = 8'h16 == new_ptr_14_value ? ghv_22 : _GEN_1178; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1180 = 8'h17 == new_ptr_14_value ? ghv_23 : _GEN_1179; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1181 = 8'h18 == new_ptr_14_value ? ghv_24 : _GEN_1180; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1182 = 8'h19 == new_ptr_14_value ? ghv_25 : _GEN_1181; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1183 = 8'h1a == new_ptr_14_value ? ghv_26 : _GEN_1182; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1184 = 8'h1b == new_ptr_14_value ? ghv_27 : _GEN_1183; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1185 = 8'h1c == new_ptr_14_value ? ghv_28 : _GEN_1184; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1186 = 8'h1d == new_ptr_14_value ? ghv_29 : _GEN_1185; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1187 = 8'h1e == new_ptr_14_value ? ghv_30 : _GEN_1186; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1188 = 8'h1f == new_ptr_14_value ? ghv_31 : _GEN_1187; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1189 = 8'h20 == new_ptr_14_value ? ghv_32 : _GEN_1188; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1190 = 8'h21 == new_ptr_14_value ? ghv_33 : _GEN_1189; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1191 = 8'h22 == new_ptr_14_value ? ghv_34 : _GEN_1190; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1192 = 8'h23 == new_ptr_14_value ? ghv_35 : _GEN_1191; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1193 = 8'h24 == new_ptr_14_value ? ghv_36 : _GEN_1192; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1194 = 8'h25 == new_ptr_14_value ? ghv_37 : _GEN_1193; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1195 = 8'h26 == new_ptr_14_value ? ghv_38 : _GEN_1194; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1196 = 8'h27 == new_ptr_14_value ? ghv_39 : _GEN_1195; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1197 = 8'h28 == new_ptr_14_value ? ghv_40 : _GEN_1196; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1198 = 8'h29 == new_ptr_14_value ? ghv_41 : _GEN_1197; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1199 = 8'h2a == new_ptr_14_value ? ghv_42 : _GEN_1198; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1200 = 8'h2b == new_ptr_14_value ? ghv_43 : _GEN_1199; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1201 = 8'h2c == new_ptr_14_value ? ghv_44 : _GEN_1200; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1202 = 8'h2d == new_ptr_14_value ? ghv_45 : _GEN_1201; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1203 = 8'h2e == new_ptr_14_value ? ghv_46 : _GEN_1202; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1204 = 8'h2f == new_ptr_14_value ? ghv_47 : _GEN_1203; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1205 = 8'h30 == new_ptr_14_value ? ghv_48 : _GEN_1204; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1206 = 8'h31 == new_ptr_14_value ? ghv_49 : _GEN_1205; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1207 = 8'h32 == new_ptr_14_value ? ghv_50 : _GEN_1206; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1208 = 8'h33 == new_ptr_14_value ? ghv_51 : _GEN_1207; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1209 = 8'h34 == new_ptr_14_value ? ghv_52 : _GEN_1208; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1210 = 8'h35 == new_ptr_14_value ? ghv_53 : _GEN_1209; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1211 = 8'h36 == new_ptr_14_value ? ghv_54 : _GEN_1210; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1212 = 8'h37 == new_ptr_14_value ? ghv_55 : _GEN_1211; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1213 = 8'h38 == new_ptr_14_value ? ghv_56 : _GEN_1212; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1214 = 8'h39 == new_ptr_14_value ? ghv_57 : _GEN_1213; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1215 = 8'h3a == new_ptr_14_value ? ghv_58 : _GEN_1214; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1216 = 8'h3b == new_ptr_14_value ? ghv_59 : _GEN_1215; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1217 = 8'h3c == new_ptr_14_value ? ghv_60 : _GEN_1216; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1218 = 8'h3d == new_ptr_14_value ? ghv_61 : _GEN_1217; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1219 = 8'h3e == new_ptr_14_value ? ghv_62 : _GEN_1218; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1220 = 8'h3f == new_ptr_14_value ? ghv_63 : _GEN_1219; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1221 = 8'h40 == new_ptr_14_value ? ghv_64 : _GEN_1220; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1222 = 8'h41 == new_ptr_14_value ? ghv_65 : _GEN_1221; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1223 = 8'h42 == new_ptr_14_value ? ghv_66 : _GEN_1222; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1224 = 8'h43 == new_ptr_14_value ? ghv_67 : _GEN_1223; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1225 = 8'h44 == new_ptr_14_value ? ghv_68 : _GEN_1224; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1226 = 8'h45 == new_ptr_14_value ? ghv_69 : _GEN_1225; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1227 = 8'h46 == new_ptr_14_value ? ghv_70 : _GEN_1226; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1228 = 8'h47 == new_ptr_14_value ? ghv_71 : _GEN_1227; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1229 = 8'h48 == new_ptr_14_value ? ghv_72 : _GEN_1228; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1230 = 8'h49 == new_ptr_14_value ? ghv_73 : _GEN_1229; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1231 = 8'h4a == new_ptr_14_value ? ghv_74 : _GEN_1230; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1232 = 8'h4b == new_ptr_14_value ? ghv_75 : _GEN_1231; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1233 = 8'h4c == new_ptr_14_value ? ghv_76 : _GEN_1232; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1234 = 8'h4d == new_ptr_14_value ? ghv_77 : _GEN_1233; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1235 = 8'h4e == new_ptr_14_value ? ghv_78 : _GEN_1234; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1236 = 8'h4f == new_ptr_14_value ? ghv_79 : _GEN_1235; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1237 = 8'h50 == new_ptr_14_value ? ghv_80 : _GEN_1236; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1238 = 8'h51 == new_ptr_14_value ? ghv_81 : _GEN_1237; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1239 = 8'h52 == new_ptr_14_value ? ghv_82 : _GEN_1238; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1240 = 8'h53 == new_ptr_14_value ? ghv_83 : _GEN_1239; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1241 = 8'h54 == new_ptr_14_value ? ghv_84 : _GEN_1240; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1242 = 8'h55 == new_ptr_14_value ? ghv_85 : _GEN_1241; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1243 = 8'h56 == new_ptr_14_value ? ghv_86 : _GEN_1242; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1244 = 8'h57 == new_ptr_14_value ? ghv_87 : _GEN_1243; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1245 = 8'h58 == new_ptr_14_value ? ghv_88 : _GEN_1244; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1246 = 8'h59 == new_ptr_14_value ? ghv_89 : _GEN_1245; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1247 = 8'h5a == new_ptr_14_value ? ghv_90 : _GEN_1246; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1248 = 8'h5b == new_ptr_14_value ? ghv_91 : _GEN_1247; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1249 = 8'h5c == new_ptr_14_value ? ghv_92 : _GEN_1248; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1250 = 8'h5d == new_ptr_14_value ? ghv_93 : _GEN_1249; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1251 = 8'h5e == new_ptr_14_value ? ghv_94 : _GEN_1250; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1252 = 8'h5f == new_ptr_14_value ? ghv_95 : _GEN_1251; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1253 = 8'h60 == new_ptr_14_value ? ghv_96 : _GEN_1252; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1254 = 8'h61 == new_ptr_14_value ? ghv_97 : _GEN_1253; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1255 = 8'h62 == new_ptr_14_value ? ghv_98 : _GEN_1254; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1256 = 8'h63 == new_ptr_14_value ? ghv_99 : _GEN_1255; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1257 = 8'h64 == new_ptr_14_value ? ghv_100 : _GEN_1256; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1258 = 8'h65 == new_ptr_14_value ? ghv_101 : _GEN_1257; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1259 = 8'h66 == new_ptr_14_value ? ghv_102 : _GEN_1258; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1260 = 8'h67 == new_ptr_14_value ? ghv_103 : _GEN_1259; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1261 = 8'h68 == new_ptr_14_value ? ghv_104 : _GEN_1260; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1262 = 8'h69 == new_ptr_14_value ? ghv_105 : _GEN_1261; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1263 = 8'h6a == new_ptr_14_value ? ghv_106 : _GEN_1262; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1264 = 8'h6b == new_ptr_14_value ? ghv_107 : _GEN_1263; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1265 = 8'h6c == new_ptr_14_value ? ghv_108 : _GEN_1264; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1266 = 8'h6d == new_ptr_14_value ? ghv_109 : _GEN_1265; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1267 = 8'h6e == new_ptr_14_value ? ghv_110 : _GEN_1266; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1268 = 8'h6f == new_ptr_14_value ? ghv_111 : _GEN_1267; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1269 = 8'h70 == new_ptr_14_value ? ghv_112 : _GEN_1268; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1270 = 8'h71 == new_ptr_14_value ? ghv_113 : _GEN_1269; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1271 = 8'h72 == new_ptr_14_value ? ghv_114 : _GEN_1270; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1272 = 8'h73 == new_ptr_14_value ? ghv_115 : _GEN_1271; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1273 = 8'h74 == new_ptr_14_value ? ghv_116 : _GEN_1272; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1274 = 8'h75 == new_ptr_14_value ? ghv_117 : _GEN_1273; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1275 = 8'h76 == new_ptr_14_value ? ghv_118 : _GEN_1274; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1276 = 8'h77 == new_ptr_14_value ? ghv_119 : _GEN_1275; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1277 = 8'h78 == new_ptr_14_value ? ghv_120 : _GEN_1276; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1278 = 8'h79 == new_ptr_14_value ? ghv_121 : _GEN_1277; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1279 = 8'h7a == new_ptr_14_value ? ghv_122 : _GEN_1278; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1280 = 8'h7b == new_ptr_14_value ? ghv_123 : _GEN_1279; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1281 = 8'h7c == new_ptr_14_value ? ghv_124 : _GEN_1280; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1282 = 8'h7d == new_ptr_14_value ? ghv_125 : _GEN_1281; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1283 = 8'h7e == new_ptr_14_value ? ghv_126 : _GEN_1282; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1284 = 8'h7f == new_ptr_14_value ? ghv_127 : _GEN_1283; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1285 = 8'h80 == new_ptr_14_value ? ghv_128 : _GEN_1284; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1286 = 8'h81 == new_ptr_14_value ? ghv_129 : _GEN_1285; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1287 = 8'h82 == new_ptr_14_value ? ghv_130 : _GEN_1286; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1288 = 8'h83 == new_ptr_14_value ? ghv_131 : _GEN_1287; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1289 = 8'h84 == new_ptr_14_value ? ghv_132 : _GEN_1288; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1290 = 8'h85 == new_ptr_14_value ? ghv_133 : _GEN_1289; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1291 = 8'h86 == new_ptr_14_value ? ghv_134 : _GEN_1290; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1292 = 8'h87 == new_ptr_14_value ? ghv_135 : _GEN_1291; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1293 = 8'h88 == new_ptr_14_value ? ghv_136 : _GEN_1292; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1294 = 8'h89 == new_ptr_14_value ? ghv_137 : _GEN_1293; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1295 = 8'h8a == new_ptr_14_value ? ghv_138 : _GEN_1294; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1296 = 8'h8b == new_ptr_14_value ? ghv_139 : _GEN_1295; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1297 = 8'h8c == new_ptr_14_value ? ghv_140 : _GEN_1296; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1298 = 8'h8d == new_ptr_14_value ? ghv_141 : _GEN_1297; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1299 = 8'h8e == new_ptr_14_value ? ghv_142 : _GEN_1298; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_17_value = _new_ptr_value_T_35[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_1302 = 8'h1 == new_ptr_17_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1303 = 8'h2 == new_ptr_17_value ? ghv_2 : _GEN_1302; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1304 = 8'h3 == new_ptr_17_value ? ghv_3 : _GEN_1303; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1305 = 8'h4 == new_ptr_17_value ? ghv_4 : _GEN_1304; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1306 = 8'h5 == new_ptr_17_value ? ghv_5 : _GEN_1305; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1307 = 8'h6 == new_ptr_17_value ? ghv_6 : _GEN_1306; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1308 = 8'h7 == new_ptr_17_value ? ghv_7 : _GEN_1307; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1309 = 8'h8 == new_ptr_17_value ? ghv_8 : _GEN_1308; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1310 = 8'h9 == new_ptr_17_value ? ghv_9 : _GEN_1309; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1311 = 8'ha == new_ptr_17_value ? ghv_10 : _GEN_1310; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1312 = 8'hb == new_ptr_17_value ? ghv_11 : _GEN_1311; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1313 = 8'hc == new_ptr_17_value ? ghv_12 : _GEN_1312; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1314 = 8'hd == new_ptr_17_value ? ghv_13 : _GEN_1313; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1315 = 8'he == new_ptr_17_value ? ghv_14 : _GEN_1314; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1316 = 8'hf == new_ptr_17_value ? ghv_15 : _GEN_1315; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1317 = 8'h10 == new_ptr_17_value ? ghv_16 : _GEN_1316; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1318 = 8'h11 == new_ptr_17_value ? ghv_17 : _GEN_1317; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1319 = 8'h12 == new_ptr_17_value ? ghv_18 : _GEN_1318; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1320 = 8'h13 == new_ptr_17_value ? ghv_19 : _GEN_1319; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1321 = 8'h14 == new_ptr_17_value ? ghv_20 : _GEN_1320; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1322 = 8'h15 == new_ptr_17_value ? ghv_21 : _GEN_1321; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1323 = 8'h16 == new_ptr_17_value ? ghv_22 : _GEN_1322; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1324 = 8'h17 == new_ptr_17_value ? ghv_23 : _GEN_1323; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1325 = 8'h18 == new_ptr_17_value ? ghv_24 : _GEN_1324; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1326 = 8'h19 == new_ptr_17_value ? ghv_25 : _GEN_1325; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1327 = 8'h1a == new_ptr_17_value ? ghv_26 : _GEN_1326; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1328 = 8'h1b == new_ptr_17_value ? ghv_27 : _GEN_1327; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1329 = 8'h1c == new_ptr_17_value ? ghv_28 : _GEN_1328; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1330 = 8'h1d == new_ptr_17_value ? ghv_29 : _GEN_1329; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1331 = 8'h1e == new_ptr_17_value ? ghv_30 : _GEN_1330; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1332 = 8'h1f == new_ptr_17_value ? ghv_31 : _GEN_1331; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1333 = 8'h20 == new_ptr_17_value ? ghv_32 : _GEN_1332; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1334 = 8'h21 == new_ptr_17_value ? ghv_33 : _GEN_1333; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1335 = 8'h22 == new_ptr_17_value ? ghv_34 : _GEN_1334; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1336 = 8'h23 == new_ptr_17_value ? ghv_35 : _GEN_1335; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1337 = 8'h24 == new_ptr_17_value ? ghv_36 : _GEN_1336; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1338 = 8'h25 == new_ptr_17_value ? ghv_37 : _GEN_1337; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1339 = 8'h26 == new_ptr_17_value ? ghv_38 : _GEN_1338; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1340 = 8'h27 == new_ptr_17_value ? ghv_39 : _GEN_1339; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1341 = 8'h28 == new_ptr_17_value ? ghv_40 : _GEN_1340; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1342 = 8'h29 == new_ptr_17_value ? ghv_41 : _GEN_1341; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1343 = 8'h2a == new_ptr_17_value ? ghv_42 : _GEN_1342; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1344 = 8'h2b == new_ptr_17_value ? ghv_43 : _GEN_1343; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1345 = 8'h2c == new_ptr_17_value ? ghv_44 : _GEN_1344; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1346 = 8'h2d == new_ptr_17_value ? ghv_45 : _GEN_1345; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1347 = 8'h2e == new_ptr_17_value ? ghv_46 : _GEN_1346; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1348 = 8'h2f == new_ptr_17_value ? ghv_47 : _GEN_1347; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1349 = 8'h30 == new_ptr_17_value ? ghv_48 : _GEN_1348; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1350 = 8'h31 == new_ptr_17_value ? ghv_49 : _GEN_1349; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1351 = 8'h32 == new_ptr_17_value ? ghv_50 : _GEN_1350; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1352 = 8'h33 == new_ptr_17_value ? ghv_51 : _GEN_1351; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1353 = 8'h34 == new_ptr_17_value ? ghv_52 : _GEN_1352; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1354 = 8'h35 == new_ptr_17_value ? ghv_53 : _GEN_1353; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1355 = 8'h36 == new_ptr_17_value ? ghv_54 : _GEN_1354; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1356 = 8'h37 == new_ptr_17_value ? ghv_55 : _GEN_1355; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1357 = 8'h38 == new_ptr_17_value ? ghv_56 : _GEN_1356; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1358 = 8'h39 == new_ptr_17_value ? ghv_57 : _GEN_1357; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1359 = 8'h3a == new_ptr_17_value ? ghv_58 : _GEN_1358; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1360 = 8'h3b == new_ptr_17_value ? ghv_59 : _GEN_1359; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1361 = 8'h3c == new_ptr_17_value ? ghv_60 : _GEN_1360; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1362 = 8'h3d == new_ptr_17_value ? ghv_61 : _GEN_1361; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1363 = 8'h3e == new_ptr_17_value ? ghv_62 : _GEN_1362; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1364 = 8'h3f == new_ptr_17_value ? ghv_63 : _GEN_1363; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1365 = 8'h40 == new_ptr_17_value ? ghv_64 : _GEN_1364; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1366 = 8'h41 == new_ptr_17_value ? ghv_65 : _GEN_1365; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1367 = 8'h42 == new_ptr_17_value ? ghv_66 : _GEN_1366; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1368 = 8'h43 == new_ptr_17_value ? ghv_67 : _GEN_1367; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1369 = 8'h44 == new_ptr_17_value ? ghv_68 : _GEN_1368; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1370 = 8'h45 == new_ptr_17_value ? ghv_69 : _GEN_1369; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1371 = 8'h46 == new_ptr_17_value ? ghv_70 : _GEN_1370; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1372 = 8'h47 == new_ptr_17_value ? ghv_71 : _GEN_1371; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1373 = 8'h48 == new_ptr_17_value ? ghv_72 : _GEN_1372; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1374 = 8'h49 == new_ptr_17_value ? ghv_73 : _GEN_1373; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1375 = 8'h4a == new_ptr_17_value ? ghv_74 : _GEN_1374; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1376 = 8'h4b == new_ptr_17_value ? ghv_75 : _GEN_1375; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1377 = 8'h4c == new_ptr_17_value ? ghv_76 : _GEN_1376; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1378 = 8'h4d == new_ptr_17_value ? ghv_77 : _GEN_1377; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1379 = 8'h4e == new_ptr_17_value ? ghv_78 : _GEN_1378; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1380 = 8'h4f == new_ptr_17_value ? ghv_79 : _GEN_1379; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1381 = 8'h50 == new_ptr_17_value ? ghv_80 : _GEN_1380; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1382 = 8'h51 == new_ptr_17_value ? ghv_81 : _GEN_1381; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1383 = 8'h52 == new_ptr_17_value ? ghv_82 : _GEN_1382; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1384 = 8'h53 == new_ptr_17_value ? ghv_83 : _GEN_1383; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1385 = 8'h54 == new_ptr_17_value ? ghv_84 : _GEN_1384; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1386 = 8'h55 == new_ptr_17_value ? ghv_85 : _GEN_1385; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1387 = 8'h56 == new_ptr_17_value ? ghv_86 : _GEN_1386; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1388 = 8'h57 == new_ptr_17_value ? ghv_87 : _GEN_1387; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1389 = 8'h58 == new_ptr_17_value ? ghv_88 : _GEN_1388; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1390 = 8'h59 == new_ptr_17_value ? ghv_89 : _GEN_1389; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1391 = 8'h5a == new_ptr_17_value ? ghv_90 : _GEN_1390; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1392 = 8'h5b == new_ptr_17_value ? ghv_91 : _GEN_1391; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1393 = 8'h5c == new_ptr_17_value ? ghv_92 : _GEN_1392; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1394 = 8'h5d == new_ptr_17_value ? ghv_93 : _GEN_1393; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1395 = 8'h5e == new_ptr_17_value ? ghv_94 : _GEN_1394; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1396 = 8'h5f == new_ptr_17_value ? ghv_95 : _GEN_1395; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1397 = 8'h60 == new_ptr_17_value ? ghv_96 : _GEN_1396; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1398 = 8'h61 == new_ptr_17_value ? ghv_97 : _GEN_1397; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1399 = 8'h62 == new_ptr_17_value ? ghv_98 : _GEN_1398; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1400 = 8'h63 == new_ptr_17_value ? ghv_99 : _GEN_1399; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1401 = 8'h64 == new_ptr_17_value ? ghv_100 : _GEN_1400; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1402 = 8'h65 == new_ptr_17_value ? ghv_101 : _GEN_1401; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1403 = 8'h66 == new_ptr_17_value ? ghv_102 : _GEN_1402; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1404 = 8'h67 == new_ptr_17_value ? ghv_103 : _GEN_1403; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1405 = 8'h68 == new_ptr_17_value ? ghv_104 : _GEN_1404; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1406 = 8'h69 == new_ptr_17_value ? ghv_105 : _GEN_1405; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1407 = 8'h6a == new_ptr_17_value ? ghv_106 : _GEN_1406; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1408 = 8'h6b == new_ptr_17_value ? ghv_107 : _GEN_1407; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1409 = 8'h6c == new_ptr_17_value ? ghv_108 : _GEN_1408; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1410 = 8'h6d == new_ptr_17_value ? ghv_109 : _GEN_1409; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1411 = 8'h6e == new_ptr_17_value ? ghv_110 : _GEN_1410; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1412 = 8'h6f == new_ptr_17_value ? ghv_111 : _GEN_1411; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1413 = 8'h70 == new_ptr_17_value ? ghv_112 : _GEN_1412; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1414 = 8'h71 == new_ptr_17_value ? ghv_113 : _GEN_1413; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1415 = 8'h72 == new_ptr_17_value ? ghv_114 : _GEN_1414; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1416 = 8'h73 == new_ptr_17_value ? ghv_115 : _GEN_1415; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1417 = 8'h74 == new_ptr_17_value ? ghv_116 : _GEN_1416; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1418 = 8'h75 == new_ptr_17_value ? ghv_117 : _GEN_1417; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1419 = 8'h76 == new_ptr_17_value ? ghv_118 : _GEN_1418; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1420 = 8'h77 == new_ptr_17_value ? ghv_119 : _GEN_1419; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1421 = 8'h78 == new_ptr_17_value ? ghv_120 : _GEN_1420; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1422 = 8'h79 == new_ptr_17_value ? ghv_121 : _GEN_1421; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1423 = 8'h7a == new_ptr_17_value ? ghv_122 : _GEN_1422; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1424 = 8'h7b == new_ptr_17_value ? ghv_123 : _GEN_1423; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1425 = 8'h7c == new_ptr_17_value ? ghv_124 : _GEN_1424; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1426 = 8'h7d == new_ptr_17_value ? ghv_125 : _GEN_1425; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1427 = 8'h7e == new_ptr_17_value ? ghv_126 : _GEN_1426; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1428 = 8'h7f == new_ptr_17_value ? ghv_127 : _GEN_1427; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1429 = 8'h80 == new_ptr_17_value ? ghv_128 : _GEN_1428; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1430 = 8'h81 == new_ptr_17_value ? ghv_129 : _GEN_1429; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1431 = 8'h82 == new_ptr_17_value ? ghv_130 : _GEN_1430; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1432 = 8'h83 == new_ptr_17_value ? ghv_131 : _GEN_1431; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1433 = 8'h84 == new_ptr_17_value ? ghv_132 : _GEN_1432; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1434 = 8'h85 == new_ptr_17_value ? ghv_133 : _GEN_1433; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1435 = 8'h86 == new_ptr_17_value ? ghv_134 : _GEN_1434; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1436 = 8'h87 == new_ptr_17_value ? ghv_135 : _GEN_1435; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1437 = 8'h88 == new_ptr_17_value ? ghv_136 : _GEN_1436; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1438 = 8'h89 == new_ptr_17_value ? ghv_137 : _GEN_1437; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1439 = 8'h8a == new_ptr_17_value ? ghv_138 : _GEN_1438; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1440 = 8'h8b == new_ptr_17_value ? ghv_139 : _GEN_1439; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1441 = 8'h8c == new_ptr_17_value ? ghv_140 : _GEN_1440; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1442 = 8'h8d == new_ptr_17_value ? ghv_141 : _GEN_1441; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1443 = 8'h8e == new_ptr_17_value ? ghv_142 : _GEN_1442; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_4_value = _new_ptr_value_T_9[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_1446 = 8'h1 == new_ptr_4_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1447 = 8'h2 == new_ptr_4_value ? ghv_2 : _GEN_1446; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1448 = 8'h3 == new_ptr_4_value ? ghv_3 : _GEN_1447; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1449 = 8'h4 == new_ptr_4_value ? ghv_4 : _GEN_1448; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1450 = 8'h5 == new_ptr_4_value ? ghv_5 : _GEN_1449; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1451 = 8'h6 == new_ptr_4_value ? ghv_6 : _GEN_1450; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1452 = 8'h7 == new_ptr_4_value ? ghv_7 : _GEN_1451; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1453 = 8'h8 == new_ptr_4_value ? ghv_8 : _GEN_1452; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1454 = 8'h9 == new_ptr_4_value ? ghv_9 : _GEN_1453; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1455 = 8'ha == new_ptr_4_value ? ghv_10 : _GEN_1454; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1456 = 8'hb == new_ptr_4_value ? ghv_11 : _GEN_1455; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1457 = 8'hc == new_ptr_4_value ? ghv_12 : _GEN_1456; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1458 = 8'hd == new_ptr_4_value ? ghv_13 : _GEN_1457; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1459 = 8'he == new_ptr_4_value ? ghv_14 : _GEN_1458; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1460 = 8'hf == new_ptr_4_value ? ghv_15 : _GEN_1459; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1461 = 8'h10 == new_ptr_4_value ? ghv_16 : _GEN_1460; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1462 = 8'h11 == new_ptr_4_value ? ghv_17 : _GEN_1461; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1463 = 8'h12 == new_ptr_4_value ? ghv_18 : _GEN_1462; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1464 = 8'h13 == new_ptr_4_value ? ghv_19 : _GEN_1463; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1465 = 8'h14 == new_ptr_4_value ? ghv_20 : _GEN_1464; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1466 = 8'h15 == new_ptr_4_value ? ghv_21 : _GEN_1465; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1467 = 8'h16 == new_ptr_4_value ? ghv_22 : _GEN_1466; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1468 = 8'h17 == new_ptr_4_value ? ghv_23 : _GEN_1467; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1469 = 8'h18 == new_ptr_4_value ? ghv_24 : _GEN_1468; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1470 = 8'h19 == new_ptr_4_value ? ghv_25 : _GEN_1469; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1471 = 8'h1a == new_ptr_4_value ? ghv_26 : _GEN_1470; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1472 = 8'h1b == new_ptr_4_value ? ghv_27 : _GEN_1471; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1473 = 8'h1c == new_ptr_4_value ? ghv_28 : _GEN_1472; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1474 = 8'h1d == new_ptr_4_value ? ghv_29 : _GEN_1473; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1475 = 8'h1e == new_ptr_4_value ? ghv_30 : _GEN_1474; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1476 = 8'h1f == new_ptr_4_value ? ghv_31 : _GEN_1475; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1477 = 8'h20 == new_ptr_4_value ? ghv_32 : _GEN_1476; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1478 = 8'h21 == new_ptr_4_value ? ghv_33 : _GEN_1477; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1479 = 8'h22 == new_ptr_4_value ? ghv_34 : _GEN_1478; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1480 = 8'h23 == new_ptr_4_value ? ghv_35 : _GEN_1479; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1481 = 8'h24 == new_ptr_4_value ? ghv_36 : _GEN_1480; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1482 = 8'h25 == new_ptr_4_value ? ghv_37 : _GEN_1481; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1483 = 8'h26 == new_ptr_4_value ? ghv_38 : _GEN_1482; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1484 = 8'h27 == new_ptr_4_value ? ghv_39 : _GEN_1483; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1485 = 8'h28 == new_ptr_4_value ? ghv_40 : _GEN_1484; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1486 = 8'h29 == new_ptr_4_value ? ghv_41 : _GEN_1485; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1487 = 8'h2a == new_ptr_4_value ? ghv_42 : _GEN_1486; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1488 = 8'h2b == new_ptr_4_value ? ghv_43 : _GEN_1487; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1489 = 8'h2c == new_ptr_4_value ? ghv_44 : _GEN_1488; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1490 = 8'h2d == new_ptr_4_value ? ghv_45 : _GEN_1489; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1491 = 8'h2e == new_ptr_4_value ? ghv_46 : _GEN_1490; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1492 = 8'h2f == new_ptr_4_value ? ghv_47 : _GEN_1491; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1493 = 8'h30 == new_ptr_4_value ? ghv_48 : _GEN_1492; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1494 = 8'h31 == new_ptr_4_value ? ghv_49 : _GEN_1493; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1495 = 8'h32 == new_ptr_4_value ? ghv_50 : _GEN_1494; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1496 = 8'h33 == new_ptr_4_value ? ghv_51 : _GEN_1495; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1497 = 8'h34 == new_ptr_4_value ? ghv_52 : _GEN_1496; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1498 = 8'h35 == new_ptr_4_value ? ghv_53 : _GEN_1497; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1499 = 8'h36 == new_ptr_4_value ? ghv_54 : _GEN_1498; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1500 = 8'h37 == new_ptr_4_value ? ghv_55 : _GEN_1499; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1501 = 8'h38 == new_ptr_4_value ? ghv_56 : _GEN_1500; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1502 = 8'h39 == new_ptr_4_value ? ghv_57 : _GEN_1501; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1503 = 8'h3a == new_ptr_4_value ? ghv_58 : _GEN_1502; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1504 = 8'h3b == new_ptr_4_value ? ghv_59 : _GEN_1503; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1505 = 8'h3c == new_ptr_4_value ? ghv_60 : _GEN_1504; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1506 = 8'h3d == new_ptr_4_value ? ghv_61 : _GEN_1505; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1507 = 8'h3e == new_ptr_4_value ? ghv_62 : _GEN_1506; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1508 = 8'h3f == new_ptr_4_value ? ghv_63 : _GEN_1507; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1509 = 8'h40 == new_ptr_4_value ? ghv_64 : _GEN_1508; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1510 = 8'h41 == new_ptr_4_value ? ghv_65 : _GEN_1509; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1511 = 8'h42 == new_ptr_4_value ? ghv_66 : _GEN_1510; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1512 = 8'h43 == new_ptr_4_value ? ghv_67 : _GEN_1511; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1513 = 8'h44 == new_ptr_4_value ? ghv_68 : _GEN_1512; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1514 = 8'h45 == new_ptr_4_value ? ghv_69 : _GEN_1513; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1515 = 8'h46 == new_ptr_4_value ? ghv_70 : _GEN_1514; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1516 = 8'h47 == new_ptr_4_value ? ghv_71 : _GEN_1515; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1517 = 8'h48 == new_ptr_4_value ? ghv_72 : _GEN_1516; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1518 = 8'h49 == new_ptr_4_value ? ghv_73 : _GEN_1517; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1519 = 8'h4a == new_ptr_4_value ? ghv_74 : _GEN_1518; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1520 = 8'h4b == new_ptr_4_value ? ghv_75 : _GEN_1519; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1521 = 8'h4c == new_ptr_4_value ? ghv_76 : _GEN_1520; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1522 = 8'h4d == new_ptr_4_value ? ghv_77 : _GEN_1521; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1523 = 8'h4e == new_ptr_4_value ? ghv_78 : _GEN_1522; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1524 = 8'h4f == new_ptr_4_value ? ghv_79 : _GEN_1523; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1525 = 8'h50 == new_ptr_4_value ? ghv_80 : _GEN_1524; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1526 = 8'h51 == new_ptr_4_value ? ghv_81 : _GEN_1525; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1527 = 8'h52 == new_ptr_4_value ? ghv_82 : _GEN_1526; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1528 = 8'h53 == new_ptr_4_value ? ghv_83 : _GEN_1527; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1529 = 8'h54 == new_ptr_4_value ? ghv_84 : _GEN_1528; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1530 = 8'h55 == new_ptr_4_value ? ghv_85 : _GEN_1529; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1531 = 8'h56 == new_ptr_4_value ? ghv_86 : _GEN_1530; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1532 = 8'h57 == new_ptr_4_value ? ghv_87 : _GEN_1531; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1533 = 8'h58 == new_ptr_4_value ? ghv_88 : _GEN_1532; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1534 = 8'h59 == new_ptr_4_value ? ghv_89 : _GEN_1533; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1535 = 8'h5a == new_ptr_4_value ? ghv_90 : _GEN_1534; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1536 = 8'h5b == new_ptr_4_value ? ghv_91 : _GEN_1535; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1537 = 8'h5c == new_ptr_4_value ? ghv_92 : _GEN_1536; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1538 = 8'h5d == new_ptr_4_value ? ghv_93 : _GEN_1537; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1539 = 8'h5e == new_ptr_4_value ? ghv_94 : _GEN_1538; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1540 = 8'h5f == new_ptr_4_value ? ghv_95 : _GEN_1539; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1541 = 8'h60 == new_ptr_4_value ? ghv_96 : _GEN_1540; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1542 = 8'h61 == new_ptr_4_value ? ghv_97 : _GEN_1541; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1543 = 8'h62 == new_ptr_4_value ? ghv_98 : _GEN_1542; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1544 = 8'h63 == new_ptr_4_value ? ghv_99 : _GEN_1543; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1545 = 8'h64 == new_ptr_4_value ? ghv_100 : _GEN_1544; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1546 = 8'h65 == new_ptr_4_value ? ghv_101 : _GEN_1545; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1547 = 8'h66 == new_ptr_4_value ? ghv_102 : _GEN_1546; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1548 = 8'h67 == new_ptr_4_value ? ghv_103 : _GEN_1547; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1549 = 8'h68 == new_ptr_4_value ? ghv_104 : _GEN_1548; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1550 = 8'h69 == new_ptr_4_value ? ghv_105 : _GEN_1549; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1551 = 8'h6a == new_ptr_4_value ? ghv_106 : _GEN_1550; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1552 = 8'h6b == new_ptr_4_value ? ghv_107 : _GEN_1551; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1553 = 8'h6c == new_ptr_4_value ? ghv_108 : _GEN_1552; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1554 = 8'h6d == new_ptr_4_value ? ghv_109 : _GEN_1553; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1555 = 8'h6e == new_ptr_4_value ? ghv_110 : _GEN_1554; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1556 = 8'h6f == new_ptr_4_value ? ghv_111 : _GEN_1555; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1557 = 8'h70 == new_ptr_4_value ? ghv_112 : _GEN_1556; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1558 = 8'h71 == new_ptr_4_value ? ghv_113 : _GEN_1557; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1559 = 8'h72 == new_ptr_4_value ? ghv_114 : _GEN_1558; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1560 = 8'h73 == new_ptr_4_value ? ghv_115 : _GEN_1559; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1561 = 8'h74 == new_ptr_4_value ? ghv_116 : _GEN_1560; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1562 = 8'h75 == new_ptr_4_value ? ghv_117 : _GEN_1561; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1563 = 8'h76 == new_ptr_4_value ? ghv_118 : _GEN_1562; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1564 = 8'h77 == new_ptr_4_value ? ghv_119 : _GEN_1563; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1565 = 8'h78 == new_ptr_4_value ? ghv_120 : _GEN_1564; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1566 = 8'h79 == new_ptr_4_value ? ghv_121 : _GEN_1565; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1567 = 8'h7a == new_ptr_4_value ? ghv_122 : _GEN_1566; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1568 = 8'h7b == new_ptr_4_value ? ghv_123 : _GEN_1567; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1569 = 8'h7c == new_ptr_4_value ? ghv_124 : _GEN_1568; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1570 = 8'h7d == new_ptr_4_value ? ghv_125 : _GEN_1569; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1571 = 8'h7e == new_ptr_4_value ? ghv_126 : _GEN_1570; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1572 = 8'h7f == new_ptr_4_value ? ghv_127 : _GEN_1571; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1573 = 8'h80 == new_ptr_4_value ? ghv_128 : _GEN_1572; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1574 = 8'h81 == new_ptr_4_value ? ghv_129 : _GEN_1573; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1575 = 8'h82 == new_ptr_4_value ? ghv_130 : _GEN_1574; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1576 = 8'h83 == new_ptr_4_value ? ghv_131 : _GEN_1575; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1577 = 8'h84 == new_ptr_4_value ? ghv_132 : _GEN_1576; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1578 = 8'h85 == new_ptr_4_value ? ghv_133 : _GEN_1577; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1579 = 8'h86 == new_ptr_4_value ? ghv_134 : _GEN_1578; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1580 = 8'h87 == new_ptr_4_value ? ghv_135 : _GEN_1579; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1581 = 8'h88 == new_ptr_4_value ? ghv_136 : _GEN_1580; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1582 = 8'h89 == new_ptr_4_value ? ghv_137 : _GEN_1581; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1583 = 8'h8a == new_ptr_4_value ? ghv_138 : _GEN_1582; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1584 = 8'h8b == new_ptr_4_value ? ghv_139 : _GEN_1583; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1585 = 8'h8c == new_ptr_4_value ? ghv_140 : _GEN_1584; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1586 = 8'h8d == new_ptr_4_value ? ghv_141 : _GEN_1585; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1587 = 8'h8e == new_ptr_4_value ? ghv_142 : _GEN_1586; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_8_value = _new_ptr_value_T_17[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_1590 = 8'h1 == new_ptr_8_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1591 = 8'h2 == new_ptr_8_value ? ghv_2 : _GEN_1590; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1592 = 8'h3 == new_ptr_8_value ? ghv_3 : _GEN_1591; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1593 = 8'h4 == new_ptr_8_value ? ghv_4 : _GEN_1592; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1594 = 8'h5 == new_ptr_8_value ? ghv_5 : _GEN_1593; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1595 = 8'h6 == new_ptr_8_value ? ghv_6 : _GEN_1594; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1596 = 8'h7 == new_ptr_8_value ? ghv_7 : _GEN_1595; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1597 = 8'h8 == new_ptr_8_value ? ghv_8 : _GEN_1596; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1598 = 8'h9 == new_ptr_8_value ? ghv_9 : _GEN_1597; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1599 = 8'ha == new_ptr_8_value ? ghv_10 : _GEN_1598; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1600 = 8'hb == new_ptr_8_value ? ghv_11 : _GEN_1599; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1601 = 8'hc == new_ptr_8_value ? ghv_12 : _GEN_1600; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1602 = 8'hd == new_ptr_8_value ? ghv_13 : _GEN_1601; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1603 = 8'he == new_ptr_8_value ? ghv_14 : _GEN_1602; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1604 = 8'hf == new_ptr_8_value ? ghv_15 : _GEN_1603; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1605 = 8'h10 == new_ptr_8_value ? ghv_16 : _GEN_1604; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1606 = 8'h11 == new_ptr_8_value ? ghv_17 : _GEN_1605; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1607 = 8'h12 == new_ptr_8_value ? ghv_18 : _GEN_1606; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1608 = 8'h13 == new_ptr_8_value ? ghv_19 : _GEN_1607; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1609 = 8'h14 == new_ptr_8_value ? ghv_20 : _GEN_1608; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1610 = 8'h15 == new_ptr_8_value ? ghv_21 : _GEN_1609; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1611 = 8'h16 == new_ptr_8_value ? ghv_22 : _GEN_1610; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1612 = 8'h17 == new_ptr_8_value ? ghv_23 : _GEN_1611; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1613 = 8'h18 == new_ptr_8_value ? ghv_24 : _GEN_1612; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1614 = 8'h19 == new_ptr_8_value ? ghv_25 : _GEN_1613; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1615 = 8'h1a == new_ptr_8_value ? ghv_26 : _GEN_1614; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1616 = 8'h1b == new_ptr_8_value ? ghv_27 : _GEN_1615; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1617 = 8'h1c == new_ptr_8_value ? ghv_28 : _GEN_1616; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1618 = 8'h1d == new_ptr_8_value ? ghv_29 : _GEN_1617; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1619 = 8'h1e == new_ptr_8_value ? ghv_30 : _GEN_1618; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1620 = 8'h1f == new_ptr_8_value ? ghv_31 : _GEN_1619; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1621 = 8'h20 == new_ptr_8_value ? ghv_32 : _GEN_1620; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1622 = 8'h21 == new_ptr_8_value ? ghv_33 : _GEN_1621; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1623 = 8'h22 == new_ptr_8_value ? ghv_34 : _GEN_1622; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1624 = 8'h23 == new_ptr_8_value ? ghv_35 : _GEN_1623; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1625 = 8'h24 == new_ptr_8_value ? ghv_36 : _GEN_1624; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1626 = 8'h25 == new_ptr_8_value ? ghv_37 : _GEN_1625; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1627 = 8'h26 == new_ptr_8_value ? ghv_38 : _GEN_1626; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1628 = 8'h27 == new_ptr_8_value ? ghv_39 : _GEN_1627; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1629 = 8'h28 == new_ptr_8_value ? ghv_40 : _GEN_1628; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1630 = 8'h29 == new_ptr_8_value ? ghv_41 : _GEN_1629; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1631 = 8'h2a == new_ptr_8_value ? ghv_42 : _GEN_1630; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1632 = 8'h2b == new_ptr_8_value ? ghv_43 : _GEN_1631; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1633 = 8'h2c == new_ptr_8_value ? ghv_44 : _GEN_1632; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1634 = 8'h2d == new_ptr_8_value ? ghv_45 : _GEN_1633; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1635 = 8'h2e == new_ptr_8_value ? ghv_46 : _GEN_1634; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1636 = 8'h2f == new_ptr_8_value ? ghv_47 : _GEN_1635; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1637 = 8'h30 == new_ptr_8_value ? ghv_48 : _GEN_1636; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1638 = 8'h31 == new_ptr_8_value ? ghv_49 : _GEN_1637; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1639 = 8'h32 == new_ptr_8_value ? ghv_50 : _GEN_1638; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1640 = 8'h33 == new_ptr_8_value ? ghv_51 : _GEN_1639; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1641 = 8'h34 == new_ptr_8_value ? ghv_52 : _GEN_1640; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1642 = 8'h35 == new_ptr_8_value ? ghv_53 : _GEN_1641; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1643 = 8'h36 == new_ptr_8_value ? ghv_54 : _GEN_1642; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1644 = 8'h37 == new_ptr_8_value ? ghv_55 : _GEN_1643; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1645 = 8'h38 == new_ptr_8_value ? ghv_56 : _GEN_1644; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1646 = 8'h39 == new_ptr_8_value ? ghv_57 : _GEN_1645; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1647 = 8'h3a == new_ptr_8_value ? ghv_58 : _GEN_1646; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1648 = 8'h3b == new_ptr_8_value ? ghv_59 : _GEN_1647; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1649 = 8'h3c == new_ptr_8_value ? ghv_60 : _GEN_1648; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1650 = 8'h3d == new_ptr_8_value ? ghv_61 : _GEN_1649; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1651 = 8'h3e == new_ptr_8_value ? ghv_62 : _GEN_1650; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1652 = 8'h3f == new_ptr_8_value ? ghv_63 : _GEN_1651; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1653 = 8'h40 == new_ptr_8_value ? ghv_64 : _GEN_1652; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1654 = 8'h41 == new_ptr_8_value ? ghv_65 : _GEN_1653; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1655 = 8'h42 == new_ptr_8_value ? ghv_66 : _GEN_1654; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1656 = 8'h43 == new_ptr_8_value ? ghv_67 : _GEN_1655; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1657 = 8'h44 == new_ptr_8_value ? ghv_68 : _GEN_1656; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1658 = 8'h45 == new_ptr_8_value ? ghv_69 : _GEN_1657; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1659 = 8'h46 == new_ptr_8_value ? ghv_70 : _GEN_1658; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1660 = 8'h47 == new_ptr_8_value ? ghv_71 : _GEN_1659; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1661 = 8'h48 == new_ptr_8_value ? ghv_72 : _GEN_1660; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1662 = 8'h49 == new_ptr_8_value ? ghv_73 : _GEN_1661; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1663 = 8'h4a == new_ptr_8_value ? ghv_74 : _GEN_1662; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1664 = 8'h4b == new_ptr_8_value ? ghv_75 : _GEN_1663; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1665 = 8'h4c == new_ptr_8_value ? ghv_76 : _GEN_1664; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1666 = 8'h4d == new_ptr_8_value ? ghv_77 : _GEN_1665; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1667 = 8'h4e == new_ptr_8_value ? ghv_78 : _GEN_1666; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1668 = 8'h4f == new_ptr_8_value ? ghv_79 : _GEN_1667; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1669 = 8'h50 == new_ptr_8_value ? ghv_80 : _GEN_1668; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1670 = 8'h51 == new_ptr_8_value ? ghv_81 : _GEN_1669; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1671 = 8'h52 == new_ptr_8_value ? ghv_82 : _GEN_1670; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1672 = 8'h53 == new_ptr_8_value ? ghv_83 : _GEN_1671; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1673 = 8'h54 == new_ptr_8_value ? ghv_84 : _GEN_1672; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1674 = 8'h55 == new_ptr_8_value ? ghv_85 : _GEN_1673; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1675 = 8'h56 == new_ptr_8_value ? ghv_86 : _GEN_1674; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1676 = 8'h57 == new_ptr_8_value ? ghv_87 : _GEN_1675; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1677 = 8'h58 == new_ptr_8_value ? ghv_88 : _GEN_1676; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1678 = 8'h59 == new_ptr_8_value ? ghv_89 : _GEN_1677; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1679 = 8'h5a == new_ptr_8_value ? ghv_90 : _GEN_1678; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1680 = 8'h5b == new_ptr_8_value ? ghv_91 : _GEN_1679; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1681 = 8'h5c == new_ptr_8_value ? ghv_92 : _GEN_1680; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1682 = 8'h5d == new_ptr_8_value ? ghv_93 : _GEN_1681; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1683 = 8'h5e == new_ptr_8_value ? ghv_94 : _GEN_1682; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1684 = 8'h5f == new_ptr_8_value ? ghv_95 : _GEN_1683; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1685 = 8'h60 == new_ptr_8_value ? ghv_96 : _GEN_1684; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1686 = 8'h61 == new_ptr_8_value ? ghv_97 : _GEN_1685; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1687 = 8'h62 == new_ptr_8_value ? ghv_98 : _GEN_1686; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1688 = 8'h63 == new_ptr_8_value ? ghv_99 : _GEN_1687; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1689 = 8'h64 == new_ptr_8_value ? ghv_100 : _GEN_1688; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1690 = 8'h65 == new_ptr_8_value ? ghv_101 : _GEN_1689; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1691 = 8'h66 == new_ptr_8_value ? ghv_102 : _GEN_1690; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1692 = 8'h67 == new_ptr_8_value ? ghv_103 : _GEN_1691; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1693 = 8'h68 == new_ptr_8_value ? ghv_104 : _GEN_1692; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1694 = 8'h69 == new_ptr_8_value ? ghv_105 : _GEN_1693; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1695 = 8'h6a == new_ptr_8_value ? ghv_106 : _GEN_1694; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1696 = 8'h6b == new_ptr_8_value ? ghv_107 : _GEN_1695; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1697 = 8'h6c == new_ptr_8_value ? ghv_108 : _GEN_1696; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1698 = 8'h6d == new_ptr_8_value ? ghv_109 : _GEN_1697; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1699 = 8'h6e == new_ptr_8_value ? ghv_110 : _GEN_1698; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1700 = 8'h6f == new_ptr_8_value ? ghv_111 : _GEN_1699; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1701 = 8'h70 == new_ptr_8_value ? ghv_112 : _GEN_1700; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1702 = 8'h71 == new_ptr_8_value ? ghv_113 : _GEN_1701; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1703 = 8'h72 == new_ptr_8_value ? ghv_114 : _GEN_1702; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1704 = 8'h73 == new_ptr_8_value ? ghv_115 : _GEN_1703; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1705 = 8'h74 == new_ptr_8_value ? ghv_116 : _GEN_1704; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1706 = 8'h75 == new_ptr_8_value ? ghv_117 : _GEN_1705; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1707 = 8'h76 == new_ptr_8_value ? ghv_118 : _GEN_1706; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1708 = 8'h77 == new_ptr_8_value ? ghv_119 : _GEN_1707; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1709 = 8'h78 == new_ptr_8_value ? ghv_120 : _GEN_1708; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1710 = 8'h79 == new_ptr_8_value ? ghv_121 : _GEN_1709; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1711 = 8'h7a == new_ptr_8_value ? ghv_122 : _GEN_1710; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1712 = 8'h7b == new_ptr_8_value ? ghv_123 : _GEN_1711; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1713 = 8'h7c == new_ptr_8_value ? ghv_124 : _GEN_1712; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1714 = 8'h7d == new_ptr_8_value ? ghv_125 : _GEN_1713; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1715 = 8'h7e == new_ptr_8_value ? ghv_126 : _GEN_1714; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1716 = 8'h7f == new_ptr_8_value ? ghv_127 : _GEN_1715; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1717 = 8'h80 == new_ptr_8_value ? ghv_128 : _GEN_1716; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1718 = 8'h81 == new_ptr_8_value ? ghv_129 : _GEN_1717; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1719 = 8'h82 == new_ptr_8_value ? ghv_130 : _GEN_1718; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1720 = 8'h83 == new_ptr_8_value ? ghv_131 : _GEN_1719; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1721 = 8'h84 == new_ptr_8_value ? ghv_132 : _GEN_1720; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1722 = 8'h85 == new_ptr_8_value ? ghv_133 : _GEN_1721; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1723 = 8'h86 == new_ptr_8_value ? ghv_134 : _GEN_1722; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1724 = 8'h87 == new_ptr_8_value ? ghv_135 : _GEN_1723; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1725 = 8'h88 == new_ptr_8_value ? ghv_136 : _GEN_1724; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1726 = 8'h89 == new_ptr_8_value ? ghv_137 : _GEN_1725; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1727 = 8'h8a == new_ptr_8_value ? ghv_138 : _GEN_1726; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1728 = 8'h8b == new_ptr_8_value ? ghv_139 : _GEN_1727; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1729 = 8'h8c == new_ptr_8_value ? ghv_140 : _GEN_1728; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1730 = 8'h8d == new_ptr_8_value ? ghv_141 : _GEN_1729; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1731 = 8'h8e == new_ptr_8_value ? ghv_142 : _GEN_1730; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_19_value = _new_ptr_value_T_39[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_1734 = 8'h1 == new_ptr_19_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1735 = 8'h2 == new_ptr_19_value ? ghv_2 : _GEN_1734; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1736 = 8'h3 == new_ptr_19_value ? ghv_3 : _GEN_1735; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1737 = 8'h4 == new_ptr_19_value ? ghv_4 : _GEN_1736; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1738 = 8'h5 == new_ptr_19_value ? ghv_5 : _GEN_1737; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1739 = 8'h6 == new_ptr_19_value ? ghv_6 : _GEN_1738; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1740 = 8'h7 == new_ptr_19_value ? ghv_7 : _GEN_1739; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1741 = 8'h8 == new_ptr_19_value ? ghv_8 : _GEN_1740; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1742 = 8'h9 == new_ptr_19_value ? ghv_9 : _GEN_1741; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1743 = 8'ha == new_ptr_19_value ? ghv_10 : _GEN_1742; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1744 = 8'hb == new_ptr_19_value ? ghv_11 : _GEN_1743; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1745 = 8'hc == new_ptr_19_value ? ghv_12 : _GEN_1744; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1746 = 8'hd == new_ptr_19_value ? ghv_13 : _GEN_1745; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1747 = 8'he == new_ptr_19_value ? ghv_14 : _GEN_1746; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1748 = 8'hf == new_ptr_19_value ? ghv_15 : _GEN_1747; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1749 = 8'h10 == new_ptr_19_value ? ghv_16 : _GEN_1748; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1750 = 8'h11 == new_ptr_19_value ? ghv_17 : _GEN_1749; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1751 = 8'h12 == new_ptr_19_value ? ghv_18 : _GEN_1750; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1752 = 8'h13 == new_ptr_19_value ? ghv_19 : _GEN_1751; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1753 = 8'h14 == new_ptr_19_value ? ghv_20 : _GEN_1752; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1754 = 8'h15 == new_ptr_19_value ? ghv_21 : _GEN_1753; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1755 = 8'h16 == new_ptr_19_value ? ghv_22 : _GEN_1754; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1756 = 8'h17 == new_ptr_19_value ? ghv_23 : _GEN_1755; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1757 = 8'h18 == new_ptr_19_value ? ghv_24 : _GEN_1756; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1758 = 8'h19 == new_ptr_19_value ? ghv_25 : _GEN_1757; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1759 = 8'h1a == new_ptr_19_value ? ghv_26 : _GEN_1758; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1760 = 8'h1b == new_ptr_19_value ? ghv_27 : _GEN_1759; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1761 = 8'h1c == new_ptr_19_value ? ghv_28 : _GEN_1760; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1762 = 8'h1d == new_ptr_19_value ? ghv_29 : _GEN_1761; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1763 = 8'h1e == new_ptr_19_value ? ghv_30 : _GEN_1762; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1764 = 8'h1f == new_ptr_19_value ? ghv_31 : _GEN_1763; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1765 = 8'h20 == new_ptr_19_value ? ghv_32 : _GEN_1764; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1766 = 8'h21 == new_ptr_19_value ? ghv_33 : _GEN_1765; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1767 = 8'h22 == new_ptr_19_value ? ghv_34 : _GEN_1766; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1768 = 8'h23 == new_ptr_19_value ? ghv_35 : _GEN_1767; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1769 = 8'h24 == new_ptr_19_value ? ghv_36 : _GEN_1768; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1770 = 8'h25 == new_ptr_19_value ? ghv_37 : _GEN_1769; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1771 = 8'h26 == new_ptr_19_value ? ghv_38 : _GEN_1770; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1772 = 8'h27 == new_ptr_19_value ? ghv_39 : _GEN_1771; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1773 = 8'h28 == new_ptr_19_value ? ghv_40 : _GEN_1772; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1774 = 8'h29 == new_ptr_19_value ? ghv_41 : _GEN_1773; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1775 = 8'h2a == new_ptr_19_value ? ghv_42 : _GEN_1774; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1776 = 8'h2b == new_ptr_19_value ? ghv_43 : _GEN_1775; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1777 = 8'h2c == new_ptr_19_value ? ghv_44 : _GEN_1776; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1778 = 8'h2d == new_ptr_19_value ? ghv_45 : _GEN_1777; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1779 = 8'h2e == new_ptr_19_value ? ghv_46 : _GEN_1778; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1780 = 8'h2f == new_ptr_19_value ? ghv_47 : _GEN_1779; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1781 = 8'h30 == new_ptr_19_value ? ghv_48 : _GEN_1780; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1782 = 8'h31 == new_ptr_19_value ? ghv_49 : _GEN_1781; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1783 = 8'h32 == new_ptr_19_value ? ghv_50 : _GEN_1782; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1784 = 8'h33 == new_ptr_19_value ? ghv_51 : _GEN_1783; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1785 = 8'h34 == new_ptr_19_value ? ghv_52 : _GEN_1784; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1786 = 8'h35 == new_ptr_19_value ? ghv_53 : _GEN_1785; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1787 = 8'h36 == new_ptr_19_value ? ghv_54 : _GEN_1786; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1788 = 8'h37 == new_ptr_19_value ? ghv_55 : _GEN_1787; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1789 = 8'h38 == new_ptr_19_value ? ghv_56 : _GEN_1788; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1790 = 8'h39 == new_ptr_19_value ? ghv_57 : _GEN_1789; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1791 = 8'h3a == new_ptr_19_value ? ghv_58 : _GEN_1790; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1792 = 8'h3b == new_ptr_19_value ? ghv_59 : _GEN_1791; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1793 = 8'h3c == new_ptr_19_value ? ghv_60 : _GEN_1792; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1794 = 8'h3d == new_ptr_19_value ? ghv_61 : _GEN_1793; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1795 = 8'h3e == new_ptr_19_value ? ghv_62 : _GEN_1794; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1796 = 8'h3f == new_ptr_19_value ? ghv_63 : _GEN_1795; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1797 = 8'h40 == new_ptr_19_value ? ghv_64 : _GEN_1796; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1798 = 8'h41 == new_ptr_19_value ? ghv_65 : _GEN_1797; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1799 = 8'h42 == new_ptr_19_value ? ghv_66 : _GEN_1798; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1800 = 8'h43 == new_ptr_19_value ? ghv_67 : _GEN_1799; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1801 = 8'h44 == new_ptr_19_value ? ghv_68 : _GEN_1800; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1802 = 8'h45 == new_ptr_19_value ? ghv_69 : _GEN_1801; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1803 = 8'h46 == new_ptr_19_value ? ghv_70 : _GEN_1802; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1804 = 8'h47 == new_ptr_19_value ? ghv_71 : _GEN_1803; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1805 = 8'h48 == new_ptr_19_value ? ghv_72 : _GEN_1804; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1806 = 8'h49 == new_ptr_19_value ? ghv_73 : _GEN_1805; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1807 = 8'h4a == new_ptr_19_value ? ghv_74 : _GEN_1806; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1808 = 8'h4b == new_ptr_19_value ? ghv_75 : _GEN_1807; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1809 = 8'h4c == new_ptr_19_value ? ghv_76 : _GEN_1808; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1810 = 8'h4d == new_ptr_19_value ? ghv_77 : _GEN_1809; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1811 = 8'h4e == new_ptr_19_value ? ghv_78 : _GEN_1810; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1812 = 8'h4f == new_ptr_19_value ? ghv_79 : _GEN_1811; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1813 = 8'h50 == new_ptr_19_value ? ghv_80 : _GEN_1812; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1814 = 8'h51 == new_ptr_19_value ? ghv_81 : _GEN_1813; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1815 = 8'h52 == new_ptr_19_value ? ghv_82 : _GEN_1814; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1816 = 8'h53 == new_ptr_19_value ? ghv_83 : _GEN_1815; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1817 = 8'h54 == new_ptr_19_value ? ghv_84 : _GEN_1816; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1818 = 8'h55 == new_ptr_19_value ? ghv_85 : _GEN_1817; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1819 = 8'h56 == new_ptr_19_value ? ghv_86 : _GEN_1818; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1820 = 8'h57 == new_ptr_19_value ? ghv_87 : _GEN_1819; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1821 = 8'h58 == new_ptr_19_value ? ghv_88 : _GEN_1820; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1822 = 8'h59 == new_ptr_19_value ? ghv_89 : _GEN_1821; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1823 = 8'h5a == new_ptr_19_value ? ghv_90 : _GEN_1822; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1824 = 8'h5b == new_ptr_19_value ? ghv_91 : _GEN_1823; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1825 = 8'h5c == new_ptr_19_value ? ghv_92 : _GEN_1824; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1826 = 8'h5d == new_ptr_19_value ? ghv_93 : _GEN_1825; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1827 = 8'h5e == new_ptr_19_value ? ghv_94 : _GEN_1826; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1828 = 8'h5f == new_ptr_19_value ? ghv_95 : _GEN_1827; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1829 = 8'h60 == new_ptr_19_value ? ghv_96 : _GEN_1828; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1830 = 8'h61 == new_ptr_19_value ? ghv_97 : _GEN_1829; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1831 = 8'h62 == new_ptr_19_value ? ghv_98 : _GEN_1830; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1832 = 8'h63 == new_ptr_19_value ? ghv_99 : _GEN_1831; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1833 = 8'h64 == new_ptr_19_value ? ghv_100 : _GEN_1832; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1834 = 8'h65 == new_ptr_19_value ? ghv_101 : _GEN_1833; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1835 = 8'h66 == new_ptr_19_value ? ghv_102 : _GEN_1834; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1836 = 8'h67 == new_ptr_19_value ? ghv_103 : _GEN_1835; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1837 = 8'h68 == new_ptr_19_value ? ghv_104 : _GEN_1836; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1838 = 8'h69 == new_ptr_19_value ? ghv_105 : _GEN_1837; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1839 = 8'h6a == new_ptr_19_value ? ghv_106 : _GEN_1838; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1840 = 8'h6b == new_ptr_19_value ? ghv_107 : _GEN_1839; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1841 = 8'h6c == new_ptr_19_value ? ghv_108 : _GEN_1840; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1842 = 8'h6d == new_ptr_19_value ? ghv_109 : _GEN_1841; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1843 = 8'h6e == new_ptr_19_value ? ghv_110 : _GEN_1842; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1844 = 8'h6f == new_ptr_19_value ? ghv_111 : _GEN_1843; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1845 = 8'h70 == new_ptr_19_value ? ghv_112 : _GEN_1844; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1846 = 8'h71 == new_ptr_19_value ? ghv_113 : _GEN_1845; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1847 = 8'h72 == new_ptr_19_value ? ghv_114 : _GEN_1846; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1848 = 8'h73 == new_ptr_19_value ? ghv_115 : _GEN_1847; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1849 = 8'h74 == new_ptr_19_value ? ghv_116 : _GEN_1848; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1850 = 8'h75 == new_ptr_19_value ? ghv_117 : _GEN_1849; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1851 = 8'h76 == new_ptr_19_value ? ghv_118 : _GEN_1850; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1852 = 8'h77 == new_ptr_19_value ? ghv_119 : _GEN_1851; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1853 = 8'h78 == new_ptr_19_value ? ghv_120 : _GEN_1852; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1854 = 8'h79 == new_ptr_19_value ? ghv_121 : _GEN_1853; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1855 = 8'h7a == new_ptr_19_value ? ghv_122 : _GEN_1854; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1856 = 8'h7b == new_ptr_19_value ? ghv_123 : _GEN_1855; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1857 = 8'h7c == new_ptr_19_value ? ghv_124 : _GEN_1856; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1858 = 8'h7d == new_ptr_19_value ? ghv_125 : _GEN_1857; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1859 = 8'h7e == new_ptr_19_value ? ghv_126 : _GEN_1858; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1860 = 8'h7f == new_ptr_19_value ? ghv_127 : _GEN_1859; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1861 = 8'h80 == new_ptr_19_value ? ghv_128 : _GEN_1860; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1862 = 8'h81 == new_ptr_19_value ? ghv_129 : _GEN_1861; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1863 = 8'h82 == new_ptr_19_value ? ghv_130 : _GEN_1862; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1864 = 8'h83 == new_ptr_19_value ? ghv_131 : _GEN_1863; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1865 = 8'h84 == new_ptr_19_value ? ghv_132 : _GEN_1864; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1866 = 8'h85 == new_ptr_19_value ? ghv_133 : _GEN_1865; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1867 = 8'h86 == new_ptr_19_value ? ghv_134 : _GEN_1866; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1868 = 8'h87 == new_ptr_19_value ? ghv_135 : _GEN_1867; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1869 = 8'h88 == new_ptr_19_value ? ghv_136 : _GEN_1868; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1870 = 8'h89 == new_ptr_19_value ? ghv_137 : _GEN_1869; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1871 = 8'h8a == new_ptr_19_value ? ghv_138 : _GEN_1870; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1872 = 8'h8b == new_ptr_19_value ? ghv_139 : _GEN_1871; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1873 = 8'h8c == new_ptr_19_value ? ghv_140 : _GEN_1872; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1874 = 8'h8d == new_ptr_19_value ? ghv_141 : _GEN_1873; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1875 = 8'h8e == new_ptr_19_value ? ghv_142 : _GEN_1874; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_3_value = _new_ptr_value_T_7[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_1878 = 8'h1 == new_ptr_3_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1879 = 8'h2 == new_ptr_3_value ? ghv_2 : _GEN_1878; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1880 = 8'h3 == new_ptr_3_value ? ghv_3 : _GEN_1879; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1881 = 8'h4 == new_ptr_3_value ? ghv_4 : _GEN_1880; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1882 = 8'h5 == new_ptr_3_value ? ghv_5 : _GEN_1881; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1883 = 8'h6 == new_ptr_3_value ? ghv_6 : _GEN_1882; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1884 = 8'h7 == new_ptr_3_value ? ghv_7 : _GEN_1883; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1885 = 8'h8 == new_ptr_3_value ? ghv_8 : _GEN_1884; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1886 = 8'h9 == new_ptr_3_value ? ghv_9 : _GEN_1885; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1887 = 8'ha == new_ptr_3_value ? ghv_10 : _GEN_1886; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1888 = 8'hb == new_ptr_3_value ? ghv_11 : _GEN_1887; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1889 = 8'hc == new_ptr_3_value ? ghv_12 : _GEN_1888; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1890 = 8'hd == new_ptr_3_value ? ghv_13 : _GEN_1889; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1891 = 8'he == new_ptr_3_value ? ghv_14 : _GEN_1890; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1892 = 8'hf == new_ptr_3_value ? ghv_15 : _GEN_1891; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1893 = 8'h10 == new_ptr_3_value ? ghv_16 : _GEN_1892; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1894 = 8'h11 == new_ptr_3_value ? ghv_17 : _GEN_1893; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1895 = 8'h12 == new_ptr_3_value ? ghv_18 : _GEN_1894; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1896 = 8'h13 == new_ptr_3_value ? ghv_19 : _GEN_1895; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1897 = 8'h14 == new_ptr_3_value ? ghv_20 : _GEN_1896; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1898 = 8'h15 == new_ptr_3_value ? ghv_21 : _GEN_1897; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1899 = 8'h16 == new_ptr_3_value ? ghv_22 : _GEN_1898; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1900 = 8'h17 == new_ptr_3_value ? ghv_23 : _GEN_1899; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1901 = 8'h18 == new_ptr_3_value ? ghv_24 : _GEN_1900; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1902 = 8'h19 == new_ptr_3_value ? ghv_25 : _GEN_1901; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1903 = 8'h1a == new_ptr_3_value ? ghv_26 : _GEN_1902; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1904 = 8'h1b == new_ptr_3_value ? ghv_27 : _GEN_1903; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1905 = 8'h1c == new_ptr_3_value ? ghv_28 : _GEN_1904; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1906 = 8'h1d == new_ptr_3_value ? ghv_29 : _GEN_1905; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1907 = 8'h1e == new_ptr_3_value ? ghv_30 : _GEN_1906; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1908 = 8'h1f == new_ptr_3_value ? ghv_31 : _GEN_1907; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1909 = 8'h20 == new_ptr_3_value ? ghv_32 : _GEN_1908; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1910 = 8'h21 == new_ptr_3_value ? ghv_33 : _GEN_1909; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1911 = 8'h22 == new_ptr_3_value ? ghv_34 : _GEN_1910; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1912 = 8'h23 == new_ptr_3_value ? ghv_35 : _GEN_1911; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1913 = 8'h24 == new_ptr_3_value ? ghv_36 : _GEN_1912; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1914 = 8'h25 == new_ptr_3_value ? ghv_37 : _GEN_1913; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1915 = 8'h26 == new_ptr_3_value ? ghv_38 : _GEN_1914; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1916 = 8'h27 == new_ptr_3_value ? ghv_39 : _GEN_1915; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1917 = 8'h28 == new_ptr_3_value ? ghv_40 : _GEN_1916; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1918 = 8'h29 == new_ptr_3_value ? ghv_41 : _GEN_1917; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1919 = 8'h2a == new_ptr_3_value ? ghv_42 : _GEN_1918; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1920 = 8'h2b == new_ptr_3_value ? ghv_43 : _GEN_1919; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1921 = 8'h2c == new_ptr_3_value ? ghv_44 : _GEN_1920; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1922 = 8'h2d == new_ptr_3_value ? ghv_45 : _GEN_1921; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1923 = 8'h2e == new_ptr_3_value ? ghv_46 : _GEN_1922; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1924 = 8'h2f == new_ptr_3_value ? ghv_47 : _GEN_1923; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1925 = 8'h30 == new_ptr_3_value ? ghv_48 : _GEN_1924; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1926 = 8'h31 == new_ptr_3_value ? ghv_49 : _GEN_1925; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1927 = 8'h32 == new_ptr_3_value ? ghv_50 : _GEN_1926; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1928 = 8'h33 == new_ptr_3_value ? ghv_51 : _GEN_1927; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1929 = 8'h34 == new_ptr_3_value ? ghv_52 : _GEN_1928; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1930 = 8'h35 == new_ptr_3_value ? ghv_53 : _GEN_1929; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1931 = 8'h36 == new_ptr_3_value ? ghv_54 : _GEN_1930; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1932 = 8'h37 == new_ptr_3_value ? ghv_55 : _GEN_1931; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1933 = 8'h38 == new_ptr_3_value ? ghv_56 : _GEN_1932; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1934 = 8'h39 == new_ptr_3_value ? ghv_57 : _GEN_1933; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1935 = 8'h3a == new_ptr_3_value ? ghv_58 : _GEN_1934; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1936 = 8'h3b == new_ptr_3_value ? ghv_59 : _GEN_1935; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1937 = 8'h3c == new_ptr_3_value ? ghv_60 : _GEN_1936; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1938 = 8'h3d == new_ptr_3_value ? ghv_61 : _GEN_1937; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1939 = 8'h3e == new_ptr_3_value ? ghv_62 : _GEN_1938; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1940 = 8'h3f == new_ptr_3_value ? ghv_63 : _GEN_1939; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1941 = 8'h40 == new_ptr_3_value ? ghv_64 : _GEN_1940; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1942 = 8'h41 == new_ptr_3_value ? ghv_65 : _GEN_1941; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1943 = 8'h42 == new_ptr_3_value ? ghv_66 : _GEN_1942; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1944 = 8'h43 == new_ptr_3_value ? ghv_67 : _GEN_1943; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1945 = 8'h44 == new_ptr_3_value ? ghv_68 : _GEN_1944; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1946 = 8'h45 == new_ptr_3_value ? ghv_69 : _GEN_1945; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1947 = 8'h46 == new_ptr_3_value ? ghv_70 : _GEN_1946; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1948 = 8'h47 == new_ptr_3_value ? ghv_71 : _GEN_1947; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1949 = 8'h48 == new_ptr_3_value ? ghv_72 : _GEN_1948; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1950 = 8'h49 == new_ptr_3_value ? ghv_73 : _GEN_1949; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1951 = 8'h4a == new_ptr_3_value ? ghv_74 : _GEN_1950; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1952 = 8'h4b == new_ptr_3_value ? ghv_75 : _GEN_1951; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1953 = 8'h4c == new_ptr_3_value ? ghv_76 : _GEN_1952; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1954 = 8'h4d == new_ptr_3_value ? ghv_77 : _GEN_1953; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1955 = 8'h4e == new_ptr_3_value ? ghv_78 : _GEN_1954; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1956 = 8'h4f == new_ptr_3_value ? ghv_79 : _GEN_1955; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1957 = 8'h50 == new_ptr_3_value ? ghv_80 : _GEN_1956; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1958 = 8'h51 == new_ptr_3_value ? ghv_81 : _GEN_1957; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1959 = 8'h52 == new_ptr_3_value ? ghv_82 : _GEN_1958; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1960 = 8'h53 == new_ptr_3_value ? ghv_83 : _GEN_1959; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1961 = 8'h54 == new_ptr_3_value ? ghv_84 : _GEN_1960; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1962 = 8'h55 == new_ptr_3_value ? ghv_85 : _GEN_1961; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1963 = 8'h56 == new_ptr_3_value ? ghv_86 : _GEN_1962; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1964 = 8'h57 == new_ptr_3_value ? ghv_87 : _GEN_1963; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1965 = 8'h58 == new_ptr_3_value ? ghv_88 : _GEN_1964; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1966 = 8'h59 == new_ptr_3_value ? ghv_89 : _GEN_1965; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1967 = 8'h5a == new_ptr_3_value ? ghv_90 : _GEN_1966; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1968 = 8'h5b == new_ptr_3_value ? ghv_91 : _GEN_1967; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1969 = 8'h5c == new_ptr_3_value ? ghv_92 : _GEN_1968; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1970 = 8'h5d == new_ptr_3_value ? ghv_93 : _GEN_1969; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1971 = 8'h5e == new_ptr_3_value ? ghv_94 : _GEN_1970; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1972 = 8'h5f == new_ptr_3_value ? ghv_95 : _GEN_1971; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1973 = 8'h60 == new_ptr_3_value ? ghv_96 : _GEN_1972; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1974 = 8'h61 == new_ptr_3_value ? ghv_97 : _GEN_1973; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1975 = 8'h62 == new_ptr_3_value ? ghv_98 : _GEN_1974; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1976 = 8'h63 == new_ptr_3_value ? ghv_99 : _GEN_1975; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1977 = 8'h64 == new_ptr_3_value ? ghv_100 : _GEN_1976; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1978 = 8'h65 == new_ptr_3_value ? ghv_101 : _GEN_1977; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1979 = 8'h66 == new_ptr_3_value ? ghv_102 : _GEN_1978; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1980 = 8'h67 == new_ptr_3_value ? ghv_103 : _GEN_1979; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1981 = 8'h68 == new_ptr_3_value ? ghv_104 : _GEN_1980; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1982 = 8'h69 == new_ptr_3_value ? ghv_105 : _GEN_1981; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1983 = 8'h6a == new_ptr_3_value ? ghv_106 : _GEN_1982; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1984 = 8'h6b == new_ptr_3_value ? ghv_107 : _GEN_1983; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1985 = 8'h6c == new_ptr_3_value ? ghv_108 : _GEN_1984; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1986 = 8'h6d == new_ptr_3_value ? ghv_109 : _GEN_1985; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1987 = 8'h6e == new_ptr_3_value ? ghv_110 : _GEN_1986; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1988 = 8'h6f == new_ptr_3_value ? ghv_111 : _GEN_1987; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1989 = 8'h70 == new_ptr_3_value ? ghv_112 : _GEN_1988; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1990 = 8'h71 == new_ptr_3_value ? ghv_113 : _GEN_1989; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1991 = 8'h72 == new_ptr_3_value ? ghv_114 : _GEN_1990; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1992 = 8'h73 == new_ptr_3_value ? ghv_115 : _GEN_1991; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1993 = 8'h74 == new_ptr_3_value ? ghv_116 : _GEN_1992; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1994 = 8'h75 == new_ptr_3_value ? ghv_117 : _GEN_1993; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1995 = 8'h76 == new_ptr_3_value ? ghv_118 : _GEN_1994; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1996 = 8'h77 == new_ptr_3_value ? ghv_119 : _GEN_1995; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1997 = 8'h78 == new_ptr_3_value ? ghv_120 : _GEN_1996; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1998 = 8'h79 == new_ptr_3_value ? ghv_121 : _GEN_1997; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_1999 = 8'h7a == new_ptr_3_value ? ghv_122 : _GEN_1998; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2000 = 8'h7b == new_ptr_3_value ? ghv_123 : _GEN_1999; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2001 = 8'h7c == new_ptr_3_value ? ghv_124 : _GEN_2000; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2002 = 8'h7d == new_ptr_3_value ? ghv_125 : _GEN_2001; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2003 = 8'h7e == new_ptr_3_value ? ghv_126 : _GEN_2002; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2004 = 8'h7f == new_ptr_3_value ? ghv_127 : _GEN_2003; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2005 = 8'h80 == new_ptr_3_value ? ghv_128 : _GEN_2004; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2006 = 8'h81 == new_ptr_3_value ? ghv_129 : _GEN_2005; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2007 = 8'h82 == new_ptr_3_value ? ghv_130 : _GEN_2006; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2008 = 8'h83 == new_ptr_3_value ? ghv_131 : _GEN_2007; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2009 = 8'h84 == new_ptr_3_value ? ghv_132 : _GEN_2008; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2010 = 8'h85 == new_ptr_3_value ? ghv_133 : _GEN_2009; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2011 = 8'h86 == new_ptr_3_value ? ghv_134 : _GEN_2010; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2012 = 8'h87 == new_ptr_3_value ? ghv_135 : _GEN_2011; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2013 = 8'h88 == new_ptr_3_value ? ghv_136 : _GEN_2012; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2014 = 8'h89 == new_ptr_3_value ? ghv_137 : _GEN_2013; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2015 = 8'h8a == new_ptr_3_value ? ghv_138 : _GEN_2014; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2016 = 8'h8b == new_ptr_3_value ? ghv_139 : _GEN_2015; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2017 = 8'h8c == new_ptr_3_value ? ghv_140 : _GEN_2016; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2018 = 8'h8d == new_ptr_3_value ? ghv_141 : _GEN_2017; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2019 = 8'h8e == new_ptr_3_value ? ghv_142 : _GEN_2018; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_10_value = _new_ptr_value_T_21[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_2022 = 8'h1 == new_ptr_10_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2023 = 8'h2 == new_ptr_10_value ? ghv_2 : _GEN_2022; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2024 = 8'h3 == new_ptr_10_value ? ghv_3 : _GEN_2023; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2025 = 8'h4 == new_ptr_10_value ? ghv_4 : _GEN_2024; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2026 = 8'h5 == new_ptr_10_value ? ghv_5 : _GEN_2025; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2027 = 8'h6 == new_ptr_10_value ? ghv_6 : _GEN_2026; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2028 = 8'h7 == new_ptr_10_value ? ghv_7 : _GEN_2027; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2029 = 8'h8 == new_ptr_10_value ? ghv_8 : _GEN_2028; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2030 = 8'h9 == new_ptr_10_value ? ghv_9 : _GEN_2029; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2031 = 8'ha == new_ptr_10_value ? ghv_10 : _GEN_2030; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2032 = 8'hb == new_ptr_10_value ? ghv_11 : _GEN_2031; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2033 = 8'hc == new_ptr_10_value ? ghv_12 : _GEN_2032; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2034 = 8'hd == new_ptr_10_value ? ghv_13 : _GEN_2033; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2035 = 8'he == new_ptr_10_value ? ghv_14 : _GEN_2034; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2036 = 8'hf == new_ptr_10_value ? ghv_15 : _GEN_2035; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2037 = 8'h10 == new_ptr_10_value ? ghv_16 : _GEN_2036; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2038 = 8'h11 == new_ptr_10_value ? ghv_17 : _GEN_2037; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2039 = 8'h12 == new_ptr_10_value ? ghv_18 : _GEN_2038; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2040 = 8'h13 == new_ptr_10_value ? ghv_19 : _GEN_2039; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2041 = 8'h14 == new_ptr_10_value ? ghv_20 : _GEN_2040; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2042 = 8'h15 == new_ptr_10_value ? ghv_21 : _GEN_2041; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2043 = 8'h16 == new_ptr_10_value ? ghv_22 : _GEN_2042; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2044 = 8'h17 == new_ptr_10_value ? ghv_23 : _GEN_2043; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2045 = 8'h18 == new_ptr_10_value ? ghv_24 : _GEN_2044; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2046 = 8'h19 == new_ptr_10_value ? ghv_25 : _GEN_2045; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2047 = 8'h1a == new_ptr_10_value ? ghv_26 : _GEN_2046; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2048 = 8'h1b == new_ptr_10_value ? ghv_27 : _GEN_2047; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2049 = 8'h1c == new_ptr_10_value ? ghv_28 : _GEN_2048; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2050 = 8'h1d == new_ptr_10_value ? ghv_29 : _GEN_2049; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2051 = 8'h1e == new_ptr_10_value ? ghv_30 : _GEN_2050; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2052 = 8'h1f == new_ptr_10_value ? ghv_31 : _GEN_2051; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2053 = 8'h20 == new_ptr_10_value ? ghv_32 : _GEN_2052; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2054 = 8'h21 == new_ptr_10_value ? ghv_33 : _GEN_2053; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2055 = 8'h22 == new_ptr_10_value ? ghv_34 : _GEN_2054; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2056 = 8'h23 == new_ptr_10_value ? ghv_35 : _GEN_2055; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2057 = 8'h24 == new_ptr_10_value ? ghv_36 : _GEN_2056; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2058 = 8'h25 == new_ptr_10_value ? ghv_37 : _GEN_2057; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2059 = 8'h26 == new_ptr_10_value ? ghv_38 : _GEN_2058; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2060 = 8'h27 == new_ptr_10_value ? ghv_39 : _GEN_2059; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2061 = 8'h28 == new_ptr_10_value ? ghv_40 : _GEN_2060; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2062 = 8'h29 == new_ptr_10_value ? ghv_41 : _GEN_2061; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2063 = 8'h2a == new_ptr_10_value ? ghv_42 : _GEN_2062; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2064 = 8'h2b == new_ptr_10_value ? ghv_43 : _GEN_2063; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2065 = 8'h2c == new_ptr_10_value ? ghv_44 : _GEN_2064; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2066 = 8'h2d == new_ptr_10_value ? ghv_45 : _GEN_2065; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2067 = 8'h2e == new_ptr_10_value ? ghv_46 : _GEN_2066; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2068 = 8'h2f == new_ptr_10_value ? ghv_47 : _GEN_2067; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2069 = 8'h30 == new_ptr_10_value ? ghv_48 : _GEN_2068; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2070 = 8'h31 == new_ptr_10_value ? ghv_49 : _GEN_2069; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2071 = 8'h32 == new_ptr_10_value ? ghv_50 : _GEN_2070; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2072 = 8'h33 == new_ptr_10_value ? ghv_51 : _GEN_2071; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2073 = 8'h34 == new_ptr_10_value ? ghv_52 : _GEN_2072; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2074 = 8'h35 == new_ptr_10_value ? ghv_53 : _GEN_2073; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2075 = 8'h36 == new_ptr_10_value ? ghv_54 : _GEN_2074; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2076 = 8'h37 == new_ptr_10_value ? ghv_55 : _GEN_2075; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2077 = 8'h38 == new_ptr_10_value ? ghv_56 : _GEN_2076; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2078 = 8'h39 == new_ptr_10_value ? ghv_57 : _GEN_2077; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2079 = 8'h3a == new_ptr_10_value ? ghv_58 : _GEN_2078; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2080 = 8'h3b == new_ptr_10_value ? ghv_59 : _GEN_2079; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2081 = 8'h3c == new_ptr_10_value ? ghv_60 : _GEN_2080; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2082 = 8'h3d == new_ptr_10_value ? ghv_61 : _GEN_2081; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2083 = 8'h3e == new_ptr_10_value ? ghv_62 : _GEN_2082; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2084 = 8'h3f == new_ptr_10_value ? ghv_63 : _GEN_2083; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2085 = 8'h40 == new_ptr_10_value ? ghv_64 : _GEN_2084; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2086 = 8'h41 == new_ptr_10_value ? ghv_65 : _GEN_2085; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2087 = 8'h42 == new_ptr_10_value ? ghv_66 : _GEN_2086; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2088 = 8'h43 == new_ptr_10_value ? ghv_67 : _GEN_2087; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2089 = 8'h44 == new_ptr_10_value ? ghv_68 : _GEN_2088; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2090 = 8'h45 == new_ptr_10_value ? ghv_69 : _GEN_2089; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2091 = 8'h46 == new_ptr_10_value ? ghv_70 : _GEN_2090; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2092 = 8'h47 == new_ptr_10_value ? ghv_71 : _GEN_2091; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2093 = 8'h48 == new_ptr_10_value ? ghv_72 : _GEN_2092; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2094 = 8'h49 == new_ptr_10_value ? ghv_73 : _GEN_2093; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2095 = 8'h4a == new_ptr_10_value ? ghv_74 : _GEN_2094; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2096 = 8'h4b == new_ptr_10_value ? ghv_75 : _GEN_2095; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2097 = 8'h4c == new_ptr_10_value ? ghv_76 : _GEN_2096; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2098 = 8'h4d == new_ptr_10_value ? ghv_77 : _GEN_2097; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2099 = 8'h4e == new_ptr_10_value ? ghv_78 : _GEN_2098; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2100 = 8'h4f == new_ptr_10_value ? ghv_79 : _GEN_2099; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2101 = 8'h50 == new_ptr_10_value ? ghv_80 : _GEN_2100; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2102 = 8'h51 == new_ptr_10_value ? ghv_81 : _GEN_2101; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2103 = 8'h52 == new_ptr_10_value ? ghv_82 : _GEN_2102; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2104 = 8'h53 == new_ptr_10_value ? ghv_83 : _GEN_2103; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2105 = 8'h54 == new_ptr_10_value ? ghv_84 : _GEN_2104; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2106 = 8'h55 == new_ptr_10_value ? ghv_85 : _GEN_2105; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2107 = 8'h56 == new_ptr_10_value ? ghv_86 : _GEN_2106; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2108 = 8'h57 == new_ptr_10_value ? ghv_87 : _GEN_2107; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2109 = 8'h58 == new_ptr_10_value ? ghv_88 : _GEN_2108; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2110 = 8'h59 == new_ptr_10_value ? ghv_89 : _GEN_2109; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2111 = 8'h5a == new_ptr_10_value ? ghv_90 : _GEN_2110; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2112 = 8'h5b == new_ptr_10_value ? ghv_91 : _GEN_2111; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2113 = 8'h5c == new_ptr_10_value ? ghv_92 : _GEN_2112; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2114 = 8'h5d == new_ptr_10_value ? ghv_93 : _GEN_2113; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2115 = 8'h5e == new_ptr_10_value ? ghv_94 : _GEN_2114; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2116 = 8'h5f == new_ptr_10_value ? ghv_95 : _GEN_2115; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2117 = 8'h60 == new_ptr_10_value ? ghv_96 : _GEN_2116; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2118 = 8'h61 == new_ptr_10_value ? ghv_97 : _GEN_2117; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2119 = 8'h62 == new_ptr_10_value ? ghv_98 : _GEN_2118; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2120 = 8'h63 == new_ptr_10_value ? ghv_99 : _GEN_2119; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2121 = 8'h64 == new_ptr_10_value ? ghv_100 : _GEN_2120; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2122 = 8'h65 == new_ptr_10_value ? ghv_101 : _GEN_2121; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2123 = 8'h66 == new_ptr_10_value ? ghv_102 : _GEN_2122; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2124 = 8'h67 == new_ptr_10_value ? ghv_103 : _GEN_2123; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2125 = 8'h68 == new_ptr_10_value ? ghv_104 : _GEN_2124; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2126 = 8'h69 == new_ptr_10_value ? ghv_105 : _GEN_2125; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2127 = 8'h6a == new_ptr_10_value ? ghv_106 : _GEN_2126; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2128 = 8'h6b == new_ptr_10_value ? ghv_107 : _GEN_2127; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2129 = 8'h6c == new_ptr_10_value ? ghv_108 : _GEN_2128; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2130 = 8'h6d == new_ptr_10_value ? ghv_109 : _GEN_2129; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2131 = 8'h6e == new_ptr_10_value ? ghv_110 : _GEN_2130; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2132 = 8'h6f == new_ptr_10_value ? ghv_111 : _GEN_2131; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2133 = 8'h70 == new_ptr_10_value ? ghv_112 : _GEN_2132; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2134 = 8'h71 == new_ptr_10_value ? ghv_113 : _GEN_2133; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2135 = 8'h72 == new_ptr_10_value ? ghv_114 : _GEN_2134; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2136 = 8'h73 == new_ptr_10_value ? ghv_115 : _GEN_2135; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2137 = 8'h74 == new_ptr_10_value ? ghv_116 : _GEN_2136; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2138 = 8'h75 == new_ptr_10_value ? ghv_117 : _GEN_2137; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2139 = 8'h76 == new_ptr_10_value ? ghv_118 : _GEN_2138; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2140 = 8'h77 == new_ptr_10_value ? ghv_119 : _GEN_2139; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2141 = 8'h78 == new_ptr_10_value ? ghv_120 : _GEN_2140; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2142 = 8'h79 == new_ptr_10_value ? ghv_121 : _GEN_2141; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2143 = 8'h7a == new_ptr_10_value ? ghv_122 : _GEN_2142; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2144 = 8'h7b == new_ptr_10_value ? ghv_123 : _GEN_2143; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2145 = 8'h7c == new_ptr_10_value ? ghv_124 : _GEN_2144; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2146 = 8'h7d == new_ptr_10_value ? ghv_125 : _GEN_2145; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2147 = 8'h7e == new_ptr_10_value ? ghv_126 : _GEN_2146; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2148 = 8'h7f == new_ptr_10_value ? ghv_127 : _GEN_2147; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2149 = 8'h80 == new_ptr_10_value ? ghv_128 : _GEN_2148; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2150 = 8'h81 == new_ptr_10_value ? ghv_129 : _GEN_2149; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2151 = 8'h82 == new_ptr_10_value ? ghv_130 : _GEN_2150; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2152 = 8'h83 == new_ptr_10_value ? ghv_131 : _GEN_2151; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2153 = 8'h84 == new_ptr_10_value ? ghv_132 : _GEN_2152; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2154 = 8'h85 == new_ptr_10_value ? ghv_133 : _GEN_2153; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2155 = 8'h86 == new_ptr_10_value ? ghv_134 : _GEN_2154; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2156 = 8'h87 == new_ptr_10_value ? ghv_135 : _GEN_2155; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2157 = 8'h88 == new_ptr_10_value ? ghv_136 : _GEN_2156; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2158 = 8'h89 == new_ptr_10_value ? ghv_137 : _GEN_2157; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2159 = 8'h8a == new_ptr_10_value ? ghv_138 : _GEN_2158; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2160 = 8'h8b == new_ptr_10_value ? ghv_139 : _GEN_2159; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2161 = 8'h8c == new_ptr_10_value ? ghv_140 : _GEN_2160; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2162 = 8'h8d == new_ptr_10_value ? ghv_141 : _GEN_2161; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2163 = 8'h8e == new_ptr_10_value ? ghv_142 : _GEN_2162; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_1_value = _new_ptr_value_T_3[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_2166 = 8'h1 == new_ptr_1_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2167 = 8'h2 == new_ptr_1_value ? ghv_2 : _GEN_2166; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2168 = 8'h3 == new_ptr_1_value ? ghv_3 : _GEN_2167; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2169 = 8'h4 == new_ptr_1_value ? ghv_4 : _GEN_2168; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2170 = 8'h5 == new_ptr_1_value ? ghv_5 : _GEN_2169; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2171 = 8'h6 == new_ptr_1_value ? ghv_6 : _GEN_2170; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2172 = 8'h7 == new_ptr_1_value ? ghv_7 : _GEN_2171; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2173 = 8'h8 == new_ptr_1_value ? ghv_8 : _GEN_2172; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2174 = 8'h9 == new_ptr_1_value ? ghv_9 : _GEN_2173; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2175 = 8'ha == new_ptr_1_value ? ghv_10 : _GEN_2174; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2176 = 8'hb == new_ptr_1_value ? ghv_11 : _GEN_2175; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2177 = 8'hc == new_ptr_1_value ? ghv_12 : _GEN_2176; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2178 = 8'hd == new_ptr_1_value ? ghv_13 : _GEN_2177; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2179 = 8'he == new_ptr_1_value ? ghv_14 : _GEN_2178; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2180 = 8'hf == new_ptr_1_value ? ghv_15 : _GEN_2179; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2181 = 8'h10 == new_ptr_1_value ? ghv_16 : _GEN_2180; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2182 = 8'h11 == new_ptr_1_value ? ghv_17 : _GEN_2181; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2183 = 8'h12 == new_ptr_1_value ? ghv_18 : _GEN_2182; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2184 = 8'h13 == new_ptr_1_value ? ghv_19 : _GEN_2183; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2185 = 8'h14 == new_ptr_1_value ? ghv_20 : _GEN_2184; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2186 = 8'h15 == new_ptr_1_value ? ghv_21 : _GEN_2185; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2187 = 8'h16 == new_ptr_1_value ? ghv_22 : _GEN_2186; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2188 = 8'h17 == new_ptr_1_value ? ghv_23 : _GEN_2187; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2189 = 8'h18 == new_ptr_1_value ? ghv_24 : _GEN_2188; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2190 = 8'h19 == new_ptr_1_value ? ghv_25 : _GEN_2189; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2191 = 8'h1a == new_ptr_1_value ? ghv_26 : _GEN_2190; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2192 = 8'h1b == new_ptr_1_value ? ghv_27 : _GEN_2191; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2193 = 8'h1c == new_ptr_1_value ? ghv_28 : _GEN_2192; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2194 = 8'h1d == new_ptr_1_value ? ghv_29 : _GEN_2193; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2195 = 8'h1e == new_ptr_1_value ? ghv_30 : _GEN_2194; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2196 = 8'h1f == new_ptr_1_value ? ghv_31 : _GEN_2195; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2197 = 8'h20 == new_ptr_1_value ? ghv_32 : _GEN_2196; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2198 = 8'h21 == new_ptr_1_value ? ghv_33 : _GEN_2197; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2199 = 8'h22 == new_ptr_1_value ? ghv_34 : _GEN_2198; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2200 = 8'h23 == new_ptr_1_value ? ghv_35 : _GEN_2199; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2201 = 8'h24 == new_ptr_1_value ? ghv_36 : _GEN_2200; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2202 = 8'h25 == new_ptr_1_value ? ghv_37 : _GEN_2201; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2203 = 8'h26 == new_ptr_1_value ? ghv_38 : _GEN_2202; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2204 = 8'h27 == new_ptr_1_value ? ghv_39 : _GEN_2203; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2205 = 8'h28 == new_ptr_1_value ? ghv_40 : _GEN_2204; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2206 = 8'h29 == new_ptr_1_value ? ghv_41 : _GEN_2205; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2207 = 8'h2a == new_ptr_1_value ? ghv_42 : _GEN_2206; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2208 = 8'h2b == new_ptr_1_value ? ghv_43 : _GEN_2207; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2209 = 8'h2c == new_ptr_1_value ? ghv_44 : _GEN_2208; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2210 = 8'h2d == new_ptr_1_value ? ghv_45 : _GEN_2209; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2211 = 8'h2e == new_ptr_1_value ? ghv_46 : _GEN_2210; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2212 = 8'h2f == new_ptr_1_value ? ghv_47 : _GEN_2211; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2213 = 8'h30 == new_ptr_1_value ? ghv_48 : _GEN_2212; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2214 = 8'h31 == new_ptr_1_value ? ghv_49 : _GEN_2213; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2215 = 8'h32 == new_ptr_1_value ? ghv_50 : _GEN_2214; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2216 = 8'h33 == new_ptr_1_value ? ghv_51 : _GEN_2215; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2217 = 8'h34 == new_ptr_1_value ? ghv_52 : _GEN_2216; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2218 = 8'h35 == new_ptr_1_value ? ghv_53 : _GEN_2217; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2219 = 8'h36 == new_ptr_1_value ? ghv_54 : _GEN_2218; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2220 = 8'h37 == new_ptr_1_value ? ghv_55 : _GEN_2219; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2221 = 8'h38 == new_ptr_1_value ? ghv_56 : _GEN_2220; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2222 = 8'h39 == new_ptr_1_value ? ghv_57 : _GEN_2221; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2223 = 8'h3a == new_ptr_1_value ? ghv_58 : _GEN_2222; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2224 = 8'h3b == new_ptr_1_value ? ghv_59 : _GEN_2223; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2225 = 8'h3c == new_ptr_1_value ? ghv_60 : _GEN_2224; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2226 = 8'h3d == new_ptr_1_value ? ghv_61 : _GEN_2225; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2227 = 8'h3e == new_ptr_1_value ? ghv_62 : _GEN_2226; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2228 = 8'h3f == new_ptr_1_value ? ghv_63 : _GEN_2227; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2229 = 8'h40 == new_ptr_1_value ? ghv_64 : _GEN_2228; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2230 = 8'h41 == new_ptr_1_value ? ghv_65 : _GEN_2229; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2231 = 8'h42 == new_ptr_1_value ? ghv_66 : _GEN_2230; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2232 = 8'h43 == new_ptr_1_value ? ghv_67 : _GEN_2231; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2233 = 8'h44 == new_ptr_1_value ? ghv_68 : _GEN_2232; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2234 = 8'h45 == new_ptr_1_value ? ghv_69 : _GEN_2233; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2235 = 8'h46 == new_ptr_1_value ? ghv_70 : _GEN_2234; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2236 = 8'h47 == new_ptr_1_value ? ghv_71 : _GEN_2235; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2237 = 8'h48 == new_ptr_1_value ? ghv_72 : _GEN_2236; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2238 = 8'h49 == new_ptr_1_value ? ghv_73 : _GEN_2237; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2239 = 8'h4a == new_ptr_1_value ? ghv_74 : _GEN_2238; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2240 = 8'h4b == new_ptr_1_value ? ghv_75 : _GEN_2239; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2241 = 8'h4c == new_ptr_1_value ? ghv_76 : _GEN_2240; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2242 = 8'h4d == new_ptr_1_value ? ghv_77 : _GEN_2241; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2243 = 8'h4e == new_ptr_1_value ? ghv_78 : _GEN_2242; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2244 = 8'h4f == new_ptr_1_value ? ghv_79 : _GEN_2243; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2245 = 8'h50 == new_ptr_1_value ? ghv_80 : _GEN_2244; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2246 = 8'h51 == new_ptr_1_value ? ghv_81 : _GEN_2245; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2247 = 8'h52 == new_ptr_1_value ? ghv_82 : _GEN_2246; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2248 = 8'h53 == new_ptr_1_value ? ghv_83 : _GEN_2247; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2249 = 8'h54 == new_ptr_1_value ? ghv_84 : _GEN_2248; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2250 = 8'h55 == new_ptr_1_value ? ghv_85 : _GEN_2249; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2251 = 8'h56 == new_ptr_1_value ? ghv_86 : _GEN_2250; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2252 = 8'h57 == new_ptr_1_value ? ghv_87 : _GEN_2251; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2253 = 8'h58 == new_ptr_1_value ? ghv_88 : _GEN_2252; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2254 = 8'h59 == new_ptr_1_value ? ghv_89 : _GEN_2253; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2255 = 8'h5a == new_ptr_1_value ? ghv_90 : _GEN_2254; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2256 = 8'h5b == new_ptr_1_value ? ghv_91 : _GEN_2255; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2257 = 8'h5c == new_ptr_1_value ? ghv_92 : _GEN_2256; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2258 = 8'h5d == new_ptr_1_value ? ghv_93 : _GEN_2257; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2259 = 8'h5e == new_ptr_1_value ? ghv_94 : _GEN_2258; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2260 = 8'h5f == new_ptr_1_value ? ghv_95 : _GEN_2259; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2261 = 8'h60 == new_ptr_1_value ? ghv_96 : _GEN_2260; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2262 = 8'h61 == new_ptr_1_value ? ghv_97 : _GEN_2261; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2263 = 8'h62 == new_ptr_1_value ? ghv_98 : _GEN_2262; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2264 = 8'h63 == new_ptr_1_value ? ghv_99 : _GEN_2263; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2265 = 8'h64 == new_ptr_1_value ? ghv_100 : _GEN_2264; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2266 = 8'h65 == new_ptr_1_value ? ghv_101 : _GEN_2265; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2267 = 8'h66 == new_ptr_1_value ? ghv_102 : _GEN_2266; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2268 = 8'h67 == new_ptr_1_value ? ghv_103 : _GEN_2267; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2269 = 8'h68 == new_ptr_1_value ? ghv_104 : _GEN_2268; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2270 = 8'h69 == new_ptr_1_value ? ghv_105 : _GEN_2269; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2271 = 8'h6a == new_ptr_1_value ? ghv_106 : _GEN_2270; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2272 = 8'h6b == new_ptr_1_value ? ghv_107 : _GEN_2271; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2273 = 8'h6c == new_ptr_1_value ? ghv_108 : _GEN_2272; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2274 = 8'h6d == new_ptr_1_value ? ghv_109 : _GEN_2273; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2275 = 8'h6e == new_ptr_1_value ? ghv_110 : _GEN_2274; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2276 = 8'h6f == new_ptr_1_value ? ghv_111 : _GEN_2275; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2277 = 8'h70 == new_ptr_1_value ? ghv_112 : _GEN_2276; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2278 = 8'h71 == new_ptr_1_value ? ghv_113 : _GEN_2277; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2279 = 8'h72 == new_ptr_1_value ? ghv_114 : _GEN_2278; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2280 = 8'h73 == new_ptr_1_value ? ghv_115 : _GEN_2279; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2281 = 8'h74 == new_ptr_1_value ? ghv_116 : _GEN_2280; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2282 = 8'h75 == new_ptr_1_value ? ghv_117 : _GEN_2281; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2283 = 8'h76 == new_ptr_1_value ? ghv_118 : _GEN_2282; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2284 = 8'h77 == new_ptr_1_value ? ghv_119 : _GEN_2283; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2285 = 8'h78 == new_ptr_1_value ? ghv_120 : _GEN_2284; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2286 = 8'h79 == new_ptr_1_value ? ghv_121 : _GEN_2285; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2287 = 8'h7a == new_ptr_1_value ? ghv_122 : _GEN_2286; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2288 = 8'h7b == new_ptr_1_value ? ghv_123 : _GEN_2287; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2289 = 8'h7c == new_ptr_1_value ? ghv_124 : _GEN_2288; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2290 = 8'h7d == new_ptr_1_value ? ghv_125 : _GEN_2289; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2291 = 8'h7e == new_ptr_1_value ? ghv_126 : _GEN_2290; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2292 = 8'h7f == new_ptr_1_value ? ghv_127 : _GEN_2291; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2293 = 8'h80 == new_ptr_1_value ? ghv_128 : _GEN_2292; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2294 = 8'h81 == new_ptr_1_value ? ghv_129 : _GEN_2293; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2295 = 8'h82 == new_ptr_1_value ? ghv_130 : _GEN_2294; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2296 = 8'h83 == new_ptr_1_value ? ghv_131 : _GEN_2295; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2297 = 8'h84 == new_ptr_1_value ? ghv_132 : _GEN_2296; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2298 = 8'h85 == new_ptr_1_value ? ghv_133 : _GEN_2297; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2299 = 8'h86 == new_ptr_1_value ? ghv_134 : _GEN_2298; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2300 = 8'h87 == new_ptr_1_value ? ghv_135 : _GEN_2299; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2301 = 8'h88 == new_ptr_1_value ? ghv_136 : _GEN_2300; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2302 = 8'h89 == new_ptr_1_value ? ghv_137 : _GEN_2301; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2303 = 8'h8a == new_ptr_1_value ? ghv_138 : _GEN_2302; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2304 = 8'h8b == new_ptr_1_value ? ghv_139 : _GEN_2303; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2305 = 8'h8c == new_ptr_1_value ? ghv_140 : _GEN_2304; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2306 = 8'h8d == new_ptr_1_value ? ghv_141 : _GEN_2305; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2307 = 8'h8e == new_ptr_1_value ? ghv_142 : _GEN_2306; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_18_value = _new_ptr_value_T_37[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_2310 = 8'h1 == new_ptr_18_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2311 = 8'h2 == new_ptr_18_value ? ghv_2 : _GEN_2310; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2312 = 8'h3 == new_ptr_18_value ? ghv_3 : _GEN_2311; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2313 = 8'h4 == new_ptr_18_value ? ghv_4 : _GEN_2312; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2314 = 8'h5 == new_ptr_18_value ? ghv_5 : _GEN_2313; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2315 = 8'h6 == new_ptr_18_value ? ghv_6 : _GEN_2314; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2316 = 8'h7 == new_ptr_18_value ? ghv_7 : _GEN_2315; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2317 = 8'h8 == new_ptr_18_value ? ghv_8 : _GEN_2316; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2318 = 8'h9 == new_ptr_18_value ? ghv_9 : _GEN_2317; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2319 = 8'ha == new_ptr_18_value ? ghv_10 : _GEN_2318; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2320 = 8'hb == new_ptr_18_value ? ghv_11 : _GEN_2319; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2321 = 8'hc == new_ptr_18_value ? ghv_12 : _GEN_2320; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2322 = 8'hd == new_ptr_18_value ? ghv_13 : _GEN_2321; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2323 = 8'he == new_ptr_18_value ? ghv_14 : _GEN_2322; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2324 = 8'hf == new_ptr_18_value ? ghv_15 : _GEN_2323; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2325 = 8'h10 == new_ptr_18_value ? ghv_16 : _GEN_2324; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2326 = 8'h11 == new_ptr_18_value ? ghv_17 : _GEN_2325; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2327 = 8'h12 == new_ptr_18_value ? ghv_18 : _GEN_2326; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2328 = 8'h13 == new_ptr_18_value ? ghv_19 : _GEN_2327; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2329 = 8'h14 == new_ptr_18_value ? ghv_20 : _GEN_2328; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2330 = 8'h15 == new_ptr_18_value ? ghv_21 : _GEN_2329; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2331 = 8'h16 == new_ptr_18_value ? ghv_22 : _GEN_2330; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2332 = 8'h17 == new_ptr_18_value ? ghv_23 : _GEN_2331; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2333 = 8'h18 == new_ptr_18_value ? ghv_24 : _GEN_2332; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2334 = 8'h19 == new_ptr_18_value ? ghv_25 : _GEN_2333; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2335 = 8'h1a == new_ptr_18_value ? ghv_26 : _GEN_2334; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2336 = 8'h1b == new_ptr_18_value ? ghv_27 : _GEN_2335; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2337 = 8'h1c == new_ptr_18_value ? ghv_28 : _GEN_2336; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2338 = 8'h1d == new_ptr_18_value ? ghv_29 : _GEN_2337; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2339 = 8'h1e == new_ptr_18_value ? ghv_30 : _GEN_2338; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2340 = 8'h1f == new_ptr_18_value ? ghv_31 : _GEN_2339; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2341 = 8'h20 == new_ptr_18_value ? ghv_32 : _GEN_2340; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2342 = 8'h21 == new_ptr_18_value ? ghv_33 : _GEN_2341; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2343 = 8'h22 == new_ptr_18_value ? ghv_34 : _GEN_2342; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2344 = 8'h23 == new_ptr_18_value ? ghv_35 : _GEN_2343; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2345 = 8'h24 == new_ptr_18_value ? ghv_36 : _GEN_2344; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2346 = 8'h25 == new_ptr_18_value ? ghv_37 : _GEN_2345; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2347 = 8'h26 == new_ptr_18_value ? ghv_38 : _GEN_2346; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2348 = 8'h27 == new_ptr_18_value ? ghv_39 : _GEN_2347; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2349 = 8'h28 == new_ptr_18_value ? ghv_40 : _GEN_2348; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2350 = 8'h29 == new_ptr_18_value ? ghv_41 : _GEN_2349; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2351 = 8'h2a == new_ptr_18_value ? ghv_42 : _GEN_2350; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2352 = 8'h2b == new_ptr_18_value ? ghv_43 : _GEN_2351; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2353 = 8'h2c == new_ptr_18_value ? ghv_44 : _GEN_2352; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2354 = 8'h2d == new_ptr_18_value ? ghv_45 : _GEN_2353; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2355 = 8'h2e == new_ptr_18_value ? ghv_46 : _GEN_2354; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2356 = 8'h2f == new_ptr_18_value ? ghv_47 : _GEN_2355; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2357 = 8'h30 == new_ptr_18_value ? ghv_48 : _GEN_2356; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2358 = 8'h31 == new_ptr_18_value ? ghv_49 : _GEN_2357; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2359 = 8'h32 == new_ptr_18_value ? ghv_50 : _GEN_2358; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2360 = 8'h33 == new_ptr_18_value ? ghv_51 : _GEN_2359; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2361 = 8'h34 == new_ptr_18_value ? ghv_52 : _GEN_2360; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2362 = 8'h35 == new_ptr_18_value ? ghv_53 : _GEN_2361; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2363 = 8'h36 == new_ptr_18_value ? ghv_54 : _GEN_2362; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2364 = 8'h37 == new_ptr_18_value ? ghv_55 : _GEN_2363; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2365 = 8'h38 == new_ptr_18_value ? ghv_56 : _GEN_2364; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2366 = 8'h39 == new_ptr_18_value ? ghv_57 : _GEN_2365; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2367 = 8'h3a == new_ptr_18_value ? ghv_58 : _GEN_2366; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2368 = 8'h3b == new_ptr_18_value ? ghv_59 : _GEN_2367; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2369 = 8'h3c == new_ptr_18_value ? ghv_60 : _GEN_2368; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2370 = 8'h3d == new_ptr_18_value ? ghv_61 : _GEN_2369; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2371 = 8'h3e == new_ptr_18_value ? ghv_62 : _GEN_2370; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2372 = 8'h3f == new_ptr_18_value ? ghv_63 : _GEN_2371; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2373 = 8'h40 == new_ptr_18_value ? ghv_64 : _GEN_2372; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2374 = 8'h41 == new_ptr_18_value ? ghv_65 : _GEN_2373; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2375 = 8'h42 == new_ptr_18_value ? ghv_66 : _GEN_2374; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2376 = 8'h43 == new_ptr_18_value ? ghv_67 : _GEN_2375; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2377 = 8'h44 == new_ptr_18_value ? ghv_68 : _GEN_2376; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2378 = 8'h45 == new_ptr_18_value ? ghv_69 : _GEN_2377; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2379 = 8'h46 == new_ptr_18_value ? ghv_70 : _GEN_2378; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2380 = 8'h47 == new_ptr_18_value ? ghv_71 : _GEN_2379; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2381 = 8'h48 == new_ptr_18_value ? ghv_72 : _GEN_2380; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2382 = 8'h49 == new_ptr_18_value ? ghv_73 : _GEN_2381; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2383 = 8'h4a == new_ptr_18_value ? ghv_74 : _GEN_2382; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2384 = 8'h4b == new_ptr_18_value ? ghv_75 : _GEN_2383; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2385 = 8'h4c == new_ptr_18_value ? ghv_76 : _GEN_2384; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2386 = 8'h4d == new_ptr_18_value ? ghv_77 : _GEN_2385; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2387 = 8'h4e == new_ptr_18_value ? ghv_78 : _GEN_2386; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2388 = 8'h4f == new_ptr_18_value ? ghv_79 : _GEN_2387; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2389 = 8'h50 == new_ptr_18_value ? ghv_80 : _GEN_2388; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2390 = 8'h51 == new_ptr_18_value ? ghv_81 : _GEN_2389; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2391 = 8'h52 == new_ptr_18_value ? ghv_82 : _GEN_2390; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2392 = 8'h53 == new_ptr_18_value ? ghv_83 : _GEN_2391; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2393 = 8'h54 == new_ptr_18_value ? ghv_84 : _GEN_2392; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2394 = 8'h55 == new_ptr_18_value ? ghv_85 : _GEN_2393; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2395 = 8'h56 == new_ptr_18_value ? ghv_86 : _GEN_2394; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2396 = 8'h57 == new_ptr_18_value ? ghv_87 : _GEN_2395; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2397 = 8'h58 == new_ptr_18_value ? ghv_88 : _GEN_2396; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2398 = 8'h59 == new_ptr_18_value ? ghv_89 : _GEN_2397; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2399 = 8'h5a == new_ptr_18_value ? ghv_90 : _GEN_2398; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2400 = 8'h5b == new_ptr_18_value ? ghv_91 : _GEN_2399; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2401 = 8'h5c == new_ptr_18_value ? ghv_92 : _GEN_2400; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2402 = 8'h5d == new_ptr_18_value ? ghv_93 : _GEN_2401; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2403 = 8'h5e == new_ptr_18_value ? ghv_94 : _GEN_2402; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2404 = 8'h5f == new_ptr_18_value ? ghv_95 : _GEN_2403; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2405 = 8'h60 == new_ptr_18_value ? ghv_96 : _GEN_2404; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2406 = 8'h61 == new_ptr_18_value ? ghv_97 : _GEN_2405; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2407 = 8'h62 == new_ptr_18_value ? ghv_98 : _GEN_2406; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2408 = 8'h63 == new_ptr_18_value ? ghv_99 : _GEN_2407; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2409 = 8'h64 == new_ptr_18_value ? ghv_100 : _GEN_2408; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2410 = 8'h65 == new_ptr_18_value ? ghv_101 : _GEN_2409; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2411 = 8'h66 == new_ptr_18_value ? ghv_102 : _GEN_2410; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2412 = 8'h67 == new_ptr_18_value ? ghv_103 : _GEN_2411; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2413 = 8'h68 == new_ptr_18_value ? ghv_104 : _GEN_2412; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2414 = 8'h69 == new_ptr_18_value ? ghv_105 : _GEN_2413; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2415 = 8'h6a == new_ptr_18_value ? ghv_106 : _GEN_2414; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2416 = 8'h6b == new_ptr_18_value ? ghv_107 : _GEN_2415; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2417 = 8'h6c == new_ptr_18_value ? ghv_108 : _GEN_2416; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2418 = 8'h6d == new_ptr_18_value ? ghv_109 : _GEN_2417; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2419 = 8'h6e == new_ptr_18_value ? ghv_110 : _GEN_2418; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2420 = 8'h6f == new_ptr_18_value ? ghv_111 : _GEN_2419; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2421 = 8'h70 == new_ptr_18_value ? ghv_112 : _GEN_2420; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2422 = 8'h71 == new_ptr_18_value ? ghv_113 : _GEN_2421; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2423 = 8'h72 == new_ptr_18_value ? ghv_114 : _GEN_2422; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2424 = 8'h73 == new_ptr_18_value ? ghv_115 : _GEN_2423; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2425 = 8'h74 == new_ptr_18_value ? ghv_116 : _GEN_2424; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2426 = 8'h75 == new_ptr_18_value ? ghv_117 : _GEN_2425; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2427 = 8'h76 == new_ptr_18_value ? ghv_118 : _GEN_2426; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2428 = 8'h77 == new_ptr_18_value ? ghv_119 : _GEN_2427; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2429 = 8'h78 == new_ptr_18_value ? ghv_120 : _GEN_2428; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2430 = 8'h79 == new_ptr_18_value ? ghv_121 : _GEN_2429; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2431 = 8'h7a == new_ptr_18_value ? ghv_122 : _GEN_2430; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2432 = 8'h7b == new_ptr_18_value ? ghv_123 : _GEN_2431; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2433 = 8'h7c == new_ptr_18_value ? ghv_124 : _GEN_2432; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2434 = 8'h7d == new_ptr_18_value ? ghv_125 : _GEN_2433; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2435 = 8'h7e == new_ptr_18_value ? ghv_126 : _GEN_2434; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2436 = 8'h7f == new_ptr_18_value ? ghv_127 : _GEN_2435; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2437 = 8'h80 == new_ptr_18_value ? ghv_128 : _GEN_2436; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2438 = 8'h81 == new_ptr_18_value ? ghv_129 : _GEN_2437; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2439 = 8'h82 == new_ptr_18_value ? ghv_130 : _GEN_2438; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2440 = 8'h83 == new_ptr_18_value ? ghv_131 : _GEN_2439; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2441 = 8'h84 == new_ptr_18_value ? ghv_132 : _GEN_2440; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2442 = 8'h85 == new_ptr_18_value ? ghv_133 : _GEN_2441; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2443 = 8'h86 == new_ptr_18_value ? ghv_134 : _GEN_2442; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2444 = 8'h87 == new_ptr_18_value ? ghv_135 : _GEN_2443; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2445 = 8'h88 == new_ptr_18_value ? ghv_136 : _GEN_2444; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2446 = 8'h89 == new_ptr_18_value ? ghv_137 : _GEN_2445; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2447 = 8'h8a == new_ptr_18_value ? ghv_138 : _GEN_2446; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2448 = 8'h8b == new_ptr_18_value ? ghv_139 : _GEN_2447; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2449 = 8'h8c == new_ptr_18_value ? ghv_140 : _GEN_2448; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2450 = 8'h8d == new_ptr_18_value ? ghv_141 : _GEN_2449; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2451 = 8'h8e == new_ptr_18_value ? ghv_142 : _GEN_2450; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_11_value = _new_ptr_value_T_23[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_2454 = 8'h1 == new_ptr_11_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2455 = 8'h2 == new_ptr_11_value ? ghv_2 : _GEN_2454; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2456 = 8'h3 == new_ptr_11_value ? ghv_3 : _GEN_2455; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2457 = 8'h4 == new_ptr_11_value ? ghv_4 : _GEN_2456; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2458 = 8'h5 == new_ptr_11_value ? ghv_5 : _GEN_2457; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2459 = 8'h6 == new_ptr_11_value ? ghv_6 : _GEN_2458; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2460 = 8'h7 == new_ptr_11_value ? ghv_7 : _GEN_2459; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2461 = 8'h8 == new_ptr_11_value ? ghv_8 : _GEN_2460; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2462 = 8'h9 == new_ptr_11_value ? ghv_9 : _GEN_2461; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2463 = 8'ha == new_ptr_11_value ? ghv_10 : _GEN_2462; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2464 = 8'hb == new_ptr_11_value ? ghv_11 : _GEN_2463; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2465 = 8'hc == new_ptr_11_value ? ghv_12 : _GEN_2464; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2466 = 8'hd == new_ptr_11_value ? ghv_13 : _GEN_2465; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2467 = 8'he == new_ptr_11_value ? ghv_14 : _GEN_2466; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2468 = 8'hf == new_ptr_11_value ? ghv_15 : _GEN_2467; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2469 = 8'h10 == new_ptr_11_value ? ghv_16 : _GEN_2468; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2470 = 8'h11 == new_ptr_11_value ? ghv_17 : _GEN_2469; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2471 = 8'h12 == new_ptr_11_value ? ghv_18 : _GEN_2470; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2472 = 8'h13 == new_ptr_11_value ? ghv_19 : _GEN_2471; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2473 = 8'h14 == new_ptr_11_value ? ghv_20 : _GEN_2472; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2474 = 8'h15 == new_ptr_11_value ? ghv_21 : _GEN_2473; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2475 = 8'h16 == new_ptr_11_value ? ghv_22 : _GEN_2474; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2476 = 8'h17 == new_ptr_11_value ? ghv_23 : _GEN_2475; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2477 = 8'h18 == new_ptr_11_value ? ghv_24 : _GEN_2476; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2478 = 8'h19 == new_ptr_11_value ? ghv_25 : _GEN_2477; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2479 = 8'h1a == new_ptr_11_value ? ghv_26 : _GEN_2478; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2480 = 8'h1b == new_ptr_11_value ? ghv_27 : _GEN_2479; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2481 = 8'h1c == new_ptr_11_value ? ghv_28 : _GEN_2480; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2482 = 8'h1d == new_ptr_11_value ? ghv_29 : _GEN_2481; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2483 = 8'h1e == new_ptr_11_value ? ghv_30 : _GEN_2482; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2484 = 8'h1f == new_ptr_11_value ? ghv_31 : _GEN_2483; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2485 = 8'h20 == new_ptr_11_value ? ghv_32 : _GEN_2484; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2486 = 8'h21 == new_ptr_11_value ? ghv_33 : _GEN_2485; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2487 = 8'h22 == new_ptr_11_value ? ghv_34 : _GEN_2486; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2488 = 8'h23 == new_ptr_11_value ? ghv_35 : _GEN_2487; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2489 = 8'h24 == new_ptr_11_value ? ghv_36 : _GEN_2488; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2490 = 8'h25 == new_ptr_11_value ? ghv_37 : _GEN_2489; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2491 = 8'h26 == new_ptr_11_value ? ghv_38 : _GEN_2490; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2492 = 8'h27 == new_ptr_11_value ? ghv_39 : _GEN_2491; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2493 = 8'h28 == new_ptr_11_value ? ghv_40 : _GEN_2492; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2494 = 8'h29 == new_ptr_11_value ? ghv_41 : _GEN_2493; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2495 = 8'h2a == new_ptr_11_value ? ghv_42 : _GEN_2494; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2496 = 8'h2b == new_ptr_11_value ? ghv_43 : _GEN_2495; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2497 = 8'h2c == new_ptr_11_value ? ghv_44 : _GEN_2496; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2498 = 8'h2d == new_ptr_11_value ? ghv_45 : _GEN_2497; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2499 = 8'h2e == new_ptr_11_value ? ghv_46 : _GEN_2498; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2500 = 8'h2f == new_ptr_11_value ? ghv_47 : _GEN_2499; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2501 = 8'h30 == new_ptr_11_value ? ghv_48 : _GEN_2500; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2502 = 8'h31 == new_ptr_11_value ? ghv_49 : _GEN_2501; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2503 = 8'h32 == new_ptr_11_value ? ghv_50 : _GEN_2502; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2504 = 8'h33 == new_ptr_11_value ? ghv_51 : _GEN_2503; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2505 = 8'h34 == new_ptr_11_value ? ghv_52 : _GEN_2504; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2506 = 8'h35 == new_ptr_11_value ? ghv_53 : _GEN_2505; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2507 = 8'h36 == new_ptr_11_value ? ghv_54 : _GEN_2506; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2508 = 8'h37 == new_ptr_11_value ? ghv_55 : _GEN_2507; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2509 = 8'h38 == new_ptr_11_value ? ghv_56 : _GEN_2508; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2510 = 8'h39 == new_ptr_11_value ? ghv_57 : _GEN_2509; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2511 = 8'h3a == new_ptr_11_value ? ghv_58 : _GEN_2510; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2512 = 8'h3b == new_ptr_11_value ? ghv_59 : _GEN_2511; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2513 = 8'h3c == new_ptr_11_value ? ghv_60 : _GEN_2512; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2514 = 8'h3d == new_ptr_11_value ? ghv_61 : _GEN_2513; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2515 = 8'h3e == new_ptr_11_value ? ghv_62 : _GEN_2514; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2516 = 8'h3f == new_ptr_11_value ? ghv_63 : _GEN_2515; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2517 = 8'h40 == new_ptr_11_value ? ghv_64 : _GEN_2516; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2518 = 8'h41 == new_ptr_11_value ? ghv_65 : _GEN_2517; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2519 = 8'h42 == new_ptr_11_value ? ghv_66 : _GEN_2518; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2520 = 8'h43 == new_ptr_11_value ? ghv_67 : _GEN_2519; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2521 = 8'h44 == new_ptr_11_value ? ghv_68 : _GEN_2520; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2522 = 8'h45 == new_ptr_11_value ? ghv_69 : _GEN_2521; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2523 = 8'h46 == new_ptr_11_value ? ghv_70 : _GEN_2522; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2524 = 8'h47 == new_ptr_11_value ? ghv_71 : _GEN_2523; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2525 = 8'h48 == new_ptr_11_value ? ghv_72 : _GEN_2524; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2526 = 8'h49 == new_ptr_11_value ? ghv_73 : _GEN_2525; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2527 = 8'h4a == new_ptr_11_value ? ghv_74 : _GEN_2526; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2528 = 8'h4b == new_ptr_11_value ? ghv_75 : _GEN_2527; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2529 = 8'h4c == new_ptr_11_value ? ghv_76 : _GEN_2528; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2530 = 8'h4d == new_ptr_11_value ? ghv_77 : _GEN_2529; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2531 = 8'h4e == new_ptr_11_value ? ghv_78 : _GEN_2530; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2532 = 8'h4f == new_ptr_11_value ? ghv_79 : _GEN_2531; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2533 = 8'h50 == new_ptr_11_value ? ghv_80 : _GEN_2532; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2534 = 8'h51 == new_ptr_11_value ? ghv_81 : _GEN_2533; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2535 = 8'h52 == new_ptr_11_value ? ghv_82 : _GEN_2534; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2536 = 8'h53 == new_ptr_11_value ? ghv_83 : _GEN_2535; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2537 = 8'h54 == new_ptr_11_value ? ghv_84 : _GEN_2536; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2538 = 8'h55 == new_ptr_11_value ? ghv_85 : _GEN_2537; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2539 = 8'h56 == new_ptr_11_value ? ghv_86 : _GEN_2538; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2540 = 8'h57 == new_ptr_11_value ? ghv_87 : _GEN_2539; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2541 = 8'h58 == new_ptr_11_value ? ghv_88 : _GEN_2540; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2542 = 8'h59 == new_ptr_11_value ? ghv_89 : _GEN_2541; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2543 = 8'h5a == new_ptr_11_value ? ghv_90 : _GEN_2542; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2544 = 8'h5b == new_ptr_11_value ? ghv_91 : _GEN_2543; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2545 = 8'h5c == new_ptr_11_value ? ghv_92 : _GEN_2544; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2546 = 8'h5d == new_ptr_11_value ? ghv_93 : _GEN_2545; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2547 = 8'h5e == new_ptr_11_value ? ghv_94 : _GEN_2546; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2548 = 8'h5f == new_ptr_11_value ? ghv_95 : _GEN_2547; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2549 = 8'h60 == new_ptr_11_value ? ghv_96 : _GEN_2548; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2550 = 8'h61 == new_ptr_11_value ? ghv_97 : _GEN_2549; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2551 = 8'h62 == new_ptr_11_value ? ghv_98 : _GEN_2550; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2552 = 8'h63 == new_ptr_11_value ? ghv_99 : _GEN_2551; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2553 = 8'h64 == new_ptr_11_value ? ghv_100 : _GEN_2552; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2554 = 8'h65 == new_ptr_11_value ? ghv_101 : _GEN_2553; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2555 = 8'h66 == new_ptr_11_value ? ghv_102 : _GEN_2554; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2556 = 8'h67 == new_ptr_11_value ? ghv_103 : _GEN_2555; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2557 = 8'h68 == new_ptr_11_value ? ghv_104 : _GEN_2556; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2558 = 8'h69 == new_ptr_11_value ? ghv_105 : _GEN_2557; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2559 = 8'h6a == new_ptr_11_value ? ghv_106 : _GEN_2558; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2560 = 8'h6b == new_ptr_11_value ? ghv_107 : _GEN_2559; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2561 = 8'h6c == new_ptr_11_value ? ghv_108 : _GEN_2560; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2562 = 8'h6d == new_ptr_11_value ? ghv_109 : _GEN_2561; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2563 = 8'h6e == new_ptr_11_value ? ghv_110 : _GEN_2562; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2564 = 8'h6f == new_ptr_11_value ? ghv_111 : _GEN_2563; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2565 = 8'h70 == new_ptr_11_value ? ghv_112 : _GEN_2564; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2566 = 8'h71 == new_ptr_11_value ? ghv_113 : _GEN_2565; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2567 = 8'h72 == new_ptr_11_value ? ghv_114 : _GEN_2566; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2568 = 8'h73 == new_ptr_11_value ? ghv_115 : _GEN_2567; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2569 = 8'h74 == new_ptr_11_value ? ghv_116 : _GEN_2568; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2570 = 8'h75 == new_ptr_11_value ? ghv_117 : _GEN_2569; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2571 = 8'h76 == new_ptr_11_value ? ghv_118 : _GEN_2570; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2572 = 8'h77 == new_ptr_11_value ? ghv_119 : _GEN_2571; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2573 = 8'h78 == new_ptr_11_value ? ghv_120 : _GEN_2572; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2574 = 8'h79 == new_ptr_11_value ? ghv_121 : _GEN_2573; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2575 = 8'h7a == new_ptr_11_value ? ghv_122 : _GEN_2574; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2576 = 8'h7b == new_ptr_11_value ? ghv_123 : _GEN_2575; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2577 = 8'h7c == new_ptr_11_value ? ghv_124 : _GEN_2576; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2578 = 8'h7d == new_ptr_11_value ? ghv_125 : _GEN_2577; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2579 = 8'h7e == new_ptr_11_value ? ghv_126 : _GEN_2578; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2580 = 8'h7f == new_ptr_11_value ? ghv_127 : _GEN_2579; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2581 = 8'h80 == new_ptr_11_value ? ghv_128 : _GEN_2580; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2582 = 8'h81 == new_ptr_11_value ? ghv_129 : _GEN_2581; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2583 = 8'h82 == new_ptr_11_value ? ghv_130 : _GEN_2582; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2584 = 8'h83 == new_ptr_11_value ? ghv_131 : _GEN_2583; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2585 = 8'h84 == new_ptr_11_value ? ghv_132 : _GEN_2584; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2586 = 8'h85 == new_ptr_11_value ? ghv_133 : _GEN_2585; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2587 = 8'h86 == new_ptr_11_value ? ghv_134 : _GEN_2586; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2588 = 8'h87 == new_ptr_11_value ? ghv_135 : _GEN_2587; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2589 = 8'h88 == new_ptr_11_value ? ghv_136 : _GEN_2588; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2590 = 8'h89 == new_ptr_11_value ? ghv_137 : _GEN_2589; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2591 = 8'h8a == new_ptr_11_value ? ghv_138 : _GEN_2590; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2592 = 8'h8b == new_ptr_11_value ? ghv_139 : _GEN_2591; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2593 = 8'h8c == new_ptr_11_value ? ghv_140 : _GEN_2592; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2594 = 8'h8d == new_ptr_11_value ? ghv_141 : _GEN_2593; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2595 = 8'h8e == new_ptr_11_value ? ghv_142 : _GEN_2594; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_7_value = _new_ptr_value_T_15[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_2598 = 8'h1 == new_ptr_7_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2599 = 8'h2 == new_ptr_7_value ? ghv_2 : _GEN_2598; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2600 = 8'h3 == new_ptr_7_value ? ghv_3 : _GEN_2599; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2601 = 8'h4 == new_ptr_7_value ? ghv_4 : _GEN_2600; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2602 = 8'h5 == new_ptr_7_value ? ghv_5 : _GEN_2601; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2603 = 8'h6 == new_ptr_7_value ? ghv_6 : _GEN_2602; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2604 = 8'h7 == new_ptr_7_value ? ghv_7 : _GEN_2603; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2605 = 8'h8 == new_ptr_7_value ? ghv_8 : _GEN_2604; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2606 = 8'h9 == new_ptr_7_value ? ghv_9 : _GEN_2605; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2607 = 8'ha == new_ptr_7_value ? ghv_10 : _GEN_2606; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2608 = 8'hb == new_ptr_7_value ? ghv_11 : _GEN_2607; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2609 = 8'hc == new_ptr_7_value ? ghv_12 : _GEN_2608; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2610 = 8'hd == new_ptr_7_value ? ghv_13 : _GEN_2609; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2611 = 8'he == new_ptr_7_value ? ghv_14 : _GEN_2610; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2612 = 8'hf == new_ptr_7_value ? ghv_15 : _GEN_2611; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2613 = 8'h10 == new_ptr_7_value ? ghv_16 : _GEN_2612; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2614 = 8'h11 == new_ptr_7_value ? ghv_17 : _GEN_2613; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2615 = 8'h12 == new_ptr_7_value ? ghv_18 : _GEN_2614; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2616 = 8'h13 == new_ptr_7_value ? ghv_19 : _GEN_2615; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2617 = 8'h14 == new_ptr_7_value ? ghv_20 : _GEN_2616; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2618 = 8'h15 == new_ptr_7_value ? ghv_21 : _GEN_2617; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2619 = 8'h16 == new_ptr_7_value ? ghv_22 : _GEN_2618; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2620 = 8'h17 == new_ptr_7_value ? ghv_23 : _GEN_2619; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2621 = 8'h18 == new_ptr_7_value ? ghv_24 : _GEN_2620; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2622 = 8'h19 == new_ptr_7_value ? ghv_25 : _GEN_2621; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2623 = 8'h1a == new_ptr_7_value ? ghv_26 : _GEN_2622; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2624 = 8'h1b == new_ptr_7_value ? ghv_27 : _GEN_2623; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2625 = 8'h1c == new_ptr_7_value ? ghv_28 : _GEN_2624; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2626 = 8'h1d == new_ptr_7_value ? ghv_29 : _GEN_2625; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2627 = 8'h1e == new_ptr_7_value ? ghv_30 : _GEN_2626; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2628 = 8'h1f == new_ptr_7_value ? ghv_31 : _GEN_2627; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2629 = 8'h20 == new_ptr_7_value ? ghv_32 : _GEN_2628; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2630 = 8'h21 == new_ptr_7_value ? ghv_33 : _GEN_2629; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2631 = 8'h22 == new_ptr_7_value ? ghv_34 : _GEN_2630; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2632 = 8'h23 == new_ptr_7_value ? ghv_35 : _GEN_2631; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2633 = 8'h24 == new_ptr_7_value ? ghv_36 : _GEN_2632; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2634 = 8'h25 == new_ptr_7_value ? ghv_37 : _GEN_2633; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2635 = 8'h26 == new_ptr_7_value ? ghv_38 : _GEN_2634; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2636 = 8'h27 == new_ptr_7_value ? ghv_39 : _GEN_2635; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2637 = 8'h28 == new_ptr_7_value ? ghv_40 : _GEN_2636; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2638 = 8'h29 == new_ptr_7_value ? ghv_41 : _GEN_2637; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2639 = 8'h2a == new_ptr_7_value ? ghv_42 : _GEN_2638; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2640 = 8'h2b == new_ptr_7_value ? ghv_43 : _GEN_2639; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2641 = 8'h2c == new_ptr_7_value ? ghv_44 : _GEN_2640; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2642 = 8'h2d == new_ptr_7_value ? ghv_45 : _GEN_2641; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2643 = 8'h2e == new_ptr_7_value ? ghv_46 : _GEN_2642; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2644 = 8'h2f == new_ptr_7_value ? ghv_47 : _GEN_2643; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2645 = 8'h30 == new_ptr_7_value ? ghv_48 : _GEN_2644; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2646 = 8'h31 == new_ptr_7_value ? ghv_49 : _GEN_2645; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2647 = 8'h32 == new_ptr_7_value ? ghv_50 : _GEN_2646; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2648 = 8'h33 == new_ptr_7_value ? ghv_51 : _GEN_2647; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2649 = 8'h34 == new_ptr_7_value ? ghv_52 : _GEN_2648; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2650 = 8'h35 == new_ptr_7_value ? ghv_53 : _GEN_2649; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2651 = 8'h36 == new_ptr_7_value ? ghv_54 : _GEN_2650; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2652 = 8'h37 == new_ptr_7_value ? ghv_55 : _GEN_2651; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2653 = 8'h38 == new_ptr_7_value ? ghv_56 : _GEN_2652; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2654 = 8'h39 == new_ptr_7_value ? ghv_57 : _GEN_2653; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2655 = 8'h3a == new_ptr_7_value ? ghv_58 : _GEN_2654; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2656 = 8'h3b == new_ptr_7_value ? ghv_59 : _GEN_2655; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2657 = 8'h3c == new_ptr_7_value ? ghv_60 : _GEN_2656; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2658 = 8'h3d == new_ptr_7_value ? ghv_61 : _GEN_2657; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2659 = 8'h3e == new_ptr_7_value ? ghv_62 : _GEN_2658; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2660 = 8'h3f == new_ptr_7_value ? ghv_63 : _GEN_2659; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2661 = 8'h40 == new_ptr_7_value ? ghv_64 : _GEN_2660; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2662 = 8'h41 == new_ptr_7_value ? ghv_65 : _GEN_2661; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2663 = 8'h42 == new_ptr_7_value ? ghv_66 : _GEN_2662; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2664 = 8'h43 == new_ptr_7_value ? ghv_67 : _GEN_2663; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2665 = 8'h44 == new_ptr_7_value ? ghv_68 : _GEN_2664; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2666 = 8'h45 == new_ptr_7_value ? ghv_69 : _GEN_2665; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2667 = 8'h46 == new_ptr_7_value ? ghv_70 : _GEN_2666; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2668 = 8'h47 == new_ptr_7_value ? ghv_71 : _GEN_2667; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2669 = 8'h48 == new_ptr_7_value ? ghv_72 : _GEN_2668; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2670 = 8'h49 == new_ptr_7_value ? ghv_73 : _GEN_2669; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2671 = 8'h4a == new_ptr_7_value ? ghv_74 : _GEN_2670; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2672 = 8'h4b == new_ptr_7_value ? ghv_75 : _GEN_2671; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2673 = 8'h4c == new_ptr_7_value ? ghv_76 : _GEN_2672; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2674 = 8'h4d == new_ptr_7_value ? ghv_77 : _GEN_2673; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2675 = 8'h4e == new_ptr_7_value ? ghv_78 : _GEN_2674; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2676 = 8'h4f == new_ptr_7_value ? ghv_79 : _GEN_2675; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2677 = 8'h50 == new_ptr_7_value ? ghv_80 : _GEN_2676; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2678 = 8'h51 == new_ptr_7_value ? ghv_81 : _GEN_2677; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2679 = 8'h52 == new_ptr_7_value ? ghv_82 : _GEN_2678; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2680 = 8'h53 == new_ptr_7_value ? ghv_83 : _GEN_2679; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2681 = 8'h54 == new_ptr_7_value ? ghv_84 : _GEN_2680; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2682 = 8'h55 == new_ptr_7_value ? ghv_85 : _GEN_2681; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2683 = 8'h56 == new_ptr_7_value ? ghv_86 : _GEN_2682; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2684 = 8'h57 == new_ptr_7_value ? ghv_87 : _GEN_2683; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2685 = 8'h58 == new_ptr_7_value ? ghv_88 : _GEN_2684; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2686 = 8'h59 == new_ptr_7_value ? ghv_89 : _GEN_2685; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2687 = 8'h5a == new_ptr_7_value ? ghv_90 : _GEN_2686; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2688 = 8'h5b == new_ptr_7_value ? ghv_91 : _GEN_2687; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2689 = 8'h5c == new_ptr_7_value ? ghv_92 : _GEN_2688; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2690 = 8'h5d == new_ptr_7_value ? ghv_93 : _GEN_2689; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2691 = 8'h5e == new_ptr_7_value ? ghv_94 : _GEN_2690; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2692 = 8'h5f == new_ptr_7_value ? ghv_95 : _GEN_2691; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2693 = 8'h60 == new_ptr_7_value ? ghv_96 : _GEN_2692; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2694 = 8'h61 == new_ptr_7_value ? ghv_97 : _GEN_2693; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2695 = 8'h62 == new_ptr_7_value ? ghv_98 : _GEN_2694; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2696 = 8'h63 == new_ptr_7_value ? ghv_99 : _GEN_2695; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2697 = 8'h64 == new_ptr_7_value ? ghv_100 : _GEN_2696; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2698 = 8'h65 == new_ptr_7_value ? ghv_101 : _GEN_2697; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2699 = 8'h66 == new_ptr_7_value ? ghv_102 : _GEN_2698; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2700 = 8'h67 == new_ptr_7_value ? ghv_103 : _GEN_2699; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2701 = 8'h68 == new_ptr_7_value ? ghv_104 : _GEN_2700; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2702 = 8'h69 == new_ptr_7_value ? ghv_105 : _GEN_2701; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2703 = 8'h6a == new_ptr_7_value ? ghv_106 : _GEN_2702; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2704 = 8'h6b == new_ptr_7_value ? ghv_107 : _GEN_2703; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2705 = 8'h6c == new_ptr_7_value ? ghv_108 : _GEN_2704; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2706 = 8'h6d == new_ptr_7_value ? ghv_109 : _GEN_2705; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2707 = 8'h6e == new_ptr_7_value ? ghv_110 : _GEN_2706; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2708 = 8'h6f == new_ptr_7_value ? ghv_111 : _GEN_2707; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2709 = 8'h70 == new_ptr_7_value ? ghv_112 : _GEN_2708; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2710 = 8'h71 == new_ptr_7_value ? ghv_113 : _GEN_2709; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2711 = 8'h72 == new_ptr_7_value ? ghv_114 : _GEN_2710; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2712 = 8'h73 == new_ptr_7_value ? ghv_115 : _GEN_2711; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2713 = 8'h74 == new_ptr_7_value ? ghv_116 : _GEN_2712; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2714 = 8'h75 == new_ptr_7_value ? ghv_117 : _GEN_2713; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2715 = 8'h76 == new_ptr_7_value ? ghv_118 : _GEN_2714; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2716 = 8'h77 == new_ptr_7_value ? ghv_119 : _GEN_2715; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2717 = 8'h78 == new_ptr_7_value ? ghv_120 : _GEN_2716; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2718 = 8'h79 == new_ptr_7_value ? ghv_121 : _GEN_2717; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2719 = 8'h7a == new_ptr_7_value ? ghv_122 : _GEN_2718; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2720 = 8'h7b == new_ptr_7_value ? ghv_123 : _GEN_2719; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2721 = 8'h7c == new_ptr_7_value ? ghv_124 : _GEN_2720; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2722 = 8'h7d == new_ptr_7_value ? ghv_125 : _GEN_2721; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2723 = 8'h7e == new_ptr_7_value ? ghv_126 : _GEN_2722; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2724 = 8'h7f == new_ptr_7_value ? ghv_127 : _GEN_2723; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2725 = 8'h80 == new_ptr_7_value ? ghv_128 : _GEN_2724; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2726 = 8'h81 == new_ptr_7_value ? ghv_129 : _GEN_2725; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2727 = 8'h82 == new_ptr_7_value ? ghv_130 : _GEN_2726; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2728 = 8'h83 == new_ptr_7_value ? ghv_131 : _GEN_2727; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2729 = 8'h84 == new_ptr_7_value ? ghv_132 : _GEN_2728; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2730 = 8'h85 == new_ptr_7_value ? ghv_133 : _GEN_2729; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2731 = 8'h86 == new_ptr_7_value ? ghv_134 : _GEN_2730; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2732 = 8'h87 == new_ptr_7_value ? ghv_135 : _GEN_2731; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2733 = 8'h88 == new_ptr_7_value ? ghv_136 : _GEN_2732; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2734 = 8'h89 == new_ptr_7_value ? ghv_137 : _GEN_2733; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2735 = 8'h8a == new_ptr_7_value ? ghv_138 : _GEN_2734; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2736 = 8'h8b == new_ptr_7_value ? ghv_139 : _GEN_2735; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2737 = 8'h8c == new_ptr_7_value ? ghv_140 : _GEN_2736; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2738 = 8'h8d == new_ptr_7_value ? ghv_141 : _GEN_2737; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2739 = 8'h8e == new_ptr_7_value ? ghv_142 : _GEN_2738; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_5_value = _new_ptr_value_T_11[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_2742 = 8'h1 == new_ptr_5_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2743 = 8'h2 == new_ptr_5_value ? ghv_2 : _GEN_2742; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2744 = 8'h3 == new_ptr_5_value ? ghv_3 : _GEN_2743; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2745 = 8'h4 == new_ptr_5_value ? ghv_4 : _GEN_2744; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2746 = 8'h5 == new_ptr_5_value ? ghv_5 : _GEN_2745; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2747 = 8'h6 == new_ptr_5_value ? ghv_6 : _GEN_2746; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2748 = 8'h7 == new_ptr_5_value ? ghv_7 : _GEN_2747; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2749 = 8'h8 == new_ptr_5_value ? ghv_8 : _GEN_2748; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2750 = 8'h9 == new_ptr_5_value ? ghv_9 : _GEN_2749; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2751 = 8'ha == new_ptr_5_value ? ghv_10 : _GEN_2750; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2752 = 8'hb == new_ptr_5_value ? ghv_11 : _GEN_2751; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2753 = 8'hc == new_ptr_5_value ? ghv_12 : _GEN_2752; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2754 = 8'hd == new_ptr_5_value ? ghv_13 : _GEN_2753; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2755 = 8'he == new_ptr_5_value ? ghv_14 : _GEN_2754; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2756 = 8'hf == new_ptr_5_value ? ghv_15 : _GEN_2755; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2757 = 8'h10 == new_ptr_5_value ? ghv_16 : _GEN_2756; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2758 = 8'h11 == new_ptr_5_value ? ghv_17 : _GEN_2757; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2759 = 8'h12 == new_ptr_5_value ? ghv_18 : _GEN_2758; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2760 = 8'h13 == new_ptr_5_value ? ghv_19 : _GEN_2759; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2761 = 8'h14 == new_ptr_5_value ? ghv_20 : _GEN_2760; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2762 = 8'h15 == new_ptr_5_value ? ghv_21 : _GEN_2761; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2763 = 8'h16 == new_ptr_5_value ? ghv_22 : _GEN_2762; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2764 = 8'h17 == new_ptr_5_value ? ghv_23 : _GEN_2763; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2765 = 8'h18 == new_ptr_5_value ? ghv_24 : _GEN_2764; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2766 = 8'h19 == new_ptr_5_value ? ghv_25 : _GEN_2765; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2767 = 8'h1a == new_ptr_5_value ? ghv_26 : _GEN_2766; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2768 = 8'h1b == new_ptr_5_value ? ghv_27 : _GEN_2767; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2769 = 8'h1c == new_ptr_5_value ? ghv_28 : _GEN_2768; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2770 = 8'h1d == new_ptr_5_value ? ghv_29 : _GEN_2769; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2771 = 8'h1e == new_ptr_5_value ? ghv_30 : _GEN_2770; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2772 = 8'h1f == new_ptr_5_value ? ghv_31 : _GEN_2771; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2773 = 8'h20 == new_ptr_5_value ? ghv_32 : _GEN_2772; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2774 = 8'h21 == new_ptr_5_value ? ghv_33 : _GEN_2773; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2775 = 8'h22 == new_ptr_5_value ? ghv_34 : _GEN_2774; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2776 = 8'h23 == new_ptr_5_value ? ghv_35 : _GEN_2775; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2777 = 8'h24 == new_ptr_5_value ? ghv_36 : _GEN_2776; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2778 = 8'h25 == new_ptr_5_value ? ghv_37 : _GEN_2777; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2779 = 8'h26 == new_ptr_5_value ? ghv_38 : _GEN_2778; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2780 = 8'h27 == new_ptr_5_value ? ghv_39 : _GEN_2779; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2781 = 8'h28 == new_ptr_5_value ? ghv_40 : _GEN_2780; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2782 = 8'h29 == new_ptr_5_value ? ghv_41 : _GEN_2781; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2783 = 8'h2a == new_ptr_5_value ? ghv_42 : _GEN_2782; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2784 = 8'h2b == new_ptr_5_value ? ghv_43 : _GEN_2783; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2785 = 8'h2c == new_ptr_5_value ? ghv_44 : _GEN_2784; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2786 = 8'h2d == new_ptr_5_value ? ghv_45 : _GEN_2785; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2787 = 8'h2e == new_ptr_5_value ? ghv_46 : _GEN_2786; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2788 = 8'h2f == new_ptr_5_value ? ghv_47 : _GEN_2787; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2789 = 8'h30 == new_ptr_5_value ? ghv_48 : _GEN_2788; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2790 = 8'h31 == new_ptr_5_value ? ghv_49 : _GEN_2789; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2791 = 8'h32 == new_ptr_5_value ? ghv_50 : _GEN_2790; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2792 = 8'h33 == new_ptr_5_value ? ghv_51 : _GEN_2791; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2793 = 8'h34 == new_ptr_5_value ? ghv_52 : _GEN_2792; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2794 = 8'h35 == new_ptr_5_value ? ghv_53 : _GEN_2793; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2795 = 8'h36 == new_ptr_5_value ? ghv_54 : _GEN_2794; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2796 = 8'h37 == new_ptr_5_value ? ghv_55 : _GEN_2795; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2797 = 8'h38 == new_ptr_5_value ? ghv_56 : _GEN_2796; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2798 = 8'h39 == new_ptr_5_value ? ghv_57 : _GEN_2797; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2799 = 8'h3a == new_ptr_5_value ? ghv_58 : _GEN_2798; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2800 = 8'h3b == new_ptr_5_value ? ghv_59 : _GEN_2799; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2801 = 8'h3c == new_ptr_5_value ? ghv_60 : _GEN_2800; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2802 = 8'h3d == new_ptr_5_value ? ghv_61 : _GEN_2801; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2803 = 8'h3e == new_ptr_5_value ? ghv_62 : _GEN_2802; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2804 = 8'h3f == new_ptr_5_value ? ghv_63 : _GEN_2803; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2805 = 8'h40 == new_ptr_5_value ? ghv_64 : _GEN_2804; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2806 = 8'h41 == new_ptr_5_value ? ghv_65 : _GEN_2805; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2807 = 8'h42 == new_ptr_5_value ? ghv_66 : _GEN_2806; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2808 = 8'h43 == new_ptr_5_value ? ghv_67 : _GEN_2807; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2809 = 8'h44 == new_ptr_5_value ? ghv_68 : _GEN_2808; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2810 = 8'h45 == new_ptr_5_value ? ghv_69 : _GEN_2809; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2811 = 8'h46 == new_ptr_5_value ? ghv_70 : _GEN_2810; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2812 = 8'h47 == new_ptr_5_value ? ghv_71 : _GEN_2811; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2813 = 8'h48 == new_ptr_5_value ? ghv_72 : _GEN_2812; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2814 = 8'h49 == new_ptr_5_value ? ghv_73 : _GEN_2813; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2815 = 8'h4a == new_ptr_5_value ? ghv_74 : _GEN_2814; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2816 = 8'h4b == new_ptr_5_value ? ghv_75 : _GEN_2815; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2817 = 8'h4c == new_ptr_5_value ? ghv_76 : _GEN_2816; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2818 = 8'h4d == new_ptr_5_value ? ghv_77 : _GEN_2817; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2819 = 8'h4e == new_ptr_5_value ? ghv_78 : _GEN_2818; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2820 = 8'h4f == new_ptr_5_value ? ghv_79 : _GEN_2819; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2821 = 8'h50 == new_ptr_5_value ? ghv_80 : _GEN_2820; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2822 = 8'h51 == new_ptr_5_value ? ghv_81 : _GEN_2821; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2823 = 8'h52 == new_ptr_5_value ? ghv_82 : _GEN_2822; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2824 = 8'h53 == new_ptr_5_value ? ghv_83 : _GEN_2823; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2825 = 8'h54 == new_ptr_5_value ? ghv_84 : _GEN_2824; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2826 = 8'h55 == new_ptr_5_value ? ghv_85 : _GEN_2825; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2827 = 8'h56 == new_ptr_5_value ? ghv_86 : _GEN_2826; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2828 = 8'h57 == new_ptr_5_value ? ghv_87 : _GEN_2827; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2829 = 8'h58 == new_ptr_5_value ? ghv_88 : _GEN_2828; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2830 = 8'h59 == new_ptr_5_value ? ghv_89 : _GEN_2829; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2831 = 8'h5a == new_ptr_5_value ? ghv_90 : _GEN_2830; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2832 = 8'h5b == new_ptr_5_value ? ghv_91 : _GEN_2831; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2833 = 8'h5c == new_ptr_5_value ? ghv_92 : _GEN_2832; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2834 = 8'h5d == new_ptr_5_value ? ghv_93 : _GEN_2833; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2835 = 8'h5e == new_ptr_5_value ? ghv_94 : _GEN_2834; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2836 = 8'h5f == new_ptr_5_value ? ghv_95 : _GEN_2835; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2837 = 8'h60 == new_ptr_5_value ? ghv_96 : _GEN_2836; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2838 = 8'h61 == new_ptr_5_value ? ghv_97 : _GEN_2837; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2839 = 8'h62 == new_ptr_5_value ? ghv_98 : _GEN_2838; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2840 = 8'h63 == new_ptr_5_value ? ghv_99 : _GEN_2839; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2841 = 8'h64 == new_ptr_5_value ? ghv_100 : _GEN_2840; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2842 = 8'h65 == new_ptr_5_value ? ghv_101 : _GEN_2841; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2843 = 8'h66 == new_ptr_5_value ? ghv_102 : _GEN_2842; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2844 = 8'h67 == new_ptr_5_value ? ghv_103 : _GEN_2843; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2845 = 8'h68 == new_ptr_5_value ? ghv_104 : _GEN_2844; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2846 = 8'h69 == new_ptr_5_value ? ghv_105 : _GEN_2845; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2847 = 8'h6a == new_ptr_5_value ? ghv_106 : _GEN_2846; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2848 = 8'h6b == new_ptr_5_value ? ghv_107 : _GEN_2847; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2849 = 8'h6c == new_ptr_5_value ? ghv_108 : _GEN_2848; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2850 = 8'h6d == new_ptr_5_value ? ghv_109 : _GEN_2849; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2851 = 8'h6e == new_ptr_5_value ? ghv_110 : _GEN_2850; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2852 = 8'h6f == new_ptr_5_value ? ghv_111 : _GEN_2851; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2853 = 8'h70 == new_ptr_5_value ? ghv_112 : _GEN_2852; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2854 = 8'h71 == new_ptr_5_value ? ghv_113 : _GEN_2853; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2855 = 8'h72 == new_ptr_5_value ? ghv_114 : _GEN_2854; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2856 = 8'h73 == new_ptr_5_value ? ghv_115 : _GEN_2855; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2857 = 8'h74 == new_ptr_5_value ? ghv_116 : _GEN_2856; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2858 = 8'h75 == new_ptr_5_value ? ghv_117 : _GEN_2857; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2859 = 8'h76 == new_ptr_5_value ? ghv_118 : _GEN_2858; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2860 = 8'h77 == new_ptr_5_value ? ghv_119 : _GEN_2859; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2861 = 8'h78 == new_ptr_5_value ? ghv_120 : _GEN_2860; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2862 = 8'h79 == new_ptr_5_value ? ghv_121 : _GEN_2861; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2863 = 8'h7a == new_ptr_5_value ? ghv_122 : _GEN_2862; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2864 = 8'h7b == new_ptr_5_value ? ghv_123 : _GEN_2863; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2865 = 8'h7c == new_ptr_5_value ? ghv_124 : _GEN_2864; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2866 = 8'h7d == new_ptr_5_value ? ghv_125 : _GEN_2865; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2867 = 8'h7e == new_ptr_5_value ? ghv_126 : _GEN_2866; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2868 = 8'h7f == new_ptr_5_value ? ghv_127 : _GEN_2867; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2869 = 8'h80 == new_ptr_5_value ? ghv_128 : _GEN_2868; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2870 = 8'h81 == new_ptr_5_value ? ghv_129 : _GEN_2869; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2871 = 8'h82 == new_ptr_5_value ? ghv_130 : _GEN_2870; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2872 = 8'h83 == new_ptr_5_value ? ghv_131 : _GEN_2871; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2873 = 8'h84 == new_ptr_5_value ? ghv_132 : _GEN_2872; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2874 = 8'h85 == new_ptr_5_value ? ghv_133 : _GEN_2873; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2875 = 8'h86 == new_ptr_5_value ? ghv_134 : _GEN_2874; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2876 = 8'h87 == new_ptr_5_value ? ghv_135 : _GEN_2875; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2877 = 8'h88 == new_ptr_5_value ? ghv_136 : _GEN_2876; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2878 = 8'h89 == new_ptr_5_value ? ghv_137 : _GEN_2877; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2879 = 8'h8a == new_ptr_5_value ? ghv_138 : _GEN_2878; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2880 = 8'h8b == new_ptr_5_value ? ghv_139 : _GEN_2879; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2881 = 8'h8c == new_ptr_5_value ? ghv_140 : _GEN_2880; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2882 = 8'h8d == new_ptr_5_value ? ghv_141 : _GEN_2881; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2883 = 8'h8e == new_ptr_5_value ? ghv_142 : _GEN_2882; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_value = _new_ptr_value_T_1[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_2886 = 8'h1 == new_ptr_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2887 = 8'h2 == new_ptr_value ? ghv_2 : _GEN_2886; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2888 = 8'h3 == new_ptr_value ? ghv_3 : _GEN_2887; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2889 = 8'h4 == new_ptr_value ? ghv_4 : _GEN_2888; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2890 = 8'h5 == new_ptr_value ? ghv_5 : _GEN_2889; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2891 = 8'h6 == new_ptr_value ? ghv_6 : _GEN_2890; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2892 = 8'h7 == new_ptr_value ? ghv_7 : _GEN_2891; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2893 = 8'h8 == new_ptr_value ? ghv_8 : _GEN_2892; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2894 = 8'h9 == new_ptr_value ? ghv_9 : _GEN_2893; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2895 = 8'ha == new_ptr_value ? ghv_10 : _GEN_2894; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2896 = 8'hb == new_ptr_value ? ghv_11 : _GEN_2895; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2897 = 8'hc == new_ptr_value ? ghv_12 : _GEN_2896; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2898 = 8'hd == new_ptr_value ? ghv_13 : _GEN_2897; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2899 = 8'he == new_ptr_value ? ghv_14 : _GEN_2898; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2900 = 8'hf == new_ptr_value ? ghv_15 : _GEN_2899; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2901 = 8'h10 == new_ptr_value ? ghv_16 : _GEN_2900; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2902 = 8'h11 == new_ptr_value ? ghv_17 : _GEN_2901; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2903 = 8'h12 == new_ptr_value ? ghv_18 : _GEN_2902; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2904 = 8'h13 == new_ptr_value ? ghv_19 : _GEN_2903; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2905 = 8'h14 == new_ptr_value ? ghv_20 : _GEN_2904; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2906 = 8'h15 == new_ptr_value ? ghv_21 : _GEN_2905; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2907 = 8'h16 == new_ptr_value ? ghv_22 : _GEN_2906; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2908 = 8'h17 == new_ptr_value ? ghv_23 : _GEN_2907; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2909 = 8'h18 == new_ptr_value ? ghv_24 : _GEN_2908; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2910 = 8'h19 == new_ptr_value ? ghv_25 : _GEN_2909; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2911 = 8'h1a == new_ptr_value ? ghv_26 : _GEN_2910; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2912 = 8'h1b == new_ptr_value ? ghv_27 : _GEN_2911; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2913 = 8'h1c == new_ptr_value ? ghv_28 : _GEN_2912; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2914 = 8'h1d == new_ptr_value ? ghv_29 : _GEN_2913; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2915 = 8'h1e == new_ptr_value ? ghv_30 : _GEN_2914; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2916 = 8'h1f == new_ptr_value ? ghv_31 : _GEN_2915; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2917 = 8'h20 == new_ptr_value ? ghv_32 : _GEN_2916; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2918 = 8'h21 == new_ptr_value ? ghv_33 : _GEN_2917; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2919 = 8'h22 == new_ptr_value ? ghv_34 : _GEN_2918; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2920 = 8'h23 == new_ptr_value ? ghv_35 : _GEN_2919; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2921 = 8'h24 == new_ptr_value ? ghv_36 : _GEN_2920; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2922 = 8'h25 == new_ptr_value ? ghv_37 : _GEN_2921; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2923 = 8'h26 == new_ptr_value ? ghv_38 : _GEN_2922; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2924 = 8'h27 == new_ptr_value ? ghv_39 : _GEN_2923; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2925 = 8'h28 == new_ptr_value ? ghv_40 : _GEN_2924; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2926 = 8'h29 == new_ptr_value ? ghv_41 : _GEN_2925; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2927 = 8'h2a == new_ptr_value ? ghv_42 : _GEN_2926; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2928 = 8'h2b == new_ptr_value ? ghv_43 : _GEN_2927; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2929 = 8'h2c == new_ptr_value ? ghv_44 : _GEN_2928; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2930 = 8'h2d == new_ptr_value ? ghv_45 : _GEN_2929; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2931 = 8'h2e == new_ptr_value ? ghv_46 : _GEN_2930; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2932 = 8'h2f == new_ptr_value ? ghv_47 : _GEN_2931; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2933 = 8'h30 == new_ptr_value ? ghv_48 : _GEN_2932; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2934 = 8'h31 == new_ptr_value ? ghv_49 : _GEN_2933; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2935 = 8'h32 == new_ptr_value ? ghv_50 : _GEN_2934; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2936 = 8'h33 == new_ptr_value ? ghv_51 : _GEN_2935; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2937 = 8'h34 == new_ptr_value ? ghv_52 : _GEN_2936; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2938 = 8'h35 == new_ptr_value ? ghv_53 : _GEN_2937; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2939 = 8'h36 == new_ptr_value ? ghv_54 : _GEN_2938; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2940 = 8'h37 == new_ptr_value ? ghv_55 : _GEN_2939; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2941 = 8'h38 == new_ptr_value ? ghv_56 : _GEN_2940; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2942 = 8'h39 == new_ptr_value ? ghv_57 : _GEN_2941; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2943 = 8'h3a == new_ptr_value ? ghv_58 : _GEN_2942; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2944 = 8'h3b == new_ptr_value ? ghv_59 : _GEN_2943; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2945 = 8'h3c == new_ptr_value ? ghv_60 : _GEN_2944; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2946 = 8'h3d == new_ptr_value ? ghv_61 : _GEN_2945; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2947 = 8'h3e == new_ptr_value ? ghv_62 : _GEN_2946; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2948 = 8'h3f == new_ptr_value ? ghv_63 : _GEN_2947; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2949 = 8'h40 == new_ptr_value ? ghv_64 : _GEN_2948; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2950 = 8'h41 == new_ptr_value ? ghv_65 : _GEN_2949; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2951 = 8'h42 == new_ptr_value ? ghv_66 : _GEN_2950; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2952 = 8'h43 == new_ptr_value ? ghv_67 : _GEN_2951; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2953 = 8'h44 == new_ptr_value ? ghv_68 : _GEN_2952; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2954 = 8'h45 == new_ptr_value ? ghv_69 : _GEN_2953; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2955 = 8'h46 == new_ptr_value ? ghv_70 : _GEN_2954; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2956 = 8'h47 == new_ptr_value ? ghv_71 : _GEN_2955; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2957 = 8'h48 == new_ptr_value ? ghv_72 : _GEN_2956; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2958 = 8'h49 == new_ptr_value ? ghv_73 : _GEN_2957; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2959 = 8'h4a == new_ptr_value ? ghv_74 : _GEN_2958; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2960 = 8'h4b == new_ptr_value ? ghv_75 : _GEN_2959; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2961 = 8'h4c == new_ptr_value ? ghv_76 : _GEN_2960; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2962 = 8'h4d == new_ptr_value ? ghv_77 : _GEN_2961; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2963 = 8'h4e == new_ptr_value ? ghv_78 : _GEN_2962; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2964 = 8'h4f == new_ptr_value ? ghv_79 : _GEN_2963; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2965 = 8'h50 == new_ptr_value ? ghv_80 : _GEN_2964; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2966 = 8'h51 == new_ptr_value ? ghv_81 : _GEN_2965; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2967 = 8'h52 == new_ptr_value ? ghv_82 : _GEN_2966; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2968 = 8'h53 == new_ptr_value ? ghv_83 : _GEN_2967; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2969 = 8'h54 == new_ptr_value ? ghv_84 : _GEN_2968; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2970 = 8'h55 == new_ptr_value ? ghv_85 : _GEN_2969; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2971 = 8'h56 == new_ptr_value ? ghv_86 : _GEN_2970; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2972 = 8'h57 == new_ptr_value ? ghv_87 : _GEN_2971; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2973 = 8'h58 == new_ptr_value ? ghv_88 : _GEN_2972; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2974 = 8'h59 == new_ptr_value ? ghv_89 : _GEN_2973; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2975 = 8'h5a == new_ptr_value ? ghv_90 : _GEN_2974; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2976 = 8'h5b == new_ptr_value ? ghv_91 : _GEN_2975; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2977 = 8'h5c == new_ptr_value ? ghv_92 : _GEN_2976; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2978 = 8'h5d == new_ptr_value ? ghv_93 : _GEN_2977; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2979 = 8'h5e == new_ptr_value ? ghv_94 : _GEN_2978; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2980 = 8'h5f == new_ptr_value ? ghv_95 : _GEN_2979; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2981 = 8'h60 == new_ptr_value ? ghv_96 : _GEN_2980; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2982 = 8'h61 == new_ptr_value ? ghv_97 : _GEN_2981; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2983 = 8'h62 == new_ptr_value ? ghv_98 : _GEN_2982; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2984 = 8'h63 == new_ptr_value ? ghv_99 : _GEN_2983; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2985 = 8'h64 == new_ptr_value ? ghv_100 : _GEN_2984; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2986 = 8'h65 == new_ptr_value ? ghv_101 : _GEN_2985; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2987 = 8'h66 == new_ptr_value ? ghv_102 : _GEN_2986; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2988 = 8'h67 == new_ptr_value ? ghv_103 : _GEN_2987; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2989 = 8'h68 == new_ptr_value ? ghv_104 : _GEN_2988; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2990 = 8'h69 == new_ptr_value ? ghv_105 : _GEN_2989; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2991 = 8'h6a == new_ptr_value ? ghv_106 : _GEN_2990; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2992 = 8'h6b == new_ptr_value ? ghv_107 : _GEN_2991; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2993 = 8'h6c == new_ptr_value ? ghv_108 : _GEN_2992; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2994 = 8'h6d == new_ptr_value ? ghv_109 : _GEN_2993; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2995 = 8'h6e == new_ptr_value ? ghv_110 : _GEN_2994; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2996 = 8'h6f == new_ptr_value ? ghv_111 : _GEN_2995; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2997 = 8'h70 == new_ptr_value ? ghv_112 : _GEN_2996; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2998 = 8'h71 == new_ptr_value ? ghv_113 : _GEN_2997; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_2999 = 8'h72 == new_ptr_value ? ghv_114 : _GEN_2998; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3000 = 8'h73 == new_ptr_value ? ghv_115 : _GEN_2999; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3001 = 8'h74 == new_ptr_value ? ghv_116 : _GEN_3000; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3002 = 8'h75 == new_ptr_value ? ghv_117 : _GEN_3001; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3003 = 8'h76 == new_ptr_value ? ghv_118 : _GEN_3002; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3004 = 8'h77 == new_ptr_value ? ghv_119 : _GEN_3003; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3005 = 8'h78 == new_ptr_value ? ghv_120 : _GEN_3004; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3006 = 8'h79 == new_ptr_value ? ghv_121 : _GEN_3005; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3007 = 8'h7a == new_ptr_value ? ghv_122 : _GEN_3006; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3008 = 8'h7b == new_ptr_value ? ghv_123 : _GEN_3007; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3009 = 8'h7c == new_ptr_value ? ghv_124 : _GEN_3008; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3010 = 8'h7d == new_ptr_value ? ghv_125 : _GEN_3009; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3011 = 8'h7e == new_ptr_value ? ghv_126 : _GEN_3010; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3012 = 8'h7f == new_ptr_value ? ghv_127 : _GEN_3011; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3013 = 8'h80 == new_ptr_value ? ghv_128 : _GEN_3012; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3014 = 8'h81 == new_ptr_value ? ghv_129 : _GEN_3013; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3015 = 8'h82 == new_ptr_value ? ghv_130 : _GEN_3014; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3016 = 8'h83 == new_ptr_value ? ghv_131 : _GEN_3015; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3017 = 8'h84 == new_ptr_value ? ghv_132 : _GEN_3016; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3018 = 8'h85 == new_ptr_value ? ghv_133 : _GEN_3017; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3019 = 8'h86 == new_ptr_value ? ghv_134 : _GEN_3018; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3020 = 8'h87 == new_ptr_value ? ghv_135 : _GEN_3019; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3021 = 8'h88 == new_ptr_value ? ghv_136 : _GEN_3020; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3022 = 8'h89 == new_ptr_value ? ghv_137 : _GEN_3021; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3023 = 8'h8a == new_ptr_value ? ghv_138 : _GEN_3022; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3024 = 8'h8b == new_ptr_value ? ghv_139 : _GEN_3023; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3025 = 8'h8c == new_ptr_value ? ghv_140 : _GEN_3024; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3026 = 8'h8d == new_ptr_value ? ghv_141 : _GEN_3025; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3027 = 8'h8e == new_ptr_value ? ghv_142 : _GEN_3026; // @[FrontendBundle.scala 329:{20,20}]
  wire [9:0] s1_ghv_wens_diff = 10'sh0 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag = $signed(s1_ghv_wens_diff) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T = 10'sh0 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_1 = s1_ghv_wens_reverse_flag ? _s1_ghv_wens_new_ptr_value_T : 10'h0; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_value = _s1_ghv_wens_new_ptr_value_T_1[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_26 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_0_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_value & _s1_predicted_ghist_ptr_WIRE__0 & s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_1 = 10'sh1 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_1 = $signed(s1_ghv_wens_diff_1) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_2 = 10'sh1 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_3 = s1_ghv_wens_reverse_flag_1 ? _s1_ghv_wens_new_ptr_value_T_2 : 10'h1; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_1_value = _s1_ghv_wens_new_ptr_value_T_3[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_53 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_1_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_0_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_1_value & _s1_predicted_ghist_ptr_T_45 & s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_80 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_1_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_1_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_1_value & _s1_predicted_ghist_ptr_WIRE__0 & s1_valid
    ; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_3 = 10'sh2 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_3 = $signed(s1_ghv_wens_diff_3) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_6 = 10'sh2 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_7 = s1_ghv_wens_reverse_flag_3 ? _s1_ghv_wens_new_ptr_value_T_6 : 10'h2; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_3_value = _s1_ghv_wens_new_ptr_value_T_7[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_107 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_3_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_1_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_3_value & _s1_predicted_ghist_ptr_T_45 & s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_134 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_3_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_2_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_3_value & _s1_predicted_ghist_ptr_WIRE__0 & s1_valid
    ; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_5 = 10'sh3 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_5 = $signed(s1_ghv_wens_diff_5) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_10 = 10'sh3 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_11 = s1_ghv_wens_reverse_flag_5 ? _s1_ghv_wens_new_ptr_value_T_10 : 10'h3; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_5_value = _s1_ghv_wens_new_ptr_value_T_11[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_161 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_5_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_2_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_5_value & _s1_predicted_ghist_ptr_T_45 & s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_188 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_5_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_3_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_5_value & _s1_predicted_ghist_ptr_WIRE__0 & s1_valid
    ; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_7 = 10'sh4 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_7 = $signed(s1_ghv_wens_diff_7) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_14 = 10'sh4 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_15 = s1_ghv_wens_reverse_flag_7 ? _s1_ghv_wens_new_ptr_value_T_14 : 10'h4; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_7_value = _s1_ghv_wens_new_ptr_value_T_15[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_215 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_7_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_3_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_7_value & _s1_predicted_ghist_ptr_T_45 & s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_242 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_7_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_4_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_7_value & _s1_predicted_ghist_ptr_WIRE__0 & s1_valid
    ; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_9 = 10'sh5 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_9 = $signed(s1_ghv_wens_diff_9) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_18 = 10'sh5 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_19 = s1_ghv_wens_reverse_flag_9 ? _s1_ghv_wens_new_ptr_value_T_18 : 10'h5; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_9_value = _s1_ghv_wens_new_ptr_value_T_19[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_269 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_9_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_4_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_9_value & _s1_predicted_ghist_ptr_T_45 & s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_296 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_9_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_5_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_9_value & _s1_predicted_ghist_ptr_WIRE__0 & s1_valid
    ; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_11 = 10'sh6 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_11 = $signed(s1_ghv_wens_diff_11) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_22 = 10'sh6 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_23 = s1_ghv_wens_reverse_flag_11 ? _s1_ghv_wens_new_ptr_value_T_22 : 10'h6; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_11_value = _s1_ghv_wens_new_ptr_value_T_23[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_323 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_11_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_5_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_11_value & _s1_predicted_ghist_ptr_T_45 & s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_350 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_11_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_6_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_11_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_13 = 10'sh7 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_13 = $signed(s1_ghv_wens_diff_13) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_26 = 10'sh7 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_27 = s1_ghv_wens_reverse_flag_13 ? _s1_ghv_wens_new_ptr_value_T_26 : 10'h7; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_13_value = _s1_ghv_wens_new_ptr_value_T_27[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_377 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_13_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_6_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_13_value & _s1_predicted_ghist_ptr_T_45 & s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_404 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_13_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_7_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_13_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_15 = 10'sh8 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_15 = $signed(s1_ghv_wens_diff_15) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_30 = 10'sh8 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_31 = s1_ghv_wens_reverse_flag_15 ? _s1_ghv_wens_new_ptr_value_T_30 : 10'h8; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_15_value = _s1_ghv_wens_new_ptr_value_T_31[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_431 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_15_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_7_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_15_value & _s1_predicted_ghist_ptr_T_45 & s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_458 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_15_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_8_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_15_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_17 = 10'sh9 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_17 = $signed(s1_ghv_wens_diff_17) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_34 = 10'sh9 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_35 = s1_ghv_wens_reverse_flag_17 ? _s1_ghv_wens_new_ptr_value_T_34 : 10'h9; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_17_value = _s1_ghv_wens_new_ptr_value_T_35[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_485 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_17_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_8_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_17_value & _s1_predicted_ghist_ptr_T_45 & s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_512 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_17_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_9_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_17_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_19 = 10'sha - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_19 = $signed(s1_ghv_wens_diff_19) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_38 = 10'sha - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_39 = s1_ghv_wens_reverse_flag_19 ? _s1_ghv_wens_new_ptr_value_T_38 : 10'ha; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_19_value = _s1_ghv_wens_new_ptr_value_T_39[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_539 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_19_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_9_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_19_value & _s1_predicted_ghist_ptr_T_45 & s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_566 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_19_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_10_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_19_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_21 = 10'shb - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_21 = $signed(s1_ghv_wens_diff_21) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_42 = 10'shb - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_43 = s1_ghv_wens_reverse_flag_21 ? _s1_ghv_wens_new_ptr_value_T_42 : 10'hb; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_21_value = _s1_ghv_wens_new_ptr_value_T_43[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_593 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_21_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_10_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_21_value & _s1_predicted_ghist_ptr_T_45 & s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_620 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_21_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_11_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_21_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_23 = 10'shc - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_23 = $signed(s1_ghv_wens_diff_23) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_46 = 10'shc - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_47 = s1_ghv_wens_reverse_flag_23 ? _s1_ghv_wens_new_ptr_value_T_46 : 10'hc; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_23_value = _s1_ghv_wens_new_ptr_value_T_47[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_647 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_23_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_11_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_23_value & _s1_predicted_ghist_ptr_T_45 & s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_674 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_23_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_12_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_23_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_25 = 10'shd - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_25 = $signed(s1_ghv_wens_diff_25) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_50 = 10'shd - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_51 = s1_ghv_wens_reverse_flag_25 ? _s1_ghv_wens_new_ptr_value_T_50 : 10'hd; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_25_value = _s1_ghv_wens_new_ptr_value_T_51[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_701 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_25_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_12_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_25_value & _s1_predicted_ghist_ptr_T_45 & s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_728 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_25_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_13_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_25_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_27 = 10'she - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_27 = $signed(s1_ghv_wens_diff_27) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_54 = 10'she - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_55 = s1_ghv_wens_reverse_flag_27 ? _s1_ghv_wens_new_ptr_value_T_54 : 10'he; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_27_value = _s1_ghv_wens_new_ptr_value_T_55[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_755 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_27_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_13_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_27_value & _s1_predicted_ghist_ptr_T_45 & s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_782 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_27_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_14_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_27_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_29 = 10'shf - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_29 = $signed(s1_ghv_wens_diff_29) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_58 = 10'shf - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_59 = s1_ghv_wens_reverse_flag_29 ? _s1_ghv_wens_new_ptr_value_T_58 : 10'hf; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_29_value = _s1_ghv_wens_new_ptr_value_T_59[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_809 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_29_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_14_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_29_value & _s1_predicted_ghist_ptr_T_45 & s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_836 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_29_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_15_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_29_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_31 = 10'sh10 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_31 = $signed(s1_ghv_wens_diff_31) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_62 = 10'sh10 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_63 = s1_ghv_wens_reverse_flag_31 ? _s1_ghv_wens_new_ptr_value_T_62 : 10'h10; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_31_value = _s1_ghv_wens_new_ptr_value_T_63[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_863 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_31_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_15_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_31_value & _s1_predicted_ghist_ptr_T_45 & s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_890 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_31_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_16_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_31_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_33 = 10'sh11 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_33 = $signed(s1_ghv_wens_diff_33) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_66 = 10'sh11 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_67 = s1_ghv_wens_reverse_flag_33 ? _s1_ghv_wens_new_ptr_value_T_66 : 10'h11; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_33_value = _s1_ghv_wens_new_ptr_value_T_67[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_917 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_33_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_16_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_33_value & _s1_predicted_ghist_ptr_T_45 & s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_944 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_33_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_17_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_33_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_35 = 10'sh12 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_35 = $signed(s1_ghv_wens_diff_35) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_70 = 10'sh12 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_71 = s1_ghv_wens_reverse_flag_35 ? _s1_ghv_wens_new_ptr_value_T_70 : 10'h12; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_35_value = _s1_ghv_wens_new_ptr_value_T_71[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_971 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_35_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_17_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_35_value & _s1_predicted_ghist_ptr_T_45 & s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_998 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_35_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_18_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_35_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_37 = 10'sh13 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_37 = $signed(s1_ghv_wens_diff_37) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_74 = 10'sh13 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_75 = s1_ghv_wens_reverse_flag_37 ? _s1_ghv_wens_new_ptr_value_T_74 : 10'h13; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_37_value = _s1_ghv_wens_new_ptr_value_T_75[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_1025 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_37_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_18_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_37_value & _s1_predicted_ghist_ptr_T_45 & s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_1052 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_37_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_19_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_37_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_39 = 10'sh14 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_39 = $signed(s1_ghv_wens_diff_39) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_78 = 10'sh14 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_79 = s1_ghv_wens_reverse_flag_39 ? _s1_ghv_wens_new_ptr_value_T_78 : 10'h14; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_39_value = _s1_ghv_wens_new_ptr_value_T_79[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_1079 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_39_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_19_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_39_value & _s1_predicted_ghist_ptr_T_45 & s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_1106 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_39_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_20_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_39_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_41 = 10'sh15 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_41 = $signed(s1_ghv_wens_diff_41) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_82 = 10'sh15 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_83 = s1_ghv_wens_reverse_flag_41 ? _s1_ghv_wens_new_ptr_value_T_82 : 10'h15; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_41_value = _s1_ghv_wens_new_ptr_value_T_83[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_1133 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_41_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_20_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_41_value & _s1_predicted_ghist_ptr_T_45 & s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_1160 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_41_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_21_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_41_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_43 = 10'sh16 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_43 = $signed(s1_ghv_wens_diff_43) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_86 = 10'sh16 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_87 = s1_ghv_wens_reverse_flag_43 ? _s1_ghv_wens_new_ptr_value_T_86 : 10'h16; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_43_value = _s1_ghv_wens_new_ptr_value_T_87[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_1187 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_43_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_21_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_43_value & _s1_predicted_ghist_ptr_T_45 & s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_1214 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_43_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_22_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_43_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_45 = 10'sh17 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_45 = $signed(s1_ghv_wens_diff_45) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_90 = 10'sh17 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_91 = s1_ghv_wens_reverse_flag_45 ? _s1_ghv_wens_new_ptr_value_T_90 : 10'h17; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_45_value = _s1_ghv_wens_new_ptr_value_T_91[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_1241 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_45_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_22_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_45_value & _s1_predicted_ghist_ptr_T_45 & s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_1268 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_45_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_23_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_45_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_47 = 10'sh18 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_47 = $signed(s1_ghv_wens_diff_47) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_94 = 10'sh18 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_95 = s1_ghv_wens_reverse_flag_47 ? _s1_ghv_wens_new_ptr_value_T_94 : 10'h18; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_47_value = _s1_ghv_wens_new_ptr_value_T_95[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_1295 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_47_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_23_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_47_value & _s1_predicted_ghist_ptr_T_45 & s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_1322 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_47_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_24_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_47_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_49 = 10'sh19 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_49 = $signed(s1_ghv_wens_diff_49) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_98 = 10'sh19 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_99 = s1_ghv_wens_reverse_flag_49 ? _s1_ghv_wens_new_ptr_value_T_98 : 10'h19; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_49_value = _s1_ghv_wens_new_ptr_value_T_99[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_1349 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_49_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_24_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_49_value & _s1_predicted_ghist_ptr_T_45 & s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_1376 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_49_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_25_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_49_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_51 = 10'sh1a - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_51 = $signed(s1_ghv_wens_diff_51) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_102 = 10'sh1a - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_103 = s1_ghv_wens_reverse_flag_51 ? _s1_ghv_wens_new_ptr_value_T_102 : 10'h1a; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_51_value = _s1_ghv_wens_new_ptr_value_T_103[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_1403 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_51_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_25_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_51_value & _s1_predicted_ghist_ptr_T_45 & s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_1430 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_51_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_26_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_51_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_53 = 10'sh1b - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_53 = $signed(s1_ghv_wens_diff_53) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_106 = 10'sh1b - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_107 = s1_ghv_wens_reverse_flag_53 ? _s1_ghv_wens_new_ptr_value_T_106 : 10'h1b; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_53_value = _s1_ghv_wens_new_ptr_value_T_107[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_1457 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_53_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_26_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_53_value & _s1_predicted_ghist_ptr_T_45 & s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_1484 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_53_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_27_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_53_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_55 = 10'sh1c - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_55 = $signed(s1_ghv_wens_diff_55) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_110 = 10'sh1c - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_111 = s1_ghv_wens_reverse_flag_55 ? _s1_ghv_wens_new_ptr_value_T_110 : 10'h1c; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_55_value = _s1_ghv_wens_new_ptr_value_T_111[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_1511 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_55_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_27_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_55_value & _s1_predicted_ghist_ptr_T_45 & s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_1538 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_55_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_28_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_55_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_57 = 10'sh1d - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_57 = $signed(s1_ghv_wens_diff_57) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_114 = 10'sh1d - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_115 = s1_ghv_wens_reverse_flag_57 ? _s1_ghv_wens_new_ptr_value_T_114 : 10'h1d; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_57_value = _s1_ghv_wens_new_ptr_value_T_115[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_1565 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_57_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_28_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_57_value & _s1_predicted_ghist_ptr_T_45 & s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_1592 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_57_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_29_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_57_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_59 = 10'sh1e - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_59 = $signed(s1_ghv_wens_diff_59) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_118 = 10'sh1e - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_119 = s1_ghv_wens_reverse_flag_59 ? _s1_ghv_wens_new_ptr_value_T_118 : 10'h1e; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_59_value = _s1_ghv_wens_new_ptr_value_T_119[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_1619 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_59_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_29_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_59_value & _s1_predicted_ghist_ptr_T_45 & s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_1646 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_59_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_30_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_59_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_61 = 10'sh1f - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_61 = $signed(s1_ghv_wens_diff_61) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_122 = 10'sh1f - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_123 = s1_ghv_wens_reverse_flag_61 ? _s1_ghv_wens_new_ptr_value_T_122 : 10'h1f; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_61_value = _s1_ghv_wens_new_ptr_value_T_123[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_1673 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_61_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_30_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_61_value & _s1_predicted_ghist_ptr_T_45 & s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_1700 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_61_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_31_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_61_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_63 = 10'sh20 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_63 = $signed(s1_ghv_wens_diff_63) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_126 = 10'sh20 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_127 = s1_ghv_wens_reverse_flag_63 ? _s1_ghv_wens_new_ptr_value_T_126 : 10'h20; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_63_value = _s1_ghv_wens_new_ptr_value_T_127[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_1727 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_63_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_31_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_63_value & _s1_predicted_ghist_ptr_T_45 & s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_1754 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_63_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_32_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_63_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_65 = 10'sh21 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_65 = $signed(s1_ghv_wens_diff_65) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_130 = 10'sh21 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_131 = s1_ghv_wens_reverse_flag_65 ? _s1_ghv_wens_new_ptr_value_T_130 : 10'h21; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_65_value = _s1_ghv_wens_new_ptr_value_T_131[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_1781 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_65_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_32_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_65_value & _s1_predicted_ghist_ptr_T_45 & s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_1808 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_65_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_33_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_65_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_67 = 10'sh22 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_67 = $signed(s1_ghv_wens_diff_67) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_134 = 10'sh22 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_135 = s1_ghv_wens_reverse_flag_67 ? _s1_ghv_wens_new_ptr_value_T_134 : 10'h22; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_67_value = _s1_ghv_wens_new_ptr_value_T_135[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_1835 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_67_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_33_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_67_value & _s1_predicted_ghist_ptr_T_45 & s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_1862 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_67_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_34_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_67_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_69 = 10'sh23 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_69 = $signed(s1_ghv_wens_diff_69) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_138 = 10'sh23 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_139 = s1_ghv_wens_reverse_flag_69 ? _s1_ghv_wens_new_ptr_value_T_138 : 10'h23; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_69_value = _s1_ghv_wens_new_ptr_value_T_139[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_1889 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_69_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_34_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_69_value & _s1_predicted_ghist_ptr_T_45 & s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_1916 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_69_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_35_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_69_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_71 = 10'sh24 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_71 = $signed(s1_ghv_wens_diff_71) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_142 = 10'sh24 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_143 = s1_ghv_wens_reverse_flag_71 ? _s1_ghv_wens_new_ptr_value_T_142 : 10'h24; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_71_value = _s1_ghv_wens_new_ptr_value_T_143[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_1943 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_71_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_35_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_71_value & _s1_predicted_ghist_ptr_T_45 & s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_1970 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_71_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_36_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_71_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_73 = 10'sh25 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_73 = $signed(s1_ghv_wens_diff_73) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_146 = 10'sh25 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_147 = s1_ghv_wens_reverse_flag_73 ? _s1_ghv_wens_new_ptr_value_T_146 : 10'h25; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_73_value = _s1_ghv_wens_new_ptr_value_T_147[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_1997 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_73_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_36_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_73_value & _s1_predicted_ghist_ptr_T_45 & s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_2024 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_73_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_37_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_73_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_75 = 10'sh26 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_75 = $signed(s1_ghv_wens_diff_75) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_150 = 10'sh26 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_151 = s1_ghv_wens_reverse_flag_75 ? _s1_ghv_wens_new_ptr_value_T_150 : 10'h26; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_75_value = _s1_ghv_wens_new_ptr_value_T_151[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_2051 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_75_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_37_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_75_value & _s1_predicted_ghist_ptr_T_45 & s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_2078 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_75_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_38_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_75_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_77 = 10'sh27 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_77 = $signed(s1_ghv_wens_diff_77) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_154 = 10'sh27 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_155 = s1_ghv_wens_reverse_flag_77 ? _s1_ghv_wens_new_ptr_value_T_154 : 10'h27; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_77_value = _s1_ghv_wens_new_ptr_value_T_155[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_2105 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_77_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_38_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_77_value & _s1_predicted_ghist_ptr_T_45 & s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_2132 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_77_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_39_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_77_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_79 = 10'sh28 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_79 = $signed(s1_ghv_wens_diff_79) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_158 = 10'sh28 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_159 = s1_ghv_wens_reverse_flag_79 ? _s1_ghv_wens_new_ptr_value_T_158 : 10'h28; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_79_value = _s1_ghv_wens_new_ptr_value_T_159[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_2159 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_79_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_39_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_79_value & _s1_predicted_ghist_ptr_T_45 & s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_2186 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_79_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_40_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_79_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_81 = 10'sh29 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_81 = $signed(s1_ghv_wens_diff_81) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_162 = 10'sh29 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_163 = s1_ghv_wens_reverse_flag_81 ? _s1_ghv_wens_new_ptr_value_T_162 : 10'h29; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_81_value = _s1_ghv_wens_new_ptr_value_T_163[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_2213 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_81_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_40_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_81_value & _s1_predicted_ghist_ptr_T_45 & s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_2240 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_81_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_41_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_81_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_83 = 10'sh2a - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_83 = $signed(s1_ghv_wens_diff_83) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_166 = 10'sh2a - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_167 = s1_ghv_wens_reverse_flag_83 ? _s1_ghv_wens_new_ptr_value_T_166 : 10'h2a; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_83_value = _s1_ghv_wens_new_ptr_value_T_167[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_2267 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_83_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_41_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_83_value & _s1_predicted_ghist_ptr_T_45 & s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_2294 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_83_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_42_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_83_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_85 = 10'sh2b - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_85 = $signed(s1_ghv_wens_diff_85) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_170 = 10'sh2b - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_171 = s1_ghv_wens_reverse_flag_85 ? _s1_ghv_wens_new_ptr_value_T_170 : 10'h2b; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_85_value = _s1_ghv_wens_new_ptr_value_T_171[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_2321 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_85_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_42_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_85_value & _s1_predicted_ghist_ptr_T_45 & s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_2348 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_85_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_43_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_85_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_87 = 10'sh2c - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_87 = $signed(s1_ghv_wens_diff_87) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_174 = 10'sh2c - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_175 = s1_ghv_wens_reverse_flag_87 ? _s1_ghv_wens_new_ptr_value_T_174 : 10'h2c; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_87_value = _s1_ghv_wens_new_ptr_value_T_175[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_2375 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_87_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_43_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_87_value & _s1_predicted_ghist_ptr_T_45 & s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_2402 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_87_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_44_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_87_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_89 = 10'sh2d - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_89 = $signed(s1_ghv_wens_diff_89) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_178 = 10'sh2d - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_179 = s1_ghv_wens_reverse_flag_89 ? _s1_ghv_wens_new_ptr_value_T_178 : 10'h2d; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_89_value = _s1_ghv_wens_new_ptr_value_T_179[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_2429 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_89_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_44_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_89_value & _s1_predicted_ghist_ptr_T_45 & s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_2456 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_89_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_45_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_89_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_91 = 10'sh2e - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_91 = $signed(s1_ghv_wens_diff_91) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_182 = 10'sh2e - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_183 = s1_ghv_wens_reverse_flag_91 ? _s1_ghv_wens_new_ptr_value_T_182 : 10'h2e; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_91_value = _s1_ghv_wens_new_ptr_value_T_183[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_2483 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_91_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_45_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_91_value & _s1_predicted_ghist_ptr_T_45 & s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_2510 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_91_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_46_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_91_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_93 = 10'sh2f - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_93 = $signed(s1_ghv_wens_diff_93) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_186 = 10'sh2f - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_187 = s1_ghv_wens_reverse_flag_93 ? _s1_ghv_wens_new_ptr_value_T_186 : 10'h2f; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_93_value = _s1_ghv_wens_new_ptr_value_T_187[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_2537 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_93_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_46_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_93_value & _s1_predicted_ghist_ptr_T_45 & s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_2564 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_93_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_47_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_93_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_95 = 10'sh30 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_95 = $signed(s1_ghv_wens_diff_95) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_190 = 10'sh30 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_191 = s1_ghv_wens_reverse_flag_95 ? _s1_ghv_wens_new_ptr_value_T_190 : 10'h30; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_95_value = _s1_ghv_wens_new_ptr_value_T_191[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_2591 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_95_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_47_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_95_value & _s1_predicted_ghist_ptr_T_45 & s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_2618 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_95_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_48_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_95_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_97 = 10'sh31 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_97 = $signed(s1_ghv_wens_diff_97) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_194 = 10'sh31 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_195 = s1_ghv_wens_reverse_flag_97 ? _s1_ghv_wens_new_ptr_value_T_194 : 10'h31; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_97_value = _s1_ghv_wens_new_ptr_value_T_195[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_2645 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_97_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_48_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_97_value & _s1_predicted_ghist_ptr_T_45 & s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_2672 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_97_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_49_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_97_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_99 = 10'sh32 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_99 = $signed(s1_ghv_wens_diff_99) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_198 = 10'sh32 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_199 = s1_ghv_wens_reverse_flag_99 ? _s1_ghv_wens_new_ptr_value_T_198 : 10'h32; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_99_value = _s1_ghv_wens_new_ptr_value_T_199[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_2699 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_99_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_49_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_99_value & _s1_predicted_ghist_ptr_T_45 & s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_2726 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_99_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_50_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_99_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_101 = 10'sh33 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_101 = $signed(s1_ghv_wens_diff_101) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_202 = 10'sh33 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_203 = s1_ghv_wens_reverse_flag_101 ? _s1_ghv_wens_new_ptr_value_T_202 : 10'h33
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_101_value = _s1_ghv_wens_new_ptr_value_T_203[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_2753 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_101_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_50_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_101_value & _s1_predicted_ghist_ptr_T_45 & s1_valid
    ; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_2780 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_101_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_51_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_101_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_103 = 10'sh34 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_103 = $signed(s1_ghv_wens_diff_103) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_206 = 10'sh34 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_207 = s1_ghv_wens_reverse_flag_103 ? _s1_ghv_wens_new_ptr_value_T_206 : 10'h34
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_103_value = _s1_ghv_wens_new_ptr_value_T_207[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_2807 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_103_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_51_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_103_value & _s1_predicted_ghist_ptr_T_45 & s1_valid
    ; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_2834 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_103_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_52_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_103_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_105 = 10'sh35 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_105 = $signed(s1_ghv_wens_diff_105) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_210 = 10'sh35 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_211 = s1_ghv_wens_reverse_flag_105 ? _s1_ghv_wens_new_ptr_value_T_210 : 10'h35
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_105_value = _s1_ghv_wens_new_ptr_value_T_211[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_2861 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_105_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_52_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_105_value & _s1_predicted_ghist_ptr_T_45 & s1_valid
    ; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_2888 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_105_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_53_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_105_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_107 = 10'sh36 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_107 = $signed(s1_ghv_wens_diff_107) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_214 = 10'sh36 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_215 = s1_ghv_wens_reverse_flag_107 ? _s1_ghv_wens_new_ptr_value_T_214 : 10'h36
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_107_value = _s1_ghv_wens_new_ptr_value_T_215[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_2915 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_107_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_53_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_107_value & _s1_predicted_ghist_ptr_T_45 & s1_valid
    ; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_2942 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_107_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_54_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_107_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_109 = 10'sh37 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_109 = $signed(s1_ghv_wens_diff_109) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_218 = 10'sh37 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_219 = s1_ghv_wens_reverse_flag_109 ? _s1_ghv_wens_new_ptr_value_T_218 : 10'h37
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_109_value = _s1_ghv_wens_new_ptr_value_T_219[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_2969 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_109_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_54_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_109_value & _s1_predicted_ghist_ptr_T_45 & s1_valid
    ; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_2996 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_109_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_55_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_109_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_111 = 10'sh38 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_111 = $signed(s1_ghv_wens_diff_111) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_222 = 10'sh38 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_223 = s1_ghv_wens_reverse_flag_111 ? _s1_ghv_wens_new_ptr_value_T_222 : 10'h38
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_111_value = _s1_ghv_wens_new_ptr_value_T_223[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_3023 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_111_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_55_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_111_value & _s1_predicted_ghist_ptr_T_45 & s1_valid
    ; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_3050 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_111_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_56_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_111_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_113 = 10'sh39 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_113 = $signed(s1_ghv_wens_diff_113) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_226 = 10'sh39 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_227 = s1_ghv_wens_reverse_flag_113 ? _s1_ghv_wens_new_ptr_value_T_226 : 10'h39
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_113_value = _s1_ghv_wens_new_ptr_value_T_227[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_3077 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_113_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_56_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_113_value & _s1_predicted_ghist_ptr_T_45 & s1_valid
    ; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_3104 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_113_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_57_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_113_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_115 = 10'sh3a - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_115 = $signed(s1_ghv_wens_diff_115) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_230 = 10'sh3a - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_231 = s1_ghv_wens_reverse_flag_115 ? _s1_ghv_wens_new_ptr_value_T_230 : 10'h3a
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_115_value = _s1_ghv_wens_new_ptr_value_T_231[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_3131 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_115_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_57_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_115_value & _s1_predicted_ghist_ptr_T_45 & s1_valid
    ; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_3158 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_115_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_58_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_115_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_117 = 10'sh3b - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_117 = $signed(s1_ghv_wens_diff_117) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_234 = 10'sh3b - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_235 = s1_ghv_wens_reverse_flag_117 ? _s1_ghv_wens_new_ptr_value_T_234 : 10'h3b
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_117_value = _s1_ghv_wens_new_ptr_value_T_235[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_3185 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_117_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_58_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_117_value & _s1_predicted_ghist_ptr_T_45 & s1_valid
    ; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_3212 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_117_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_59_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_117_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_119 = 10'sh3c - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_119 = $signed(s1_ghv_wens_diff_119) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_238 = 10'sh3c - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_239 = s1_ghv_wens_reverse_flag_119 ? _s1_ghv_wens_new_ptr_value_T_238 : 10'h3c
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_119_value = _s1_ghv_wens_new_ptr_value_T_239[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_3239 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_119_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_59_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_119_value & _s1_predicted_ghist_ptr_T_45 & s1_valid
    ; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_3266 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_119_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_60_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_119_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_121 = 10'sh3d - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_121 = $signed(s1_ghv_wens_diff_121) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_242 = 10'sh3d - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_243 = s1_ghv_wens_reverse_flag_121 ? _s1_ghv_wens_new_ptr_value_T_242 : 10'h3d
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_121_value = _s1_ghv_wens_new_ptr_value_T_243[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_3293 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_121_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_60_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_121_value & _s1_predicted_ghist_ptr_T_45 & s1_valid
    ; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_3320 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_121_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_61_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_121_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_123 = 10'sh3e - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_123 = $signed(s1_ghv_wens_diff_123) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_246 = 10'sh3e - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_247 = s1_ghv_wens_reverse_flag_123 ? _s1_ghv_wens_new_ptr_value_T_246 : 10'h3e
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_123_value = _s1_ghv_wens_new_ptr_value_T_247[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_3347 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_123_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_61_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_123_value & _s1_predicted_ghist_ptr_T_45 & s1_valid
    ; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_3374 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_123_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_62_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_123_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_125 = 10'sh3f - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_125 = $signed(s1_ghv_wens_diff_125) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_250 = 10'sh3f - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_251 = s1_ghv_wens_reverse_flag_125 ? _s1_ghv_wens_new_ptr_value_T_250 : 10'h3f
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_125_value = _s1_ghv_wens_new_ptr_value_T_251[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_3401 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_125_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_62_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_125_value & _s1_predicted_ghist_ptr_T_45 & s1_valid
    ; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_3428 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_125_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_63_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_125_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_127 = 10'sh40 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_127 = $signed(s1_ghv_wens_diff_127) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_254 = 10'sh40 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_255 = s1_ghv_wens_reverse_flag_127 ? _s1_ghv_wens_new_ptr_value_T_254 : 10'h40
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_127_value = _s1_ghv_wens_new_ptr_value_T_255[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_3455 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_127_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_63_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_127_value & _s1_predicted_ghist_ptr_T_45 & s1_valid
    ; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_3482 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_127_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_64_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_127_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_129 = 10'sh41 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_129 = $signed(s1_ghv_wens_diff_129) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_258 = 10'sh41 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_259 = s1_ghv_wens_reverse_flag_129 ? _s1_ghv_wens_new_ptr_value_T_258 : 10'h41
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_129_value = _s1_ghv_wens_new_ptr_value_T_259[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_3509 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_129_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_64_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_129_value & _s1_predicted_ghist_ptr_T_45 & s1_valid
    ; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_3536 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_129_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_65_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_129_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_131 = 10'sh42 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_131 = $signed(s1_ghv_wens_diff_131) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_262 = 10'sh42 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_263 = s1_ghv_wens_reverse_flag_131 ? _s1_ghv_wens_new_ptr_value_T_262 : 10'h42
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_131_value = _s1_ghv_wens_new_ptr_value_T_263[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_3563 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_131_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_65_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_131_value & _s1_predicted_ghist_ptr_T_45 & s1_valid
    ; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_3590 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_131_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_66_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_131_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_133 = 10'sh43 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_133 = $signed(s1_ghv_wens_diff_133) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_266 = 10'sh43 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_267 = s1_ghv_wens_reverse_flag_133 ? _s1_ghv_wens_new_ptr_value_T_266 : 10'h43
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_133_value = _s1_ghv_wens_new_ptr_value_T_267[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_3617 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_133_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_66_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_133_value & _s1_predicted_ghist_ptr_T_45 & s1_valid
    ; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_3644 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_133_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_67_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_133_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_135 = 10'sh44 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_135 = $signed(s1_ghv_wens_diff_135) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_270 = 10'sh44 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_271 = s1_ghv_wens_reverse_flag_135 ? _s1_ghv_wens_new_ptr_value_T_270 : 10'h44
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_135_value = _s1_ghv_wens_new_ptr_value_T_271[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_3671 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_135_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_67_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_135_value & _s1_predicted_ghist_ptr_T_45 & s1_valid
    ; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_3698 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_135_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_68_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_135_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_137 = 10'sh45 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_137 = $signed(s1_ghv_wens_diff_137) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_274 = 10'sh45 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_275 = s1_ghv_wens_reverse_flag_137 ? _s1_ghv_wens_new_ptr_value_T_274 : 10'h45
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_137_value = _s1_ghv_wens_new_ptr_value_T_275[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_3725 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_137_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_68_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_137_value & _s1_predicted_ghist_ptr_T_45 & s1_valid
    ; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_3752 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_137_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_69_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_137_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_139 = 10'sh46 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_139 = $signed(s1_ghv_wens_diff_139) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_278 = 10'sh46 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_279 = s1_ghv_wens_reverse_flag_139 ? _s1_ghv_wens_new_ptr_value_T_278 : 10'h46
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_139_value = _s1_ghv_wens_new_ptr_value_T_279[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_3779 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_139_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_69_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_139_value & _s1_predicted_ghist_ptr_T_45 & s1_valid
    ; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_3806 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_139_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_70_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_139_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_141 = 10'sh47 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_141 = $signed(s1_ghv_wens_diff_141) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_282 = 10'sh47 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_283 = s1_ghv_wens_reverse_flag_141 ? _s1_ghv_wens_new_ptr_value_T_282 : 10'h47
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_141_value = _s1_ghv_wens_new_ptr_value_T_283[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_3833 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_141_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_70_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_141_value & _s1_predicted_ghist_ptr_T_45 & s1_valid
    ; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_3860 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_141_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_71_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_141_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_143 = 10'sh48 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_143 = $signed(s1_ghv_wens_diff_143) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_286 = 10'sh48 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_287 = s1_ghv_wens_reverse_flag_143 ? _s1_ghv_wens_new_ptr_value_T_286 : 10'h48
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_143_value = _s1_ghv_wens_new_ptr_value_T_287[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_3887 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_143_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_71_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_143_value & _s1_predicted_ghist_ptr_T_45 & s1_valid
    ; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_3914 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_143_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_72_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_143_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_145 = 10'sh49 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_145 = $signed(s1_ghv_wens_diff_145) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_290 = 10'sh49 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_291 = s1_ghv_wens_reverse_flag_145 ? _s1_ghv_wens_new_ptr_value_T_290 : 10'h49
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_145_value = _s1_ghv_wens_new_ptr_value_T_291[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_3941 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_145_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_72_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_145_value & _s1_predicted_ghist_ptr_T_45 & s1_valid
    ; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_3968 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_145_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_73_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_145_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_147 = 10'sh4a - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_147 = $signed(s1_ghv_wens_diff_147) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_294 = 10'sh4a - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_295 = s1_ghv_wens_reverse_flag_147 ? _s1_ghv_wens_new_ptr_value_T_294 : 10'h4a
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_147_value = _s1_ghv_wens_new_ptr_value_T_295[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_3995 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_147_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_73_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_147_value & _s1_predicted_ghist_ptr_T_45 & s1_valid
    ; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_4022 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_147_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_74_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_147_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_149 = 10'sh4b - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_149 = $signed(s1_ghv_wens_diff_149) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_298 = 10'sh4b - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_299 = s1_ghv_wens_reverse_flag_149 ? _s1_ghv_wens_new_ptr_value_T_298 : 10'h4b
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_149_value = _s1_ghv_wens_new_ptr_value_T_299[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_4049 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_149_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_74_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_149_value & _s1_predicted_ghist_ptr_T_45 & s1_valid
    ; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_4076 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_149_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_75_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_149_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_151 = 10'sh4c - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_151 = $signed(s1_ghv_wens_diff_151) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_302 = 10'sh4c - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_303 = s1_ghv_wens_reverse_flag_151 ? _s1_ghv_wens_new_ptr_value_T_302 : 10'h4c
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_151_value = _s1_ghv_wens_new_ptr_value_T_303[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_4103 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_151_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_75_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_151_value & _s1_predicted_ghist_ptr_T_45 & s1_valid
    ; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_4130 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_151_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_76_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_151_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_153 = 10'sh4d - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_153 = $signed(s1_ghv_wens_diff_153) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_306 = 10'sh4d - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_307 = s1_ghv_wens_reverse_flag_153 ? _s1_ghv_wens_new_ptr_value_T_306 : 10'h4d
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_153_value = _s1_ghv_wens_new_ptr_value_T_307[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_4157 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_153_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_76_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_153_value & _s1_predicted_ghist_ptr_T_45 & s1_valid
    ; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_4184 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_153_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_77_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_153_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_155 = 10'sh4e - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_155 = $signed(s1_ghv_wens_diff_155) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_310 = 10'sh4e - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_311 = s1_ghv_wens_reverse_flag_155 ? _s1_ghv_wens_new_ptr_value_T_310 : 10'h4e
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_155_value = _s1_ghv_wens_new_ptr_value_T_311[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_4211 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_155_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_77_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_155_value & _s1_predicted_ghist_ptr_T_45 & s1_valid
    ; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_4238 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_155_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_78_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_155_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_157 = 10'sh4f - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_157 = $signed(s1_ghv_wens_diff_157) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_314 = 10'sh4f - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_315 = s1_ghv_wens_reverse_flag_157 ? _s1_ghv_wens_new_ptr_value_T_314 : 10'h4f
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_157_value = _s1_ghv_wens_new_ptr_value_T_315[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_4265 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_157_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_78_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_157_value & _s1_predicted_ghist_ptr_T_45 & s1_valid
    ; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_4292 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_157_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_79_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_157_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_159 = 10'sh50 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_159 = $signed(s1_ghv_wens_diff_159) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_318 = 10'sh50 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_319 = s1_ghv_wens_reverse_flag_159 ? _s1_ghv_wens_new_ptr_value_T_318 : 10'h50
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_159_value = _s1_ghv_wens_new_ptr_value_T_319[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_4319 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_159_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_79_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_159_value & _s1_predicted_ghist_ptr_T_45 & s1_valid
    ; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_4346 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_159_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_80_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_159_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_161 = 10'sh51 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_161 = $signed(s1_ghv_wens_diff_161) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_322 = 10'sh51 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_323 = s1_ghv_wens_reverse_flag_161 ? _s1_ghv_wens_new_ptr_value_T_322 : 10'h51
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_161_value = _s1_ghv_wens_new_ptr_value_T_323[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_4373 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_161_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_80_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_161_value & _s1_predicted_ghist_ptr_T_45 & s1_valid
    ; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_4400 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_161_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_81_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_161_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_163 = 10'sh52 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_163 = $signed(s1_ghv_wens_diff_163) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_326 = 10'sh52 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_327 = s1_ghv_wens_reverse_flag_163 ? _s1_ghv_wens_new_ptr_value_T_326 : 10'h52
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_163_value = _s1_ghv_wens_new_ptr_value_T_327[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_4427 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_163_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_81_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_163_value & _s1_predicted_ghist_ptr_T_45 & s1_valid
    ; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_4454 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_163_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_82_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_163_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_165 = 10'sh53 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_165 = $signed(s1_ghv_wens_diff_165) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_330 = 10'sh53 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_331 = s1_ghv_wens_reverse_flag_165 ? _s1_ghv_wens_new_ptr_value_T_330 : 10'h53
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_165_value = _s1_ghv_wens_new_ptr_value_T_331[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_4481 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_165_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_82_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_165_value & _s1_predicted_ghist_ptr_T_45 & s1_valid
    ; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_4508 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_165_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_83_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_165_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_167 = 10'sh54 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_167 = $signed(s1_ghv_wens_diff_167) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_334 = 10'sh54 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_335 = s1_ghv_wens_reverse_flag_167 ? _s1_ghv_wens_new_ptr_value_T_334 : 10'h54
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_167_value = _s1_ghv_wens_new_ptr_value_T_335[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_4535 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_167_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_83_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_167_value & _s1_predicted_ghist_ptr_T_45 & s1_valid
    ; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_4562 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_167_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_84_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_167_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_169 = 10'sh55 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_169 = $signed(s1_ghv_wens_diff_169) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_338 = 10'sh55 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_339 = s1_ghv_wens_reverse_flag_169 ? _s1_ghv_wens_new_ptr_value_T_338 : 10'h55
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_169_value = _s1_ghv_wens_new_ptr_value_T_339[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_4589 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_169_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_84_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_169_value & _s1_predicted_ghist_ptr_T_45 & s1_valid
    ; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_4616 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_169_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_85_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_169_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_171 = 10'sh56 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_171 = $signed(s1_ghv_wens_diff_171) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_342 = 10'sh56 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_343 = s1_ghv_wens_reverse_flag_171 ? _s1_ghv_wens_new_ptr_value_T_342 : 10'h56
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_171_value = _s1_ghv_wens_new_ptr_value_T_343[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_4643 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_171_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_85_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_171_value & _s1_predicted_ghist_ptr_T_45 & s1_valid
    ; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_4670 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_171_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_86_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_171_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_173 = 10'sh57 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_173 = $signed(s1_ghv_wens_diff_173) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_346 = 10'sh57 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_347 = s1_ghv_wens_reverse_flag_173 ? _s1_ghv_wens_new_ptr_value_T_346 : 10'h57
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_173_value = _s1_ghv_wens_new_ptr_value_T_347[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_4697 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_173_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_86_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_173_value & _s1_predicted_ghist_ptr_T_45 & s1_valid
    ; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_4724 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_173_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_87_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_173_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_175 = 10'sh58 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_175 = $signed(s1_ghv_wens_diff_175) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_350 = 10'sh58 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_351 = s1_ghv_wens_reverse_flag_175 ? _s1_ghv_wens_new_ptr_value_T_350 : 10'h58
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_175_value = _s1_ghv_wens_new_ptr_value_T_351[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_4751 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_175_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_87_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_175_value & _s1_predicted_ghist_ptr_T_45 & s1_valid
    ; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_4778 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_175_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_88_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_175_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_177 = 10'sh59 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_177 = $signed(s1_ghv_wens_diff_177) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_354 = 10'sh59 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_355 = s1_ghv_wens_reverse_flag_177 ? _s1_ghv_wens_new_ptr_value_T_354 : 10'h59
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_177_value = _s1_ghv_wens_new_ptr_value_T_355[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_4805 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_177_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_88_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_177_value & _s1_predicted_ghist_ptr_T_45 & s1_valid
    ; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_4832 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_177_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_89_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_177_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_179 = 10'sh5a - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_179 = $signed(s1_ghv_wens_diff_179) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_358 = 10'sh5a - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_359 = s1_ghv_wens_reverse_flag_179 ? _s1_ghv_wens_new_ptr_value_T_358 : 10'h5a
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_179_value = _s1_ghv_wens_new_ptr_value_T_359[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_4859 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_179_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_89_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_179_value & _s1_predicted_ghist_ptr_T_45 & s1_valid
    ; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_4886 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_179_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_90_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_179_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_181 = 10'sh5b - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_181 = $signed(s1_ghv_wens_diff_181) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_362 = 10'sh5b - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_363 = s1_ghv_wens_reverse_flag_181 ? _s1_ghv_wens_new_ptr_value_T_362 : 10'h5b
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_181_value = _s1_ghv_wens_new_ptr_value_T_363[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_4913 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_181_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_90_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_181_value & _s1_predicted_ghist_ptr_T_45 & s1_valid
    ; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_4940 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_181_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_91_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_181_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_183 = 10'sh5c - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_183 = $signed(s1_ghv_wens_diff_183) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_366 = 10'sh5c - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_367 = s1_ghv_wens_reverse_flag_183 ? _s1_ghv_wens_new_ptr_value_T_366 : 10'h5c
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_183_value = _s1_ghv_wens_new_ptr_value_T_367[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_4967 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_183_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_91_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_183_value & _s1_predicted_ghist_ptr_T_45 & s1_valid
    ; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_4994 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_183_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_92_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_183_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_185 = 10'sh5d - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_185 = $signed(s1_ghv_wens_diff_185) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_370 = 10'sh5d - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_371 = s1_ghv_wens_reverse_flag_185 ? _s1_ghv_wens_new_ptr_value_T_370 : 10'h5d
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_185_value = _s1_ghv_wens_new_ptr_value_T_371[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_5021 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_185_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_92_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_185_value & _s1_predicted_ghist_ptr_T_45 & s1_valid
    ; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_5048 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_185_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_93_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_185_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_187 = 10'sh5e - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_187 = $signed(s1_ghv_wens_diff_187) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_374 = 10'sh5e - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_375 = s1_ghv_wens_reverse_flag_187 ? _s1_ghv_wens_new_ptr_value_T_374 : 10'h5e
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_187_value = _s1_ghv_wens_new_ptr_value_T_375[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_5075 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_187_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_93_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_187_value & _s1_predicted_ghist_ptr_T_45 & s1_valid
    ; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_5102 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_187_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_94_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_187_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_189 = 10'sh5f - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_189 = $signed(s1_ghv_wens_diff_189) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_378 = 10'sh5f - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_379 = s1_ghv_wens_reverse_flag_189 ? _s1_ghv_wens_new_ptr_value_T_378 : 10'h5f
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_189_value = _s1_ghv_wens_new_ptr_value_T_379[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_5129 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_189_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_94_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_189_value & _s1_predicted_ghist_ptr_T_45 & s1_valid
    ; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_5156 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_189_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_95_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_189_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_191 = 10'sh60 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_191 = $signed(s1_ghv_wens_diff_191) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_382 = 10'sh60 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_383 = s1_ghv_wens_reverse_flag_191 ? _s1_ghv_wens_new_ptr_value_T_382 : 10'h60
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_191_value = _s1_ghv_wens_new_ptr_value_T_383[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_5183 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_191_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_95_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_191_value & _s1_predicted_ghist_ptr_T_45 & s1_valid
    ; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_5210 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_191_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_96_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_191_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_193 = 10'sh61 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_193 = $signed(s1_ghv_wens_diff_193) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_386 = 10'sh61 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_387 = s1_ghv_wens_reverse_flag_193 ? _s1_ghv_wens_new_ptr_value_T_386 : 10'h61
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_193_value = _s1_ghv_wens_new_ptr_value_T_387[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_5237 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_193_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_96_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_193_value & _s1_predicted_ghist_ptr_T_45 & s1_valid
    ; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_5264 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_193_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_97_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_193_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_195 = 10'sh62 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_195 = $signed(s1_ghv_wens_diff_195) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_390 = 10'sh62 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_391 = s1_ghv_wens_reverse_flag_195 ? _s1_ghv_wens_new_ptr_value_T_390 : 10'h62
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_195_value = _s1_ghv_wens_new_ptr_value_T_391[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_5291 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_195_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_97_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_195_value & _s1_predicted_ghist_ptr_T_45 & s1_valid
    ; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_5318 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_195_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_98_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_195_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_197 = 10'sh63 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_197 = $signed(s1_ghv_wens_diff_197) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_394 = 10'sh63 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_395 = s1_ghv_wens_reverse_flag_197 ? _s1_ghv_wens_new_ptr_value_T_394 : 10'h63
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_197_value = _s1_ghv_wens_new_ptr_value_T_395[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_5345 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_197_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_98_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_197_value & _s1_predicted_ghist_ptr_T_45 & s1_valid
    ; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_5372 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_197_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_99_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_197_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_199 = 10'sh64 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_199 = $signed(s1_ghv_wens_diff_199) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_398 = 10'sh64 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_399 = s1_ghv_wens_reverse_flag_199 ? _s1_ghv_wens_new_ptr_value_T_398 : 10'h64
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_199_value = _s1_ghv_wens_new_ptr_value_T_399[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_5399 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_199_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_99_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_199_value & _s1_predicted_ghist_ptr_T_45 & s1_valid
    ; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_5426 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_199_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_100_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_199_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_201 = 10'sh65 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_201 = $signed(s1_ghv_wens_diff_201) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_402 = 10'sh65 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_403 = s1_ghv_wens_reverse_flag_201 ? _s1_ghv_wens_new_ptr_value_T_402 : 10'h65
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_201_value = _s1_ghv_wens_new_ptr_value_T_403[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_5453 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_201_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_100_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_201_value & _s1_predicted_ghist_ptr_T_45 &
    s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_5480 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_201_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_101_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_201_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_203 = 10'sh66 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_203 = $signed(s1_ghv_wens_diff_203) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_406 = 10'sh66 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_407 = s1_ghv_wens_reverse_flag_203 ? _s1_ghv_wens_new_ptr_value_T_406 : 10'h66
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_203_value = _s1_ghv_wens_new_ptr_value_T_407[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_5507 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_203_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_101_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_203_value & _s1_predicted_ghist_ptr_T_45 &
    s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_5534 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_203_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_102_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_203_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_205 = 10'sh67 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_205 = $signed(s1_ghv_wens_diff_205) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_410 = 10'sh67 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_411 = s1_ghv_wens_reverse_flag_205 ? _s1_ghv_wens_new_ptr_value_T_410 : 10'h67
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_205_value = _s1_ghv_wens_new_ptr_value_T_411[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_5561 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_205_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_102_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_205_value & _s1_predicted_ghist_ptr_T_45 &
    s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_5588 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_205_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_103_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_205_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_207 = 10'sh68 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_207 = $signed(s1_ghv_wens_diff_207) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_414 = 10'sh68 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_415 = s1_ghv_wens_reverse_flag_207 ? _s1_ghv_wens_new_ptr_value_T_414 : 10'h68
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_207_value = _s1_ghv_wens_new_ptr_value_T_415[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_5615 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_207_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_103_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_207_value & _s1_predicted_ghist_ptr_T_45 &
    s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_5642 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_207_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_104_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_207_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_209 = 10'sh69 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_209 = $signed(s1_ghv_wens_diff_209) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_418 = 10'sh69 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_419 = s1_ghv_wens_reverse_flag_209 ? _s1_ghv_wens_new_ptr_value_T_418 : 10'h69
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_209_value = _s1_ghv_wens_new_ptr_value_T_419[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_5669 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_209_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_104_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_209_value & _s1_predicted_ghist_ptr_T_45 &
    s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_5696 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_209_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_105_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_209_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_211 = 10'sh6a - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_211 = $signed(s1_ghv_wens_diff_211) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_422 = 10'sh6a - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_423 = s1_ghv_wens_reverse_flag_211 ? _s1_ghv_wens_new_ptr_value_T_422 : 10'h6a
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_211_value = _s1_ghv_wens_new_ptr_value_T_423[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_5723 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_211_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_105_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_211_value & _s1_predicted_ghist_ptr_T_45 &
    s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_5750 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_211_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_106_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_211_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_213 = 10'sh6b - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_213 = $signed(s1_ghv_wens_diff_213) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_426 = 10'sh6b - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_427 = s1_ghv_wens_reverse_flag_213 ? _s1_ghv_wens_new_ptr_value_T_426 : 10'h6b
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_213_value = _s1_ghv_wens_new_ptr_value_T_427[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_5777 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_213_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_106_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_213_value & _s1_predicted_ghist_ptr_T_45 &
    s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_5804 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_213_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_107_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_213_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_215 = 10'sh6c - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_215 = $signed(s1_ghv_wens_diff_215) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_430 = 10'sh6c - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_431 = s1_ghv_wens_reverse_flag_215 ? _s1_ghv_wens_new_ptr_value_T_430 : 10'h6c
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_215_value = _s1_ghv_wens_new_ptr_value_T_431[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_5831 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_215_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_107_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_215_value & _s1_predicted_ghist_ptr_T_45 &
    s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_5858 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_215_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_108_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_215_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_217 = 10'sh6d - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_217 = $signed(s1_ghv_wens_diff_217) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_434 = 10'sh6d - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_435 = s1_ghv_wens_reverse_flag_217 ? _s1_ghv_wens_new_ptr_value_T_434 : 10'h6d
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_217_value = _s1_ghv_wens_new_ptr_value_T_435[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_5885 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_217_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_108_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_217_value & _s1_predicted_ghist_ptr_T_45 &
    s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_5912 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_217_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_109_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_217_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_219 = 10'sh6e - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_219 = $signed(s1_ghv_wens_diff_219) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_438 = 10'sh6e - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_439 = s1_ghv_wens_reverse_flag_219 ? _s1_ghv_wens_new_ptr_value_T_438 : 10'h6e
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_219_value = _s1_ghv_wens_new_ptr_value_T_439[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_5939 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_219_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_109_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_219_value & _s1_predicted_ghist_ptr_T_45 &
    s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_5966 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_219_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_110_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_219_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_221 = 10'sh6f - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_221 = $signed(s1_ghv_wens_diff_221) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_442 = 10'sh6f - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_443 = s1_ghv_wens_reverse_flag_221 ? _s1_ghv_wens_new_ptr_value_T_442 : 10'h6f
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_221_value = _s1_ghv_wens_new_ptr_value_T_443[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_5993 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_221_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_110_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_221_value & _s1_predicted_ghist_ptr_T_45 &
    s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_6020 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_221_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_111_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_221_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_223 = 10'sh70 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_223 = $signed(s1_ghv_wens_diff_223) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_446 = 10'sh70 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_447 = s1_ghv_wens_reverse_flag_223 ? _s1_ghv_wens_new_ptr_value_T_446 : 10'h70
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_223_value = _s1_ghv_wens_new_ptr_value_T_447[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_6047 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_223_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_111_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_223_value & _s1_predicted_ghist_ptr_T_45 &
    s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_6074 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_223_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_112_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_223_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_225 = 10'sh71 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_225 = $signed(s1_ghv_wens_diff_225) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_450 = 10'sh71 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_451 = s1_ghv_wens_reverse_flag_225 ? _s1_ghv_wens_new_ptr_value_T_450 : 10'h71
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_225_value = _s1_ghv_wens_new_ptr_value_T_451[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_6101 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_225_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_112_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_225_value & _s1_predicted_ghist_ptr_T_45 &
    s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_6128 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_225_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_113_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_225_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_227 = 10'sh72 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_227 = $signed(s1_ghv_wens_diff_227) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_454 = 10'sh72 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_455 = s1_ghv_wens_reverse_flag_227 ? _s1_ghv_wens_new_ptr_value_T_454 : 10'h72
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_227_value = _s1_ghv_wens_new_ptr_value_T_455[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_6155 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_227_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_113_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_227_value & _s1_predicted_ghist_ptr_T_45 &
    s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_6182 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_227_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_114_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_227_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_229 = 10'sh73 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_229 = $signed(s1_ghv_wens_diff_229) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_458 = 10'sh73 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_459 = s1_ghv_wens_reverse_flag_229 ? _s1_ghv_wens_new_ptr_value_T_458 : 10'h73
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_229_value = _s1_ghv_wens_new_ptr_value_T_459[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_6209 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_229_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_114_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_229_value & _s1_predicted_ghist_ptr_T_45 &
    s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_6236 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_229_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_115_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_229_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_231 = 10'sh74 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_231 = $signed(s1_ghv_wens_diff_231) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_462 = 10'sh74 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_463 = s1_ghv_wens_reverse_flag_231 ? _s1_ghv_wens_new_ptr_value_T_462 : 10'h74
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_231_value = _s1_ghv_wens_new_ptr_value_T_463[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_6263 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_231_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_115_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_231_value & _s1_predicted_ghist_ptr_T_45 &
    s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_6290 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_231_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_116_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_231_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_233 = 10'sh75 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_233 = $signed(s1_ghv_wens_diff_233) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_466 = 10'sh75 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_467 = s1_ghv_wens_reverse_flag_233 ? _s1_ghv_wens_new_ptr_value_T_466 : 10'h75
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_233_value = _s1_ghv_wens_new_ptr_value_T_467[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_6317 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_233_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_116_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_233_value & _s1_predicted_ghist_ptr_T_45 &
    s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_6344 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_233_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_117_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_233_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_235 = 10'sh76 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_235 = $signed(s1_ghv_wens_diff_235) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_470 = 10'sh76 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_471 = s1_ghv_wens_reverse_flag_235 ? _s1_ghv_wens_new_ptr_value_T_470 : 10'h76
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_235_value = _s1_ghv_wens_new_ptr_value_T_471[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_6371 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_235_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_117_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_235_value & _s1_predicted_ghist_ptr_T_45 &
    s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_6398 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_235_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_118_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_235_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_237 = 10'sh77 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_237 = $signed(s1_ghv_wens_diff_237) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_474 = 10'sh77 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_475 = s1_ghv_wens_reverse_flag_237 ? _s1_ghv_wens_new_ptr_value_T_474 : 10'h77
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_237_value = _s1_ghv_wens_new_ptr_value_T_475[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_6425 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_237_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_118_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_237_value & _s1_predicted_ghist_ptr_T_45 &
    s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_6452 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_237_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_119_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_237_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_239 = 10'sh78 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_239 = $signed(s1_ghv_wens_diff_239) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_478 = 10'sh78 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_479 = s1_ghv_wens_reverse_flag_239 ? _s1_ghv_wens_new_ptr_value_T_478 : 10'h78
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_239_value = _s1_ghv_wens_new_ptr_value_T_479[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_6479 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_239_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_119_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_239_value & _s1_predicted_ghist_ptr_T_45 &
    s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_6506 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_239_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_120_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_239_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_241 = 10'sh79 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_241 = $signed(s1_ghv_wens_diff_241) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_482 = 10'sh79 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_483 = s1_ghv_wens_reverse_flag_241 ? _s1_ghv_wens_new_ptr_value_T_482 : 10'h79
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_241_value = _s1_ghv_wens_new_ptr_value_T_483[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_6533 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_241_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_120_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_241_value & _s1_predicted_ghist_ptr_T_45 &
    s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_6560 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_241_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_121_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_241_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_243 = 10'sh7a - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_243 = $signed(s1_ghv_wens_diff_243) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_486 = 10'sh7a - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_487 = s1_ghv_wens_reverse_flag_243 ? _s1_ghv_wens_new_ptr_value_T_486 : 10'h7a
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_243_value = _s1_ghv_wens_new_ptr_value_T_487[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_6587 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_243_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_121_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_243_value & _s1_predicted_ghist_ptr_T_45 &
    s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_6614 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_243_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_122_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_243_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_245 = 10'sh7b - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_245 = $signed(s1_ghv_wens_diff_245) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_490 = 10'sh7b - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_491 = s1_ghv_wens_reverse_flag_245 ? _s1_ghv_wens_new_ptr_value_T_490 : 10'h7b
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_245_value = _s1_ghv_wens_new_ptr_value_T_491[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_6641 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_245_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_122_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_245_value & _s1_predicted_ghist_ptr_T_45 &
    s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_6668 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_245_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_123_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_245_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_247 = 10'sh7c - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_247 = $signed(s1_ghv_wens_diff_247) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_494 = 10'sh7c - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_495 = s1_ghv_wens_reverse_flag_247 ? _s1_ghv_wens_new_ptr_value_T_494 : 10'h7c
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_247_value = _s1_ghv_wens_new_ptr_value_T_495[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_6695 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_247_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_123_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_247_value & _s1_predicted_ghist_ptr_T_45 &
    s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_6722 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_247_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_124_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_247_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_249 = 10'sh7d - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_249 = $signed(s1_ghv_wens_diff_249) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_498 = 10'sh7d - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_499 = s1_ghv_wens_reverse_flag_249 ? _s1_ghv_wens_new_ptr_value_T_498 : 10'h7d
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_249_value = _s1_ghv_wens_new_ptr_value_T_499[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_6749 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_249_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_124_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_249_value & _s1_predicted_ghist_ptr_T_45 &
    s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_6776 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_249_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_125_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_249_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_251 = 10'sh7e - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_251 = $signed(s1_ghv_wens_diff_251) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_502 = 10'sh7e - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_503 = s1_ghv_wens_reverse_flag_251 ? _s1_ghv_wens_new_ptr_value_T_502 : 10'h7e
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_251_value = _s1_ghv_wens_new_ptr_value_T_503[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_6803 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_251_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_125_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_251_value & _s1_predicted_ghist_ptr_T_45 &
    s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_6830 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_251_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_126_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_251_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_253 = 10'sh7f - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_253 = $signed(s1_ghv_wens_diff_253) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_506 = 10'sh7f - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_507 = s1_ghv_wens_reverse_flag_253 ? _s1_ghv_wens_new_ptr_value_T_506 : 10'h7f
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_253_value = _s1_ghv_wens_new_ptr_value_T_507[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_6857 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_253_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_126_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_253_value & _s1_predicted_ghist_ptr_T_45 &
    s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_6884 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_253_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_127_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_253_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_255 = 10'sh80 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_255 = $signed(s1_ghv_wens_diff_255) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_510 = 10'sh80 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_511 = s1_ghv_wens_reverse_flag_255 ? _s1_ghv_wens_new_ptr_value_T_510 : 10'h80
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_255_value = _s1_ghv_wens_new_ptr_value_T_511[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_6911 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_255_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_127_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_255_value & _s1_predicted_ghist_ptr_T_45 &
    s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_6938 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_255_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_128_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_255_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_257 = 10'sh81 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_257 = $signed(s1_ghv_wens_diff_257) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_514 = 10'sh81 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_515 = s1_ghv_wens_reverse_flag_257 ? _s1_ghv_wens_new_ptr_value_T_514 : 10'h81
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_257_value = _s1_ghv_wens_new_ptr_value_T_515[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_6965 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_257_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_128_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_257_value & _s1_predicted_ghist_ptr_T_45 &
    s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_6992 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_257_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_129_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_257_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_259 = 10'sh82 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_259 = $signed(s1_ghv_wens_diff_259) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_518 = 10'sh82 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_519 = s1_ghv_wens_reverse_flag_259 ? _s1_ghv_wens_new_ptr_value_T_518 : 10'h82
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_259_value = _s1_ghv_wens_new_ptr_value_T_519[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_7019 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_259_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_129_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_259_value & _s1_predicted_ghist_ptr_T_45 &
    s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_7046 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_259_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_130_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_259_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_261 = 10'sh83 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_261 = $signed(s1_ghv_wens_diff_261) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_522 = 10'sh83 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_523 = s1_ghv_wens_reverse_flag_261 ? _s1_ghv_wens_new_ptr_value_T_522 : 10'h83
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_261_value = _s1_ghv_wens_new_ptr_value_T_523[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_7073 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_261_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_130_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_261_value & _s1_predicted_ghist_ptr_T_45 &
    s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_7100 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_261_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_131_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_261_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_263 = 10'sh84 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_263 = $signed(s1_ghv_wens_diff_263) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_526 = 10'sh84 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_527 = s1_ghv_wens_reverse_flag_263 ? _s1_ghv_wens_new_ptr_value_T_526 : 10'h84
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_263_value = _s1_ghv_wens_new_ptr_value_T_527[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_7127 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_263_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_131_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_263_value & _s1_predicted_ghist_ptr_T_45 &
    s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_7154 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_263_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_132_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_263_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_265 = 10'sh85 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_265 = $signed(s1_ghv_wens_diff_265) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_530 = 10'sh85 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_531 = s1_ghv_wens_reverse_flag_265 ? _s1_ghv_wens_new_ptr_value_T_530 : 10'h85
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_265_value = _s1_ghv_wens_new_ptr_value_T_531[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_7181 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_265_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_132_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_265_value & _s1_predicted_ghist_ptr_T_45 &
    s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_7208 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_265_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_133_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_265_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_267 = 10'sh86 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_267 = $signed(s1_ghv_wens_diff_267) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_534 = 10'sh86 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_535 = s1_ghv_wens_reverse_flag_267 ? _s1_ghv_wens_new_ptr_value_T_534 : 10'h86
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_267_value = _s1_ghv_wens_new_ptr_value_T_535[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_7235 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_267_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_133_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_267_value & _s1_predicted_ghist_ptr_T_45 &
    s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_7262 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_267_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_134_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_267_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_269 = 10'sh87 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_269 = $signed(s1_ghv_wens_diff_269) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_538 = 10'sh87 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_539 = s1_ghv_wens_reverse_flag_269 ? _s1_ghv_wens_new_ptr_value_T_538 : 10'h87
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_269_value = _s1_ghv_wens_new_ptr_value_T_539[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_7289 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_269_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_134_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_269_value & _s1_predicted_ghist_ptr_T_45 &
    s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_7316 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_269_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_135_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_269_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_271 = 10'sh88 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_271 = $signed(s1_ghv_wens_diff_271) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_542 = 10'sh88 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_543 = s1_ghv_wens_reverse_flag_271 ? _s1_ghv_wens_new_ptr_value_T_542 : 10'h88
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_271_value = _s1_ghv_wens_new_ptr_value_T_543[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_7343 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_271_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_135_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_271_value & _s1_predicted_ghist_ptr_T_45 &
    s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_7370 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_271_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_136_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_271_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_273 = 10'sh89 - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_273 = $signed(s1_ghv_wens_diff_273) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_546 = 10'sh89 - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_547 = s1_ghv_wens_reverse_flag_273 ? _s1_ghv_wens_new_ptr_value_T_546 : 10'h89
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_273_value = _s1_ghv_wens_new_ptr_value_T_547[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_7397 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_273_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_136_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_273_value & _s1_predicted_ghist_ptr_T_45 &
    s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_7424 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_273_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_137_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_273_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_275 = 10'sh8a - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_275 = $signed(s1_ghv_wens_diff_275) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_550 = 10'sh8a - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_551 = s1_ghv_wens_reverse_flag_275 ? _s1_ghv_wens_new_ptr_value_T_550 : 10'h8a
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_275_value = _s1_ghv_wens_new_ptr_value_T_551[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_7451 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_275_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_137_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_275_value & _s1_predicted_ghist_ptr_T_45 &
    s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_7478 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_275_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_138_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_275_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_277 = 10'sh8b - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_277 = $signed(s1_ghv_wens_diff_277) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_554 = 10'sh8b - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_555 = s1_ghv_wens_reverse_flag_277 ? _s1_ghv_wens_new_ptr_value_T_554 : 10'h8b
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_277_value = _s1_ghv_wens_new_ptr_value_T_555[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_7505 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_277_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_138_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_277_value & _s1_predicted_ghist_ptr_T_45 &
    s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_7532 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_277_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_139_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_277_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_279 = 10'sh8c - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_279 = $signed(s1_ghv_wens_diff_279) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_558 = 10'sh8c - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_559 = s1_ghv_wens_reverse_flag_279 ? _s1_ghv_wens_new_ptr_value_T_558 : 10'h8c
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_279_value = _s1_ghv_wens_new_ptr_value_T_559[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_7559 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_279_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_139_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_279_value & _s1_predicted_ghist_ptr_T_45 &
    s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_7586 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_279_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_140_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_279_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_281 = 10'sh8d - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_281 = $signed(s1_ghv_wens_diff_281) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_562 = 10'sh8d - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_563 = s1_ghv_wens_reverse_flag_281 ? _s1_ghv_wens_new_ptr_value_T_562 : 10'h8d
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_281_value = _s1_ghv_wens_new_ptr_value_T_563[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_7613 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_281_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_140_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_281_value & _s1_predicted_ghist_ptr_T_45 &
    s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_7640 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_281_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_141_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_281_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_283 = 10'sh8e - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_283 = $signed(s1_ghv_wens_diff_283) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_566 = 10'sh8e - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_567 = s1_ghv_wens_reverse_flag_283 ? _s1_ghv_wens_new_ptr_value_T_566 : 10'h8e
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_283_value = _s1_ghv_wens_new_ptr_value_T_567[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_7667 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_283_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_141_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_283_value & _s1_predicted_ghist_ptr_T_45 &
    s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_7694 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_283_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_142_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_283_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire [9:0] s1_ghv_wens_diff_285 = 10'sh8f - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s1_ghv_wens_reverse_flag_285 = $signed(s1_ghv_wens_diff_285) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_570 = 10'sh8f - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s1_ghv_wens_new_ptr_value_T_571 = s1_ghv_wens_reverse_flag_285 ? _s1_ghv_wens_new_ptr_value_T_570 : 10'h8f
    ; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] s1_ghv_wens_new_ptr_285_value = _s1_ghv_wens_new_ptr_value_T_571[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _s1_ghv_wens_T_7721 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_285_value & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_142_1 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_285_value & _s1_predicted_ghist_ptr_T_45 &
    s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_7748 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_285_value & _s1_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_143_0 = s1_ghist_ptr_value == s1_ghv_wens_new_ptr_285_value & _s1_predicted_ghist_ptr_WIRE__0 &
    s1_valid; // @[BPU.scala 422:119]
  wire  _s1_ghv_wens_T_7775 = s1_ghist_ptr_value == 8'h0 & _s1_predicted_ghist_ptr_T_45; // @[BPU.scala 422:90]
  wire  s1_ghv_wens_143_1 = s1_ghist_ptr_value == 8'h0 & _s1_predicted_ghist_ptr_T_45 & s1_valid; // @[BPU.scala 422:119]
  wire [38:0] targetVec_3 = predictors_io_out_s1_pc + 39'h10; // @[FrontendBundle.scala 473:55]
  wire  selVecOH_1 = ~_s1_predicted_ghist_ptr_T_6 & _s1_predicted_ghist_ptr_T_10 & predictors_io_out_s1_full_pred_hit; // @[FrontendBundle.scala 476:80]
  wire [1:0] _selVecOH_T_5 = {_s1_predicted_ghist_ptr_T_10,_s1_predicted_ghist_ptr_T_6}; // @[FrontendBundle.scala 477:12]
  wire  selVecOH_2 = ~(|_selVecOH_T_5) & predictors_io_out_s1_full_pred_hit; // @[FrontendBundle.scala 477:23]
  wire [38:0] _T_54 = _s1_predicted_ghist_ptr_T_11 ? predictors_io_out_s1_full_pred_targets_0 : 39'h0; // @[Mux.scala 27:73]
  wire [38:0] _T_55 = selVecOH_1 ? predictors_io_out_s1_full_pred_targets_1 : 39'h0; // @[Mux.scala 27:73]
  wire [38:0] _T_56 = selVecOH_2 ? predictors_io_out_s1_full_pred_fallThroughAddr : 39'h0; // @[Mux.scala 27:73]
  wire [38:0] _T_57 = _s1_predicted_ghist_ptr_T ? targetVec_3 : 39'h0; // @[Mux.scala 27:73]
  wire [38:0] _T_58 = _T_54 | _T_55; // @[Mux.scala 27:73]
  wire [38:0] _T_59 = _T_58 | _T_56; // @[Mux.scala 27:73]
  wire [38:0] _T_60 = _T_59 | _T_57; // @[Mux.scala 27:73]
  wire [1:0] hi = {_s1_predicted_ghist_ptr_T_60,_s1_predicted_ghist_ptr_T_32}; // @[BPU.scala 435:57]
  wire [2:0] _T_122 = {_s1_predicted_ghist_ptr_T_60,_s1_predicted_ghist_ptr_T_32,_s1_predicted_ghist_ptr_T_4}; // @[BPU.scala 435:57]
  wire  _T_123 = s1_ghv_wens_0_0 | s1_ghv_wens_0_1; // @[BPU.scala 438:26]
  wire  _T_124 = s1_ghv_wens_1_0 | s1_ghv_wens_1_1; // @[BPU.scala 438:26]
  wire  _T_125 = s1_ghv_wens_2_0 | s1_ghv_wens_2_1; // @[BPU.scala 438:26]
  wire  _T_126 = s1_ghv_wens_3_0 | s1_ghv_wens_3_1; // @[BPU.scala 438:26]
  wire  _T_127 = s1_ghv_wens_4_0 | s1_ghv_wens_4_1; // @[BPU.scala 438:26]
  wire  _T_128 = s1_ghv_wens_5_0 | s1_ghv_wens_5_1; // @[BPU.scala 438:26]
  wire  _T_129 = s1_ghv_wens_6_0 | s1_ghv_wens_6_1; // @[BPU.scala 438:26]
  wire  _T_130 = s1_ghv_wens_7_0 | s1_ghv_wens_7_1; // @[BPU.scala 438:26]
  wire  _T_131 = s1_ghv_wens_8_0 | s1_ghv_wens_8_1; // @[BPU.scala 438:26]
  wire  _T_132 = s1_ghv_wens_9_0 | s1_ghv_wens_9_1; // @[BPU.scala 438:26]
  wire  _T_133 = s1_ghv_wens_10_0 | s1_ghv_wens_10_1; // @[BPU.scala 438:26]
  wire  _T_134 = s1_ghv_wens_11_0 | s1_ghv_wens_11_1; // @[BPU.scala 438:26]
  wire  _T_135 = s1_ghv_wens_12_0 | s1_ghv_wens_12_1; // @[BPU.scala 438:26]
  wire  _T_136 = s1_ghv_wens_13_0 | s1_ghv_wens_13_1; // @[BPU.scala 438:26]
  wire  _T_137 = s1_ghv_wens_14_0 | s1_ghv_wens_14_1; // @[BPU.scala 438:26]
  wire  _T_138 = s1_ghv_wens_15_0 | s1_ghv_wens_15_1; // @[BPU.scala 438:26]
  wire  _T_139 = s1_ghv_wens_16_0 | s1_ghv_wens_16_1; // @[BPU.scala 438:26]
  wire  _T_140 = s1_ghv_wens_17_0 | s1_ghv_wens_17_1; // @[BPU.scala 438:26]
  wire  _T_141 = s1_ghv_wens_18_0 | s1_ghv_wens_18_1; // @[BPU.scala 438:26]
  wire  _T_142 = s1_ghv_wens_19_0 | s1_ghv_wens_19_1; // @[BPU.scala 438:26]
  wire  _T_143 = s1_ghv_wens_20_0 | s1_ghv_wens_20_1; // @[BPU.scala 438:26]
  wire  _T_144 = s1_ghv_wens_21_0 | s1_ghv_wens_21_1; // @[BPU.scala 438:26]
  wire  _T_145 = s1_ghv_wens_22_0 | s1_ghv_wens_22_1; // @[BPU.scala 438:26]
  wire  _T_146 = s1_ghv_wens_23_0 | s1_ghv_wens_23_1; // @[BPU.scala 438:26]
  wire  _T_147 = s1_ghv_wens_24_0 | s1_ghv_wens_24_1; // @[BPU.scala 438:26]
  wire  _T_148 = s1_ghv_wens_25_0 | s1_ghv_wens_25_1; // @[BPU.scala 438:26]
  wire  _T_149 = s1_ghv_wens_26_0 | s1_ghv_wens_26_1; // @[BPU.scala 438:26]
  wire  _T_150 = s1_ghv_wens_27_0 | s1_ghv_wens_27_1; // @[BPU.scala 438:26]
  wire  _T_151 = s1_ghv_wens_28_0 | s1_ghv_wens_28_1; // @[BPU.scala 438:26]
  wire  _T_152 = s1_ghv_wens_29_0 | s1_ghv_wens_29_1; // @[BPU.scala 438:26]
  wire  _T_153 = s1_ghv_wens_30_0 | s1_ghv_wens_30_1; // @[BPU.scala 438:26]
  wire  _T_154 = s1_ghv_wens_31_0 | s1_ghv_wens_31_1; // @[BPU.scala 438:26]
  wire  _T_155 = s1_ghv_wens_32_0 | s1_ghv_wens_32_1; // @[BPU.scala 438:26]
  wire  _T_156 = s1_ghv_wens_33_0 | s1_ghv_wens_33_1; // @[BPU.scala 438:26]
  wire  _T_157 = s1_ghv_wens_34_0 | s1_ghv_wens_34_1; // @[BPU.scala 438:26]
  wire  _T_158 = s1_ghv_wens_35_0 | s1_ghv_wens_35_1; // @[BPU.scala 438:26]
  wire  _T_159 = s1_ghv_wens_36_0 | s1_ghv_wens_36_1; // @[BPU.scala 438:26]
  wire  _T_160 = s1_ghv_wens_37_0 | s1_ghv_wens_37_1; // @[BPU.scala 438:26]
  wire  _T_161 = s1_ghv_wens_38_0 | s1_ghv_wens_38_1; // @[BPU.scala 438:26]
  wire  _T_162 = s1_ghv_wens_39_0 | s1_ghv_wens_39_1; // @[BPU.scala 438:26]
  wire  _T_163 = s1_ghv_wens_40_0 | s1_ghv_wens_40_1; // @[BPU.scala 438:26]
  wire  _T_164 = s1_ghv_wens_41_0 | s1_ghv_wens_41_1; // @[BPU.scala 438:26]
  wire  _T_165 = s1_ghv_wens_42_0 | s1_ghv_wens_42_1; // @[BPU.scala 438:26]
  wire  _T_166 = s1_ghv_wens_43_0 | s1_ghv_wens_43_1; // @[BPU.scala 438:26]
  wire  _T_167 = s1_ghv_wens_44_0 | s1_ghv_wens_44_1; // @[BPU.scala 438:26]
  wire  _T_168 = s1_ghv_wens_45_0 | s1_ghv_wens_45_1; // @[BPU.scala 438:26]
  wire  _T_169 = s1_ghv_wens_46_0 | s1_ghv_wens_46_1; // @[BPU.scala 438:26]
  wire  _T_170 = s1_ghv_wens_47_0 | s1_ghv_wens_47_1; // @[BPU.scala 438:26]
  wire  _T_171 = s1_ghv_wens_48_0 | s1_ghv_wens_48_1; // @[BPU.scala 438:26]
  wire  _T_172 = s1_ghv_wens_49_0 | s1_ghv_wens_49_1; // @[BPU.scala 438:26]
  wire  _T_173 = s1_ghv_wens_50_0 | s1_ghv_wens_50_1; // @[BPU.scala 438:26]
  wire  _T_174 = s1_ghv_wens_51_0 | s1_ghv_wens_51_1; // @[BPU.scala 438:26]
  wire  _T_175 = s1_ghv_wens_52_0 | s1_ghv_wens_52_1; // @[BPU.scala 438:26]
  wire  _T_176 = s1_ghv_wens_53_0 | s1_ghv_wens_53_1; // @[BPU.scala 438:26]
  wire  _T_177 = s1_ghv_wens_54_0 | s1_ghv_wens_54_1; // @[BPU.scala 438:26]
  wire  _T_178 = s1_ghv_wens_55_0 | s1_ghv_wens_55_1; // @[BPU.scala 438:26]
  wire  _T_179 = s1_ghv_wens_56_0 | s1_ghv_wens_56_1; // @[BPU.scala 438:26]
  wire  _T_180 = s1_ghv_wens_57_0 | s1_ghv_wens_57_1; // @[BPU.scala 438:26]
  wire  _T_181 = s1_ghv_wens_58_0 | s1_ghv_wens_58_1; // @[BPU.scala 438:26]
  wire  _T_182 = s1_ghv_wens_59_0 | s1_ghv_wens_59_1; // @[BPU.scala 438:26]
  wire  _T_183 = s1_ghv_wens_60_0 | s1_ghv_wens_60_1; // @[BPU.scala 438:26]
  wire  _T_184 = s1_ghv_wens_61_0 | s1_ghv_wens_61_1; // @[BPU.scala 438:26]
  wire  _T_185 = s1_ghv_wens_62_0 | s1_ghv_wens_62_1; // @[BPU.scala 438:26]
  wire  _T_186 = s1_ghv_wens_63_0 | s1_ghv_wens_63_1; // @[BPU.scala 438:26]
  wire  _T_187 = s1_ghv_wens_64_0 | s1_ghv_wens_64_1; // @[BPU.scala 438:26]
  wire  _T_188 = s1_ghv_wens_65_0 | s1_ghv_wens_65_1; // @[BPU.scala 438:26]
  wire  _T_189 = s1_ghv_wens_66_0 | s1_ghv_wens_66_1; // @[BPU.scala 438:26]
  wire  _T_190 = s1_ghv_wens_67_0 | s1_ghv_wens_67_1; // @[BPU.scala 438:26]
  wire  _T_191 = s1_ghv_wens_68_0 | s1_ghv_wens_68_1; // @[BPU.scala 438:26]
  wire  _T_192 = s1_ghv_wens_69_0 | s1_ghv_wens_69_1; // @[BPU.scala 438:26]
  wire  _T_193 = s1_ghv_wens_70_0 | s1_ghv_wens_70_1; // @[BPU.scala 438:26]
  wire  _T_194 = s1_ghv_wens_71_0 | s1_ghv_wens_71_1; // @[BPU.scala 438:26]
  wire  _T_195 = s1_ghv_wens_72_0 | s1_ghv_wens_72_1; // @[BPU.scala 438:26]
  wire  _T_196 = s1_ghv_wens_73_0 | s1_ghv_wens_73_1; // @[BPU.scala 438:26]
  wire  _T_197 = s1_ghv_wens_74_0 | s1_ghv_wens_74_1; // @[BPU.scala 438:26]
  wire  _T_198 = s1_ghv_wens_75_0 | s1_ghv_wens_75_1; // @[BPU.scala 438:26]
  wire  _T_199 = s1_ghv_wens_76_0 | s1_ghv_wens_76_1; // @[BPU.scala 438:26]
  wire  _T_200 = s1_ghv_wens_77_0 | s1_ghv_wens_77_1; // @[BPU.scala 438:26]
  wire  _T_201 = s1_ghv_wens_78_0 | s1_ghv_wens_78_1; // @[BPU.scala 438:26]
  wire  _T_202 = s1_ghv_wens_79_0 | s1_ghv_wens_79_1; // @[BPU.scala 438:26]
  wire  _T_203 = s1_ghv_wens_80_0 | s1_ghv_wens_80_1; // @[BPU.scala 438:26]
  wire  _T_204 = s1_ghv_wens_81_0 | s1_ghv_wens_81_1; // @[BPU.scala 438:26]
  wire  _T_205 = s1_ghv_wens_82_0 | s1_ghv_wens_82_1; // @[BPU.scala 438:26]
  wire  _T_206 = s1_ghv_wens_83_0 | s1_ghv_wens_83_1; // @[BPU.scala 438:26]
  wire  _T_207 = s1_ghv_wens_84_0 | s1_ghv_wens_84_1; // @[BPU.scala 438:26]
  wire  _T_208 = s1_ghv_wens_85_0 | s1_ghv_wens_85_1; // @[BPU.scala 438:26]
  wire  _T_209 = s1_ghv_wens_86_0 | s1_ghv_wens_86_1; // @[BPU.scala 438:26]
  wire  _T_210 = s1_ghv_wens_87_0 | s1_ghv_wens_87_1; // @[BPU.scala 438:26]
  wire  _T_211 = s1_ghv_wens_88_0 | s1_ghv_wens_88_1; // @[BPU.scala 438:26]
  wire  _T_212 = s1_ghv_wens_89_0 | s1_ghv_wens_89_1; // @[BPU.scala 438:26]
  wire  _T_213 = s1_ghv_wens_90_0 | s1_ghv_wens_90_1; // @[BPU.scala 438:26]
  wire  _T_214 = s1_ghv_wens_91_0 | s1_ghv_wens_91_1; // @[BPU.scala 438:26]
  wire  _T_215 = s1_ghv_wens_92_0 | s1_ghv_wens_92_1; // @[BPU.scala 438:26]
  wire  _T_216 = s1_ghv_wens_93_0 | s1_ghv_wens_93_1; // @[BPU.scala 438:26]
  wire  _T_217 = s1_ghv_wens_94_0 | s1_ghv_wens_94_1; // @[BPU.scala 438:26]
  wire  _T_218 = s1_ghv_wens_95_0 | s1_ghv_wens_95_1; // @[BPU.scala 438:26]
  wire  _T_219 = s1_ghv_wens_96_0 | s1_ghv_wens_96_1; // @[BPU.scala 438:26]
  wire  _T_220 = s1_ghv_wens_97_0 | s1_ghv_wens_97_1; // @[BPU.scala 438:26]
  wire  _T_221 = s1_ghv_wens_98_0 | s1_ghv_wens_98_1; // @[BPU.scala 438:26]
  wire  _T_222 = s1_ghv_wens_99_0 | s1_ghv_wens_99_1; // @[BPU.scala 438:26]
  wire  _T_223 = s1_ghv_wens_100_0 | s1_ghv_wens_100_1; // @[BPU.scala 438:26]
  wire  _T_224 = s1_ghv_wens_101_0 | s1_ghv_wens_101_1; // @[BPU.scala 438:26]
  wire  _T_225 = s1_ghv_wens_102_0 | s1_ghv_wens_102_1; // @[BPU.scala 438:26]
  wire  _T_226 = s1_ghv_wens_103_0 | s1_ghv_wens_103_1; // @[BPU.scala 438:26]
  wire  _T_227 = s1_ghv_wens_104_0 | s1_ghv_wens_104_1; // @[BPU.scala 438:26]
  wire  _T_228 = s1_ghv_wens_105_0 | s1_ghv_wens_105_1; // @[BPU.scala 438:26]
  wire  _T_229 = s1_ghv_wens_106_0 | s1_ghv_wens_106_1; // @[BPU.scala 438:26]
  wire  _T_230 = s1_ghv_wens_107_0 | s1_ghv_wens_107_1; // @[BPU.scala 438:26]
  wire  _T_231 = s1_ghv_wens_108_0 | s1_ghv_wens_108_1; // @[BPU.scala 438:26]
  wire  _T_232 = s1_ghv_wens_109_0 | s1_ghv_wens_109_1; // @[BPU.scala 438:26]
  wire  _T_233 = s1_ghv_wens_110_0 | s1_ghv_wens_110_1; // @[BPU.scala 438:26]
  wire  _T_234 = s1_ghv_wens_111_0 | s1_ghv_wens_111_1; // @[BPU.scala 438:26]
  wire  _T_235 = s1_ghv_wens_112_0 | s1_ghv_wens_112_1; // @[BPU.scala 438:26]
  wire  _T_236 = s1_ghv_wens_113_0 | s1_ghv_wens_113_1; // @[BPU.scala 438:26]
  wire  _T_237 = s1_ghv_wens_114_0 | s1_ghv_wens_114_1; // @[BPU.scala 438:26]
  wire  _T_238 = s1_ghv_wens_115_0 | s1_ghv_wens_115_1; // @[BPU.scala 438:26]
  wire  _T_239 = s1_ghv_wens_116_0 | s1_ghv_wens_116_1; // @[BPU.scala 438:26]
  wire  _T_240 = s1_ghv_wens_117_0 | s1_ghv_wens_117_1; // @[BPU.scala 438:26]
  wire  _T_241 = s1_ghv_wens_118_0 | s1_ghv_wens_118_1; // @[BPU.scala 438:26]
  wire  _T_242 = s1_ghv_wens_119_0 | s1_ghv_wens_119_1; // @[BPU.scala 438:26]
  wire  _T_243 = s1_ghv_wens_120_0 | s1_ghv_wens_120_1; // @[BPU.scala 438:26]
  wire  _T_244 = s1_ghv_wens_121_0 | s1_ghv_wens_121_1; // @[BPU.scala 438:26]
  wire  _T_245 = s1_ghv_wens_122_0 | s1_ghv_wens_122_1; // @[BPU.scala 438:26]
  wire  _T_246 = s1_ghv_wens_123_0 | s1_ghv_wens_123_1; // @[BPU.scala 438:26]
  wire  _T_247 = s1_ghv_wens_124_0 | s1_ghv_wens_124_1; // @[BPU.scala 438:26]
  wire  _T_248 = s1_ghv_wens_125_0 | s1_ghv_wens_125_1; // @[BPU.scala 438:26]
  wire  _T_249 = s1_ghv_wens_126_0 | s1_ghv_wens_126_1; // @[BPU.scala 438:26]
  wire  _T_250 = s1_ghv_wens_127_0 | s1_ghv_wens_127_1; // @[BPU.scala 438:26]
  wire  _T_251 = s1_ghv_wens_128_0 | s1_ghv_wens_128_1; // @[BPU.scala 438:26]
  wire  _T_252 = s1_ghv_wens_129_0 | s1_ghv_wens_129_1; // @[BPU.scala 438:26]
  wire  _T_253 = s1_ghv_wens_130_0 | s1_ghv_wens_130_1; // @[BPU.scala 438:26]
  wire  _T_254 = s1_ghv_wens_131_0 | s1_ghv_wens_131_1; // @[BPU.scala 438:26]
  wire  _T_255 = s1_ghv_wens_132_0 | s1_ghv_wens_132_1; // @[BPU.scala 438:26]
  wire  _T_256 = s1_ghv_wens_133_0 | s1_ghv_wens_133_1; // @[BPU.scala 438:26]
  wire  _T_257 = s1_ghv_wens_134_0 | s1_ghv_wens_134_1; // @[BPU.scala 438:26]
  wire  _T_258 = s1_ghv_wens_135_0 | s1_ghv_wens_135_1; // @[BPU.scala 438:26]
  wire  _T_259 = s1_ghv_wens_136_0 | s1_ghv_wens_136_1; // @[BPU.scala 438:26]
  wire  _T_260 = s1_ghv_wens_137_0 | s1_ghv_wens_137_1; // @[BPU.scala 438:26]
  wire  _T_261 = s1_ghv_wens_138_0 | s1_ghv_wens_138_1; // @[BPU.scala 438:26]
  wire  _T_262 = s1_ghv_wens_139_0 | s1_ghv_wens_139_1; // @[BPU.scala 438:26]
  wire  _T_263 = s1_ghv_wens_140_0 | s1_ghv_wens_140_1; // @[BPU.scala 438:26]
  wire  _T_264 = s1_ghv_wens_141_0 | s1_ghv_wens_141_1; // @[BPU.scala 438:26]
  wire  _T_265 = s1_ghv_wens_142_0 | s1_ghv_wens_142_1; // @[BPU.scala 438:26]
  wire  _T_266 = s1_ghv_wens_143_0 | s1_ghv_wens_143_1; // @[BPU.scala 438:26]
  wire [8:0] s2_possible_predicted_ghist_ptrs_flipped_new_ptr_new_value = s2_ghist_ptr_value +
    _s1_possible_predicted_ghist_ptrs_flipped_new_ptr_T_1; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _s2_possible_predicted_ghist_ptrs_flipped_new_ptr_diff_T_1 = {1'h0,
    s2_possible_predicted_ghist_ptrs_flipped_new_ptr_new_value}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] s2_possible_predicted_ghist_ptrs_flipped_new_ptr_diff = $signed(
    _s2_possible_predicted_ghist_ptrs_flipped_new_ptr_diff_T_1) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s2_possible_predicted_ghist_ptrs_flipped_new_ptr_reverse_flag = $signed(
    s2_possible_predicted_ghist_ptrs_flipped_new_ptr_diff) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire  s2_possible_predicted_ghist_ptrs_flipped_new_ptr_flag =
    s2_possible_predicted_ghist_ptrs_flipped_new_ptr_reverse_flag ? ~s2_ghist_ptr_flag : s2_ghist_ptr_flag; // @[CircularQueuePtr.scala 44:26]
  wire [9:0] _s2_possible_predicted_ghist_ptrs_flipped_new_ptr_new_ptr_value_T = $signed(
    _s2_possible_predicted_ghist_ptrs_flipped_new_ptr_diff_T_1) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s2_possible_predicted_ghist_ptrs_flipped_new_ptr_new_ptr_value_T_1 =
    s2_possible_predicted_ghist_ptrs_flipped_new_ptr_reverse_flag ?
    _s2_possible_predicted_ghist_ptrs_flipped_new_ptr_new_ptr_value_T : {{1'd0},
    s2_possible_predicted_ghist_ptrs_flipped_new_ptr_new_value}; // @[CircularQueuePtr.scala 45:27]
  wire  s2_possible_predicted_ghist_ptrs_0_flag = ~s2_possible_predicted_ghist_ptrs_flipped_new_ptr_flag; // @[CircularQueuePtr.scala 56:21]
  wire [8:0] s2_possible_predicted_ghist_ptrs_flipped_new_ptr_new_value_1 = s2_ghist_ptr_value +
    _s1_possible_predicted_ghist_ptrs_flipped_new_ptr_T_3; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _s2_possible_predicted_ghist_ptrs_flipped_new_ptr_diff_T_7 = {1'h0,
    s2_possible_predicted_ghist_ptrs_flipped_new_ptr_new_value_1}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] s2_possible_predicted_ghist_ptrs_flipped_new_ptr_diff_1 = $signed(
    _s2_possible_predicted_ghist_ptrs_flipped_new_ptr_diff_T_7) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s2_possible_predicted_ghist_ptrs_flipped_new_ptr_reverse_flag_1 = $signed(
    s2_possible_predicted_ghist_ptrs_flipped_new_ptr_diff_1) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire  s2_possible_predicted_ghist_ptrs_flipped_new_ptr_1_flag =
    s2_possible_predicted_ghist_ptrs_flipped_new_ptr_reverse_flag_1 ? ~s2_ghist_ptr_flag : s2_ghist_ptr_flag; // @[CircularQueuePtr.scala 44:26]
  wire [9:0] _s2_possible_predicted_ghist_ptrs_flipped_new_ptr_new_ptr_value_T_2 = $signed(
    _s2_possible_predicted_ghist_ptrs_flipped_new_ptr_diff_T_7) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s2_possible_predicted_ghist_ptrs_flipped_new_ptr_new_ptr_value_T_3 =
    s2_possible_predicted_ghist_ptrs_flipped_new_ptr_reverse_flag_1 ?
    _s2_possible_predicted_ghist_ptrs_flipped_new_ptr_new_ptr_value_T_2 : {{1'd0},
    s2_possible_predicted_ghist_ptrs_flipped_new_ptr_new_value_1}; // @[CircularQueuePtr.scala 45:27]
  wire  s2_possible_predicted_ghist_ptrs_1_flag = ~s2_possible_predicted_ghist_ptrs_flipped_new_ptr_1_flag; // @[CircularQueuePtr.scala 56:21]
  wire [8:0] s2_possible_predicted_ghist_ptrs_flipped_new_ptr_new_value_2 = s2_ghist_ptr_value +
    _s1_possible_predicted_ghist_ptrs_flipped_new_ptr_T_5; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _s2_possible_predicted_ghist_ptrs_flipped_new_ptr_diff_T_13 = {1'h0,
    s2_possible_predicted_ghist_ptrs_flipped_new_ptr_new_value_2}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] s2_possible_predicted_ghist_ptrs_flipped_new_ptr_diff_2 = $signed(
    _s2_possible_predicted_ghist_ptrs_flipped_new_ptr_diff_T_13) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s2_possible_predicted_ghist_ptrs_flipped_new_ptr_reverse_flag_2 = $signed(
    s2_possible_predicted_ghist_ptrs_flipped_new_ptr_diff_2) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire  s2_possible_predicted_ghist_ptrs_flipped_new_ptr_2_flag =
    s2_possible_predicted_ghist_ptrs_flipped_new_ptr_reverse_flag_2 ? ~s2_ghist_ptr_flag : s2_ghist_ptr_flag; // @[CircularQueuePtr.scala 44:26]
  wire [9:0] _s2_possible_predicted_ghist_ptrs_flipped_new_ptr_new_ptr_value_T_4 = $signed(
    _s2_possible_predicted_ghist_ptrs_flipped_new_ptr_diff_T_13) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s2_possible_predicted_ghist_ptrs_flipped_new_ptr_new_ptr_value_T_5 =
    s2_possible_predicted_ghist_ptrs_flipped_new_ptr_reverse_flag_2 ?
    _s2_possible_predicted_ghist_ptrs_flipped_new_ptr_new_ptr_value_T_4 : {{1'd0},
    s2_possible_predicted_ghist_ptrs_flipped_new_ptr_new_value_2}; // @[CircularQueuePtr.scala 45:27]
  wire  s2_possible_predicted_ghist_ptrs_2_flag = ~s2_possible_predicted_ghist_ptrs_flipped_new_ptr_2_flag; // @[CircularQueuePtr.scala 56:21]
  wire [7:0] s2_possible_predicted_ghist_ptrs_flipped_new_ptr_value =
    _s2_possible_predicted_ghist_ptrs_flipped_new_ptr_new_ptr_value_T_1[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire [7:0] _s2_predicted_ghist_ptr_T_61 = _s2_redirect_s1_last_pred_vec_T_12 ?
    s2_possible_predicted_ghist_ptrs_flipped_new_ptr_value : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] s2_possible_predicted_ghist_ptrs_flipped_new_ptr_1_value =
    _s2_possible_predicted_ghist_ptrs_flipped_new_ptr_new_ptr_value_T_3[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire [7:0] _s2_predicted_ghist_ptr_T_62 = _s2_redirect_s1_last_pred_vec_T_40 ?
    s2_possible_predicted_ghist_ptrs_flipped_new_ptr_1_value : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] s2_possible_predicted_ghist_ptrs_flipped_new_ptr_2_value =
    _s2_possible_predicted_ghist_ptrs_flipped_new_ptr_new_ptr_value_T_5[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire [7:0] _s2_predicted_ghist_ptr_T_63 = _s2_redirect_s1_last_pred_vec_T_68 ?
    s2_possible_predicted_ghist_ptrs_flipped_new_ptr_2_value : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _s2_predicted_ghist_ptr_T_64 = _s2_predicted_ghist_ptr_T_61 | _s2_predicted_ghist_ptr_T_62; // @[Mux.scala 27:73]
  wire  s2_possible_predicted_fhs_ob__0 = s2_last_br_num_oh[0] & s2_ahead_fh_oldest_bits_afhob_3_bits_0 |
    s2_last_br_num_oh[1] & s2_ahead_fh_oldest_bits_afhob_3_bits_1 | s2_last_br_num_oh[2] &
    s2_ahead_fh_oldest_bits_afhob_3_bits_2; // @[Mux.scala 27:73]
  wire  s2_possible_predicted_fhs_ob__1 = s2_last_br_num_oh[0] & s2_ahead_fh_oldest_bits_afhob_3_bits_1 |
    s2_last_br_num_oh[1] & s2_ahead_fh_oldest_bits_afhob_3_bits_2 | s2_last_br_num_oh[2] &
    s2_ahead_fh_oldest_bits_afhob_3_bits_3; // @[Mux.scala 27:73]
  wire  s2_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__0 = s2_folded_gh_hist_0_folded_hist[0
    ]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__1 = s2_folded_gh_hist_0_folded_hist[1
    ]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__2 = s2_folded_gh_hist_0_folded_hist[2
    ]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__3 = s2_folded_gh_hist_0_folded_hist[3
    ]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__4 = s2_folded_gh_hist_0_folded_hist[4
    ]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__5 = s2_folded_gh_hist_0_folded_hist[5
    ]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__6 = s2_folded_gh_hist_0_folded_hist[6
    ]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__7 = s2_folded_gh_hist_0_folded_hist[7
    ]; // @[FrontendBundle.scala 280:54]
  wire [7:0] s2_possible_predicted_fhs_res_hist_0_new_folded_hist_xored = {
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__7,
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__6,
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__5,
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__4,
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__3,
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__1,
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [15:0] s2_possible_predicted_fhs_res_hist_0_new_folded_hist_src_doubled = {
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__7,
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__6,
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__5,
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__4,
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__3,
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__1,
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__0,
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_xored}; // @[Cat.scala 31:58]
  wire [7:0] s2_possible_predicted_fhs_res_hist_0_new_folded_hist =
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_src_doubled[15:8]; // @[FrontendBundle.scala 221:30]
  wire  s2_possible_predicted_fhs_ob_1_0 = s2_last_br_num_oh[0] & s2_ahead_fh_oldest_bits_afhob_2_bits_0 |
    s2_last_br_num_oh[1] & s2_ahead_fh_oldest_bits_afhob_2_bits_1 | s2_last_br_num_oh[2] &
    s2_ahead_fh_oldest_bits_afhob_2_bits_2; // @[Mux.scala 27:73]
  wire  s2_possible_predicted_fhs_ob_1_1 = s2_last_br_num_oh[0] & s2_ahead_fh_oldest_bits_afhob_2_bits_1 |
    s2_last_br_num_oh[1] & s2_ahead_fh_oldest_bits_afhob_2_bits_2 | s2_last_br_num_oh[2] &
    s2_ahead_fh_oldest_bits_afhob_2_bits_3; // @[Mux.scala 27:73]
  wire  s2_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__0 = s2_folded_gh_hist_1_folded_hist[0
    ]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__1 = s2_folded_gh_hist_1_folded_hist[1
    ]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__2 = s2_folded_gh_hist_1_folded_hist[2
    ]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__3 = s2_folded_gh_hist_1_folded_hist[3
    ]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__4 = s2_folded_gh_hist_1_folded_hist[4
    ]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__5 = s2_folded_gh_hist_1_folded_hist[5
    ]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__6 = s2_folded_gh_hist_1_folded_hist[6
    ]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__7 = s2_folded_gh_hist_1_folded_hist[7
    ]; // @[FrontendBundle.scala 280:54]
  wire [7:0] s2_possible_predicted_fhs_res_hist_1_new_folded_hist_xored = {
    s2_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__7,
    s2_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__6,
    s2_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__5,
    s2_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__4,
    s2_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__3,
    s2_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__1,
    s2_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [15:0] s2_possible_predicted_fhs_res_hist_1_new_folded_hist_src_doubled = {
    s2_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__7,
    s2_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__6,
    s2_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__5,
    s2_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__4,
    s2_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__3,
    s2_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__1,
    s2_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__0,
    s2_possible_predicted_fhs_res_hist_1_new_folded_hist_xored}; // @[Cat.scala 31:58]
  wire [7:0] s2_possible_predicted_fhs_res_hist_1_new_folded_hist =
    s2_possible_predicted_fhs_res_hist_1_new_folded_hist_src_doubled[15:8]; // @[FrontendBundle.scala 221:30]
  wire  s2_possible_predicted_fhs_ob_2_0 = s2_last_br_num_oh[0] & s2_ahead_fh_oldest_bits_afhob_5_bits_0 |
    s2_last_br_num_oh[1] & s2_ahead_fh_oldest_bits_afhob_5_bits_1 | s2_last_br_num_oh[2] &
    s2_ahead_fh_oldest_bits_afhob_5_bits_2; // @[Mux.scala 27:73]
  wire  s2_possible_predicted_fhs_ob_2_1 = s2_last_br_num_oh[0] & s2_ahead_fh_oldest_bits_afhob_5_bits_1 |
    s2_last_br_num_oh[1] & s2_ahead_fh_oldest_bits_afhob_5_bits_2 | s2_last_br_num_oh[2] &
    s2_ahead_fh_oldest_bits_afhob_5_bits_3; // @[Mux.scala 27:73]
  wire  s2_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__0 = s2_folded_gh_hist_2_folded_hist[0
    ]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__1 = s2_folded_gh_hist_2_folded_hist[1
    ]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__2 = s2_folded_gh_hist_2_folded_hist[2
    ]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__3 = s2_folded_gh_hist_2_folded_hist[3
    ]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__4 = s2_folded_gh_hist_2_folded_hist[4
    ]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__5 = s2_folded_gh_hist_2_folded_hist[5
    ]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__6 = s2_folded_gh_hist_2_folded_hist[6
    ]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__7 = s2_folded_gh_hist_2_folded_hist[7
    ]; // @[FrontendBundle.scala 280:54]
  wire [7:0] s2_possible_predicted_fhs_res_hist_2_new_folded_hist_xored = {
    s2_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__7,
    s2_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__6,
    s2_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__5,
    s2_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__4,
    s2_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__3,
    s2_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__1,
    s2_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [15:0] s2_possible_predicted_fhs_res_hist_2_new_folded_hist_src_doubled = {
    s2_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__7,
    s2_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__6,
    s2_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__5,
    s2_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__4,
    s2_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__3,
    s2_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__1,
    s2_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__0,
    s2_possible_predicted_fhs_res_hist_2_new_folded_hist_xored}; // @[Cat.scala 31:58]
  wire [7:0] s2_possible_predicted_fhs_res_hist_2_new_folded_hist =
    s2_possible_predicted_fhs_res_hist_2_new_folded_hist_src_doubled[15:8]; // @[FrontendBundle.scala 221:30]
  wire  s2_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__0 = s2_folded_gh_hist_3_folded_hist[0
    ]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__1 = s2_folded_gh_hist_3_folded_hist[1
    ]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__2 = s2_folded_gh_hist_3_folded_hist[2
    ]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__3 = s2_folded_gh_hist_3_folded_hist[3
    ]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__4 = s2_folded_gh_hist_3_folded_hist[4
    ]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__5 = s2_folded_gh_hist_3_folded_hist[5
    ]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__6 = s2_folded_gh_hist_3_folded_hist[6
    ]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__7 = s2_folded_gh_hist_3_folded_hist[7
    ]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__8 = s2_folded_gh_hist_3_folded_hist[8
    ]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__9 = s2_folded_gh_hist_3_folded_hist[9
    ]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__10 = s2_folded_gh_hist_3_folded_hist[
    10]; // @[FrontendBundle.scala 280:54]
  wire [4:0] s2_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_lo = {
    s2_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__4,
    s2_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__3,
    s2_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__1,
    s2_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [10:0] s2_possible_predicted_fhs_res_hist_3_new_folded_hist_xored = {
    s2_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__10,
    s2_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__9,
    s2_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__8,
    s2_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__7,
    s2_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__6,
    s2_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__5,
    s2_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_lo}; // @[FrontendBundle.scala 258:11]
  wire [21:0] s2_possible_predicted_fhs_res_hist_3_new_folded_hist_src_doubled = {
    s2_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__10,
    s2_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__9,
    s2_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__8,
    s2_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__7,
    s2_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__6,
    s2_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__5,
    s2_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_lo,
    s2_possible_predicted_fhs_res_hist_3_new_folded_hist_xored}; // @[Cat.scala 31:58]
  wire [10:0] s2_possible_predicted_fhs_res_hist_3_new_folded_hist =
    s2_possible_predicted_fhs_res_hist_3_new_folded_hist_src_doubled[21:11]; // @[FrontendBundle.scala 221:30]
  wire  s2_possible_predicted_fhs_ob_4_0 = s2_last_br_num_oh[0] & s2_ahead_fh_oldest_bits_afhob_1_bits_0 |
    s2_last_br_num_oh[1] & s2_ahead_fh_oldest_bits_afhob_1_bits_1 | s2_last_br_num_oh[2] &
    s2_ahead_fh_oldest_bits_afhob_1_bits_2; // @[Mux.scala 27:73]
  wire  s2_possible_predicted_fhs_ob_4_1 = s2_last_br_num_oh[0] & s2_ahead_fh_oldest_bits_afhob_1_bits_1 |
    s2_last_br_num_oh[1] & s2_ahead_fh_oldest_bits_afhob_1_bits_2 | s2_last_br_num_oh[2] &
    s2_ahead_fh_oldest_bits_afhob_1_bits_3; // @[Mux.scala 27:73]
  wire  s2_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__0 = s2_folded_gh_hist_5_folded_hist[0
    ]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__1 = s2_folded_gh_hist_5_folded_hist[1
    ]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__2 = s2_folded_gh_hist_5_folded_hist[2
    ]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__3 = s2_folded_gh_hist_5_folded_hist[3
    ]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__4 = s2_folded_gh_hist_5_folded_hist[4
    ]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__5 = s2_folded_gh_hist_5_folded_hist[5
    ]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__6 = s2_folded_gh_hist_5_folded_hist[6
    ]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__7 = s2_folded_gh_hist_5_folded_hist[7
    ]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__8 = s2_folded_gh_hist_5_folded_hist[8
    ]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__9 = s2_folded_gh_hist_5_folded_hist[9
    ]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__10 = s2_folded_gh_hist_5_folded_hist[
    10]; // @[FrontendBundle.scala 280:54]
  wire [4:0] s2_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_lo = {
    s2_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__4,
    s2_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__3,
    s2_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__1,
    s2_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [10:0] s2_possible_predicted_fhs_res_hist_5_new_folded_hist_xored = {
    s2_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__10,
    s2_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__9,
    s2_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__8,
    s2_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__7,
    s2_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__6,
    s2_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__5,
    s2_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_lo}; // @[FrontendBundle.scala 258:11]
  wire [21:0] s2_possible_predicted_fhs_res_hist_5_new_folded_hist_src_doubled = {
    s2_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__10,
    s2_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__9,
    s2_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__8,
    s2_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__7,
    s2_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__6,
    s2_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__5,
    s2_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_lo,
    s2_possible_predicted_fhs_res_hist_5_new_folded_hist_xored}; // @[Cat.scala 31:58]
  wire [10:0] s2_possible_predicted_fhs_res_hist_5_new_folded_hist =
    s2_possible_predicted_fhs_res_hist_5_new_folded_hist_src_doubled[21:11]; // @[FrontendBundle.scala 221:30]
  wire  s2_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__0 = s2_folded_gh_hist_6_folded_hist[0
    ]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__1 = s2_folded_gh_hist_6_folded_hist[1
    ]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__2 = s2_folded_gh_hist_6_folded_hist[2
    ]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__3 = s2_folded_gh_hist_6_folded_hist[3
    ]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__4 = s2_folded_gh_hist_6_folded_hist[4
    ]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__5 = s2_folded_gh_hist_6_folded_hist[5
    ]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__6 = s2_folded_gh_hist_6_folded_hist[6
    ]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__7 = s2_folded_gh_hist_6_folded_hist[7
    ]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__8 = s2_folded_gh_hist_6_folded_hist[8
    ]; // @[FrontendBundle.scala 280:54]
  wire [8:0] s2_possible_predicted_fhs_res_hist_6_new_folded_hist_xored = {
    s2_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__8,
    s2_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__7,
    s2_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__6,
    s2_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__5,
    s2_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__4,
    s2_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__3,
    s2_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__1,
    s2_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [17:0] s2_possible_predicted_fhs_res_hist_6_new_folded_hist_src_doubled = {
    s2_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__8,
    s2_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__7,
    s2_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__6,
    s2_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__5,
    s2_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__4,
    s2_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__3,
    s2_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__1,
    s2_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__0,
    s2_possible_predicted_fhs_res_hist_6_new_folded_hist_xored}; // @[Cat.scala 31:58]
  wire [8:0] s2_possible_predicted_fhs_res_hist_6_new_folded_hist =
    s2_possible_predicted_fhs_res_hist_6_new_folded_hist_src_doubled[17:9]; // @[FrontendBundle.scala 221:30]
  wire  s2_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__0 = s2_folded_gh_hist_7_folded_hist[0
    ]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__1 = s2_folded_gh_hist_7_folded_hist[1
    ]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__2 = s2_folded_gh_hist_7_folded_hist[2
    ]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__3 = s2_folded_gh_hist_7_folded_hist[3
    ]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__4 = s2_folded_gh_hist_7_folded_hist[4
    ]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__5 = s2_folded_gh_hist_7_folded_hist[5
    ]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__6 = s2_folded_gh_hist_7_folded_hist[6
    ]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__7 = s2_folded_gh_hist_7_folded_hist[7
    ]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__8 = s2_folded_gh_hist_7_folded_hist[8
    ]; // @[FrontendBundle.scala 280:54]
  wire [8:0] s2_possible_predicted_fhs_res_hist_7_new_folded_hist_xored = {
    s2_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__8,
    s2_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__7,
    s2_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__6,
    s2_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__5,
    s2_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__4,
    s2_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__3,
    s2_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__1,
    s2_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [17:0] s2_possible_predicted_fhs_res_hist_7_new_folded_hist_src_doubled = {
    s2_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__8,
    s2_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__7,
    s2_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__6,
    s2_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__5,
    s2_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__4,
    s2_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__3,
    s2_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__1,
    s2_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__0,
    s2_possible_predicted_fhs_res_hist_7_new_folded_hist_xored}; // @[Cat.scala 31:58]
  wire [8:0] s2_possible_predicted_fhs_res_hist_7_new_folded_hist =
    s2_possible_predicted_fhs_res_hist_7_new_folded_hist_src_doubled[17:9]; // @[FrontendBundle.scala 221:30]
  wire  s2_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__0 = s2_folded_gh_hist_9_folded_hist[0
    ]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__1 = s2_folded_gh_hist_9_folded_hist[1
    ]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__2 = s2_folded_gh_hist_9_folded_hist[2
    ]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__3 = s2_folded_gh_hist_9_folded_hist[3
    ]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__4 = s2_folded_gh_hist_9_folded_hist[4
    ]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__5 = s2_folded_gh_hist_9_folded_hist[5
    ]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__6 = s2_folded_gh_hist_9_folded_hist[6
    ]; // @[FrontendBundle.scala 280:54]
  wire [6:0] s2_possible_predicted_fhs_res_hist_9_new_folded_hist_xored = {
    s2_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__6,
    s2_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__5,
    s2_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__4,
    s2_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__3,
    s2_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__1,
    s2_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [13:0] s2_possible_predicted_fhs_res_hist_9_new_folded_hist_src_doubled = {
    s2_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__6,
    s2_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__5,
    s2_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__4,
    s2_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__3,
    s2_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__1,
    s2_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__0,
    s2_possible_predicted_fhs_res_hist_9_new_folded_hist_xored}; // @[Cat.scala 31:58]
  wire [6:0] s2_possible_predicted_fhs_res_hist_9_new_folded_hist =
    s2_possible_predicted_fhs_res_hist_9_new_folded_hist_src_doubled[13:7]; // @[FrontendBundle.scala 221:30]
  wire  s2_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__0 = s2_folded_gh_hist_10_folded_hist
    [0]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__1 = s2_folded_gh_hist_10_folded_hist
    [1]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__2 = s2_folded_gh_hist_10_folded_hist
    [2]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__3 = s2_folded_gh_hist_10_folded_hist
    [3]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__4 = s2_folded_gh_hist_10_folded_hist
    [4]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__5 = s2_folded_gh_hist_10_folded_hist
    [5]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__6 = s2_folded_gh_hist_10_folded_hist
    [6]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__7 = s2_folded_gh_hist_10_folded_hist
    [7]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__8 = s2_folded_gh_hist_10_folded_hist
    [8]; // @[FrontendBundle.scala 280:54]
  wire [8:0] s2_possible_predicted_fhs_res_hist_10_new_folded_hist_xored = {
    s2_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__8,
    s2_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__7,
    s2_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__6,
    s2_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__5,
    s2_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__4,
    s2_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__3,
    s2_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__1,
    s2_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [17:0] s2_possible_predicted_fhs_res_hist_10_new_folded_hist_src_doubled = {
    s2_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__8,
    s2_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__7,
    s2_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__6,
    s2_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__5,
    s2_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__4,
    s2_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__3,
    s2_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__1,
    s2_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__0,
    s2_possible_predicted_fhs_res_hist_10_new_folded_hist_xored}; // @[Cat.scala 31:58]
  wire [8:0] s2_possible_predicted_fhs_res_hist_10_new_folded_hist =
    s2_possible_predicted_fhs_res_hist_10_new_folded_hist_src_doubled[17:9]; // @[FrontendBundle.scala 221:30]
  wire  s2_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__0 = s2_folded_gh_hist_12_folded_hist
    [0]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__1 = s2_folded_gh_hist_12_folded_hist
    [1]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__2 = s2_folded_gh_hist_12_folded_hist
    [2]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__3 = s2_folded_gh_hist_12_folded_hist
    [3]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__4 = s2_folded_gh_hist_12_folded_hist
    [4]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__5 = s2_folded_gh_hist_12_folded_hist
    [5]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__6 = s2_folded_gh_hist_12_folded_hist
    [6]; // @[FrontendBundle.scala 280:54]
  wire [6:0] s2_possible_predicted_fhs_res_hist_12_new_folded_hist_xored = {
    s2_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__6,
    s2_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__5,
    s2_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__4,
    s2_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__3,
    s2_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__1,
    s2_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [13:0] s2_possible_predicted_fhs_res_hist_12_new_folded_hist_src_doubled = {
    s2_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__6,
    s2_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__5,
    s2_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__4,
    s2_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__3,
    s2_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__1,
    s2_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__0,
    s2_possible_predicted_fhs_res_hist_12_new_folded_hist_xored}; // @[Cat.scala 31:58]
  wire [6:0] s2_possible_predicted_fhs_res_hist_12_new_folded_hist =
    s2_possible_predicted_fhs_res_hist_12_new_folded_hist_src_doubled[13:7]; // @[FrontendBundle.scala 221:30]
  wire  s2_possible_predicted_fhs_ob_10_0 = s2_last_br_num_oh[0] & s2_ahead_fh_oldest_bits_afhob_4_bits_0 |
    s2_last_br_num_oh[1] & s2_ahead_fh_oldest_bits_afhob_4_bits_1 | s2_last_br_num_oh[2] &
    s2_ahead_fh_oldest_bits_afhob_4_bits_2; // @[Mux.scala 27:73]
  wire  s2_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__0 = s2_folded_gh_hist_13_folded_hist
    [0]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__1 = s2_folded_gh_hist_13_folded_hist
    [1]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__2 = s2_folded_gh_hist_13_folded_hist
    [2]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__3 = s2_folded_gh_hist_13_folded_hist
    [3]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__4 = s2_folded_gh_hist_13_folded_hist
    [4]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__5 = s2_folded_gh_hist_13_folded_hist
    [5]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__6 = s2_folded_gh_hist_13_folded_hist
    [6]; // @[FrontendBundle.scala 280:54]
  wire [6:0] s2_possible_predicted_fhs_res_hist_13_new_folded_hist_xored = {
    s2_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__6,
    s2_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__5,
    s2_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__4,
    s2_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__3,
    s2_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__1,
    s2_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [13:0] s2_possible_predicted_fhs_res_hist_13_new_folded_hist_src_doubled = {
    s2_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__6,
    s2_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__5,
    s2_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__4,
    s2_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__3,
    s2_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__1,
    s2_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__0,
    s2_possible_predicted_fhs_res_hist_13_new_folded_hist_xored}; // @[Cat.scala 31:58]
  wire [6:0] s2_possible_predicted_fhs_res_hist_13_new_folded_hist =
    s2_possible_predicted_fhs_res_hist_13_new_folded_hist_src_doubled[13:7]; // @[FrontendBundle.scala 221:30]
  wire  s2_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__0 = s2_folded_gh_hist_14_folded_hist
    [0]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__1 = s2_folded_gh_hist_14_folded_hist
    [1]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__2 = s2_folded_gh_hist_14_folded_hist
    [2]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__3 = s2_folded_gh_hist_14_folded_hist
    [3]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__4 = s2_folded_gh_hist_14_folded_hist
    [4]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__5 = s2_folded_gh_hist_14_folded_hist
    [5]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__6 = s2_folded_gh_hist_14_folded_hist
    [6]; // @[FrontendBundle.scala 280:54]
  wire [6:0] s2_possible_predicted_fhs_res_hist_14_new_folded_hist_xored = {
    s2_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__6,
    s2_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__5,
    s2_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__4,
    s2_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__3,
    s2_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__1,
    s2_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [13:0] s2_possible_predicted_fhs_res_hist_14_new_folded_hist_src_doubled = {
    s2_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__6,
    s2_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__5,
    s2_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__4,
    s2_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__3,
    s2_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__1,
    s2_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__0,
    s2_possible_predicted_fhs_res_hist_14_new_folded_hist_xored}; // @[Cat.scala 31:58]
  wire [6:0] s2_possible_predicted_fhs_res_hist_14_new_folded_hist =
    s2_possible_predicted_fhs_res_hist_14_new_folded_hist_src_doubled[13:7]; // @[FrontendBundle.scala 221:30]
  wire  s2_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__0 = s2_folded_gh_hist_15_folded_hist
    [0]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__1 = s2_folded_gh_hist_15_folded_hist
    [1]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__2 = s2_folded_gh_hist_15_folded_hist
    [2]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__3 = s2_folded_gh_hist_15_folded_hist
    [3]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__4 = s2_folded_gh_hist_15_folded_hist
    [4]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__5 = s2_folded_gh_hist_15_folded_hist
    [5]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__6 = s2_folded_gh_hist_15_folded_hist
    [6]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__7 = s2_folded_gh_hist_15_folded_hist
    [7]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__8 = s2_folded_gh_hist_15_folded_hist
    [8]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__9 = s2_folded_gh_hist_15_folded_hist
    [9]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__10 =
    s2_folded_gh_hist_15_folded_hist[10]; // @[FrontendBundle.scala 280:54]
  wire [4:0] s2_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_lo = {
    s2_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__4,
    s2_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__3,
    s2_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__1,
    s2_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [10:0] s2_possible_predicted_fhs_res_hist_15_new_folded_hist_xored = {
    s2_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__10,
    s2_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__9,
    s2_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__8,
    s2_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__7,
    s2_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__6,
    s2_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__5,
    s2_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_lo}; // @[FrontendBundle.scala 258:11]
  wire [21:0] s2_possible_predicted_fhs_res_hist_15_new_folded_hist_src_doubled = {
    s2_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__10,
    s2_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__9,
    s2_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__8,
    s2_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__7,
    s2_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__6,
    s2_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__5,
    s2_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_lo,
    s2_possible_predicted_fhs_res_hist_15_new_folded_hist_xored}; // @[Cat.scala 31:58]
  wire [10:0] s2_possible_predicted_fhs_res_hist_15_new_folded_hist =
    s2_possible_predicted_fhs_res_hist_15_new_folded_hist_src_doubled[21:11]; // @[FrontendBundle.scala 221:30]
  wire  s2_possible_predicted_fhs_ob_13_0 = s2_last_br_num_oh[0] & s2_ahead_fh_oldest_bits_afhob_0_bits_0 |
    s2_last_br_num_oh[1] & s2_ahead_fh_oldest_bits_afhob_0_bits_1 | s2_last_br_num_oh[2] &
    s2_ahead_fh_oldest_bits_afhob_0_bits_2; // @[Mux.scala 27:73]
  wire  s2_possible_predicted_fhs_ob_13_1 = s2_last_br_num_oh[0] & s2_ahead_fh_oldest_bits_afhob_0_bits_1 |
    s2_last_br_num_oh[1] & s2_ahead_fh_oldest_bits_afhob_0_bits_2 | s2_last_br_num_oh[2] &
    s2_ahead_fh_oldest_bits_afhob_0_bits_3; // @[Mux.scala 27:73]
  wire  s2_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__0 = s2_folded_gh_hist_16_folded_hist
    [0]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__1 = s2_folded_gh_hist_16_folded_hist
    [1]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__2 = s2_folded_gh_hist_16_folded_hist
    [2]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__3 = s2_folded_gh_hist_16_folded_hist
    [3]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__4 = s2_folded_gh_hist_16_folded_hist
    [4]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__5 = s2_folded_gh_hist_16_folded_hist
    [5]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__6 = s2_folded_gh_hist_16_folded_hist
    [6]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__7 = s2_folded_gh_hist_16_folded_hist
    [7]; // @[FrontendBundle.scala 280:54]
  wire [7:0] s2_possible_predicted_fhs_res_hist_16_new_folded_hist_xored = {
    s2_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__7,
    s2_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__6,
    s2_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__5,
    s2_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__4,
    s2_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__3,
    s2_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__1,
    s2_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [15:0] s2_possible_predicted_fhs_res_hist_16_new_folded_hist_src_doubled = {
    s2_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__7,
    s2_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__6,
    s2_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__5,
    s2_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__4,
    s2_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__3,
    s2_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__1,
    s2_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__0,
    s2_possible_predicted_fhs_res_hist_16_new_folded_hist_xored}; // @[Cat.scala 31:58]
  wire [7:0] s2_possible_predicted_fhs_res_hist_16_new_folded_hist =
    s2_possible_predicted_fhs_res_hist_16_new_folded_hist_src_doubled[15:8]; // @[FrontendBundle.scala 221:30]
  wire  s2_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__0 = s2_folded_gh_hist_17_folded_hist
    [0]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__1 = s2_folded_gh_hist_17_folded_hist
    [1]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__2 = s2_folded_gh_hist_17_folded_hist
    [2]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__3 = s2_folded_gh_hist_17_folded_hist
    [3]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__4 = s2_folded_gh_hist_17_folded_hist
    [4]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__5 = s2_folded_gh_hist_17_folded_hist
    [5]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__6 = s2_folded_gh_hist_17_folded_hist
    [6]; // @[FrontendBundle.scala 280:54]
  wire  s2_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__7 = s2_folded_gh_hist_17_folded_hist
    [7]; // @[FrontendBundle.scala 280:54]
  wire [7:0] s2_possible_predicted_fhs_res_hist_17_new_folded_hist_xored = {
    s2_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__7,
    s2_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__6,
    s2_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__5,
    s2_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__4,
    s2_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__3,
    s2_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__1,
    s2_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [15:0] s2_possible_predicted_fhs_res_hist_17_new_folded_hist_src_doubled = {
    s2_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__7,
    s2_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__6,
    s2_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__5,
    s2_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__4,
    s2_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__3,
    s2_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__1,
    s2_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__0,
    s2_possible_predicted_fhs_res_hist_17_new_folded_hist_xored}; // @[Cat.scala 31:58]
  wire [7:0] s2_possible_predicted_fhs_res_hist_17_new_folded_hist =
    s2_possible_predicted_fhs_res_hist_17_new_folded_hist_src_doubled[15:8]; // @[FrontendBundle.scala 221:30]
  wire  _s2_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_T_2 =
    predictors_io_out_s2_full_pred_br_taken_mask_0; // @[FrontendBundle.scala 274:80]
  wire [1:0] s2_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1 = {1'h0,
    _s2_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_T_2}; // @[FrontendBundle.scala 274:102]
  wire  s2_possible_predicted_fhs_res_hist_0_new_folded_hist_xored_res_1_6 =
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[1] ^
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__6; // @[FrontendBundle.scala 256:48]
  wire  s2_possible_predicted_fhs_res_hist_0_new_folded_hist_xored_res_1_7 =
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[0] ^ s2_possible_predicted_fhs_ob__0 ^
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__7; // @[FrontendBundle.scala 256:48]
  wire [7:0] s2_possible_predicted_fhs_res_hist_0_new_folded_hist_xored_1 = {
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_xored_res_1_7,
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_xored_res_1_6,
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__5,
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__4,
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__3,
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__1,
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [15:0] s2_possible_predicted_fhs_res_hist_0_new_folded_hist_src_doubled_1 = {
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_xored_res_1_7,
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_xored_res_1_6,
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__5,
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__4,
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__3,
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__1,
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__0,
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_xored_1}; // @[Cat.scala 31:58]
  wire [7:0] s2_possible_predicted_fhs_res_hist_0_new_folded_hist_1 =
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_src_doubled_1[14:7]; // @[FrontendBundle.scala 221:30]
  wire  s2_possible_predicted_fhs_res_hist_1_new_folded_hist_xored_res_1_6 =
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[1] ^
    s2_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__6; // @[FrontendBundle.scala 256:48]
  wire  s2_possible_predicted_fhs_res_hist_1_new_folded_hist_xored_res_1_7 =
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[0] ^ s2_possible_predicted_fhs_ob_1_0 ^
    s2_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__7; // @[FrontendBundle.scala 256:48]
  wire [7:0] s2_possible_predicted_fhs_res_hist_1_new_folded_hist_xored_1 = {
    s2_possible_predicted_fhs_res_hist_1_new_folded_hist_xored_res_1_7,
    s2_possible_predicted_fhs_res_hist_1_new_folded_hist_xored_res_1_6,
    s2_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__5,
    s2_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__4,
    s2_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__3,
    s2_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__1,
    s2_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [15:0] s2_possible_predicted_fhs_res_hist_1_new_folded_hist_src_doubled_1 = {
    s2_possible_predicted_fhs_res_hist_1_new_folded_hist_xored_res_1_7,
    s2_possible_predicted_fhs_res_hist_1_new_folded_hist_xored_res_1_6,
    s2_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__5,
    s2_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__4,
    s2_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__3,
    s2_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__1,
    s2_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__0,
    s2_possible_predicted_fhs_res_hist_1_new_folded_hist_xored_1}; // @[Cat.scala 31:58]
  wire [7:0] s2_possible_predicted_fhs_res_hist_1_new_folded_hist_1 =
    s2_possible_predicted_fhs_res_hist_1_new_folded_hist_src_doubled_1[14:7]; // @[FrontendBundle.scala 221:30]
  wire  s2_possible_predicted_fhs_res_hist_2_new_folded_hist_xored_res_1_6 =
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[1] ^ s2_possible_predicted_fhs_ob_2_0 ^
    s2_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__6; // @[FrontendBundle.scala 256:48]
  wire  s2_possible_predicted_fhs_res_hist_2_new_folded_hist_xored_res_1_7 =
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[0] ^
    s2_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__7; // @[FrontendBundle.scala 256:48]
  wire [7:0] s2_possible_predicted_fhs_res_hist_2_new_folded_hist_xored_1 = {
    s2_possible_predicted_fhs_res_hist_2_new_folded_hist_xored_res_1_7,
    s2_possible_predicted_fhs_res_hist_2_new_folded_hist_xored_res_1_6,
    s2_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__5,
    s2_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__4,
    s2_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__3,
    s2_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__1,
    s2_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [15:0] s2_possible_predicted_fhs_res_hist_2_new_folded_hist_src_doubled_1 = {
    s2_possible_predicted_fhs_res_hist_2_new_folded_hist_xored_res_1_7,
    s2_possible_predicted_fhs_res_hist_2_new_folded_hist_xored_res_1_6,
    s2_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__5,
    s2_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__4,
    s2_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__3,
    s2_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__1,
    s2_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__0,
    s2_possible_predicted_fhs_res_hist_2_new_folded_hist_xored_1}; // @[Cat.scala 31:58]
  wire [7:0] s2_possible_predicted_fhs_res_hist_2_new_folded_hist_1 =
    s2_possible_predicted_fhs_res_hist_2_new_folded_hist_src_doubled_1[14:7]; // @[FrontendBundle.scala 221:30]
  wire  s2_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_res_1_9 =
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[1] ^ s2_possible_predicted_fhs_ob_1_0 ^
    s2_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__9; // @[FrontendBundle.scala 256:48]
  wire  s2_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_res_1_10 =
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[0] ^
    s2_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__10; // @[FrontendBundle.scala 256:48]
  wire [10:0] s2_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_1 = {
    s2_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_res_1_10,
    s2_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_res_1_9,
    s2_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__8,
    s2_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__7,
    s2_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__6,
    s2_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__5,
    s2_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_lo}; // @[FrontendBundle.scala 258:11]
  wire [21:0] s2_possible_predicted_fhs_res_hist_3_new_folded_hist_src_doubled_1 = {
    s2_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_res_1_10,
    s2_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_res_1_9,
    s2_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__8,
    s2_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__7,
    s2_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__6,
    s2_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__5,
    s2_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_lo,
    s2_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_1}; // @[Cat.scala 31:58]
  wire [10:0] s2_possible_predicted_fhs_res_hist_3_new_folded_hist_1 =
    s2_possible_predicted_fhs_res_hist_3_new_folded_hist_src_doubled_1[20:10]; // @[FrontendBundle.scala 221:30]
  wire [4:0] _s2_possible_predicted_fhs_res_hist_4_new_folded_hist_T_2 = {s2_folded_gh_hist_4_folded_hist, 1'h0}; // @[FrontendBundle.scala 290:21]
  wire [4:0] _GEN_11919 = {{4'd0}, predictors_io_out_s2_full_pred_br_taken_mask_0}; // @[FrontendBundle.scala 290:29]
  wire [4:0] _s2_possible_predicted_fhs_res_hist_4_new_folded_hist_T_3 =
    _s2_possible_predicted_fhs_res_hist_4_new_folded_hist_T_2 | _GEN_11919; // @[FrontendBundle.scala 290:29]
  wire [3:0] s2_possible_predicted_fhs_res_hist_4_new_folded_hist_1 =
    _s2_possible_predicted_fhs_res_hist_4_new_folded_hist_T_3[3:0]; // @[FrontendBundle.scala 290:37]
  wire  s2_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_res_1_1 = s2_possible_predicted_fhs_ob_4_0 ^
    s2_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__1; // @[FrontendBundle.scala 256:48]
  wire  s2_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_res_1_9 =
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[1] ^
    s2_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__9; // @[FrontendBundle.scala 256:48]
  wire  s2_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_res_1_10 =
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[0] ^
    s2_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__10; // @[FrontendBundle.scala 256:48]
  wire [4:0] s2_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_lo_1 = {
    s2_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__4,
    s2_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__3,
    s2_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_res_1_1,
    s2_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [10:0] s2_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_1 = {
    s2_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_res_1_10,
    s2_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_res_1_9,
    s2_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__8,
    s2_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__7,
    s2_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__6,
    s2_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__5,
    s2_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_lo_1}; // @[FrontendBundle.scala 258:11]
  wire [21:0] s2_possible_predicted_fhs_res_hist_5_new_folded_hist_src_doubled_1 = {
    s2_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_res_1_10,
    s2_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_res_1_9,
    s2_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__8,
    s2_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__7,
    s2_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__6,
    s2_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__5,
    s2_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_lo_1,
    s2_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_1}; // @[Cat.scala 31:58]
  wire [10:0] s2_possible_predicted_fhs_res_hist_5_new_folded_hist_1 =
    s2_possible_predicted_fhs_res_hist_5_new_folded_hist_src_doubled_1[20:10]; // @[FrontendBundle.scala 221:30]
  wire  s2_possible_predicted_fhs_res_hist_6_new_folded_hist_xored_res_1_3 = s2_possible_predicted_fhs_ob_4_0 ^
    s2_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__3; // @[FrontendBundle.scala 256:48]
  wire  s2_possible_predicted_fhs_res_hist_6_new_folded_hist_xored_res_1_7 =
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[1] ^
    s2_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__7; // @[FrontendBundle.scala 256:48]
  wire  s2_possible_predicted_fhs_res_hist_6_new_folded_hist_xored_res_1_8 =
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[0] ^
    s2_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__8; // @[FrontendBundle.scala 256:48]
  wire [8:0] s2_possible_predicted_fhs_res_hist_6_new_folded_hist_xored_1 = {
    s2_possible_predicted_fhs_res_hist_6_new_folded_hist_xored_res_1_8,
    s2_possible_predicted_fhs_res_hist_6_new_folded_hist_xored_res_1_7,
    s2_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__6,
    s2_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__5,
    s2_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__4,
    s2_possible_predicted_fhs_res_hist_6_new_folded_hist_xored_res_1_3,
    s2_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__1,
    s2_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [17:0] s2_possible_predicted_fhs_res_hist_6_new_folded_hist_src_doubled_1 = {
    s2_possible_predicted_fhs_res_hist_6_new_folded_hist_xored_res_1_8,
    s2_possible_predicted_fhs_res_hist_6_new_folded_hist_xored_res_1_7,
    s2_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__6,
    s2_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__5,
    s2_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__4,
    s2_possible_predicted_fhs_res_hist_6_new_folded_hist_xored_res_1_3,
    s2_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__1,
    s2_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__0,
    s2_possible_predicted_fhs_res_hist_6_new_folded_hist_xored_1}; // @[Cat.scala 31:58]
  wire [8:0] s2_possible_predicted_fhs_res_hist_6_new_folded_hist_1 =
    s2_possible_predicted_fhs_res_hist_6_new_folded_hist_src_doubled_1[16:8]; // @[FrontendBundle.scala 221:30]
  wire  s2_possible_predicted_fhs_res_hist_7_new_folded_hist_xored_res_1_6 = s2_possible_predicted_fhs_ob__0 ^
    s2_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__6; // @[FrontendBundle.scala 256:48]
  wire  s2_possible_predicted_fhs_res_hist_7_new_folded_hist_xored_res_1_7 =
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[1] ^
    s2_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__7; // @[FrontendBundle.scala 256:48]
  wire  s2_possible_predicted_fhs_res_hist_7_new_folded_hist_xored_res_1_8 =
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[0] ^
    s2_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__8; // @[FrontendBundle.scala 256:48]
  wire [8:0] s2_possible_predicted_fhs_res_hist_7_new_folded_hist_xored_1 = {
    s2_possible_predicted_fhs_res_hist_7_new_folded_hist_xored_res_1_8,
    s2_possible_predicted_fhs_res_hist_7_new_folded_hist_xored_res_1_7,
    s2_possible_predicted_fhs_res_hist_7_new_folded_hist_xored_res_1_6,
    s2_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__5,
    s2_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__4,
    s2_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__3,
    s2_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__1,
    s2_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [17:0] s2_possible_predicted_fhs_res_hist_7_new_folded_hist_src_doubled_1 = {
    s2_possible_predicted_fhs_res_hist_7_new_folded_hist_xored_res_1_8,
    s2_possible_predicted_fhs_res_hist_7_new_folded_hist_xored_res_1_7,
    s2_possible_predicted_fhs_res_hist_7_new_folded_hist_xored_res_1_6,
    s2_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__5,
    s2_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__4,
    s2_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__3,
    s2_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__1,
    s2_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__0,
    s2_possible_predicted_fhs_res_hist_7_new_folded_hist_xored_1}; // @[Cat.scala 31:58]
  wire [8:0] s2_possible_predicted_fhs_res_hist_7_new_folded_hist_1 =
    s2_possible_predicted_fhs_res_hist_7_new_folded_hist_src_doubled_1[16:8]; // @[FrontendBundle.scala 221:30]
  wire [8:0] _s2_possible_predicted_fhs_res_hist_8_new_folded_hist_T_2 = {s2_folded_gh_hist_8_folded_hist, 1'h0}; // @[FrontendBundle.scala 290:21]
  wire [8:0] _GEN_11920 = {{8'd0}, predictors_io_out_s2_full_pred_br_taken_mask_0}; // @[FrontendBundle.scala 290:29]
  wire [8:0] _s2_possible_predicted_fhs_res_hist_8_new_folded_hist_T_3 =
    _s2_possible_predicted_fhs_res_hist_8_new_folded_hist_T_2 | _GEN_11920; // @[FrontendBundle.scala 290:29]
  wire [7:0] s2_possible_predicted_fhs_res_hist_8_new_folded_hist_1 =
    _s2_possible_predicted_fhs_res_hist_8_new_folded_hist_T_3[7:0]; // @[FrontendBundle.scala 290:37]
  wire  s2_possible_predicted_fhs_res_hist_9_new_folded_hist_xored_res_1_3 = s2_possible_predicted_fhs_ob_1_0 ^
    s2_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__3; // @[FrontendBundle.scala 256:48]
  wire  s2_possible_predicted_fhs_res_hist_9_new_folded_hist_xored_res_1_5 =
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[1] ^
    s2_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__5; // @[FrontendBundle.scala 256:48]
  wire  s2_possible_predicted_fhs_res_hist_9_new_folded_hist_xored_res_1_6 =
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[0] ^
    s2_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__6; // @[FrontendBundle.scala 256:48]
  wire [6:0] s2_possible_predicted_fhs_res_hist_9_new_folded_hist_xored_1 = {
    s2_possible_predicted_fhs_res_hist_9_new_folded_hist_xored_res_1_6,
    s2_possible_predicted_fhs_res_hist_9_new_folded_hist_xored_res_1_5,
    s2_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__4,
    s2_possible_predicted_fhs_res_hist_9_new_folded_hist_xored_res_1_3,
    s2_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__1,
    s2_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [13:0] s2_possible_predicted_fhs_res_hist_9_new_folded_hist_src_doubled_1 = {
    s2_possible_predicted_fhs_res_hist_9_new_folded_hist_xored_res_1_6,
    s2_possible_predicted_fhs_res_hist_9_new_folded_hist_xored_res_1_5,
    s2_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__4,
    s2_possible_predicted_fhs_res_hist_9_new_folded_hist_xored_res_1_3,
    s2_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__1,
    s2_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__0,
    s2_possible_predicted_fhs_res_hist_9_new_folded_hist_xored_1}; // @[Cat.scala 31:58]
  wire [6:0] s2_possible_predicted_fhs_res_hist_9_new_folded_hist_1 =
    s2_possible_predicted_fhs_res_hist_9_new_folded_hist_src_doubled_1[12:6]; // @[FrontendBundle.scala 221:30]
  wire  s2_possible_predicted_fhs_res_hist_10_new_folded_hist_xored_res_1_4 = s2_possible_predicted_fhs_ob_1_0 ^
    s2_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__4; // @[FrontendBundle.scala 256:48]
  wire  s2_possible_predicted_fhs_res_hist_10_new_folded_hist_xored_res_1_7 =
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[1] ^
    s2_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__7; // @[FrontendBundle.scala 256:48]
  wire  s2_possible_predicted_fhs_res_hist_10_new_folded_hist_xored_res_1_8 =
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[0] ^
    s2_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__8; // @[FrontendBundle.scala 256:48]
  wire [8:0] s2_possible_predicted_fhs_res_hist_10_new_folded_hist_xored_1 = {
    s2_possible_predicted_fhs_res_hist_10_new_folded_hist_xored_res_1_8,
    s2_possible_predicted_fhs_res_hist_10_new_folded_hist_xored_res_1_7,
    s2_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__6,
    s2_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__5,
    s2_possible_predicted_fhs_res_hist_10_new_folded_hist_xored_res_1_4,
    s2_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__3,
    s2_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__1,
    s2_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [17:0] s2_possible_predicted_fhs_res_hist_10_new_folded_hist_src_doubled_1 = {
    s2_possible_predicted_fhs_res_hist_10_new_folded_hist_xored_res_1_8,
    s2_possible_predicted_fhs_res_hist_10_new_folded_hist_xored_res_1_7,
    s2_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__6,
    s2_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__5,
    s2_possible_predicted_fhs_res_hist_10_new_folded_hist_xored_res_1_4,
    s2_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__3,
    s2_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__1,
    s2_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__0,
    s2_possible_predicted_fhs_res_hist_10_new_folded_hist_xored_1}; // @[Cat.scala 31:58]
  wire [8:0] s2_possible_predicted_fhs_res_hist_10_new_folded_hist_1 =
    s2_possible_predicted_fhs_res_hist_10_new_folded_hist_src_doubled_1[16:8]; // @[FrontendBundle.scala 221:30]
  wire [8:0] _s2_possible_predicted_fhs_res_hist_11_new_folded_hist_T_2 = {s2_folded_gh_hist_11_folded_hist, 1'h0}; // @[FrontendBundle.scala 290:21]
  wire [8:0] _s2_possible_predicted_fhs_res_hist_11_new_folded_hist_T_3 =
    _s2_possible_predicted_fhs_res_hist_11_new_folded_hist_T_2 | _GEN_11920; // @[FrontendBundle.scala 290:29]
  wire [7:0] s2_possible_predicted_fhs_res_hist_11_new_folded_hist_1 =
    _s2_possible_predicted_fhs_res_hist_11_new_folded_hist_T_3[7:0]; // @[FrontendBundle.scala 290:37]
  wire  s2_possible_predicted_fhs_res_hist_12_new_folded_hist_xored_res_1_5 =
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[1] ^ s2_possible_predicted_fhs_ob_4_0 ^
    s2_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__5; // @[FrontendBundle.scala 256:48]
  wire  s2_possible_predicted_fhs_res_hist_12_new_folded_hist_xored_res_1_6 =
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[0] ^
    s2_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__6; // @[FrontendBundle.scala 256:48]
  wire [6:0] s2_possible_predicted_fhs_res_hist_12_new_folded_hist_xored_1 = {
    s2_possible_predicted_fhs_res_hist_12_new_folded_hist_xored_res_1_6,
    s2_possible_predicted_fhs_res_hist_12_new_folded_hist_xored_res_1_5,
    s2_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__4,
    s2_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__3,
    s2_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__1,
    s2_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [13:0] s2_possible_predicted_fhs_res_hist_12_new_folded_hist_src_doubled_1 = {
    s2_possible_predicted_fhs_res_hist_12_new_folded_hist_xored_res_1_6,
    s2_possible_predicted_fhs_res_hist_12_new_folded_hist_xored_res_1_5,
    s2_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__4,
    s2_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__3,
    s2_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__1,
    s2_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__0,
    s2_possible_predicted_fhs_res_hist_12_new_folded_hist_xored_1}; // @[Cat.scala 31:58]
  wire [6:0] s2_possible_predicted_fhs_res_hist_12_new_folded_hist_1 =
    s2_possible_predicted_fhs_res_hist_12_new_folded_hist_src_doubled_1[12:6]; // @[FrontendBundle.scala 221:30]
  wire  s2_possible_predicted_fhs_res_hist_13_new_folded_hist_xored_res_1_0 = s2_possible_predicted_fhs_ob_10_0 ^
    s2_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__0; // @[FrontendBundle.scala 256:48]
  wire  s2_possible_predicted_fhs_res_hist_13_new_folded_hist_xored_res_1_5 =
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[1] ^
    s2_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__5; // @[FrontendBundle.scala 256:48]
  wire  s2_possible_predicted_fhs_res_hist_13_new_folded_hist_xored_res_1_6 =
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[0] ^
    s2_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__6; // @[FrontendBundle.scala 256:48]
  wire [6:0] s2_possible_predicted_fhs_res_hist_13_new_folded_hist_xored_1 = {
    s2_possible_predicted_fhs_res_hist_13_new_folded_hist_xored_res_1_6,
    s2_possible_predicted_fhs_res_hist_13_new_folded_hist_xored_res_1_5,
    s2_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__4,
    s2_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__3,
    s2_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__1,
    s2_possible_predicted_fhs_res_hist_13_new_folded_hist_xored_res_1_0}; // @[FrontendBundle.scala 258:11]
  wire [13:0] s2_possible_predicted_fhs_res_hist_13_new_folded_hist_src_doubled_1 = {
    s2_possible_predicted_fhs_res_hist_13_new_folded_hist_xored_res_1_6,
    s2_possible_predicted_fhs_res_hist_13_new_folded_hist_xored_res_1_5,
    s2_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__4,
    s2_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__3,
    s2_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__1,
    s2_possible_predicted_fhs_res_hist_13_new_folded_hist_xored_res_1_0,
    s2_possible_predicted_fhs_res_hist_13_new_folded_hist_xored_1}; // @[Cat.scala 31:58]
  wire [6:0] s2_possible_predicted_fhs_res_hist_13_new_folded_hist_1 =
    s2_possible_predicted_fhs_res_hist_13_new_folded_hist_src_doubled_1[12:6]; // @[FrontendBundle.scala 221:30]
  wire  s2_possible_predicted_fhs_res_hist_14_new_folded_hist_xored_res_1_5 =
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[1] ^
    s2_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__5; // @[FrontendBundle.scala 256:48]
  wire  s2_possible_predicted_fhs_res_hist_14_new_folded_hist_xored_res_1_6 =
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[0] ^ s2_possible_predicted_fhs_ob_2_0 ^
    s2_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__6; // @[FrontendBundle.scala 256:48]
  wire [6:0] s2_possible_predicted_fhs_res_hist_14_new_folded_hist_xored_1 = {
    s2_possible_predicted_fhs_res_hist_14_new_folded_hist_xored_res_1_6,
    s2_possible_predicted_fhs_res_hist_14_new_folded_hist_xored_res_1_5,
    s2_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__4,
    s2_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__3,
    s2_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__1,
    s2_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [13:0] s2_possible_predicted_fhs_res_hist_14_new_folded_hist_src_doubled_1 = {
    s2_possible_predicted_fhs_res_hist_14_new_folded_hist_xored_res_1_6,
    s2_possible_predicted_fhs_res_hist_14_new_folded_hist_xored_res_1_5,
    s2_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__4,
    s2_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__3,
    s2_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__1,
    s2_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__0,
    s2_possible_predicted_fhs_res_hist_14_new_folded_hist_xored_1}; // @[Cat.scala 31:58]
  wire [6:0] s2_possible_predicted_fhs_res_hist_14_new_folded_hist_1 =
    s2_possible_predicted_fhs_res_hist_14_new_folded_hist_src_doubled_1[12:6]; // @[FrontendBundle.scala 221:30]
  wire  s2_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_res_1_8 = s2_possible_predicted_fhs_ob_2_0 ^
    s2_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__8; // @[FrontendBundle.scala 256:48]
  wire  s2_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_res_1_9 =
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[1] ^
    s2_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__9; // @[FrontendBundle.scala 256:48]
  wire  s2_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_res_1_10 =
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[0] ^
    s2_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__10; // @[FrontendBundle.scala 256:48]
  wire [10:0] s2_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_1 = {
    s2_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_res_1_10,
    s2_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_res_1_9,
    s2_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_res_1_8,
    s2_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__7,
    s2_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__6,
    s2_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__5,
    s2_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_lo}; // @[FrontendBundle.scala 258:11]
  wire [21:0] s2_possible_predicted_fhs_res_hist_15_new_folded_hist_src_doubled_1 = {
    s2_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_res_1_10,
    s2_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_res_1_9,
    s2_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_res_1_8,
    s2_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__7,
    s2_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__6,
    s2_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__5,
    s2_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_lo,
    s2_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_1}; // @[Cat.scala 31:58]
  wire [10:0] s2_possible_predicted_fhs_res_hist_15_new_folded_hist_1 =
    s2_possible_predicted_fhs_res_hist_15_new_folded_hist_src_doubled_1[20:10]; // @[FrontendBundle.scala 221:30]
  wire  s2_possible_predicted_fhs_res_hist_16_new_folded_hist_xored_res_1_1 = s2_possible_predicted_fhs_ob_13_0 ^
    s2_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__1; // @[FrontendBundle.scala 256:48]
  wire  s2_possible_predicted_fhs_res_hist_16_new_folded_hist_xored_res_1_6 =
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[1] ^
    s2_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__6; // @[FrontendBundle.scala 256:48]
  wire  s2_possible_predicted_fhs_res_hist_16_new_folded_hist_xored_res_1_7 =
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[0] ^
    s2_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__7; // @[FrontendBundle.scala 256:48]
  wire [7:0] s2_possible_predicted_fhs_res_hist_16_new_folded_hist_xored_1 = {
    s2_possible_predicted_fhs_res_hist_16_new_folded_hist_xored_res_1_7,
    s2_possible_predicted_fhs_res_hist_16_new_folded_hist_xored_res_1_6,
    s2_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__5,
    s2_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__4,
    s2_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__3,
    s2_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_16_new_folded_hist_xored_res_1_1,
    s2_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [15:0] s2_possible_predicted_fhs_res_hist_16_new_folded_hist_src_doubled_1 = {
    s2_possible_predicted_fhs_res_hist_16_new_folded_hist_xored_res_1_7,
    s2_possible_predicted_fhs_res_hist_16_new_folded_hist_xored_res_1_6,
    s2_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__5,
    s2_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__4,
    s2_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__3,
    s2_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_16_new_folded_hist_xored_res_1_1,
    s2_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__0,
    s2_possible_predicted_fhs_res_hist_16_new_folded_hist_xored_1}; // @[Cat.scala 31:58]
  wire [7:0] s2_possible_predicted_fhs_res_hist_16_new_folded_hist_1 =
    s2_possible_predicted_fhs_res_hist_16_new_folded_hist_src_doubled_1[14:7]; // @[FrontendBundle.scala 221:30]
  wire  s2_possible_predicted_fhs_res_hist_17_new_folded_hist_xored_res_1_4 = s2_possible_predicted_fhs_ob_4_0 ^
    s2_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__4; // @[FrontendBundle.scala 256:48]
  wire  s2_possible_predicted_fhs_res_hist_17_new_folded_hist_xored_res_1_6 =
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[1] ^
    s2_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__6; // @[FrontendBundle.scala 256:48]
  wire  s2_possible_predicted_fhs_res_hist_17_new_folded_hist_xored_res_1_7 =
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[0] ^
    s2_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__7; // @[FrontendBundle.scala 256:48]
  wire [7:0] s2_possible_predicted_fhs_res_hist_17_new_folded_hist_xored_1 = {
    s2_possible_predicted_fhs_res_hist_17_new_folded_hist_xored_res_1_7,
    s2_possible_predicted_fhs_res_hist_17_new_folded_hist_xored_res_1_6,
    s2_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__5,
    s2_possible_predicted_fhs_res_hist_17_new_folded_hist_xored_res_1_4,
    s2_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__3,
    s2_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__1,
    s2_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [15:0] s2_possible_predicted_fhs_res_hist_17_new_folded_hist_src_doubled_1 = {
    s2_possible_predicted_fhs_res_hist_17_new_folded_hist_xored_res_1_7,
    s2_possible_predicted_fhs_res_hist_17_new_folded_hist_xored_res_1_6,
    s2_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__5,
    s2_possible_predicted_fhs_res_hist_17_new_folded_hist_xored_res_1_4,
    s2_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__3,
    s2_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__1,
    s2_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__0,
    s2_possible_predicted_fhs_res_hist_17_new_folded_hist_xored_1}; // @[Cat.scala 31:58]
  wire [7:0] s2_possible_predicted_fhs_res_hist_17_new_folded_hist_1 =
    s2_possible_predicted_fhs_res_hist_17_new_folded_hist_src_doubled_1[14:7]; // @[FrontendBundle.scala 221:30]
  wire  _s2_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_T_5 =
    predictors_io_out_s2_full_pred_br_taken_mask_1; // @[FrontendBundle.scala 274:80]
  wire [1:0] s2_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2 = {
    _s2_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_T_5,1'h0}; // @[FrontendBundle.scala 274:102]
  wire  s2_possible_predicted_fhs_res_hist_0_new_folded_hist_xored_res_2_6 =
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[1] ^ s2_possible_predicted_fhs_ob__1 ^
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__6; // @[FrontendBundle.scala 256:48]
  wire  s2_possible_predicted_fhs_res_hist_0_new_folded_hist_xored_res_2_7 =
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[0] ^ s2_possible_predicted_fhs_ob__0 ^
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__7; // @[FrontendBundle.scala 256:48]
  wire [7:0] s2_possible_predicted_fhs_res_hist_0_new_folded_hist_xored_2 = {
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_xored_res_2_7,
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_xored_res_2_6,
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__5,
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__4,
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__3,
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__1,
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [15:0] s2_possible_predicted_fhs_res_hist_0_new_folded_hist_src_doubled_2 = {
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_xored_res_2_7,
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_xored_res_2_6,
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__5,
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__4,
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__3,
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__1,
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__0,
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_xored_2}; // @[Cat.scala 31:58]
  wire [7:0] s2_possible_predicted_fhs_res_hist_0_new_folded_hist_2 =
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_src_doubled_2[13:6]; // @[FrontendBundle.scala 221:30]
  wire  s2_possible_predicted_fhs_res_hist_1_new_folded_hist_xored_res_2_6 =
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[1] ^ s2_possible_predicted_fhs_ob_1_1 ^
    s2_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__6; // @[FrontendBundle.scala 256:48]
  wire  s2_possible_predicted_fhs_res_hist_1_new_folded_hist_xored_res_2_7 =
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[0] ^ s2_possible_predicted_fhs_ob_1_0 ^
    s2_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__7; // @[FrontendBundle.scala 256:48]
  wire [7:0] s2_possible_predicted_fhs_res_hist_1_new_folded_hist_xored_2 = {
    s2_possible_predicted_fhs_res_hist_1_new_folded_hist_xored_res_2_7,
    s2_possible_predicted_fhs_res_hist_1_new_folded_hist_xored_res_2_6,
    s2_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__5,
    s2_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__4,
    s2_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__3,
    s2_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__1,
    s2_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [15:0] s2_possible_predicted_fhs_res_hist_1_new_folded_hist_src_doubled_2 = {
    s2_possible_predicted_fhs_res_hist_1_new_folded_hist_xored_res_2_7,
    s2_possible_predicted_fhs_res_hist_1_new_folded_hist_xored_res_2_6,
    s2_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__5,
    s2_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__4,
    s2_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__3,
    s2_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__1,
    s2_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__0,
    s2_possible_predicted_fhs_res_hist_1_new_folded_hist_xored_2}; // @[Cat.scala 31:58]
  wire [7:0] s2_possible_predicted_fhs_res_hist_1_new_folded_hist_2 =
    s2_possible_predicted_fhs_res_hist_1_new_folded_hist_src_doubled_2[13:6]; // @[FrontendBundle.scala 221:30]
  wire  s2_possible_predicted_fhs_res_hist_2_new_folded_hist_xored_res_2_5 = s2_possible_predicted_fhs_ob_2_1 ^
    s2_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__5; // @[FrontendBundle.scala 256:48]
  wire  s2_possible_predicted_fhs_res_hist_2_new_folded_hist_xored_res_2_6 =
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[1] ^ s2_possible_predicted_fhs_ob_2_0 ^
    s2_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__6; // @[FrontendBundle.scala 256:48]
  wire  s2_possible_predicted_fhs_res_hist_2_new_folded_hist_xored_res_2_7 =
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[0] ^
    s2_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__7; // @[FrontendBundle.scala 256:48]
  wire [7:0] s2_possible_predicted_fhs_res_hist_2_new_folded_hist_xored_2 = {
    s2_possible_predicted_fhs_res_hist_2_new_folded_hist_xored_res_2_7,
    s2_possible_predicted_fhs_res_hist_2_new_folded_hist_xored_res_2_6,
    s2_possible_predicted_fhs_res_hist_2_new_folded_hist_xored_res_2_5,
    s2_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__4,
    s2_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__3,
    s2_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__1,
    s2_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [15:0] s2_possible_predicted_fhs_res_hist_2_new_folded_hist_src_doubled_2 = {
    s2_possible_predicted_fhs_res_hist_2_new_folded_hist_xored_res_2_7,
    s2_possible_predicted_fhs_res_hist_2_new_folded_hist_xored_res_2_6,
    s2_possible_predicted_fhs_res_hist_2_new_folded_hist_xored_res_2_5,
    s2_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__4,
    s2_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__3,
    s2_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__1,
    s2_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__0,
    s2_possible_predicted_fhs_res_hist_2_new_folded_hist_xored_2}; // @[Cat.scala 31:58]
  wire [7:0] s2_possible_predicted_fhs_res_hist_2_new_folded_hist_2 =
    s2_possible_predicted_fhs_res_hist_2_new_folded_hist_src_doubled_2[13:6]; // @[FrontendBundle.scala 221:30]
  wire  s2_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_res_2_8 = s2_possible_predicted_fhs_ob_1_1 ^
    s2_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__8; // @[FrontendBundle.scala 256:48]
  wire  s2_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_res_2_9 =
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[1] ^ s2_possible_predicted_fhs_ob_1_0 ^
    s2_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__9; // @[FrontendBundle.scala 256:48]
  wire  s2_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_res_2_10 =
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[0] ^
    s2_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__10; // @[FrontendBundle.scala 256:48]
  wire [10:0] s2_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_2 = {
    s2_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_res_2_10,
    s2_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_res_2_9,
    s2_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_res_2_8,
    s2_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__7,
    s2_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__6,
    s2_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__5,
    s2_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_lo}; // @[FrontendBundle.scala 258:11]
  wire [21:0] s2_possible_predicted_fhs_res_hist_3_new_folded_hist_src_doubled_2 = {
    s2_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_res_2_10,
    s2_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_res_2_9,
    s2_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_res_2_8,
    s2_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__7,
    s2_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__6,
    s2_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__5,
    s2_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_lo,
    s2_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_2}; // @[Cat.scala 31:58]
  wire [10:0] s2_possible_predicted_fhs_res_hist_3_new_folded_hist_2 =
    s2_possible_predicted_fhs_res_hist_3_new_folded_hist_src_doubled_2[19:9]; // @[FrontendBundle.scala 221:30]
  wire [5:0] _s2_possible_predicted_fhs_res_hist_4_new_folded_hist_T_4 = {s2_folded_gh_hist_4_folded_hist, 2'h0}; // @[FrontendBundle.scala 290:21]
  wire [5:0] _GEN_11922 = {{5'd0}, predictors_io_out_s2_full_pred_br_taken_mask_1}; // @[FrontendBundle.scala 290:29]
  wire [5:0] _s2_possible_predicted_fhs_res_hist_4_new_folded_hist_T_5 =
    _s2_possible_predicted_fhs_res_hist_4_new_folded_hist_T_4 | _GEN_11922; // @[FrontendBundle.scala 290:29]
  wire [3:0] s2_possible_predicted_fhs_res_hist_4_new_folded_hist_2 =
    _s2_possible_predicted_fhs_res_hist_4_new_folded_hist_T_5[3:0]; // @[FrontendBundle.scala 290:37]
  wire  s2_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_res_2_0 = s2_possible_predicted_fhs_ob_4_1 ^
    s2_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__0; // @[FrontendBundle.scala 256:48]
  wire  s2_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_res_2_9 =
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[1] ^
    s2_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__9; // @[FrontendBundle.scala 256:48]
  wire  s2_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_res_2_10 =
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[0] ^
    s2_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__10; // @[FrontendBundle.scala 256:48]
  wire [4:0] s2_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_lo_2 = {
    s2_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__4,
    s2_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__3,
    s2_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_res_1_1,
    s2_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_res_2_0}; // @[FrontendBundle.scala 258:11]
  wire [10:0] s2_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_2 = {
    s2_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_res_2_10,
    s2_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_res_2_9,
    s2_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__8,
    s2_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__7,
    s2_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__6,
    s2_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__5,
    s2_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_lo_2}; // @[FrontendBundle.scala 258:11]
  wire [21:0] s2_possible_predicted_fhs_res_hist_5_new_folded_hist_src_doubled_2 = {
    s2_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_res_2_10,
    s2_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_res_2_9,
    s2_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__8,
    s2_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__7,
    s2_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__6,
    s2_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__5,
    s2_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_lo_2,
    s2_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_2}; // @[Cat.scala 31:58]
  wire [10:0] s2_possible_predicted_fhs_res_hist_5_new_folded_hist_2 =
    s2_possible_predicted_fhs_res_hist_5_new_folded_hist_src_doubled_2[19:9]; // @[FrontendBundle.scala 221:30]
  wire  s2_possible_predicted_fhs_res_hist_6_new_folded_hist_xored_res_2_2 = s2_possible_predicted_fhs_ob_4_1 ^
    s2_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__2; // @[FrontendBundle.scala 256:48]
  wire  s2_possible_predicted_fhs_res_hist_6_new_folded_hist_xored_res_2_7 =
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[1] ^
    s2_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__7; // @[FrontendBundle.scala 256:48]
  wire  s2_possible_predicted_fhs_res_hist_6_new_folded_hist_xored_res_2_8 =
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[0] ^
    s2_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__8; // @[FrontendBundle.scala 256:48]
  wire [8:0] s2_possible_predicted_fhs_res_hist_6_new_folded_hist_xored_2 = {
    s2_possible_predicted_fhs_res_hist_6_new_folded_hist_xored_res_2_8,
    s2_possible_predicted_fhs_res_hist_6_new_folded_hist_xored_res_2_7,
    s2_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__6,
    s2_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__5,
    s2_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__4,
    s2_possible_predicted_fhs_res_hist_6_new_folded_hist_xored_res_1_3,
    s2_possible_predicted_fhs_res_hist_6_new_folded_hist_xored_res_2_2,
    s2_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__1,
    s2_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [17:0] s2_possible_predicted_fhs_res_hist_6_new_folded_hist_src_doubled_2 = {
    s2_possible_predicted_fhs_res_hist_6_new_folded_hist_xored_res_2_8,
    s2_possible_predicted_fhs_res_hist_6_new_folded_hist_xored_res_2_7,
    s2_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__6,
    s2_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__5,
    s2_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__4,
    s2_possible_predicted_fhs_res_hist_6_new_folded_hist_xored_res_1_3,
    s2_possible_predicted_fhs_res_hist_6_new_folded_hist_xored_res_2_2,
    s2_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__1,
    s2_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__0,
    s2_possible_predicted_fhs_res_hist_6_new_folded_hist_xored_2}; // @[Cat.scala 31:58]
  wire [8:0] s2_possible_predicted_fhs_res_hist_6_new_folded_hist_2 =
    s2_possible_predicted_fhs_res_hist_6_new_folded_hist_src_doubled_2[15:7]; // @[FrontendBundle.scala 221:30]
  wire  s2_possible_predicted_fhs_res_hist_7_new_folded_hist_xored_res_2_5 = s2_possible_predicted_fhs_ob__1 ^
    s2_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__5; // @[FrontendBundle.scala 256:48]
  wire  s2_possible_predicted_fhs_res_hist_7_new_folded_hist_xored_res_2_7 =
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[1] ^
    s2_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__7; // @[FrontendBundle.scala 256:48]
  wire  s2_possible_predicted_fhs_res_hist_7_new_folded_hist_xored_res_2_8 =
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[0] ^
    s2_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__8; // @[FrontendBundle.scala 256:48]
  wire [8:0] s2_possible_predicted_fhs_res_hist_7_new_folded_hist_xored_2 = {
    s2_possible_predicted_fhs_res_hist_7_new_folded_hist_xored_res_2_8,
    s2_possible_predicted_fhs_res_hist_7_new_folded_hist_xored_res_2_7,
    s2_possible_predicted_fhs_res_hist_7_new_folded_hist_xored_res_1_6,
    s2_possible_predicted_fhs_res_hist_7_new_folded_hist_xored_res_2_5,
    s2_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__4,
    s2_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__3,
    s2_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__1,
    s2_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [17:0] s2_possible_predicted_fhs_res_hist_7_new_folded_hist_src_doubled_2 = {
    s2_possible_predicted_fhs_res_hist_7_new_folded_hist_xored_res_2_8,
    s2_possible_predicted_fhs_res_hist_7_new_folded_hist_xored_res_2_7,
    s2_possible_predicted_fhs_res_hist_7_new_folded_hist_xored_res_1_6,
    s2_possible_predicted_fhs_res_hist_7_new_folded_hist_xored_res_2_5,
    s2_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__4,
    s2_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__3,
    s2_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__1,
    s2_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__0,
    s2_possible_predicted_fhs_res_hist_7_new_folded_hist_xored_2}; // @[Cat.scala 31:58]
  wire [8:0] s2_possible_predicted_fhs_res_hist_7_new_folded_hist_2 =
    s2_possible_predicted_fhs_res_hist_7_new_folded_hist_src_doubled_2[15:7]; // @[FrontendBundle.scala 221:30]
  wire [9:0] _s2_possible_predicted_fhs_res_hist_8_new_folded_hist_T_4 = {s2_folded_gh_hist_8_folded_hist, 2'h0}; // @[FrontendBundle.scala 290:21]
  wire [9:0] _GEN_11923 = {{9'd0}, predictors_io_out_s2_full_pred_br_taken_mask_1}; // @[FrontendBundle.scala 290:29]
  wire [9:0] _s2_possible_predicted_fhs_res_hist_8_new_folded_hist_T_5 =
    _s2_possible_predicted_fhs_res_hist_8_new_folded_hist_T_4 | _GEN_11923; // @[FrontendBundle.scala 290:29]
  wire [7:0] s2_possible_predicted_fhs_res_hist_8_new_folded_hist_2 =
    _s2_possible_predicted_fhs_res_hist_8_new_folded_hist_T_5[7:0]; // @[FrontendBundle.scala 290:37]
  wire  s2_possible_predicted_fhs_res_hist_9_new_folded_hist_xored_res_2_2 = s2_possible_predicted_fhs_ob_1_1 ^
    s2_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__2; // @[FrontendBundle.scala 256:48]
  wire  s2_possible_predicted_fhs_res_hist_9_new_folded_hist_xored_res_2_5 =
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[1] ^
    s2_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__5; // @[FrontendBundle.scala 256:48]
  wire  s2_possible_predicted_fhs_res_hist_9_new_folded_hist_xored_res_2_6 =
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[0] ^
    s2_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__6; // @[FrontendBundle.scala 256:48]
  wire [6:0] s2_possible_predicted_fhs_res_hist_9_new_folded_hist_xored_2 = {
    s2_possible_predicted_fhs_res_hist_9_new_folded_hist_xored_res_2_6,
    s2_possible_predicted_fhs_res_hist_9_new_folded_hist_xored_res_2_5,
    s2_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__4,
    s2_possible_predicted_fhs_res_hist_9_new_folded_hist_xored_res_1_3,
    s2_possible_predicted_fhs_res_hist_9_new_folded_hist_xored_res_2_2,
    s2_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__1,
    s2_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [13:0] s2_possible_predicted_fhs_res_hist_9_new_folded_hist_src_doubled_2 = {
    s2_possible_predicted_fhs_res_hist_9_new_folded_hist_xored_res_2_6,
    s2_possible_predicted_fhs_res_hist_9_new_folded_hist_xored_res_2_5,
    s2_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__4,
    s2_possible_predicted_fhs_res_hist_9_new_folded_hist_xored_res_1_3,
    s2_possible_predicted_fhs_res_hist_9_new_folded_hist_xored_res_2_2,
    s2_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__1,
    s2_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__0,
    s2_possible_predicted_fhs_res_hist_9_new_folded_hist_xored_2}; // @[Cat.scala 31:58]
  wire [6:0] s2_possible_predicted_fhs_res_hist_9_new_folded_hist_2 =
    s2_possible_predicted_fhs_res_hist_9_new_folded_hist_src_doubled_2[11:5]; // @[FrontendBundle.scala 221:30]
  wire  s2_possible_predicted_fhs_res_hist_10_new_folded_hist_xored_res_2_3 = s2_possible_predicted_fhs_ob_1_1 ^
    s2_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__3; // @[FrontendBundle.scala 256:48]
  wire  s2_possible_predicted_fhs_res_hist_10_new_folded_hist_xored_res_2_7 =
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[1] ^
    s2_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__7; // @[FrontendBundle.scala 256:48]
  wire  s2_possible_predicted_fhs_res_hist_10_new_folded_hist_xored_res_2_8 =
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[0] ^
    s2_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__8; // @[FrontendBundle.scala 256:48]
  wire [8:0] s2_possible_predicted_fhs_res_hist_10_new_folded_hist_xored_2 = {
    s2_possible_predicted_fhs_res_hist_10_new_folded_hist_xored_res_2_8,
    s2_possible_predicted_fhs_res_hist_10_new_folded_hist_xored_res_2_7,
    s2_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__6,
    s2_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__5,
    s2_possible_predicted_fhs_res_hist_10_new_folded_hist_xored_res_1_4,
    s2_possible_predicted_fhs_res_hist_10_new_folded_hist_xored_res_2_3,
    s2_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__1,
    s2_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [17:0] s2_possible_predicted_fhs_res_hist_10_new_folded_hist_src_doubled_2 = {
    s2_possible_predicted_fhs_res_hist_10_new_folded_hist_xored_res_2_8,
    s2_possible_predicted_fhs_res_hist_10_new_folded_hist_xored_res_2_7,
    s2_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__6,
    s2_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__5,
    s2_possible_predicted_fhs_res_hist_10_new_folded_hist_xored_res_1_4,
    s2_possible_predicted_fhs_res_hist_10_new_folded_hist_xored_res_2_3,
    s2_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__1,
    s2_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__0,
    s2_possible_predicted_fhs_res_hist_10_new_folded_hist_xored_2}; // @[Cat.scala 31:58]
  wire [8:0] s2_possible_predicted_fhs_res_hist_10_new_folded_hist_2 =
    s2_possible_predicted_fhs_res_hist_10_new_folded_hist_src_doubled_2[15:7]; // @[FrontendBundle.scala 221:30]
  wire [9:0] _s2_possible_predicted_fhs_res_hist_11_new_folded_hist_T_4 = {s2_folded_gh_hist_11_folded_hist, 2'h0}; // @[FrontendBundle.scala 290:21]
  wire [9:0] _s2_possible_predicted_fhs_res_hist_11_new_folded_hist_T_5 =
    _s2_possible_predicted_fhs_res_hist_11_new_folded_hist_T_4 | _GEN_11923; // @[FrontendBundle.scala 290:29]
  wire [7:0] s2_possible_predicted_fhs_res_hist_11_new_folded_hist_2 =
    _s2_possible_predicted_fhs_res_hist_11_new_folded_hist_T_5[7:0]; // @[FrontendBundle.scala 290:37]
  wire  s2_possible_predicted_fhs_res_hist_12_new_folded_hist_xored_res_2_4 = s2_possible_predicted_fhs_ob_4_1 ^
    s2_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__4; // @[FrontendBundle.scala 256:48]
  wire  s2_possible_predicted_fhs_res_hist_12_new_folded_hist_xored_res_2_5 =
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[1] ^ s2_possible_predicted_fhs_ob_4_0 ^
    s2_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__5; // @[FrontendBundle.scala 256:48]
  wire  s2_possible_predicted_fhs_res_hist_12_new_folded_hist_xored_res_2_6 =
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[0] ^
    s2_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__6; // @[FrontendBundle.scala 256:48]
  wire [6:0] s2_possible_predicted_fhs_res_hist_12_new_folded_hist_xored_2 = {
    s2_possible_predicted_fhs_res_hist_12_new_folded_hist_xored_res_2_6,
    s2_possible_predicted_fhs_res_hist_12_new_folded_hist_xored_res_2_5,
    s2_possible_predicted_fhs_res_hist_12_new_folded_hist_xored_res_2_4,
    s2_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__3,
    s2_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__1,
    s2_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [13:0] s2_possible_predicted_fhs_res_hist_12_new_folded_hist_src_doubled_2 = {
    s2_possible_predicted_fhs_res_hist_12_new_folded_hist_xored_res_2_6,
    s2_possible_predicted_fhs_res_hist_12_new_folded_hist_xored_res_2_5,
    s2_possible_predicted_fhs_res_hist_12_new_folded_hist_xored_res_2_4,
    s2_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__3,
    s2_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__1,
    s2_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__0,
    s2_possible_predicted_fhs_res_hist_12_new_folded_hist_xored_2}; // @[Cat.scala 31:58]
  wire [6:0] s2_possible_predicted_fhs_res_hist_12_new_folded_hist_2 =
    s2_possible_predicted_fhs_res_hist_12_new_folded_hist_src_doubled_2[11:5]; // @[FrontendBundle.scala 221:30]
  wire  s2_possible_predicted_fhs_res_hist_13_new_folded_hist_xored_res_2_5 =
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[1] ^
    s2_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__5; // @[FrontendBundle.scala 256:48]
  wire [6:0] s2_possible_predicted_fhs_res_hist_13_new_folded_hist_xored_2 = {
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[0],
    s2_possible_predicted_fhs_res_hist_13_new_folded_hist_xored_res_2_5,
    s2_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__4,
    s2_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__3,
    s2_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__1,
    s2_possible_predicted_fhs_res_hist_13_new_folded_hist_xored_res_1_0}; // @[FrontendBundle.scala 258:11]
  wire [13:0] s2_possible_predicted_fhs_res_hist_13_new_folded_hist_src_doubled_2 = {
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[0],
    s2_possible_predicted_fhs_res_hist_13_new_folded_hist_xored_res_2_5,
    s2_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__4,
    s2_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__3,
    s2_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__1,
    s2_possible_predicted_fhs_res_hist_13_new_folded_hist_xored_res_1_0,
    s2_possible_predicted_fhs_res_hist_13_new_folded_hist_xored_2}; // @[Cat.scala 31:58]
  wire [6:0] s2_possible_predicted_fhs_res_hist_13_new_folded_hist_2 =
    s2_possible_predicted_fhs_res_hist_13_new_folded_hist_src_doubled_2[11:5]; // @[FrontendBundle.scala 221:30]
  wire  s2_possible_predicted_fhs_res_hist_14_new_folded_hist_xored_res_2_5 =
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[1] ^ s2_possible_predicted_fhs_ob_2_1 ^
    s2_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__5; // @[FrontendBundle.scala 256:48]
  wire  s2_possible_predicted_fhs_res_hist_14_new_folded_hist_xored_res_2_6 =
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[0] ^ s2_possible_predicted_fhs_ob_2_0 ^
    s2_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__6; // @[FrontendBundle.scala 256:48]
  wire [6:0] s2_possible_predicted_fhs_res_hist_14_new_folded_hist_xored_2 = {
    s2_possible_predicted_fhs_res_hist_14_new_folded_hist_xored_res_2_6,
    s2_possible_predicted_fhs_res_hist_14_new_folded_hist_xored_res_2_5,
    s2_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__4,
    s2_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__3,
    s2_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__1,
    s2_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [13:0] s2_possible_predicted_fhs_res_hist_14_new_folded_hist_src_doubled_2 = {
    s2_possible_predicted_fhs_res_hist_14_new_folded_hist_xored_res_2_6,
    s2_possible_predicted_fhs_res_hist_14_new_folded_hist_xored_res_2_5,
    s2_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__4,
    s2_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__3,
    s2_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__1,
    s2_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__0,
    s2_possible_predicted_fhs_res_hist_14_new_folded_hist_xored_2}; // @[Cat.scala 31:58]
  wire [6:0] s2_possible_predicted_fhs_res_hist_14_new_folded_hist_2 =
    s2_possible_predicted_fhs_res_hist_14_new_folded_hist_src_doubled_2[11:5]; // @[FrontendBundle.scala 221:30]
  wire  s2_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_res_2_7 = s2_possible_predicted_fhs_ob_2_1 ^
    s2_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__7; // @[FrontendBundle.scala 256:48]
  wire  s2_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_res_2_9 =
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[1] ^
    s2_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__9; // @[FrontendBundle.scala 256:48]
  wire  s2_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_res_2_10 =
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[0] ^
    s2_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__10; // @[FrontendBundle.scala 256:48]
  wire [10:0] s2_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_2 = {
    s2_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_res_2_10,
    s2_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_res_2_9,
    s2_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_res_1_8,
    s2_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_res_2_7,
    s2_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__6,
    s2_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__5,
    s2_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_lo}; // @[FrontendBundle.scala 258:11]
  wire [21:0] s2_possible_predicted_fhs_res_hist_15_new_folded_hist_src_doubled_2 = {
    s2_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_res_2_10,
    s2_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_res_2_9,
    s2_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_res_1_8,
    s2_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_res_2_7,
    s2_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__6,
    s2_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__5,
    s2_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_lo,
    s2_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_2}; // @[Cat.scala 31:58]
  wire [10:0] s2_possible_predicted_fhs_res_hist_15_new_folded_hist_2 =
    s2_possible_predicted_fhs_res_hist_15_new_folded_hist_src_doubled_2[19:9]; // @[FrontendBundle.scala 221:30]
  wire  s2_possible_predicted_fhs_res_hist_16_new_folded_hist_xored_res_2_0 = s2_possible_predicted_fhs_ob_13_1 ^
    s2_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__0; // @[FrontendBundle.scala 256:48]
  wire  s2_possible_predicted_fhs_res_hist_16_new_folded_hist_xored_res_2_6 =
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[1] ^
    s2_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__6; // @[FrontendBundle.scala 256:48]
  wire  s2_possible_predicted_fhs_res_hist_16_new_folded_hist_xored_res_2_7 =
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[0] ^
    s2_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__7; // @[FrontendBundle.scala 256:48]
  wire [7:0] s2_possible_predicted_fhs_res_hist_16_new_folded_hist_xored_2 = {
    s2_possible_predicted_fhs_res_hist_16_new_folded_hist_xored_res_2_7,
    s2_possible_predicted_fhs_res_hist_16_new_folded_hist_xored_res_2_6,
    s2_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__5,
    s2_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__4,
    s2_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__3,
    s2_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_16_new_folded_hist_xored_res_1_1,
    s2_possible_predicted_fhs_res_hist_16_new_folded_hist_xored_res_2_0}; // @[FrontendBundle.scala 258:11]
  wire [15:0] s2_possible_predicted_fhs_res_hist_16_new_folded_hist_src_doubled_2 = {
    s2_possible_predicted_fhs_res_hist_16_new_folded_hist_xored_res_2_7,
    s2_possible_predicted_fhs_res_hist_16_new_folded_hist_xored_res_2_6,
    s2_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__5,
    s2_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__4,
    s2_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__3,
    s2_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_16_new_folded_hist_xored_res_1_1,
    s2_possible_predicted_fhs_res_hist_16_new_folded_hist_xored_res_2_0,
    s2_possible_predicted_fhs_res_hist_16_new_folded_hist_xored_2}; // @[Cat.scala 31:58]
  wire [7:0] s2_possible_predicted_fhs_res_hist_16_new_folded_hist_2 =
    s2_possible_predicted_fhs_res_hist_16_new_folded_hist_src_doubled_2[13:6]; // @[FrontendBundle.scala 221:30]
  wire  s2_possible_predicted_fhs_res_hist_17_new_folded_hist_xored_res_2_3 = s2_possible_predicted_fhs_ob_4_1 ^
    s2_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__3; // @[FrontendBundle.scala 256:48]
  wire  s2_possible_predicted_fhs_res_hist_17_new_folded_hist_xored_res_2_6 =
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[1] ^
    s2_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__6; // @[FrontendBundle.scala 256:48]
  wire  s2_possible_predicted_fhs_res_hist_17_new_folded_hist_xored_res_2_7 =
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[0] ^
    s2_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__7; // @[FrontendBundle.scala 256:48]
  wire [7:0] s2_possible_predicted_fhs_res_hist_17_new_folded_hist_xored_2 = {
    s2_possible_predicted_fhs_res_hist_17_new_folded_hist_xored_res_2_7,
    s2_possible_predicted_fhs_res_hist_17_new_folded_hist_xored_res_2_6,
    s2_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__5,
    s2_possible_predicted_fhs_res_hist_17_new_folded_hist_xored_res_1_4,
    s2_possible_predicted_fhs_res_hist_17_new_folded_hist_xored_res_2_3,
    s2_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__1,
    s2_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [15:0] s2_possible_predicted_fhs_res_hist_17_new_folded_hist_src_doubled_2 = {
    s2_possible_predicted_fhs_res_hist_17_new_folded_hist_xored_res_2_7,
    s2_possible_predicted_fhs_res_hist_17_new_folded_hist_xored_res_2_6,
    s2_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__5,
    s2_possible_predicted_fhs_res_hist_17_new_folded_hist_xored_res_1_4,
    s2_possible_predicted_fhs_res_hist_17_new_folded_hist_xored_res_2_3,
    s2_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__2,
    s2_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__1,
    s2_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__0,
    s2_possible_predicted_fhs_res_hist_17_new_folded_hist_xored_2}; // @[Cat.scala 31:58]
  wire [7:0] s2_possible_predicted_fhs_res_hist_17_new_folded_hist_2 =
    s2_possible_predicted_fhs_res_hist_17_new_folded_hist_src_doubled_2[13:6]; // @[FrontendBundle.scala 221:30]
  wire [7:0] _s2_predicted_fh_T_61 = _s2_redirect_s1_last_pred_vec_T_12 ?
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _s2_predicted_fh_T_62 = _s2_redirect_s1_last_pred_vec_T_40 ?
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _s2_predicted_fh_T_63 = _s2_redirect_s1_last_pred_vec_T_68 ?
    s2_possible_predicted_fhs_res_hist_0_new_folded_hist_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _s2_predicted_fh_T_64 = _s2_predicted_fh_T_61 | _s2_predicted_fh_T_62; // @[Mux.scala 27:73]
  wire [7:0] _s2_predicted_fh_T_66 = _s2_redirect_s1_last_pred_vec_T_12 ?
    s2_possible_predicted_fhs_res_hist_1_new_folded_hist : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _s2_predicted_fh_T_67 = _s2_redirect_s1_last_pred_vec_T_40 ?
    s2_possible_predicted_fhs_res_hist_1_new_folded_hist_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _s2_predicted_fh_T_68 = _s2_redirect_s1_last_pred_vec_T_68 ?
    s2_possible_predicted_fhs_res_hist_1_new_folded_hist_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _s2_predicted_fh_T_69 = _s2_predicted_fh_T_66 | _s2_predicted_fh_T_67; // @[Mux.scala 27:73]
  wire [7:0] _s2_predicted_fh_T_71 = _s2_redirect_s1_last_pred_vec_T_12 ?
    s2_possible_predicted_fhs_res_hist_2_new_folded_hist : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _s2_predicted_fh_T_72 = _s2_redirect_s1_last_pred_vec_T_40 ?
    s2_possible_predicted_fhs_res_hist_2_new_folded_hist_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _s2_predicted_fh_T_73 = _s2_redirect_s1_last_pred_vec_T_68 ?
    s2_possible_predicted_fhs_res_hist_2_new_folded_hist_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _s2_predicted_fh_T_74 = _s2_predicted_fh_T_71 | _s2_predicted_fh_T_72; // @[Mux.scala 27:73]
  wire [10:0] _s2_predicted_fh_T_76 = _s2_redirect_s1_last_pred_vec_T_12 ?
    s2_possible_predicted_fhs_res_hist_3_new_folded_hist : 11'h0; // @[Mux.scala 27:73]
  wire [10:0] _s2_predicted_fh_T_77 = _s2_redirect_s1_last_pred_vec_T_40 ?
    s2_possible_predicted_fhs_res_hist_3_new_folded_hist_1 : 11'h0; // @[Mux.scala 27:73]
  wire [10:0] _s2_predicted_fh_T_78 = _s2_redirect_s1_last_pred_vec_T_68 ?
    s2_possible_predicted_fhs_res_hist_3_new_folded_hist_2 : 11'h0; // @[Mux.scala 27:73]
  wire [10:0] _s2_predicted_fh_T_79 = _s2_predicted_fh_T_76 | _s2_predicted_fh_T_77; // @[Mux.scala 27:73]
  wire [3:0] _s2_predicted_fh_T_81 = _s2_redirect_s1_last_pred_vec_T_12 ? s2_folded_gh_hist_4_folded_hist : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _s2_predicted_fh_T_82 = _s2_redirect_s1_last_pred_vec_T_40 ?
    s2_possible_predicted_fhs_res_hist_4_new_folded_hist_1 : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _s2_predicted_fh_T_83 = _s2_redirect_s1_last_pred_vec_T_68 ?
    s2_possible_predicted_fhs_res_hist_4_new_folded_hist_2 : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _s2_predicted_fh_T_84 = _s2_predicted_fh_T_81 | _s2_predicted_fh_T_82; // @[Mux.scala 27:73]
  wire [10:0] _s2_predicted_fh_T_86 = _s2_redirect_s1_last_pred_vec_T_12 ?
    s2_possible_predicted_fhs_res_hist_5_new_folded_hist : 11'h0; // @[Mux.scala 27:73]
  wire [10:0] _s2_predicted_fh_T_87 = _s2_redirect_s1_last_pred_vec_T_40 ?
    s2_possible_predicted_fhs_res_hist_5_new_folded_hist_1 : 11'h0; // @[Mux.scala 27:73]
  wire [10:0] _s2_predicted_fh_T_88 = _s2_redirect_s1_last_pred_vec_T_68 ?
    s2_possible_predicted_fhs_res_hist_5_new_folded_hist_2 : 11'h0; // @[Mux.scala 27:73]
  wire [10:0] _s2_predicted_fh_T_89 = _s2_predicted_fh_T_86 | _s2_predicted_fh_T_87; // @[Mux.scala 27:73]
  wire [8:0] _s2_predicted_fh_T_91 = _s2_redirect_s1_last_pred_vec_T_12 ?
    s2_possible_predicted_fhs_res_hist_6_new_folded_hist : 9'h0; // @[Mux.scala 27:73]
  wire [8:0] _s2_predicted_fh_T_92 = _s2_redirect_s1_last_pred_vec_T_40 ?
    s2_possible_predicted_fhs_res_hist_6_new_folded_hist_1 : 9'h0; // @[Mux.scala 27:73]
  wire [8:0] _s2_predicted_fh_T_93 = _s2_redirect_s1_last_pred_vec_T_68 ?
    s2_possible_predicted_fhs_res_hist_6_new_folded_hist_2 : 9'h0; // @[Mux.scala 27:73]
  wire [8:0] _s2_predicted_fh_T_94 = _s2_predicted_fh_T_91 | _s2_predicted_fh_T_92; // @[Mux.scala 27:73]
  wire [8:0] _s2_predicted_fh_T_96 = _s2_redirect_s1_last_pred_vec_T_12 ?
    s2_possible_predicted_fhs_res_hist_7_new_folded_hist : 9'h0; // @[Mux.scala 27:73]
  wire [8:0] _s2_predicted_fh_T_97 = _s2_redirect_s1_last_pred_vec_T_40 ?
    s2_possible_predicted_fhs_res_hist_7_new_folded_hist_1 : 9'h0; // @[Mux.scala 27:73]
  wire [8:0] _s2_predicted_fh_T_98 = _s2_redirect_s1_last_pred_vec_T_68 ?
    s2_possible_predicted_fhs_res_hist_7_new_folded_hist_2 : 9'h0; // @[Mux.scala 27:73]
  wire [8:0] _s2_predicted_fh_T_99 = _s2_predicted_fh_T_96 | _s2_predicted_fh_T_97; // @[Mux.scala 27:73]
  wire [7:0] _s2_predicted_fh_T_101 = _s2_redirect_s1_last_pred_vec_T_12 ? s2_folded_gh_hist_8_folded_hist : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _s2_predicted_fh_T_102 = _s2_redirect_s1_last_pred_vec_T_40 ?
    s2_possible_predicted_fhs_res_hist_8_new_folded_hist_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _s2_predicted_fh_T_103 = _s2_redirect_s1_last_pred_vec_T_68 ?
    s2_possible_predicted_fhs_res_hist_8_new_folded_hist_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _s2_predicted_fh_T_104 = _s2_predicted_fh_T_101 | _s2_predicted_fh_T_102; // @[Mux.scala 27:73]
  wire [6:0] _s2_predicted_fh_T_106 = _s2_redirect_s1_last_pred_vec_T_12 ?
    s2_possible_predicted_fhs_res_hist_9_new_folded_hist : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _s2_predicted_fh_T_107 = _s2_redirect_s1_last_pred_vec_T_40 ?
    s2_possible_predicted_fhs_res_hist_9_new_folded_hist_1 : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _s2_predicted_fh_T_108 = _s2_redirect_s1_last_pred_vec_T_68 ?
    s2_possible_predicted_fhs_res_hist_9_new_folded_hist_2 : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _s2_predicted_fh_T_109 = _s2_predicted_fh_T_106 | _s2_predicted_fh_T_107; // @[Mux.scala 27:73]
  wire [8:0] _s2_predicted_fh_T_111 = _s2_redirect_s1_last_pred_vec_T_12 ?
    s2_possible_predicted_fhs_res_hist_10_new_folded_hist : 9'h0; // @[Mux.scala 27:73]
  wire [8:0] _s2_predicted_fh_T_112 = _s2_redirect_s1_last_pred_vec_T_40 ?
    s2_possible_predicted_fhs_res_hist_10_new_folded_hist_1 : 9'h0; // @[Mux.scala 27:73]
  wire [8:0] _s2_predicted_fh_T_113 = _s2_redirect_s1_last_pred_vec_T_68 ?
    s2_possible_predicted_fhs_res_hist_10_new_folded_hist_2 : 9'h0; // @[Mux.scala 27:73]
  wire [8:0] _s2_predicted_fh_T_114 = _s2_predicted_fh_T_111 | _s2_predicted_fh_T_112; // @[Mux.scala 27:73]
  wire [7:0] _s2_predicted_fh_T_116 = _s2_redirect_s1_last_pred_vec_T_12 ? s2_folded_gh_hist_11_folded_hist : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _s2_predicted_fh_T_117 = _s2_redirect_s1_last_pred_vec_T_40 ?
    s2_possible_predicted_fhs_res_hist_11_new_folded_hist_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _s2_predicted_fh_T_118 = _s2_redirect_s1_last_pred_vec_T_68 ?
    s2_possible_predicted_fhs_res_hist_11_new_folded_hist_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _s2_predicted_fh_T_119 = _s2_predicted_fh_T_116 | _s2_predicted_fh_T_117; // @[Mux.scala 27:73]
  wire [6:0] _s2_predicted_fh_T_121 = _s2_redirect_s1_last_pred_vec_T_12 ?
    s2_possible_predicted_fhs_res_hist_12_new_folded_hist : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _s2_predicted_fh_T_122 = _s2_redirect_s1_last_pred_vec_T_40 ?
    s2_possible_predicted_fhs_res_hist_12_new_folded_hist_1 : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _s2_predicted_fh_T_123 = _s2_redirect_s1_last_pred_vec_T_68 ?
    s2_possible_predicted_fhs_res_hist_12_new_folded_hist_2 : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _s2_predicted_fh_T_124 = _s2_predicted_fh_T_121 | _s2_predicted_fh_T_122; // @[Mux.scala 27:73]
  wire [6:0] _s2_predicted_fh_T_126 = _s2_redirect_s1_last_pred_vec_T_12 ?
    s2_possible_predicted_fhs_res_hist_13_new_folded_hist : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _s2_predicted_fh_T_127 = _s2_redirect_s1_last_pred_vec_T_40 ?
    s2_possible_predicted_fhs_res_hist_13_new_folded_hist_1 : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _s2_predicted_fh_T_128 = _s2_redirect_s1_last_pred_vec_T_68 ?
    s2_possible_predicted_fhs_res_hist_13_new_folded_hist_2 : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _s2_predicted_fh_T_129 = _s2_predicted_fh_T_126 | _s2_predicted_fh_T_127; // @[Mux.scala 27:73]
  wire [6:0] _s2_predicted_fh_T_131 = _s2_redirect_s1_last_pred_vec_T_12 ?
    s2_possible_predicted_fhs_res_hist_14_new_folded_hist : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _s2_predicted_fh_T_132 = _s2_redirect_s1_last_pred_vec_T_40 ?
    s2_possible_predicted_fhs_res_hist_14_new_folded_hist_1 : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _s2_predicted_fh_T_133 = _s2_redirect_s1_last_pred_vec_T_68 ?
    s2_possible_predicted_fhs_res_hist_14_new_folded_hist_2 : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _s2_predicted_fh_T_134 = _s2_predicted_fh_T_131 | _s2_predicted_fh_T_132; // @[Mux.scala 27:73]
  wire [10:0] _s2_predicted_fh_T_136 = _s2_redirect_s1_last_pred_vec_T_12 ?
    s2_possible_predicted_fhs_res_hist_15_new_folded_hist : 11'h0; // @[Mux.scala 27:73]
  wire [10:0] _s2_predicted_fh_T_137 = _s2_redirect_s1_last_pred_vec_T_40 ?
    s2_possible_predicted_fhs_res_hist_15_new_folded_hist_1 : 11'h0; // @[Mux.scala 27:73]
  wire [10:0] _s2_predicted_fh_T_138 = _s2_redirect_s1_last_pred_vec_T_68 ?
    s2_possible_predicted_fhs_res_hist_15_new_folded_hist_2 : 11'h0; // @[Mux.scala 27:73]
  wire [10:0] _s2_predicted_fh_T_139 = _s2_predicted_fh_T_136 | _s2_predicted_fh_T_137; // @[Mux.scala 27:73]
  wire [7:0] _s2_predicted_fh_T_141 = _s2_redirect_s1_last_pred_vec_T_12 ?
    s2_possible_predicted_fhs_res_hist_16_new_folded_hist : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _s2_predicted_fh_T_142 = _s2_redirect_s1_last_pred_vec_T_40 ?
    s2_possible_predicted_fhs_res_hist_16_new_folded_hist_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _s2_predicted_fh_T_143 = _s2_redirect_s1_last_pred_vec_T_68 ?
    s2_possible_predicted_fhs_res_hist_16_new_folded_hist_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _s2_predicted_fh_T_144 = _s2_predicted_fh_T_141 | _s2_predicted_fh_T_142; // @[Mux.scala 27:73]
  wire [7:0] _s2_predicted_fh_T_146 = _s2_redirect_s1_last_pred_vec_T_12 ?
    s2_possible_predicted_fhs_res_hist_17_new_folded_hist : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _s2_predicted_fh_T_147 = _s2_redirect_s1_last_pred_vec_T_40 ?
    s2_possible_predicted_fhs_res_hist_17_new_folded_hist_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _s2_predicted_fh_T_148 = _s2_redirect_s1_last_pred_vec_T_68 ?
    s2_possible_predicted_fhs_res_hist_17_new_folded_hist_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _s2_predicted_fh_T_149 = _s2_predicted_fh_T_146 | _s2_predicted_fh_T_147; // @[Mux.scala 27:73]
  wire [8:0] new_value_20 = s2_ghist_ptr_value + 8'h74; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_121 = {1'h0,new_value_20}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_20 = $signed(_diff_T_121) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_20 = $signed(diff_20) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_40 = $signed(_diff_T_121) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_41 = reverse_flag_20 ? _new_ptr_value_T_40 : {{1'd0}, new_value_20}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_21 = s2_ghist_ptr_value + 8'h6; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_127 = {1'h0,new_value_21}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_21 = $signed(_diff_T_127) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_21 = $signed(diff_21) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_42 = $signed(_diff_T_127) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_43 = reverse_flag_21 ? _new_ptr_value_T_42 : {{1'd0}, new_value_21}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_22 = s2_ghist_ptr_value + 8'hb; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_133 = {1'h0,new_value_22}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_22 = $signed(_diff_T_133) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_22 = $signed(diff_22) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_44 = $signed(_diff_T_133) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_45 = reverse_flag_22 ? _new_ptr_value_T_44 : {{1'd0}, new_value_22}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_23 = s2_ghist_ptr_value + 8'hf; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_139 = {1'h0,new_value_23}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_23 = $signed(_diff_T_139) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_23 = $signed(diff_23) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_46 = $signed(_diff_T_139) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_47 = reverse_flag_23 ? _new_ptr_value_T_46 : {{1'd0}, new_value_23}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_24 = s2_ghist_ptr_value + 8'h1e; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_145 = {1'h0,new_value_24}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_24 = $signed(_diff_T_145) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_24 = $signed(diff_24) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_48 = $signed(_diff_T_145) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_49 = reverse_flag_24 ? _new_ptr_value_T_48 : {{1'd0}, new_value_24}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_25 = s2_ghist_ptr_value + 8'h75; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_151 = {1'h0,new_value_25}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_25 = $signed(_diff_T_151) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_25 = $signed(diff_25) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_50 = $signed(_diff_T_151) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_51 = reverse_flag_25 ? _new_ptr_value_T_50 : {{1'd0}, new_value_25}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_26 = s2_ghist_ptr_value + 8'h7; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_157 = {1'h0,new_value_26}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_26 = $signed(_diff_T_157) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_26 = $signed(diff_26) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_52 = $signed(_diff_T_157) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_53 = reverse_flag_26 ? _new_ptr_value_T_52 : {{1'd0}, new_value_26}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_27 = s2_ghist_ptr_value + 8'h76; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_163 = {1'h0,new_value_27}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_27 = $signed(_diff_T_163) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_27 = $signed(diff_27) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_54 = $signed(_diff_T_163) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_55 = reverse_flag_27 ? _new_ptr_value_T_54 : {{1'd0}, new_value_27}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_28 = s2_ghist_ptr_value + 8'h1d; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_169 = {1'h0,new_value_28}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_28 = $signed(_diff_T_169) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_28 = $signed(diff_28) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_56 = $signed(_diff_T_169) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_57 = reverse_flag_28 ? _new_ptr_value_T_56 : {{1'd0}, new_value_28}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_29 = s2_ghist_ptr_value + 8'ha; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_175 = {1'h0,new_value_29}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_29 = $signed(_diff_T_175) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_29 = $signed(diff_29) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_58 = $signed(_diff_T_175) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_59 = reverse_flag_29 ? _new_ptr_value_T_58 : {{1'd0}, new_value_29}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_30 = s2_ghist_ptr_value + 8'he; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_181 = {1'h0,new_value_30}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_30 = $signed(_diff_T_181) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_30 = $signed(diff_30) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_60 = $signed(_diff_T_181) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_61 = reverse_flag_30 ? _new_ptr_value_T_60 : {{1'd0}, new_value_30}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_31 = s2_ghist_ptr_value + 8'h77; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_187 = {1'h0,new_value_31}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_31 = $signed(_diff_T_187) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_31 = $signed(diff_31) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_62 = $signed(_diff_T_187) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_63 = reverse_flag_31 ? _new_ptr_value_T_62 : {{1'd0}, new_value_31}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_32 = s2_ghist_ptr_value + 8'hd; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_193 = {1'h0,new_value_32}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_32 = $signed(_diff_T_193) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_32 = $signed(diff_32) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_64 = $signed(_diff_T_193) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_65 = reverse_flag_32 ? _new_ptr_value_T_64 : {{1'd0}, new_value_32}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_33 = s2_ghist_ptr_value + 8'h8; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_199 = {1'h0,new_value_33}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_33 = $signed(_diff_T_199) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_33 = $signed(diff_33) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_66 = $signed(_diff_T_199) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_67 = reverse_flag_33 ? _new_ptr_value_T_66 : {{1'd0}, new_value_33}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_34 = s2_ghist_ptr_value + 8'h20; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_205 = {1'h0,new_value_34}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_34 = $signed(_diff_T_205) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_34 = $signed(diff_34) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_68 = $signed(_diff_T_205) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_69 = reverse_flag_34 ? _new_ptr_value_T_68 : {{1'd0}, new_value_34}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_35 = s2_ghist_ptr_value + 8'hc; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_211 = {1'h0,new_value_35}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_35 = $signed(_diff_T_211) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_35 = $signed(diff_35) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_70 = $signed(_diff_T_211) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_71 = reverse_flag_35 ? _new_ptr_value_T_70 : {{1'd0}, new_value_35}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_36 = s2_ghist_ptr_value + 8'h9; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_217 = {1'h0,new_value_36}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_36 = $signed(_diff_T_217) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_36 = $signed(diff_36) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_72 = $signed(_diff_T_217) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_73 = reverse_flag_36 ? _new_ptr_value_T_72 : {{1'd0}, new_value_36}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_37 = s2_ghist_ptr_value + 8'h1f; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_223 = {1'h0,new_value_37}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_37 = $signed(_diff_T_223) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_37 = $signed(diff_37) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_74 = $signed(_diff_T_223) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_75 = reverse_flag_37 ? _new_ptr_value_T_74 : {{1'd0}, new_value_37}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_38 = s2_ghist_ptr_value + 8'h5; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_229 = {1'h0,new_value_38}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_38 = $signed(_diff_T_229) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_38 = $signed(diff_38) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_76 = $signed(_diff_T_229) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_77 = reverse_flag_38 ? _new_ptr_value_T_76 : {{1'd0}, new_value_38}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_39 = s2_ghist_ptr_value + 8'h10; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_235 = {1'h0,new_value_39}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_39 = $signed(_diff_T_235) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_39 = $signed(diff_39) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_78 = $signed(_diff_T_235) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_79 = reverse_flag_39 ? _new_ptr_value_T_78 : {{1'd0}, new_value_39}; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] new_ptr_29_value = _new_ptr_value_T_59[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_3033 = 8'h1 == new_ptr_29_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3034 = 8'h2 == new_ptr_29_value ? ghv_2 : _GEN_3033; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3035 = 8'h3 == new_ptr_29_value ? ghv_3 : _GEN_3034; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3036 = 8'h4 == new_ptr_29_value ? ghv_4 : _GEN_3035; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3037 = 8'h5 == new_ptr_29_value ? ghv_5 : _GEN_3036; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3038 = 8'h6 == new_ptr_29_value ? ghv_6 : _GEN_3037; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3039 = 8'h7 == new_ptr_29_value ? ghv_7 : _GEN_3038; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3040 = 8'h8 == new_ptr_29_value ? ghv_8 : _GEN_3039; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3041 = 8'h9 == new_ptr_29_value ? ghv_9 : _GEN_3040; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3042 = 8'ha == new_ptr_29_value ? ghv_10 : _GEN_3041; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3043 = 8'hb == new_ptr_29_value ? ghv_11 : _GEN_3042; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3044 = 8'hc == new_ptr_29_value ? ghv_12 : _GEN_3043; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3045 = 8'hd == new_ptr_29_value ? ghv_13 : _GEN_3044; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3046 = 8'he == new_ptr_29_value ? ghv_14 : _GEN_3045; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3047 = 8'hf == new_ptr_29_value ? ghv_15 : _GEN_3046; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3048 = 8'h10 == new_ptr_29_value ? ghv_16 : _GEN_3047; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3049 = 8'h11 == new_ptr_29_value ? ghv_17 : _GEN_3048; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3050 = 8'h12 == new_ptr_29_value ? ghv_18 : _GEN_3049; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3051 = 8'h13 == new_ptr_29_value ? ghv_19 : _GEN_3050; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3052 = 8'h14 == new_ptr_29_value ? ghv_20 : _GEN_3051; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3053 = 8'h15 == new_ptr_29_value ? ghv_21 : _GEN_3052; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3054 = 8'h16 == new_ptr_29_value ? ghv_22 : _GEN_3053; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3055 = 8'h17 == new_ptr_29_value ? ghv_23 : _GEN_3054; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3056 = 8'h18 == new_ptr_29_value ? ghv_24 : _GEN_3055; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3057 = 8'h19 == new_ptr_29_value ? ghv_25 : _GEN_3056; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3058 = 8'h1a == new_ptr_29_value ? ghv_26 : _GEN_3057; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3059 = 8'h1b == new_ptr_29_value ? ghv_27 : _GEN_3058; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3060 = 8'h1c == new_ptr_29_value ? ghv_28 : _GEN_3059; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3061 = 8'h1d == new_ptr_29_value ? ghv_29 : _GEN_3060; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3062 = 8'h1e == new_ptr_29_value ? ghv_30 : _GEN_3061; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3063 = 8'h1f == new_ptr_29_value ? ghv_31 : _GEN_3062; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3064 = 8'h20 == new_ptr_29_value ? ghv_32 : _GEN_3063; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3065 = 8'h21 == new_ptr_29_value ? ghv_33 : _GEN_3064; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3066 = 8'h22 == new_ptr_29_value ? ghv_34 : _GEN_3065; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3067 = 8'h23 == new_ptr_29_value ? ghv_35 : _GEN_3066; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3068 = 8'h24 == new_ptr_29_value ? ghv_36 : _GEN_3067; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3069 = 8'h25 == new_ptr_29_value ? ghv_37 : _GEN_3068; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3070 = 8'h26 == new_ptr_29_value ? ghv_38 : _GEN_3069; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3071 = 8'h27 == new_ptr_29_value ? ghv_39 : _GEN_3070; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3072 = 8'h28 == new_ptr_29_value ? ghv_40 : _GEN_3071; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3073 = 8'h29 == new_ptr_29_value ? ghv_41 : _GEN_3072; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3074 = 8'h2a == new_ptr_29_value ? ghv_42 : _GEN_3073; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3075 = 8'h2b == new_ptr_29_value ? ghv_43 : _GEN_3074; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3076 = 8'h2c == new_ptr_29_value ? ghv_44 : _GEN_3075; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3077 = 8'h2d == new_ptr_29_value ? ghv_45 : _GEN_3076; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3078 = 8'h2e == new_ptr_29_value ? ghv_46 : _GEN_3077; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3079 = 8'h2f == new_ptr_29_value ? ghv_47 : _GEN_3078; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3080 = 8'h30 == new_ptr_29_value ? ghv_48 : _GEN_3079; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3081 = 8'h31 == new_ptr_29_value ? ghv_49 : _GEN_3080; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3082 = 8'h32 == new_ptr_29_value ? ghv_50 : _GEN_3081; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3083 = 8'h33 == new_ptr_29_value ? ghv_51 : _GEN_3082; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3084 = 8'h34 == new_ptr_29_value ? ghv_52 : _GEN_3083; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3085 = 8'h35 == new_ptr_29_value ? ghv_53 : _GEN_3084; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3086 = 8'h36 == new_ptr_29_value ? ghv_54 : _GEN_3085; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3087 = 8'h37 == new_ptr_29_value ? ghv_55 : _GEN_3086; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3088 = 8'h38 == new_ptr_29_value ? ghv_56 : _GEN_3087; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3089 = 8'h39 == new_ptr_29_value ? ghv_57 : _GEN_3088; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3090 = 8'h3a == new_ptr_29_value ? ghv_58 : _GEN_3089; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3091 = 8'h3b == new_ptr_29_value ? ghv_59 : _GEN_3090; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3092 = 8'h3c == new_ptr_29_value ? ghv_60 : _GEN_3091; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3093 = 8'h3d == new_ptr_29_value ? ghv_61 : _GEN_3092; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3094 = 8'h3e == new_ptr_29_value ? ghv_62 : _GEN_3093; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3095 = 8'h3f == new_ptr_29_value ? ghv_63 : _GEN_3094; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3096 = 8'h40 == new_ptr_29_value ? ghv_64 : _GEN_3095; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3097 = 8'h41 == new_ptr_29_value ? ghv_65 : _GEN_3096; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3098 = 8'h42 == new_ptr_29_value ? ghv_66 : _GEN_3097; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3099 = 8'h43 == new_ptr_29_value ? ghv_67 : _GEN_3098; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3100 = 8'h44 == new_ptr_29_value ? ghv_68 : _GEN_3099; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3101 = 8'h45 == new_ptr_29_value ? ghv_69 : _GEN_3100; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3102 = 8'h46 == new_ptr_29_value ? ghv_70 : _GEN_3101; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3103 = 8'h47 == new_ptr_29_value ? ghv_71 : _GEN_3102; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3104 = 8'h48 == new_ptr_29_value ? ghv_72 : _GEN_3103; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3105 = 8'h49 == new_ptr_29_value ? ghv_73 : _GEN_3104; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3106 = 8'h4a == new_ptr_29_value ? ghv_74 : _GEN_3105; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3107 = 8'h4b == new_ptr_29_value ? ghv_75 : _GEN_3106; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3108 = 8'h4c == new_ptr_29_value ? ghv_76 : _GEN_3107; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3109 = 8'h4d == new_ptr_29_value ? ghv_77 : _GEN_3108; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3110 = 8'h4e == new_ptr_29_value ? ghv_78 : _GEN_3109; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3111 = 8'h4f == new_ptr_29_value ? ghv_79 : _GEN_3110; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3112 = 8'h50 == new_ptr_29_value ? ghv_80 : _GEN_3111; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3113 = 8'h51 == new_ptr_29_value ? ghv_81 : _GEN_3112; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3114 = 8'h52 == new_ptr_29_value ? ghv_82 : _GEN_3113; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3115 = 8'h53 == new_ptr_29_value ? ghv_83 : _GEN_3114; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3116 = 8'h54 == new_ptr_29_value ? ghv_84 : _GEN_3115; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3117 = 8'h55 == new_ptr_29_value ? ghv_85 : _GEN_3116; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3118 = 8'h56 == new_ptr_29_value ? ghv_86 : _GEN_3117; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3119 = 8'h57 == new_ptr_29_value ? ghv_87 : _GEN_3118; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3120 = 8'h58 == new_ptr_29_value ? ghv_88 : _GEN_3119; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3121 = 8'h59 == new_ptr_29_value ? ghv_89 : _GEN_3120; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3122 = 8'h5a == new_ptr_29_value ? ghv_90 : _GEN_3121; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3123 = 8'h5b == new_ptr_29_value ? ghv_91 : _GEN_3122; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3124 = 8'h5c == new_ptr_29_value ? ghv_92 : _GEN_3123; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3125 = 8'h5d == new_ptr_29_value ? ghv_93 : _GEN_3124; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3126 = 8'h5e == new_ptr_29_value ? ghv_94 : _GEN_3125; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3127 = 8'h5f == new_ptr_29_value ? ghv_95 : _GEN_3126; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3128 = 8'h60 == new_ptr_29_value ? ghv_96 : _GEN_3127; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3129 = 8'h61 == new_ptr_29_value ? ghv_97 : _GEN_3128; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3130 = 8'h62 == new_ptr_29_value ? ghv_98 : _GEN_3129; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3131 = 8'h63 == new_ptr_29_value ? ghv_99 : _GEN_3130; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3132 = 8'h64 == new_ptr_29_value ? ghv_100 : _GEN_3131; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3133 = 8'h65 == new_ptr_29_value ? ghv_101 : _GEN_3132; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3134 = 8'h66 == new_ptr_29_value ? ghv_102 : _GEN_3133; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3135 = 8'h67 == new_ptr_29_value ? ghv_103 : _GEN_3134; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3136 = 8'h68 == new_ptr_29_value ? ghv_104 : _GEN_3135; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3137 = 8'h69 == new_ptr_29_value ? ghv_105 : _GEN_3136; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3138 = 8'h6a == new_ptr_29_value ? ghv_106 : _GEN_3137; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3139 = 8'h6b == new_ptr_29_value ? ghv_107 : _GEN_3138; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3140 = 8'h6c == new_ptr_29_value ? ghv_108 : _GEN_3139; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3141 = 8'h6d == new_ptr_29_value ? ghv_109 : _GEN_3140; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3142 = 8'h6e == new_ptr_29_value ? ghv_110 : _GEN_3141; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3143 = 8'h6f == new_ptr_29_value ? ghv_111 : _GEN_3142; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3144 = 8'h70 == new_ptr_29_value ? ghv_112 : _GEN_3143; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3145 = 8'h71 == new_ptr_29_value ? ghv_113 : _GEN_3144; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3146 = 8'h72 == new_ptr_29_value ? ghv_114 : _GEN_3145; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3147 = 8'h73 == new_ptr_29_value ? ghv_115 : _GEN_3146; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3148 = 8'h74 == new_ptr_29_value ? ghv_116 : _GEN_3147; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3149 = 8'h75 == new_ptr_29_value ? ghv_117 : _GEN_3148; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3150 = 8'h76 == new_ptr_29_value ? ghv_118 : _GEN_3149; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3151 = 8'h77 == new_ptr_29_value ? ghv_119 : _GEN_3150; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3152 = 8'h78 == new_ptr_29_value ? ghv_120 : _GEN_3151; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3153 = 8'h79 == new_ptr_29_value ? ghv_121 : _GEN_3152; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3154 = 8'h7a == new_ptr_29_value ? ghv_122 : _GEN_3153; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3155 = 8'h7b == new_ptr_29_value ? ghv_123 : _GEN_3154; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3156 = 8'h7c == new_ptr_29_value ? ghv_124 : _GEN_3155; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3157 = 8'h7d == new_ptr_29_value ? ghv_125 : _GEN_3156; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3158 = 8'h7e == new_ptr_29_value ? ghv_126 : _GEN_3157; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3159 = 8'h7f == new_ptr_29_value ? ghv_127 : _GEN_3158; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3160 = 8'h80 == new_ptr_29_value ? ghv_128 : _GEN_3159; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3161 = 8'h81 == new_ptr_29_value ? ghv_129 : _GEN_3160; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3162 = 8'h82 == new_ptr_29_value ? ghv_130 : _GEN_3161; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3163 = 8'h83 == new_ptr_29_value ? ghv_131 : _GEN_3162; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3164 = 8'h84 == new_ptr_29_value ? ghv_132 : _GEN_3163; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3165 = 8'h85 == new_ptr_29_value ? ghv_133 : _GEN_3164; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3166 = 8'h86 == new_ptr_29_value ? ghv_134 : _GEN_3165; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3167 = 8'h87 == new_ptr_29_value ? ghv_135 : _GEN_3166; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3168 = 8'h88 == new_ptr_29_value ? ghv_136 : _GEN_3167; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3169 = 8'h89 == new_ptr_29_value ? ghv_137 : _GEN_3168; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3170 = 8'h8a == new_ptr_29_value ? ghv_138 : _GEN_3169; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3171 = 8'h8b == new_ptr_29_value ? ghv_139 : _GEN_3170; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3172 = 8'h8c == new_ptr_29_value ? ghv_140 : _GEN_3171; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3173 = 8'h8d == new_ptr_29_value ? ghv_141 : _GEN_3172; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3174 = 8'h8e == new_ptr_29_value ? ghv_142 : _GEN_3173; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_36_value = _new_ptr_value_T_73[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_3177 = 8'h1 == new_ptr_36_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3178 = 8'h2 == new_ptr_36_value ? ghv_2 : _GEN_3177; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3179 = 8'h3 == new_ptr_36_value ? ghv_3 : _GEN_3178; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3180 = 8'h4 == new_ptr_36_value ? ghv_4 : _GEN_3179; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3181 = 8'h5 == new_ptr_36_value ? ghv_5 : _GEN_3180; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3182 = 8'h6 == new_ptr_36_value ? ghv_6 : _GEN_3181; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3183 = 8'h7 == new_ptr_36_value ? ghv_7 : _GEN_3182; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3184 = 8'h8 == new_ptr_36_value ? ghv_8 : _GEN_3183; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3185 = 8'h9 == new_ptr_36_value ? ghv_9 : _GEN_3184; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3186 = 8'ha == new_ptr_36_value ? ghv_10 : _GEN_3185; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3187 = 8'hb == new_ptr_36_value ? ghv_11 : _GEN_3186; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3188 = 8'hc == new_ptr_36_value ? ghv_12 : _GEN_3187; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3189 = 8'hd == new_ptr_36_value ? ghv_13 : _GEN_3188; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3190 = 8'he == new_ptr_36_value ? ghv_14 : _GEN_3189; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3191 = 8'hf == new_ptr_36_value ? ghv_15 : _GEN_3190; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3192 = 8'h10 == new_ptr_36_value ? ghv_16 : _GEN_3191; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3193 = 8'h11 == new_ptr_36_value ? ghv_17 : _GEN_3192; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3194 = 8'h12 == new_ptr_36_value ? ghv_18 : _GEN_3193; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3195 = 8'h13 == new_ptr_36_value ? ghv_19 : _GEN_3194; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3196 = 8'h14 == new_ptr_36_value ? ghv_20 : _GEN_3195; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3197 = 8'h15 == new_ptr_36_value ? ghv_21 : _GEN_3196; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3198 = 8'h16 == new_ptr_36_value ? ghv_22 : _GEN_3197; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3199 = 8'h17 == new_ptr_36_value ? ghv_23 : _GEN_3198; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3200 = 8'h18 == new_ptr_36_value ? ghv_24 : _GEN_3199; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3201 = 8'h19 == new_ptr_36_value ? ghv_25 : _GEN_3200; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3202 = 8'h1a == new_ptr_36_value ? ghv_26 : _GEN_3201; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3203 = 8'h1b == new_ptr_36_value ? ghv_27 : _GEN_3202; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3204 = 8'h1c == new_ptr_36_value ? ghv_28 : _GEN_3203; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3205 = 8'h1d == new_ptr_36_value ? ghv_29 : _GEN_3204; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3206 = 8'h1e == new_ptr_36_value ? ghv_30 : _GEN_3205; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3207 = 8'h1f == new_ptr_36_value ? ghv_31 : _GEN_3206; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3208 = 8'h20 == new_ptr_36_value ? ghv_32 : _GEN_3207; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3209 = 8'h21 == new_ptr_36_value ? ghv_33 : _GEN_3208; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3210 = 8'h22 == new_ptr_36_value ? ghv_34 : _GEN_3209; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3211 = 8'h23 == new_ptr_36_value ? ghv_35 : _GEN_3210; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3212 = 8'h24 == new_ptr_36_value ? ghv_36 : _GEN_3211; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3213 = 8'h25 == new_ptr_36_value ? ghv_37 : _GEN_3212; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3214 = 8'h26 == new_ptr_36_value ? ghv_38 : _GEN_3213; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3215 = 8'h27 == new_ptr_36_value ? ghv_39 : _GEN_3214; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3216 = 8'h28 == new_ptr_36_value ? ghv_40 : _GEN_3215; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3217 = 8'h29 == new_ptr_36_value ? ghv_41 : _GEN_3216; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3218 = 8'h2a == new_ptr_36_value ? ghv_42 : _GEN_3217; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3219 = 8'h2b == new_ptr_36_value ? ghv_43 : _GEN_3218; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3220 = 8'h2c == new_ptr_36_value ? ghv_44 : _GEN_3219; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3221 = 8'h2d == new_ptr_36_value ? ghv_45 : _GEN_3220; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3222 = 8'h2e == new_ptr_36_value ? ghv_46 : _GEN_3221; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3223 = 8'h2f == new_ptr_36_value ? ghv_47 : _GEN_3222; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3224 = 8'h30 == new_ptr_36_value ? ghv_48 : _GEN_3223; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3225 = 8'h31 == new_ptr_36_value ? ghv_49 : _GEN_3224; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3226 = 8'h32 == new_ptr_36_value ? ghv_50 : _GEN_3225; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3227 = 8'h33 == new_ptr_36_value ? ghv_51 : _GEN_3226; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3228 = 8'h34 == new_ptr_36_value ? ghv_52 : _GEN_3227; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3229 = 8'h35 == new_ptr_36_value ? ghv_53 : _GEN_3228; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3230 = 8'h36 == new_ptr_36_value ? ghv_54 : _GEN_3229; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3231 = 8'h37 == new_ptr_36_value ? ghv_55 : _GEN_3230; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3232 = 8'h38 == new_ptr_36_value ? ghv_56 : _GEN_3231; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3233 = 8'h39 == new_ptr_36_value ? ghv_57 : _GEN_3232; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3234 = 8'h3a == new_ptr_36_value ? ghv_58 : _GEN_3233; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3235 = 8'h3b == new_ptr_36_value ? ghv_59 : _GEN_3234; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3236 = 8'h3c == new_ptr_36_value ? ghv_60 : _GEN_3235; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3237 = 8'h3d == new_ptr_36_value ? ghv_61 : _GEN_3236; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3238 = 8'h3e == new_ptr_36_value ? ghv_62 : _GEN_3237; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3239 = 8'h3f == new_ptr_36_value ? ghv_63 : _GEN_3238; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3240 = 8'h40 == new_ptr_36_value ? ghv_64 : _GEN_3239; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3241 = 8'h41 == new_ptr_36_value ? ghv_65 : _GEN_3240; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3242 = 8'h42 == new_ptr_36_value ? ghv_66 : _GEN_3241; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3243 = 8'h43 == new_ptr_36_value ? ghv_67 : _GEN_3242; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3244 = 8'h44 == new_ptr_36_value ? ghv_68 : _GEN_3243; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3245 = 8'h45 == new_ptr_36_value ? ghv_69 : _GEN_3244; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3246 = 8'h46 == new_ptr_36_value ? ghv_70 : _GEN_3245; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3247 = 8'h47 == new_ptr_36_value ? ghv_71 : _GEN_3246; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3248 = 8'h48 == new_ptr_36_value ? ghv_72 : _GEN_3247; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3249 = 8'h49 == new_ptr_36_value ? ghv_73 : _GEN_3248; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3250 = 8'h4a == new_ptr_36_value ? ghv_74 : _GEN_3249; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3251 = 8'h4b == new_ptr_36_value ? ghv_75 : _GEN_3250; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3252 = 8'h4c == new_ptr_36_value ? ghv_76 : _GEN_3251; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3253 = 8'h4d == new_ptr_36_value ? ghv_77 : _GEN_3252; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3254 = 8'h4e == new_ptr_36_value ? ghv_78 : _GEN_3253; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3255 = 8'h4f == new_ptr_36_value ? ghv_79 : _GEN_3254; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3256 = 8'h50 == new_ptr_36_value ? ghv_80 : _GEN_3255; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3257 = 8'h51 == new_ptr_36_value ? ghv_81 : _GEN_3256; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3258 = 8'h52 == new_ptr_36_value ? ghv_82 : _GEN_3257; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3259 = 8'h53 == new_ptr_36_value ? ghv_83 : _GEN_3258; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3260 = 8'h54 == new_ptr_36_value ? ghv_84 : _GEN_3259; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3261 = 8'h55 == new_ptr_36_value ? ghv_85 : _GEN_3260; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3262 = 8'h56 == new_ptr_36_value ? ghv_86 : _GEN_3261; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3263 = 8'h57 == new_ptr_36_value ? ghv_87 : _GEN_3262; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3264 = 8'h58 == new_ptr_36_value ? ghv_88 : _GEN_3263; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3265 = 8'h59 == new_ptr_36_value ? ghv_89 : _GEN_3264; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3266 = 8'h5a == new_ptr_36_value ? ghv_90 : _GEN_3265; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3267 = 8'h5b == new_ptr_36_value ? ghv_91 : _GEN_3266; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3268 = 8'h5c == new_ptr_36_value ? ghv_92 : _GEN_3267; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3269 = 8'h5d == new_ptr_36_value ? ghv_93 : _GEN_3268; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3270 = 8'h5e == new_ptr_36_value ? ghv_94 : _GEN_3269; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3271 = 8'h5f == new_ptr_36_value ? ghv_95 : _GEN_3270; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3272 = 8'h60 == new_ptr_36_value ? ghv_96 : _GEN_3271; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3273 = 8'h61 == new_ptr_36_value ? ghv_97 : _GEN_3272; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3274 = 8'h62 == new_ptr_36_value ? ghv_98 : _GEN_3273; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3275 = 8'h63 == new_ptr_36_value ? ghv_99 : _GEN_3274; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3276 = 8'h64 == new_ptr_36_value ? ghv_100 : _GEN_3275; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3277 = 8'h65 == new_ptr_36_value ? ghv_101 : _GEN_3276; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3278 = 8'h66 == new_ptr_36_value ? ghv_102 : _GEN_3277; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3279 = 8'h67 == new_ptr_36_value ? ghv_103 : _GEN_3278; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3280 = 8'h68 == new_ptr_36_value ? ghv_104 : _GEN_3279; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3281 = 8'h69 == new_ptr_36_value ? ghv_105 : _GEN_3280; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3282 = 8'h6a == new_ptr_36_value ? ghv_106 : _GEN_3281; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3283 = 8'h6b == new_ptr_36_value ? ghv_107 : _GEN_3282; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3284 = 8'h6c == new_ptr_36_value ? ghv_108 : _GEN_3283; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3285 = 8'h6d == new_ptr_36_value ? ghv_109 : _GEN_3284; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3286 = 8'h6e == new_ptr_36_value ? ghv_110 : _GEN_3285; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3287 = 8'h6f == new_ptr_36_value ? ghv_111 : _GEN_3286; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3288 = 8'h70 == new_ptr_36_value ? ghv_112 : _GEN_3287; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3289 = 8'h71 == new_ptr_36_value ? ghv_113 : _GEN_3288; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3290 = 8'h72 == new_ptr_36_value ? ghv_114 : _GEN_3289; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3291 = 8'h73 == new_ptr_36_value ? ghv_115 : _GEN_3290; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3292 = 8'h74 == new_ptr_36_value ? ghv_116 : _GEN_3291; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3293 = 8'h75 == new_ptr_36_value ? ghv_117 : _GEN_3292; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3294 = 8'h76 == new_ptr_36_value ? ghv_118 : _GEN_3293; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3295 = 8'h77 == new_ptr_36_value ? ghv_119 : _GEN_3294; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3296 = 8'h78 == new_ptr_36_value ? ghv_120 : _GEN_3295; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3297 = 8'h79 == new_ptr_36_value ? ghv_121 : _GEN_3296; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3298 = 8'h7a == new_ptr_36_value ? ghv_122 : _GEN_3297; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3299 = 8'h7b == new_ptr_36_value ? ghv_123 : _GEN_3298; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3300 = 8'h7c == new_ptr_36_value ? ghv_124 : _GEN_3299; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3301 = 8'h7d == new_ptr_36_value ? ghv_125 : _GEN_3300; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3302 = 8'h7e == new_ptr_36_value ? ghv_126 : _GEN_3301; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3303 = 8'h7f == new_ptr_36_value ? ghv_127 : _GEN_3302; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3304 = 8'h80 == new_ptr_36_value ? ghv_128 : _GEN_3303; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3305 = 8'h81 == new_ptr_36_value ? ghv_129 : _GEN_3304; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3306 = 8'h82 == new_ptr_36_value ? ghv_130 : _GEN_3305; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3307 = 8'h83 == new_ptr_36_value ? ghv_131 : _GEN_3306; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3308 = 8'h84 == new_ptr_36_value ? ghv_132 : _GEN_3307; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3309 = 8'h85 == new_ptr_36_value ? ghv_133 : _GEN_3308; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3310 = 8'h86 == new_ptr_36_value ? ghv_134 : _GEN_3309; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3311 = 8'h87 == new_ptr_36_value ? ghv_135 : _GEN_3310; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3312 = 8'h88 == new_ptr_36_value ? ghv_136 : _GEN_3311; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3313 = 8'h89 == new_ptr_36_value ? ghv_137 : _GEN_3312; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3314 = 8'h8a == new_ptr_36_value ? ghv_138 : _GEN_3313; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3315 = 8'h8b == new_ptr_36_value ? ghv_139 : _GEN_3314; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3316 = 8'h8c == new_ptr_36_value ? ghv_140 : _GEN_3315; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3317 = 8'h8d == new_ptr_36_value ? ghv_141 : _GEN_3316; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3318 = 8'h8e == new_ptr_36_value ? ghv_142 : _GEN_3317; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_33_value = _new_ptr_value_T_67[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_3321 = 8'h1 == new_ptr_33_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3322 = 8'h2 == new_ptr_33_value ? ghv_2 : _GEN_3321; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3323 = 8'h3 == new_ptr_33_value ? ghv_3 : _GEN_3322; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3324 = 8'h4 == new_ptr_33_value ? ghv_4 : _GEN_3323; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3325 = 8'h5 == new_ptr_33_value ? ghv_5 : _GEN_3324; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3326 = 8'h6 == new_ptr_33_value ? ghv_6 : _GEN_3325; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3327 = 8'h7 == new_ptr_33_value ? ghv_7 : _GEN_3326; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3328 = 8'h8 == new_ptr_33_value ? ghv_8 : _GEN_3327; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3329 = 8'h9 == new_ptr_33_value ? ghv_9 : _GEN_3328; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3330 = 8'ha == new_ptr_33_value ? ghv_10 : _GEN_3329; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3331 = 8'hb == new_ptr_33_value ? ghv_11 : _GEN_3330; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3332 = 8'hc == new_ptr_33_value ? ghv_12 : _GEN_3331; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3333 = 8'hd == new_ptr_33_value ? ghv_13 : _GEN_3332; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3334 = 8'he == new_ptr_33_value ? ghv_14 : _GEN_3333; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3335 = 8'hf == new_ptr_33_value ? ghv_15 : _GEN_3334; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3336 = 8'h10 == new_ptr_33_value ? ghv_16 : _GEN_3335; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3337 = 8'h11 == new_ptr_33_value ? ghv_17 : _GEN_3336; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3338 = 8'h12 == new_ptr_33_value ? ghv_18 : _GEN_3337; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3339 = 8'h13 == new_ptr_33_value ? ghv_19 : _GEN_3338; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3340 = 8'h14 == new_ptr_33_value ? ghv_20 : _GEN_3339; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3341 = 8'h15 == new_ptr_33_value ? ghv_21 : _GEN_3340; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3342 = 8'h16 == new_ptr_33_value ? ghv_22 : _GEN_3341; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3343 = 8'h17 == new_ptr_33_value ? ghv_23 : _GEN_3342; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3344 = 8'h18 == new_ptr_33_value ? ghv_24 : _GEN_3343; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3345 = 8'h19 == new_ptr_33_value ? ghv_25 : _GEN_3344; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3346 = 8'h1a == new_ptr_33_value ? ghv_26 : _GEN_3345; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3347 = 8'h1b == new_ptr_33_value ? ghv_27 : _GEN_3346; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3348 = 8'h1c == new_ptr_33_value ? ghv_28 : _GEN_3347; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3349 = 8'h1d == new_ptr_33_value ? ghv_29 : _GEN_3348; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3350 = 8'h1e == new_ptr_33_value ? ghv_30 : _GEN_3349; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3351 = 8'h1f == new_ptr_33_value ? ghv_31 : _GEN_3350; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3352 = 8'h20 == new_ptr_33_value ? ghv_32 : _GEN_3351; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3353 = 8'h21 == new_ptr_33_value ? ghv_33 : _GEN_3352; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3354 = 8'h22 == new_ptr_33_value ? ghv_34 : _GEN_3353; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3355 = 8'h23 == new_ptr_33_value ? ghv_35 : _GEN_3354; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3356 = 8'h24 == new_ptr_33_value ? ghv_36 : _GEN_3355; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3357 = 8'h25 == new_ptr_33_value ? ghv_37 : _GEN_3356; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3358 = 8'h26 == new_ptr_33_value ? ghv_38 : _GEN_3357; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3359 = 8'h27 == new_ptr_33_value ? ghv_39 : _GEN_3358; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3360 = 8'h28 == new_ptr_33_value ? ghv_40 : _GEN_3359; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3361 = 8'h29 == new_ptr_33_value ? ghv_41 : _GEN_3360; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3362 = 8'h2a == new_ptr_33_value ? ghv_42 : _GEN_3361; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3363 = 8'h2b == new_ptr_33_value ? ghv_43 : _GEN_3362; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3364 = 8'h2c == new_ptr_33_value ? ghv_44 : _GEN_3363; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3365 = 8'h2d == new_ptr_33_value ? ghv_45 : _GEN_3364; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3366 = 8'h2e == new_ptr_33_value ? ghv_46 : _GEN_3365; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3367 = 8'h2f == new_ptr_33_value ? ghv_47 : _GEN_3366; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3368 = 8'h30 == new_ptr_33_value ? ghv_48 : _GEN_3367; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3369 = 8'h31 == new_ptr_33_value ? ghv_49 : _GEN_3368; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3370 = 8'h32 == new_ptr_33_value ? ghv_50 : _GEN_3369; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3371 = 8'h33 == new_ptr_33_value ? ghv_51 : _GEN_3370; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3372 = 8'h34 == new_ptr_33_value ? ghv_52 : _GEN_3371; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3373 = 8'h35 == new_ptr_33_value ? ghv_53 : _GEN_3372; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3374 = 8'h36 == new_ptr_33_value ? ghv_54 : _GEN_3373; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3375 = 8'h37 == new_ptr_33_value ? ghv_55 : _GEN_3374; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3376 = 8'h38 == new_ptr_33_value ? ghv_56 : _GEN_3375; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3377 = 8'h39 == new_ptr_33_value ? ghv_57 : _GEN_3376; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3378 = 8'h3a == new_ptr_33_value ? ghv_58 : _GEN_3377; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3379 = 8'h3b == new_ptr_33_value ? ghv_59 : _GEN_3378; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3380 = 8'h3c == new_ptr_33_value ? ghv_60 : _GEN_3379; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3381 = 8'h3d == new_ptr_33_value ? ghv_61 : _GEN_3380; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3382 = 8'h3e == new_ptr_33_value ? ghv_62 : _GEN_3381; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3383 = 8'h3f == new_ptr_33_value ? ghv_63 : _GEN_3382; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3384 = 8'h40 == new_ptr_33_value ? ghv_64 : _GEN_3383; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3385 = 8'h41 == new_ptr_33_value ? ghv_65 : _GEN_3384; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3386 = 8'h42 == new_ptr_33_value ? ghv_66 : _GEN_3385; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3387 = 8'h43 == new_ptr_33_value ? ghv_67 : _GEN_3386; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3388 = 8'h44 == new_ptr_33_value ? ghv_68 : _GEN_3387; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3389 = 8'h45 == new_ptr_33_value ? ghv_69 : _GEN_3388; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3390 = 8'h46 == new_ptr_33_value ? ghv_70 : _GEN_3389; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3391 = 8'h47 == new_ptr_33_value ? ghv_71 : _GEN_3390; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3392 = 8'h48 == new_ptr_33_value ? ghv_72 : _GEN_3391; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3393 = 8'h49 == new_ptr_33_value ? ghv_73 : _GEN_3392; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3394 = 8'h4a == new_ptr_33_value ? ghv_74 : _GEN_3393; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3395 = 8'h4b == new_ptr_33_value ? ghv_75 : _GEN_3394; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3396 = 8'h4c == new_ptr_33_value ? ghv_76 : _GEN_3395; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3397 = 8'h4d == new_ptr_33_value ? ghv_77 : _GEN_3396; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3398 = 8'h4e == new_ptr_33_value ? ghv_78 : _GEN_3397; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3399 = 8'h4f == new_ptr_33_value ? ghv_79 : _GEN_3398; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3400 = 8'h50 == new_ptr_33_value ? ghv_80 : _GEN_3399; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3401 = 8'h51 == new_ptr_33_value ? ghv_81 : _GEN_3400; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3402 = 8'h52 == new_ptr_33_value ? ghv_82 : _GEN_3401; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3403 = 8'h53 == new_ptr_33_value ? ghv_83 : _GEN_3402; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3404 = 8'h54 == new_ptr_33_value ? ghv_84 : _GEN_3403; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3405 = 8'h55 == new_ptr_33_value ? ghv_85 : _GEN_3404; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3406 = 8'h56 == new_ptr_33_value ? ghv_86 : _GEN_3405; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3407 = 8'h57 == new_ptr_33_value ? ghv_87 : _GEN_3406; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3408 = 8'h58 == new_ptr_33_value ? ghv_88 : _GEN_3407; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3409 = 8'h59 == new_ptr_33_value ? ghv_89 : _GEN_3408; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3410 = 8'h5a == new_ptr_33_value ? ghv_90 : _GEN_3409; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3411 = 8'h5b == new_ptr_33_value ? ghv_91 : _GEN_3410; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3412 = 8'h5c == new_ptr_33_value ? ghv_92 : _GEN_3411; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3413 = 8'h5d == new_ptr_33_value ? ghv_93 : _GEN_3412; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3414 = 8'h5e == new_ptr_33_value ? ghv_94 : _GEN_3413; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3415 = 8'h5f == new_ptr_33_value ? ghv_95 : _GEN_3414; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3416 = 8'h60 == new_ptr_33_value ? ghv_96 : _GEN_3415; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3417 = 8'h61 == new_ptr_33_value ? ghv_97 : _GEN_3416; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3418 = 8'h62 == new_ptr_33_value ? ghv_98 : _GEN_3417; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3419 = 8'h63 == new_ptr_33_value ? ghv_99 : _GEN_3418; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3420 = 8'h64 == new_ptr_33_value ? ghv_100 : _GEN_3419; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3421 = 8'h65 == new_ptr_33_value ? ghv_101 : _GEN_3420; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3422 = 8'h66 == new_ptr_33_value ? ghv_102 : _GEN_3421; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3423 = 8'h67 == new_ptr_33_value ? ghv_103 : _GEN_3422; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3424 = 8'h68 == new_ptr_33_value ? ghv_104 : _GEN_3423; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3425 = 8'h69 == new_ptr_33_value ? ghv_105 : _GEN_3424; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3426 = 8'h6a == new_ptr_33_value ? ghv_106 : _GEN_3425; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3427 = 8'h6b == new_ptr_33_value ? ghv_107 : _GEN_3426; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3428 = 8'h6c == new_ptr_33_value ? ghv_108 : _GEN_3427; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3429 = 8'h6d == new_ptr_33_value ? ghv_109 : _GEN_3428; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3430 = 8'h6e == new_ptr_33_value ? ghv_110 : _GEN_3429; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3431 = 8'h6f == new_ptr_33_value ? ghv_111 : _GEN_3430; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3432 = 8'h70 == new_ptr_33_value ? ghv_112 : _GEN_3431; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3433 = 8'h71 == new_ptr_33_value ? ghv_113 : _GEN_3432; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3434 = 8'h72 == new_ptr_33_value ? ghv_114 : _GEN_3433; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3435 = 8'h73 == new_ptr_33_value ? ghv_115 : _GEN_3434; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3436 = 8'h74 == new_ptr_33_value ? ghv_116 : _GEN_3435; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3437 = 8'h75 == new_ptr_33_value ? ghv_117 : _GEN_3436; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3438 = 8'h76 == new_ptr_33_value ? ghv_118 : _GEN_3437; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3439 = 8'h77 == new_ptr_33_value ? ghv_119 : _GEN_3438; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3440 = 8'h78 == new_ptr_33_value ? ghv_120 : _GEN_3439; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3441 = 8'h79 == new_ptr_33_value ? ghv_121 : _GEN_3440; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3442 = 8'h7a == new_ptr_33_value ? ghv_122 : _GEN_3441; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3443 = 8'h7b == new_ptr_33_value ? ghv_123 : _GEN_3442; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3444 = 8'h7c == new_ptr_33_value ? ghv_124 : _GEN_3443; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3445 = 8'h7d == new_ptr_33_value ? ghv_125 : _GEN_3444; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3446 = 8'h7e == new_ptr_33_value ? ghv_126 : _GEN_3445; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3447 = 8'h7f == new_ptr_33_value ? ghv_127 : _GEN_3446; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3448 = 8'h80 == new_ptr_33_value ? ghv_128 : _GEN_3447; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3449 = 8'h81 == new_ptr_33_value ? ghv_129 : _GEN_3448; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3450 = 8'h82 == new_ptr_33_value ? ghv_130 : _GEN_3449; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3451 = 8'h83 == new_ptr_33_value ? ghv_131 : _GEN_3450; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3452 = 8'h84 == new_ptr_33_value ? ghv_132 : _GEN_3451; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3453 = 8'h85 == new_ptr_33_value ? ghv_133 : _GEN_3452; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3454 = 8'h86 == new_ptr_33_value ? ghv_134 : _GEN_3453; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3455 = 8'h87 == new_ptr_33_value ? ghv_135 : _GEN_3454; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3456 = 8'h88 == new_ptr_33_value ? ghv_136 : _GEN_3455; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3457 = 8'h89 == new_ptr_33_value ? ghv_137 : _GEN_3456; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3458 = 8'h8a == new_ptr_33_value ? ghv_138 : _GEN_3457; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3459 = 8'h8b == new_ptr_33_value ? ghv_139 : _GEN_3458; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3460 = 8'h8c == new_ptr_33_value ? ghv_140 : _GEN_3459; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3461 = 8'h8d == new_ptr_33_value ? ghv_141 : _GEN_3460; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3462 = 8'h8e == new_ptr_33_value ? ghv_142 : _GEN_3461; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_26_value = _new_ptr_value_T_53[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_3465 = 8'h1 == new_ptr_26_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3466 = 8'h2 == new_ptr_26_value ? ghv_2 : _GEN_3465; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3467 = 8'h3 == new_ptr_26_value ? ghv_3 : _GEN_3466; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3468 = 8'h4 == new_ptr_26_value ? ghv_4 : _GEN_3467; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3469 = 8'h5 == new_ptr_26_value ? ghv_5 : _GEN_3468; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3470 = 8'h6 == new_ptr_26_value ? ghv_6 : _GEN_3469; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3471 = 8'h7 == new_ptr_26_value ? ghv_7 : _GEN_3470; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3472 = 8'h8 == new_ptr_26_value ? ghv_8 : _GEN_3471; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3473 = 8'h9 == new_ptr_26_value ? ghv_9 : _GEN_3472; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3474 = 8'ha == new_ptr_26_value ? ghv_10 : _GEN_3473; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3475 = 8'hb == new_ptr_26_value ? ghv_11 : _GEN_3474; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3476 = 8'hc == new_ptr_26_value ? ghv_12 : _GEN_3475; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3477 = 8'hd == new_ptr_26_value ? ghv_13 : _GEN_3476; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3478 = 8'he == new_ptr_26_value ? ghv_14 : _GEN_3477; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3479 = 8'hf == new_ptr_26_value ? ghv_15 : _GEN_3478; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3480 = 8'h10 == new_ptr_26_value ? ghv_16 : _GEN_3479; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3481 = 8'h11 == new_ptr_26_value ? ghv_17 : _GEN_3480; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3482 = 8'h12 == new_ptr_26_value ? ghv_18 : _GEN_3481; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3483 = 8'h13 == new_ptr_26_value ? ghv_19 : _GEN_3482; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3484 = 8'h14 == new_ptr_26_value ? ghv_20 : _GEN_3483; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3485 = 8'h15 == new_ptr_26_value ? ghv_21 : _GEN_3484; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3486 = 8'h16 == new_ptr_26_value ? ghv_22 : _GEN_3485; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3487 = 8'h17 == new_ptr_26_value ? ghv_23 : _GEN_3486; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3488 = 8'h18 == new_ptr_26_value ? ghv_24 : _GEN_3487; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3489 = 8'h19 == new_ptr_26_value ? ghv_25 : _GEN_3488; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3490 = 8'h1a == new_ptr_26_value ? ghv_26 : _GEN_3489; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3491 = 8'h1b == new_ptr_26_value ? ghv_27 : _GEN_3490; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3492 = 8'h1c == new_ptr_26_value ? ghv_28 : _GEN_3491; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3493 = 8'h1d == new_ptr_26_value ? ghv_29 : _GEN_3492; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3494 = 8'h1e == new_ptr_26_value ? ghv_30 : _GEN_3493; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3495 = 8'h1f == new_ptr_26_value ? ghv_31 : _GEN_3494; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3496 = 8'h20 == new_ptr_26_value ? ghv_32 : _GEN_3495; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3497 = 8'h21 == new_ptr_26_value ? ghv_33 : _GEN_3496; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3498 = 8'h22 == new_ptr_26_value ? ghv_34 : _GEN_3497; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3499 = 8'h23 == new_ptr_26_value ? ghv_35 : _GEN_3498; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3500 = 8'h24 == new_ptr_26_value ? ghv_36 : _GEN_3499; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3501 = 8'h25 == new_ptr_26_value ? ghv_37 : _GEN_3500; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3502 = 8'h26 == new_ptr_26_value ? ghv_38 : _GEN_3501; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3503 = 8'h27 == new_ptr_26_value ? ghv_39 : _GEN_3502; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3504 = 8'h28 == new_ptr_26_value ? ghv_40 : _GEN_3503; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3505 = 8'h29 == new_ptr_26_value ? ghv_41 : _GEN_3504; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3506 = 8'h2a == new_ptr_26_value ? ghv_42 : _GEN_3505; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3507 = 8'h2b == new_ptr_26_value ? ghv_43 : _GEN_3506; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3508 = 8'h2c == new_ptr_26_value ? ghv_44 : _GEN_3507; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3509 = 8'h2d == new_ptr_26_value ? ghv_45 : _GEN_3508; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3510 = 8'h2e == new_ptr_26_value ? ghv_46 : _GEN_3509; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3511 = 8'h2f == new_ptr_26_value ? ghv_47 : _GEN_3510; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3512 = 8'h30 == new_ptr_26_value ? ghv_48 : _GEN_3511; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3513 = 8'h31 == new_ptr_26_value ? ghv_49 : _GEN_3512; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3514 = 8'h32 == new_ptr_26_value ? ghv_50 : _GEN_3513; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3515 = 8'h33 == new_ptr_26_value ? ghv_51 : _GEN_3514; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3516 = 8'h34 == new_ptr_26_value ? ghv_52 : _GEN_3515; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3517 = 8'h35 == new_ptr_26_value ? ghv_53 : _GEN_3516; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3518 = 8'h36 == new_ptr_26_value ? ghv_54 : _GEN_3517; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3519 = 8'h37 == new_ptr_26_value ? ghv_55 : _GEN_3518; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3520 = 8'h38 == new_ptr_26_value ? ghv_56 : _GEN_3519; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3521 = 8'h39 == new_ptr_26_value ? ghv_57 : _GEN_3520; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3522 = 8'h3a == new_ptr_26_value ? ghv_58 : _GEN_3521; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3523 = 8'h3b == new_ptr_26_value ? ghv_59 : _GEN_3522; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3524 = 8'h3c == new_ptr_26_value ? ghv_60 : _GEN_3523; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3525 = 8'h3d == new_ptr_26_value ? ghv_61 : _GEN_3524; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3526 = 8'h3e == new_ptr_26_value ? ghv_62 : _GEN_3525; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3527 = 8'h3f == new_ptr_26_value ? ghv_63 : _GEN_3526; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3528 = 8'h40 == new_ptr_26_value ? ghv_64 : _GEN_3527; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3529 = 8'h41 == new_ptr_26_value ? ghv_65 : _GEN_3528; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3530 = 8'h42 == new_ptr_26_value ? ghv_66 : _GEN_3529; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3531 = 8'h43 == new_ptr_26_value ? ghv_67 : _GEN_3530; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3532 = 8'h44 == new_ptr_26_value ? ghv_68 : _GEN_3531; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3533 = 8'h45 == new_ptr_26_value ? ghv_69 : _GEN_3532; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3534 = 8'h46 == new_ptr_26_value ? ghv_70 : _GEN_3533; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3535 = 8'h47 == new_ptr_26_value ? ghv_71 : _GEN_3534; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3536 = 8'h48 == new_ptr_26_value ? ghv_72 : _GEN_3535; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3537 = 8'h49 == new_ptr_26_value ? ghv_73 : _GEN_3536; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3538 = 8'h4a == new_ptr_26_value ? ghv_74 : _GEN_3537; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3539 = 8'h4b == new_ptr_26_value ? ghv_75 : _GEN_3538; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3540 = 8'h4c == new_ptr_26_value ? ghv_76 : _GEN_3539; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3541 = 8'h4d == new_ptr_26_value ? ghv_77 : _GEN_3540; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3542 = 8'h4e == new_ptr_26_value ? ghv_78 : _GEN_3541; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3543 = 8'h4f == new_ptr_26_value ? ghv_79 : _GEN_3542; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3544 = 8'h50 == new_ptr_26_value ? ghv_80 : _GEN_3543; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3545 = 8'h51 == new_ptr_26_value ? ghv_81 : _GEN_3544; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3546 = 8'h52 == new_ptr_26_value ? ghv_82 : _GEN_3545; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3547 = 8'h53 == new_ptr_26_value ? ghv_83 : _GEN_3546; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3548 = 8'h54 == new_ptr_26_value ? ghv_84 : _GEN_3547; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3549 = 8'h55 == new_ptr_26_value ? ghv_85 : _GEN_3548; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3550 = 8'h56 == new_ptr_26_value ? ghv_86 : _GEN_3549; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3551 = 8'h57 == new_ptr_26_value ? ghv_87 : _GEN_3550; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3552 = 8'h58 == new_ptr_26_value ? ghv_88 : _GEN_3551; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3553 = 8'h59 == new_ptr_26_value ? ghv_89 : _GEN_3552; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3554 = 8'h5a == new_ptr_26_value ? ghv_90 : _GEN_3553; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3555 = 8'h5b == new_ptr_26_value ? ghv_91 : _GEN_3554; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3556 = 8'h5c == new_ptr_26_value ? ghv_92 : _GEN_3555; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3557 = 8'h5d == new_ptr_26_value ? ghv_93 : _GEN_3556; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3558 = 8'h5e == new_ptr_26_value ? ghv_94 : _GEN_3557; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3559 = 8'h5f == new_ptr_26_value ? ghv_95 : _GEN_3558; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3560 = 8'h60 == new_ptr_26_value ? ghv_96 : _GEN_3559; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3561 = 8'h61 == new_ptr_26_value ? ghv_97 : _GEN_3560; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3562 = 8'h62 == new_ptr_26_value ? ghv_98 : _GEN_3561; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3563 = 8'h63 == new_ptr_26_value ? ghv_99 : _GEN_3562; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3564 = 8'h64 == new_ptr_26_value ? ghv_100 : _GEN_3563; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3565 = 8'h65 == new_ptr_26_value ? ghv_101 : _GEN_3564; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3566 = 8'h66 == new_ptr_26_value ? ghv_102 : _GEN_3565; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3567 = 8'h67 == new_ptr_26_value ? ghv_103 : _GEN_3566; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3568 = 8'h68 == new_ptr_26_value ? ghv_104 : _GEN_3567; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3569 = 8'h69 == new_ptr_26_value ? ghv_105 : _GEN_3568; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3570 = 8'h6a == new_ptr_26_value ? ghv_106 : _GEN_3569; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3571 = 8'h6b == new_ptr_26_value ? ghv_107 : _GEN_3570; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3572 = 8'h6c == new_ptr_26_value ? ghv_108 : _GEN_3571; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3573 = 8'h6d == new_ptr_26_value ? ghv_109 : _GEN_3572; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3574 = 8'h6e == new_ptr_26_value ? ghv_110 : _GEN_3573; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3575 = 8'h6f == new_ptr_26_value ? ghv_111 : _GEN_3574; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3576 = 8'h70 == new_ptr_26_value ? ghv_112 : _GEN_3575; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3577 = 8'h71 == new_ptr_26_value ? ghv_113 : _GEN_3576; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3578 = 8'h72 == new_ptr_26_value ? ghv_114 : _GEN_3577; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3579 = 8'h73 == new_ptr_26_value ? ghv_115 : _GEN_3578; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3580 = 8'h74 == new_ptr_26_value ? ghv_116 : _GEN_3579; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3581 = 8'h75 == new_ptr_26_value ? ghv_117 : _GEN_3580; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3582 = 8'h76 == new_ptr_26_value ? ghv_118 : _GEN_3581; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3583 = 8'h77 == new_ptr_26_value ? ghv_119 : _GEN_3582; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3584 = 8'h78 == new_ptr_26_value ? ghv_120 : _GEN_3583; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3585 = 8'h79 == new_ptr_26_value ? ghv_121 : _GEN_3584; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3586 = 8'h7a == new_ptr_26_value ? ghv_122 : _GEN_3585; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3587 = 8'h7b == new_ptr_26_value ? ghv_123 : _GEN_3586; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3588 = 8'h7c == new_ptr_26_value ? ghv_124 : _GEN_3587; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3589 = 8'h7d == new_ptr_26_value ? ghv_125 : _GEN_3588; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3590 = 8'h7e == new_ptr_26_value ? ghv_126 : _GEN_3589; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3591 = 8'h7f == new_ptr_26_value ? ghv_127 : _GEN_3590; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3592 = 8'h80 == new_ptr_26_value ? ghv_128 : _GEN_3591; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3593 = 8'h81 == new_ptr_26_value ? ghv_129 : _GEN_3592; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3594 = 8'h82 == new_ptr_26_value ? ghv_130 : _GEN_3593; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3595 = 8'h83 == new_ptr_26_value ? ghv_131 : _GEN_3594; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3596 = 8'h84 == new_ptr_26_value ? ghv_132 : _GEN_3595; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3597 = 8'h85 == new_ptr_26_value ? ghv_133 : _GEN_3596; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3598 = 8'h86 == new_ptr_26_value ? ghv_134 : _GEN_3597; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3599 = 8'h87 == new_ptr_26_value ? ghv_135 : _GEN_3598; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3600 = 8'h88 == new_ptr_26_value ? ghv_136 : _GEN_3599; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3601 = 8'h89 == new_ptr_26_value ? ghv_137 : _GEN_3600; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3602 = 8'h8a == new_ptr_26_value ? ghv_138 : _GEN_3601; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3603 = 8'h8b == new_ptr_26_value ? ghv_139 : _GEN_3602; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3604 = 8'h8c == new_ptr_26_value ? ghv_140 : _GEN_3603; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3605 = 8'h8d == new_ptr_26_value ? ghv_141 : _GEN_3604; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3606 = 8'h8e == new_ptr_26_value ? ghv_142 : _GEN_3605; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_32_value = _new_ptr_value_T_65[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_3609 = 8'h1 == new_ptr_32_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3610 = 8'h2 == new_ptr_32_value ? ghv_2 : _GEN_3609; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3611 = 8'h3 == new_ptr_32_value ? ghv_3 : _GEN_3610; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3612 = 8'h4 == new_ptr_32_value ? ghv_4 : _GEN_3611; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3613 = 8'h5 == new_ptr_32_value ? ghv_5 : _GEN_3612; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3614 = 8'h6 == new_ptr_32_value ? ghv_6 : _GEN_3613; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3615 = 8'h7 == new_ptr_32_value ? ghv_7 : _GEN_3614; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3616 = 8'h8 == new_ptr_32_value ? ghv_8 : _GEN_3615; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3617 = 8'h9 == new_ptr_32_value ? ghv_9 : _GEN_3616; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3618 = 8'ha == new_ptr_32_value ? ghv_10 : _GEN_3617; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3619 = 8'hb == new_ptr_32_value ? ghv_11 : _GEN_3618; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3620 = 8'hc == new_ptr_32_value ? ghv_12 : _GEN_3619; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3621 = 8'hd == new_ptr_32_value ? ghv_13 : _GEN_3620; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3622 = 8'he == new_ptr_32_value ? ghv_14 : _GEN_3621; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3623 = 8'hf == new_ptr_32_value ? ghv_15 : _GEN_3622; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3624 = 8'h10 == new_ptr_32_value ? ghv_16 : _GEN_3623; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3625 = 8'h11 == new_ptr_32_value ? ghv_17 : _GEN_3624; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3626 = 8'h12 == new_ptr_32_value ? ghv_18 : _GEN_3625; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3627 = 8'h13 == new_ptr_32_value ? ghv_19 : _GEN_3626; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3628 = 8'h14 == new_ptr_32_value ? ghv_20 : _GEN_3627; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3629 = 8'h15 == new_ptr_32_value ? ghv_21 : _GEN_3628; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3630 = 8'h16 == new_ptr_32_value ? ghv_22 : _GEN_3629; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3631 = 8'h17 == new_ptr_32_value ? ghv_23 : _GEN_3630; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3632 = 8'h18 == new_ptr_32_value ? ghv_24 : _GEN_3631; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3633 = 8'h19 == new_ptr_32_value ? ghv_25 : _GEN_3632; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3634 = 8'h1a == new_ptr_32_value ? ghv_26 : _GEN_3633; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3635 = 8'h1b == new_ptr_32_value ? ghv_27 : _GEN_3634; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3636 = 8'h1c == new_ptr_32_value ? ghv_28 : _GEN_3635; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3637 = 8'h1d == new_ptr_32_value ? ghv_29 : _GEN_3636; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3638 = 8'h1e == new_ptr_32_value ? ghv_30 : _GEN_3637; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3639 = 8'h1f == new_ptr_32_value ? ghv_31 : _GEN_3638; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3640 = 8'h20 == new_ptr_32_value ? ghv_32 : _GEN_3639; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3641 = 8'h21 == new_ptr_32_value ? ghv_33 : _GEN_3640; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3642 = 8'h22 == new_ptr_32_value ? ghv_34 : _GEN_3641; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3643 = 8'h23 == new_ptr_32_value ? ghv_35 : _GEN_3642; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3644 = 8'h24 == new_ptr_32_value ? ghv_36 : _GEN_3643; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3645 = 8'h25 == new_ptr_32_value ? ghv_37 : _GEN_3644; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3646 = 8'h26 == new_ptr_32_value ? ghv_38 : _GEN_3645; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3647 = 8'h27 == new_ptr_32_value ? ghv_39 : _GEN_3646; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3648 = 8'h28 == new_ptr_32_value ? ghv_40 : _GEN_3647; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3649 = 8'h29 == new_ptr_32_value ? ghv_41 : _GEN_3648; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3650 = 8'h2a == new_ptr_32_value ? ghv_42 : _GEN_3649; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3651 = 8'h2b == new_ptr_32_value ? ghv_43 : _GEN_3650; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3652 = 8'h2c == new_ptr_32_value ? ghv_44 : _GEN_3651; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3653 = 8'h2d == new_ptr_32_value ? ghv_45 : _GEN_3652; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3654 = 8'h2e == new_ptr_32_value ? ghv_46 : _GEN_3653; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3655 = 8'h2f == new_ptr_32_value ? ghv_47 : _GEN_3654; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3656 = 8'h30 == new_ptr_32_value ? ghv_48 : _GEN_3655; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3657 = 8'h31 == new_ptr_32_value ? ghv_49 : _GEN_3656; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3658 = 8'h32 == new_ptr_32_value ? ghv_50 : _GEN_3657; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3659 = 8'h33 == new_ptr_32_value ? ghv_51 : _GEN_3658; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3660 = 8'h34 == new_ptr_32_value ? ghv_52 : _GEN_3659; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3661 = 8'h35 == new_ptr_32_value ? ghv_53 : _GEN_3660; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3662 = 8'h36 == new_ptr_32_value ? ghv_54 : _GEN_3661; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3663 = 8'h37 == new_ptr_32_value ? ghv_55 : _GEN_3662; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3664 = 8'h38 == new_ptr_32_value ? ghv_56 : _GEN_3663; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3665 = 8'h39 == new_ptr_32_value ? ghv_57 : _GEN_3664; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3666 = 8'h3a == new_ptr_32_value ? ghv_58 : _GEN_3665; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3667 = 8'h3b == new_ptr_32_value ? ghv_59 : _GEN_3666; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3668 = 8'h3c == new_ptr_32_value ? ghv_60 : _GEN_3667; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3669 = 8'h3d == new_ptr_32_value ? ghv_61 : _GEN_3668; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3670 = 8'h3e == new_ptr_32_value ? ghv_62 : _GEN_3669; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3671 = 8'h3f == new_ptr_32_value ? ghv_63 : _GEN_3670; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3672 = 8'h40 == new_ptr_32_value ? ghv_64 : _GEN_3671; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3673 = 8'h41 == new_ptr_32_value ? ghv_65 : _GEN_3672; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3674 = 8'h42 == new_ptr_32_value ? ghv_66 : _GEN_3673; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3675 = 8'h43 == new_ptr_32_value ? ghv_67 : _GEN_3674; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3676 = 8'h44 == new_ptr_32_value ? ghv_68 : _GEN_3675; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3677 = 8'h45 == new_ptr_32_value ? ghv_69 : _GEN_3676; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3678 = 8'h46 == new_ptr_32_value ? ghv_70 : _GEN_3677; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3679 = 8'h47 == new_ptr_32_value ? ghv_71 : _GEN_3678; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3680 = 8'h48 == new_ptr_32_value ? ghv_72 : _GEN_3679; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3681 = 8'h49 == new_ptr_32_value ? ghv_73 : _GEN_3680; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3682 = 8'h4a == new_ptr_32_value ? ghv_74 : _GEN_3681; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3683 = 8'h4b == new_ptr_32_value ? ghv_75 : _GEN_3682; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3684 = 8'h4c == new_ptr_32_value ? ghv_76 : _GEN_3683; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3685 = 8'h4d == new_ptr_32_value ? ghv_77 : _GEN_3684; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3686 = 8'h4e == new_ptr_32_value ? ghv_78 : _GEN_3685; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3687 = 8'h4f == new_ptr_32_value ? ghv_79 : _GEN_3686; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3688 = 8'h50 == new_ptr_32_value ? ghv_80 : _GEN_3687; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3689 = 8'h51 == new_ptr_32_value ? ghv_81 : _GEN_3688; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3690 = 8'h52 == new_ptr_32_value ? ghv_82 : _GEN_3689; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3691 = 8'h53 == new_ptr_32_value ? ghv_83 : _GEN_3690; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3692 = 8'h54 == new_ptr_32_value ? ghv_84 : _GEN_3691; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3693 = 8'h55 == new_ptr_32_value ? ghv_85 : _GEN_3692; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3694 = 8'h56 == new_ptr_32_value ? ghv_86 : _GEN_3693; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3695 = 8'h57 == new_ptr_32_value ? ghv_87 : _GEN_3694; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3696 = 8'h58 == new_ptr_32_value ? ghv_88 : _GEN_3695; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3697 = 8'h59 == new_ptr_32_value ? ghv_89 : _GEN_3696; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3698 = 8'h5a == new_ptr_32_value ? ghv_90 : _GEN_3697; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3699 = 8'h5b == new_ptr_32_value ? ghv_91 : _GEN_3698; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3700 = 8'h5c == new_ptr_32_value ? ghv_92 : _GEN_3699; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3701 = 8'h5d == new_ptr_32_value ? ghv_93 : _GEN_3700; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3702 = 8'h5e == new_ptr_32_value ? ghv_94 : _GEN_3701; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3703 = 8'h5f == new_ptr_32_value ? ghv_95 : _GEN_3702; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3704 = 8'h60 == new_ptr_32_value ? ghv_96 : _GEN_3703; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3705 = 8'h61 == new_ptr_32_value ? ghv_97 : _GEN_3704; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3706 = 8'h62 == new_ptr_32_value ? ghv_98 : _GEN_3705; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3707 = 8'h63 == new_ptr_32_value ? ghv_99 : _GEN_3706; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3708 = 8'h64 == new_ptr_32_value ? ghv_100 : _GEN_3707; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3709 = 8'h65 == new_ptr_32_value ? ghv_101 : _GEN_3708; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3710 = 8'h66 == new_ptr_32_value ? ghv_102 : _GEN_3709; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3711 = 8'h67 == new_ptr_32_value ? ghv_103 : _GEN_3710; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3712 = 8'h68 == new_ptr_32_value ? ghv_104 : _GEN_3711; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3713 = 8'h69 == new_ptr_32_value ? ghv_105 : _GEN_3712; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3714 = 8'h6a == new_ptr_32_value ? ghv_106 : _GEN_3713; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3715 = 8'h6b == new_ptr_32_value ? ghv_107 : _GEN_3714; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3716 = 8'h6c == new_ptr_32_value ? ghv_108 : _GEN_3715; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3717 = 8'h6d == new_ptr_32_value ? ghv_109 : _GEN_3716; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3718 = 8'h6e == new_ptr_32_value ? ghv_110 : _GEN_3717; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3719 = 8'h6f == new_ptr_32_value ? ghv_111 : _GEN_3718; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3720 = 8'h70 == new_ptr_32_value ? ghv_112 : _GEN_3719; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3721 = 8'h71 == new_ptr_32_value ? ghv_113 : _GEN_3720; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3722 = 8'h72 == new_ptr_32_value ? ghv_114 : _GEN_3721; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3723 = 8'h73 == new_ptr_32_value ? ghv_115 : _GEN_3722; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3724 = 8'h74 == new_ptr_32_value ? ghv_116 : _GEN_3723; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3725 = 8'h75 == new_ptr_32_value ? ghv_117 : _GEN_3724; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3726 = 8'h76 == new_ptr_32_value ? ghv_118 : _GEN_3725; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3727 = 8'h77 == new_ptr_32_value ? ghv_119 : _GEN_3726; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3728 = 8'h78 == new_ptr_32_value ? ghv_120 : _GEN_3727; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3729 = 8'h79 == new_ptr_32_value ? ghv_121 : _GEN_3728; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3730 = 8'h7a == new_ptr_32_value ? ghv_122 : _GEN_3729; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3731 = 8'h7b == new_ptr_32_value ? ghv_123 : _GEN_3730; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3732 = 8'h7c == new_ptr_32_value ? ghv_124 : _GEN_3731; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3733 = 8'h7d == new_ptr_32_value ? ghv_125 : _GEN_3732; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3734 = 8'h7e == new_ptr_32_value ? ghv_126 : _GEN_3733; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3735 = 8'h7f == new_ptr_32_value ? ghv_127 : _GEN_3734; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3736 = 8'h80 == new_ptr_32_value ? ghv_128 : _GEN_3735; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3737 = 8'h81 == new_ptr_32_value ? ghv_129 : _GEN_3736; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3738 = 8'h82 == new_ptr_32_value ? ghv_130 : _GEN_3737; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3739 = 8'h83 == new_ptr_32_value ? ghv_131 : _GEN_3738; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3740 = 8'h84 == new_ptr_32_value ? ghv_132 : _GEN_3739; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3741 = 8'h85 == new_ptr_32_value ? ghv_133 : _GEN_3740; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3742 = 8'h86 == new_ptr_32_value ? ghv_134 : _GEN_3741; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3743 = 8'h87 == new_ptr_32_value ? ghv_135 : _GEN_3742; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3744 = 8'h88 == new_ptr_32_value ? ghv_136 : _GEN_3743; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3745 = 8'h89 == new_ptr_32_value ? ghv_137 : _GEN_3744; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3746 = 8'h8a == new_ptr_32_value ? ghv_138 : _GEN_3745; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3747 = 8'h8b == new_ptr_32_value ? ghv_139 : _GEN_3746; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3748 = 8'h8c == new_ptr_32_value ? ghv_140 : _GEN_3747; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3749 = 8'h8d == new_ptr_32_value ? ghv_141 : _GEN_3748; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3750 = 8'h8e == new_ptr_32_value ? ghv_142 : _GEN_3749; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_35_value = _new_ptr_value_T_71[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_3753 = 8'h1 == new_ptr_35_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3754 = 8'h2 == new_ptr_35_value ? ghv_2 : _GEN_3753; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3755 = 8'h3 == new_ptr_35_value ? ghv_3 : _GEN_3754; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3756 = 8'h4 == new_ptr_35_value ? ghv_4 : _GEN_3755; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3757 = 8'h5 == new_ptr_35_value ? ghv_5 : _GEN_3756; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3758 = 8'h6 == new_ptr_35_value ? ghv_6 : _GEN_3757; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3759 = 8'h7 == new_ptr_35_value ? ghv_7 : _GEN_3758; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3760 = 8'h8 == new_ptr_35_value ? ghv_8 : _GEN_3759; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3761 = 8'h9 == new_ptr_35_value ? ghv_9 : _GEN_3760; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3762 = 8'ha == new_ptr_35_value ? ghv_10 : _GEN_3761; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3763 = 8'hb == new_ptr_35_value ? ghv_11 : _GEN_3762; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3764 = 8'hc == new_ptr_35_value ? ghv_12 : _GEN_3763; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3765 = 8'hd == new_ptr_35_value ? ghv_13 : _GEN_3764; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3766 = 8'he == new_ptr_35_value ? ghv_14 : _GEN_3765; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3767 = 8'hf == new_ptr_35_value ? ghv_15 : _GEN_3766; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3768 = 8'h10 == new_ptr_35_value ? ghv_16 : _GEN_3767; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3769 = 8'h11 == new_ptr_35_value ? ghv_17 : _GEN_3768; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3770 = 8'h12 == new_ptr_35_value ? ghv_18 : _GEN_3769; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3771 = 8'h13 == new_ptr_35_value ? ghv_19 : _GEN_3770; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3772 = 8'h14 == new_ptr_35_value ? ghv_20 : _GEN_3771; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3773 = 8'h15 == new_ptr_35_value ? ghv_21 : _GEN_3772; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3774 = 8'h16 == new_ptr_35_value ? ghv_22 : _GEN_3773; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3775 = 8'h17 == new_ptr_35_value ? ghv_23 : _GEN_3774; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3776 = 8'h18 == new_ptr_35_value ? ghv_24 : _GEN_3775; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3777 = 8'h19 == new_ptr_35_value ? ghv_25 : _GEN_3776; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3778 = 8'h1a == new_ptr_35_value ? ghv_26 : _GEN_3777; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3779 = 8'h1b == new_ptr_35_value ? ghv_27 : _GEN_3778; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3780 = 8'h1c == new_ptr_35_value ? ghv_28 : _GEN_3779; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3781 = 8'h1d == new_ptr_35_value ? ghv_29 : _GEN_3780; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3782 = 8'h1e == new_ptr_35_value ? ghv_30 : _GEN_3781; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3783 = 8'h1f == new_ptr_35_value ? ghv_31 : _GEN_3782; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3784 = 8'h20 == new_ptr_35_value ? ghv_32 : _GEN_3783; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3785 = 8'h21 == new_ptr_35_value ? ghv_33 : _GEN_3784; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3786 = 8'h22 == new_ptr_35_value ? ghv_34 : _GEN_3785; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3787 = 8'h23 == new_ptr_35_value ? ghv_35 : _GEN_3786; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3788 = 8'h24 == new_ptr_35_value ? ghv_36 : _GEN_3787; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3789 = 8'h25 == new_ptr_35_value ? ghv_37 : _GEN_3788; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3790 = 8'h26 == new_ptr_35_value ? ghv_38 : _GEN_3789; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3791 = 8'h27 == new_ptr_35_value ? ghv_39 : _GEN_3790; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3792 = 8'h28 == new_ptr_35_value ? ghv_40 : _GEN_3791; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3793 = 8'h29 == new_ptr_35_value ? ghv_41 : _GEN_3792; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3794 = 8'h2a == new_ptr_35_value ? ghv_42 : _GEN_3793; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3795 = 8'h2b == new_ptr_35_value ? ghv_43 : _GEN_3794; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3796 = 8'h2c == new_ptr_35_value ? ghv_44 : _GEN_3795; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3797 = 8'h2d == new_ptr_35_value ? ghv_45 : _GEN_3796; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3798 = 8'h2e == new_ptr_35_value ? ghv_46 : _GEN_3797; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3799 = 8'h2f == new_ptr_35_value ? ghv_47 : _GEN_3798; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3800 = 8'h30 == new_ptr_35_value ? ghv_48 : _GEN_3799; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3801 = 8'h31 == new_ptr_35_value ? ghv_49 : _GEN_3800; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3802 = 8'h32 == new_ptr_35_value ? ghv_50 : _GEN_3801; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3803 = 8'h33 == new_ptr_35_value ? ghv_51 : _GEN_3802; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3804 = 8'h34 == new_ptr_35_value ? ghv_52 : _GEN_3803; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3805 = 8'h35 == new_ptr_35_value ? ghv_53 : _GEN_3804; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3806 = 8'h36 == new_ptr_35_value ? ghv_54 : _GEN_3805; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3807 = 8'h37 == new_ptr_35_value ? ghv_55 : _GEN_3806; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3808 = 8'h38 == new_ptr_35_value ? ghv_56 : _GEN_3807; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3809 = 8'h39 == new_ptr_35_value ? ghv_57 : _GEN_3808; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3810 = 8'h3a == new_ptr_35_value ? ghv_58 : _GEN_3809; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3811 = 8'h3b == new_ptr_35_value ? ghv_59 : _GEN_3810; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3812 = 8'h3c == new_ptr_35_value ? ghv_60 : _GEN_3811; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3813 = 8'h3d == new_ptr_35_value ? ghv_61 : _GEN_3812; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3814 = 8'h3e == new_ptr_35_value ? ghv_62 : _GEN_3813; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3815 = 8'h3f == new_ptr_35_value ? ghv_63 : _GEN_3814; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3816 = 8'h40 == new_ptr_35_value ? ghv_64 : _GEN_3815; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3817 = 8'h41 == new_ptr_35_value ? ghv_65 : _GEN_3816; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3818 = 8'h42 == new_ptr_35_value ? ghv_66 : _GEN_3817; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3819 = 8'h43 == new_ptr_35_value ? ghv_67 : _GEN_3818; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3820 = 8'h44 == new_ptr_35_value ? ghv_68 : _GEN_3819; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3821 = 8'h45 == new_ptr_35_value ? ghv_69 : _GEN_3820; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3822 = 8'h46 == new_ptr_35_value ? ghv_70 : _GEN_3821; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3823 = 8'h47 == new_ptr_35_value ? ghv_71 : _GEN_3822; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3824 = 8'h48 == new_ptr_35_value ? ghv_72 : _GEN_3823; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3825 = 8'h49 == new_ptr_35_value ? ghv_73 : _GEN_3824; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3826 = 8'h4a == new_ptr_35_value ? ghv_74 : _GEN_3825; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3827 = 8'h4b == new_ptr_35_value ? ghv_75 : _GEN_3826; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3828 = 8'h4c == new_ptr_35_value ? ghv_76 : _GEN_3827; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3829 = 8'h4d == new_ptr_35_value ? ghv_77 : _GEN_3828; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3830 = 8'h4e == new_ptr_35_value ? ghv_78 : _GEN_3829; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3831 = 8'h4f == new_ptr_35_value ? ghv_79 : _GEN_3830; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3832 = 8'h50 == new_ptr_35_value ? ghv_80 : _GEN_3831; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3833 = 8'h51 == new_ptr_35_value ? ghv_81 : _GEN_3832; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3834 = 8'h52 == new_ptr_35_value ? ghv_82 : _GEN_3833; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3835 = 8'h53 == new_ptr_35_value ? ghv_83 : _GEN_3834; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3836 = 8'h54 == new_ptr_35_value ? ghv_84 : _GEN_3835; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3837 = 8'h55 == new_ptr_35_value ? ghv_85 : _GEN_3836; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3838 = 8'h56 == new_ptr_35_value ? ghv_86 : _GEN_3837; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3839 = 8'h57 == new_ptr_35_value ? ghv_87 : _GEN_3838; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3840 = 8'h58 == new_ptr_35_value ? ghv_88 : _GEN_3839; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3841 = 8'h59 == new_ptr_35_value ? ghv_89 : _GEN_3840; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3842 = 8'h5a == new_ptr_35_value ? ghv_90 : _GEN_3841; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3843 = 8'h5b == new_ptr_35_value ? ghv_91 : _GEN_3842; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3844 = 8'h5c == new_ptr_35_value ? ghv_92 : _GEN_3843; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3845 = 8'h5d == new_ptr_35_value ? ghv_93 : _GEN_3844; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3846 = 8'h5e == new_ptr_35_value ? ghv_94 : _GEN_3845; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3847 = 8'h5f == new_ptr_35_value ? ghv_95 : _GEN_3846; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3848 = 8'h60 == new_ptr_35_value ? ghv_96 : _GEN_3847; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3849 = 8'h61 == new_ptr_35_value ? ghv_97 : _GEN_3848; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3850 = 8'h62 == new_ptr_35_value ? ghv_98 : _GEN_3849; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3851 = 8'h63 == new_ptr_35_value ? ghv_99 : _GEN_3850; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3852 = 8'h64 == new_ptr_35_value ? ghv_100 : _GEN_3851; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3853 = 8'h65 == new_ptr_35_value ? ghv_101 : _GEN_3852; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3854 = 8'h66 == new_ptr_35_value ? ghv_102 : _GEN_3853; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3855 = 8'h67 == new_ptr_35_value ? ghv_103 : _GEN_3854; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3856 = 8'h68 == new_ptr_35_value ? ghv_104 : _GEN_3855; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3857 = 8'h69 == new_ptr_35_value ? ghv_105 : _GEN_3856; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3858 = 8'h6a == new_ptr_35_value ? ghv_106 : _GEN_3857; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3859 = 8'h6b == new_ptr_35_value ? ghv_107 : _GEN_3858; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3860 = 8'h6c == new_ptr_35_value ? ghv_108 : _GEN_3859; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3861 = 8'h6d == new_ptr_35_value ? ghv_109 : _GEN_3860; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3862 = 8'h6e == new_ptr_35_value ? ghv_110 : _GEN_3861; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3863 = 8'h6f == new_ptr_35_value ? ghv_111 : _GEN_3862; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3864 = 8'h70 == new_ptr_35_value ? ghv_112 : _GEN_3863; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3865 = 8'h71 == new_ptr_35_value ? ghv_113 : _GEN_3864; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3866 = 8'h72 == new_ptr_35_value ? ghv_114 : _GEN_3865; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3867 = 8'h73 == new_ptr_35_value ? ghv_115 : _GEN_3866; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3868 = 8'h74 == new_ptr_35_value ? ghv_116 : _GEN_3867; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3869 = 8'h75 == new_ptr_35_value ? ghv_117 : _GEN_3868; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3870 = 8'h76 == new_ptr_35_value ? ghv_118 : _GEN_3869; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3871 = 8'h77 == new_ptr_35_value ? ghv_119 : _GEN_3870; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3872 = 8'h78 == new_ptr_35_value ? ghv_120 : _GEN_3871; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3873 = 8'h79 == new_ptr_35_value ? ghv_121 : _GEN_3872; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3874 = 8'h7a == new_ptr_35_value ? ghv_122 : _GEN_3873; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3875 = 8'h7b == new_ptr_35_value ? ghv_123 : _GEN_3874; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3876 = 8'h7c == new_ptr_35_value ? ghv_124 : _GEN_3875; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3877 = 8'h7d == new_ptr_35_value ? ghv_125 : _GEN_3876; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3878 = 8'h7e == new_ptr_35_value ? ghv_126 : _GEN_3877; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3879 = 8'h7f == new_ptr_35_value ? ghv_127 : _GEN_3878; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3880 = 8'h80 == new_ptr_35_value ? ghv_128 : _GEN_3879; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3881 = 8'h81 == new_ptr_35_value ? ghv_129 : _GEN_3880; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3882 = 8'h82 == new_ptr_35_value ? ghv_130 : _GEN_3881; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3883 = 8'h83 == new_ptr_35_value ? ghv_131 : _GEN_3882; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3884 = 8'h84 == new_ptr_35_value ? ghv_132 : _GEN_3883; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3885 = 8'h85 == new_ptr_35_value ? ghv_133 : _GEN_3884; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3886 = 8'h86 == new_ptr_35_value ? ghv_134 : _GEN_3885; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3887 = 8'h87 == new_ptr_35_value ? ghv_135 : _GEN_3886; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3888 = 8'h88 == new_ptr_35_value ? ghv_136 : _GEN_3887; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3889 = 8'h89 == new_ptr_35_value ? ghv_137 : _GEN_3888; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3890 = 8'h8a == new_ptr_35_value ? ghv_138 : _GEN_3889; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3891 = 8'h8b == new_ptr_35_value ? ghv_139 : _GEN_3890; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3892 = 8'h8c == new_ptr_35_value ? ghv_140 : _GEN_3891; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3893 = 8'h8d == new_ptr_35_value ? ghv_141 : _GEN_3892; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3894 = 8'h8e == new_ptr_35_value ? ghv_142 : _GEN_3893; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_22_value = _new_ptr_value_T_45[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_3897 = 8'h1 == new_ptr_22_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3898 = 8'h2 == new_ptr_22_value ? ghv_2 : _GEN_3897; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3899 = 8'h3 == new_ptr_22_value ? ghv_3 : _GEN_3898; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3900 = 8'h4 == new_ptr_22_value ? ghv_4 : _GEN_3899; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3901 = 8'h5 == new_ptr_22_value ? ghv_5 : _GEN_3900; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3902 = 8'h6 == new_ptr_22_value ? ghv_6 : _GEN_3901; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3903 = 8'h7 == new_ptr_22_value ? ghv_7 : _GEN_3902; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3904 = 8'h8 == new_ptr_22_value ? ghv_8 : _GEN_3903; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3905 = 8'h9 == new_ptr_22_value ? ghv_9 : _GEN_3904; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3906 = 8'ha == new_ptr_22_value ? ghv_10 : _GEN_3905; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3907 = 8'hb == new_ptr_22_value ? ghv_11 : _GEN_3906; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3908 = 8'hc == new_ptr_22_value ? ghv_12 : _GEN_3907; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3909 = 8'hd == new_ptr_22_value ? ghv_13 : _GEN_3908; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3910 = 8'he == new_ptr_22_value ? ghv_14 : _GEN_3909; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3911 = 8'hf == new_ptr_22_value ? ghv_15 : _GEN_3910; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3912 = 8'h10 == new_ptr_22_value ? ghv_16 : _GEN_3911; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3913 = 8'h11 == new_ptr_22_value ? ghv_17 : _GEN_3912; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3914 = 8'h12 == new_ptr_22_value ? ghv_18 : _GEN_3913; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3915 = 8'h13 == new_ptr_22_value ? ghv_19 : _GEN_3914; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3916 = 8'h14 == new_ptr_22_value ? ghv_20 : _GEN_3915; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3917 = 8'h15 == new_ptr_22_value ? ghv_21 : _GEN_3916; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3918 = 8'h16 == new_ptr_22_value ? ghv_22 : _GEN_3917; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3919 = 8'h17 == new_ptr_22_value ? ghv_23 : _GEN_3918; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3920 = 8'h18 == new_ptr_22_value ? ghv_24 : _GEN_3919; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3921 = 8'h19 == new_ptr_22_value ? ghv_25 : _GEN_3920; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3922 = 8'h1a == new_ptr_22_value ? ghv_26 : _GEN_3921; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3923 = 8'h1b == new_ptr_22_value ? ghv_27 : _GEN_3922; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3924 = 8'h1c == new_ptr_22_value ? ghv_28 : _GEN_3923; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3925 = 8'h1d == new_ptr_22_value ? ghv_29 : _GEN_3924; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3926 = 8'h1e == new_ptr_22_value ? ghv_30 : _GEN_3925; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3927 = 8'h1f == new_ptr_22_value ? ghv_31 : _GEN_3926; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3928 = 8'h20 == new_ptr_22_value ? ghv_32 : _GEN_3927; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3929 = 8'h21 == new_ptr_22_value ? ghv_33 : _GEN_3928; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3930 = 8'h22 == new_ptr_22_value ? ghv_34 : _GEN_3929; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3931 = 8'h23 == new_ptr_22_value ? ghv_35 : _GEN_3930; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3932 = 8'h24 == new_ptr_22_value ? ghv_36 : _GEN_3931; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3933 = 8'h25 == new_ptr_22_value ? ghv_37 : _GEN_3932; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3934 = 8'h26 == new_ptr_22_value ? ghv_38 : _GEN_3933; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3935 = 8'h27 == new_ptr_22_value ? ghv_39 : _GEN_3934; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3936 = 8'h28 == new_ptr_22_value ? ghv_40 : _GEN_3935; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3937 = 8'h29 == new_ptr_22_value ? ghv_41 : _GEN_3936; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3938 = 8'h2a == new_ptr_22_value ? ghv_42 : _GEN_3937; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3939 = 8'h2b == new_ptr_22_value ? ghv_43 : _GEN_3938; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3940 = 8'h2c == new_ptr_22_value ? ghv_44 : _GEN_3939; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3941 = 8'h2d == new_ptr_22_value ? ghv_45 : _GEN_3940; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3942 = 8'h2e == new_ptr_22_value ? ghv_46 : _GEN_3941; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3943 = 8'h2f == new_ptr_22_value ? ghv_47 : _GEN_3942; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3944 = 8'h30 == new_ptr_22_value ? ghv_48 : _GEN_3943; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3945 = 8'h31 == new_ptr_22_value ? ghv_49 : _GEN_3944; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3946 = 8'h32 == new_ptr_22_value ? ghv_50 : _GEN_3945; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3947 = 8'h33 == new_ptr_22_value ? ghv_51 : _GEN_3946; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3948 = 8'h34 == new_ptr_22_value ? ghv_52 : _GEN_3947; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3949 = 8'h35 == new_ptr_22_value ? ghv_53 : _GEN_3948; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3950 = 8'h36 == new_ptr_22_value ? ghv_54 : _GEN_3949; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3951 = 8'h37 == new_ptr_22_value ? ghv_55 : _GEN_3950; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3952 = 8'h38 == new_ptr_22_value ? ghv_56 : _GEN_3951; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3953 = 8'h39 == new_ptr_22_value ? ghv_57 : _GEN_3952; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3954 = 8'h3a == new_ptr_22_value ? ghv_58 : _GEN_3953; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3955 = 8'h3b == new_ptr_22_value ? ghv_59 : _GEN_3954; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3956 = 8'h3c == new_ptr_22_value ? ghv_60 : _GEN_3955; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3957 = 8'h3d == new_ptr_22_value ? ghv_61 : _GEN_3956; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3958 = 8'h3e == new_ptr_22_value ? ghv_62 : _GEN_3957; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3959 = 8'h3f == new_ptr_22_value ? ghv_63 : _GEN_3958; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3960 = 8'h40 == new_ptr_22_value ? ghv_64 : _GEN_3959; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3961 = 8'h41 == new_ptr_22_value ? ghv_65 : _GEN_3960; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3962 = 8'h42 == new_ptr_22_value ? ghv_66 : _GEN_3961; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3963 = 8'h43 == new_ptr_22_value ? ghv_67 : _GEN_3962; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3964 = 8'h44 == new_ptr_22_value ? ghv_68 : _GEN_3963; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3965 = 8'h45 == new_ptr_22_value ? ghv_69 : _GEN_3964; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3966 = 8'h46 == new_ptr_22_value ? ghv_70 : _GEN_3965; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3967 = 8'h47 == new_ptr_22_value ? ghv_71 : _GEN_3966; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3968 = 8'h48 == new_ptr_22_value ? ghv_72 : _GEN_3967; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3969 = 8'h49 == new_ptr_22_value ? ghv_73 : _GEN_3968; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3970 = 8'h4a == new_ptr_22_value ? ghv_74 : _GEN_3969; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3971 = 8'h4b == new_ptr_22_value ? ghv_75 : _GEN_3970; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3972 = 8'h4c == new_ptr_22_value ? ghv_76 : _GEN_3971; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3973 = 8'h4d == new_ptr_22_value ? ghv_77 : _GEN_3972; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3974 = 8'h4e == new_ptr_22_value ? ghv_78 : _GEN_3973; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3975 = 8'h4f == new_ptr_22_value ? ghv_79 : _GEN_3974; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3976 = 8'h50 == new_ptr_22_value ? ghv_80 : _GEN_3975; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3977 = 8'h51 == new_ptr_22_value ? ghv_81 : _GEN_3976; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3978 = 8'h52 == new_ptr_22_value ? ghv_82 : _GEN_3977; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3979 = 8'h53 == new_ptr_22_value ? ghv_83 : _GEN_3978; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3980 = 8'h54 == new_ptr_22_value ? ghv_84 : _GEN_3979; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3981 = 8'h55 == new_ptr_22_value ? ghv_85 : _GEN_3980; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3982 = 8'h56 == new_ptr_22_value ? ghv_86 : _GEN_3981; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3983 = 8'h57 == new_ptr_22_value ? ghv_87 : _GEN_3982; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3984 = 8'h58 == new_ptr_22_value ? ghv_88 : _GEN_3983; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3985 = 8'h59 == new_ptr_22_value ? ghv_89 : _GEN_3984; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3986 = 8'h5a == new_ptr_22_value ? ghv_90 : _GEN_3985; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3987 = 8'h5b == new_ptr_22_value ? ghv_91 : _GEN_3986; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3988 = 8'h5c == new_ptr_22_value ? ghv_92 : _GEN_3987; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3989 = 8'h5d == new_ptr_22_value ? ghv_93 : _GEN_3988; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3990 = 8'h5e == new_ptr_22_value ? ghv_94 : _GEN_3989; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3991 = 8'h5f == new_ptr_22_value ? ghv_95 : _GEN_3990; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3992 = 8'h60 == new_ptr_22_value ? ghv_96 : _GEN_3991; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3993 = 8'h61 == new_ptr_22_value ? ghv_97 : _GEN_3992; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3994 = 8'h62 == new_ptr_22_value ? ghv_98 : _GEN_3993; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3995 = 8'h63 == new_ptr_22_value ? ghv_99 : _GEN_3994; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3996 = 8'h64 == new_ptr_22_value ? ghv_100 : _GEN_3995; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3997 = 8'h65 == new_ptr_22_value ? ghv_101 : _GEN_3996; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3998 = 8'h66 == new_ptr_22_value ? ghv_102 : _GEN_3997; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_3999 = 8'h67 == new_ptr_22_value ? ghv_103 : _GEN_3998; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4000 = 8'h68 == new_ptr_22_value ? ghv_104 : _GEN_3999; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4001 = 8'h69 == new_ptr_22_value ? ghv_105 : _GEN_4000; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4002 = 8'h6a == new_ptr_22_value ? ghv_106 : _GEN_4001; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4003 = 8'h6b == new_ptr_22_value ? ghv_107 : _GEN_4002; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4004 = 8'h6c == new_ptr_22_value ? ghv_108 : _GEN_4003; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4005 = 8'h6d == new_ptr_22_value ? ghv_109 : _GEN_4004; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4006 = 8'h6e == new_ptr_22_value ? ghv_110 : _GEN_4005; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4007 = 8'h6f == new_ptr_22_value ? ghv_111 : _GEN_4006; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4008 = 8'h70 == new_ptr_22_value ? ghv_112 : _GEN_4007; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4009 = 8'h71 == new_ptr_22_value ? ghv_113 : _GEN_4008; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4010 = 8'h72 == new_ptr_22_value ? ghv_114 : _GEN_4009; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4011 = 8'h73 == new_ptr_22_value ? ghv_115 : _GEN_4010; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4012 = 8'h74 == new_ptr_22_value ? ghv_116 : _GEN_4011; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4013 = 8'h75 == new_ptr_22_value ? ghv_117 : _GEN_4012; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4014 = 8'h76 == new_ptr_22_value ? ghv_118 : _GEN_4013; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4015 = 8'h77 == new_ptr_22_value ? ghv_119 : _GEN_4014; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4016 = 8'h78 == new_ptr_22_value ? ghv_120 : _GEN_4015; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4017 = 8'h79 == new_ptr_22_value ? ghv_121 : _GEN_4016; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4018 = 8'h7a == new_ptr_22_value ? ghv_122 : _GEN_4017; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4019 = 8'h7b == new_ptr_22_value ? ghv_123 : _GEN_4018; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4020 = 8'h7c == new_ptr_22_value ? ghv_124 : _GEN_4019; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4021 = 8'h7d == new_ptr_22_value ? ghv_125 : _GEN_4020; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4022 = 8'h7e == new_ptr_22_value ? ghv_126 : _GEN_4021; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4023 = 8'h7f == new_ptr_22_value ? ghv_127 : _GEN_4022; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4024 = 8'h80 == new_ptr_22_value ? ghv_128 : _GEN_4023; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4025 = 8'h81 == new_ptr_22_value ? ghv_129 : _GEN_4024; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4026 = 8'h82 == new_ptr_22_value ? ghv_130 : _GEN_4025; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4027 = 8'h83 == new_ptr_22_value ? ghv_131 : _GEN_4026; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4028 = 8'h84 == new_ptr_22_value ? ghv_132 : _GEN_4027; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4029 = 8'h85 == new_ptr_22_value ? ghv_133 : _GEN_4028; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4030 = 8'h86 == new_ptr_22_value ? ghv_134 : _GEN_4029; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4031 = 8'h87 == new_ptr_22_value ? ghv_135 : _GEN_4030; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4032 = 8'h88 == new_ptr_22_value ? ghv_136 : _GEN_4031; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4033 = 8'h89 == new_ptr_22_value ? ghv_137 : _GEN_4032; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4034 = 8'h8a == new_ptr_22_value ? ghv_138 : _GEN_4033; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4035 = 8'h8b == new_ptr_22_value ? ghv_139 : _GEN_4034; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4036 = 8'h8c == new_ptr_22_value ? ghv_140 : _GEN_4035; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4037 = 8'h8d == new_ptr_22_value ? ghv_141 : _GEN_4036; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4038 = 8'h8e == new_ptr_22_value ? ghv_142 : _GEN_4037; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_34_value = _new_ptr_value_T_69[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_4041 = 8'h1 == new_ptr_34_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4042 = 8'h2 == new_ptr_34_value ? ghv_2 : _GEN_4041; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4043 = 8'h3 == new_ptr_34_value ? ghv_3 : _GEN_4042; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4044 = 8'h4 == new_ptr_34_value ? ghv_4 : _GEN_4043; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4045 = 8'h5 == new_ptr_34_value ? ghv_5 : _GEN_4044; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4046 = 8'h6 == new_ptr_34_value ? ghv_6 : _GEN_4045; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4047 = 8'h7 == new_ptr_34_value ? ghv_7 : _GEN_4046; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4048 = 8'h8 == new_ptr_34_value ? ghv_8 : _GEN_4047; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4049 = 8'h9 == new_ptr_34_value ? ghv_9 : _GEN_4048; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4050 = 8'ha == new_ptr_34_value ? ghv_10 : _GEN_4049; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4051 = 8'hb == new_ptr_34_value ? ghv_11 : _GEN_4050; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4052 = 8'hc == new_ptr_34_value ? ghv_12 : _GEN_4051; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4053 = 8'hd == new_ptr_34_value ? ghv_13 : _GEN_4052; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4054 = 8'he == new_ptr_34_value ? ghv_14 : _GEN_4053; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4055 = 8'hf == new_ptr_34_value ? ghv_15 : _GEN_4054; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4056 = 8'h10 == new_ptr_34_value ? ghv_16 : _GEN_4055; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4057 = 8'h11 == new_ptr_34_value ? ghv_17 : _GEN_4056; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4058 = 8'h12 == new_ptr_34_value ? ghv_18 : _GEN_4057; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4059 = 8'h13 == new_ptr_34_value ? ghv_19 : _GEN_4058; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4060 = 8'h14 == new_ptr_34_value ? ghv_20 : _GEN_4059; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4061 = 8'h15 == new_ptr_34_value ? ghv_21 : _GEN_4060; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4062 = 8'h16 == new_ptr_34_value ? ghv_22 : _GEN_4061; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4063 = 8'h17 == new_ptr_34_value ? ghv_23 : _GEN_4062; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4064 = 8'h18 == new_ptr_34_value ? ghv_24 : _GEN_4063; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4065 = 8'h19 == new_ptr_34_value ? ghv_25 : _GEN_4064; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4066 = 8'h1a == new_ptr_34_value ? ghv_26 : _GEN_4065; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4067 = 8'h1b == new_ptr_34_value ? ghv_27 : _GEN_4066; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4068 = 8'h1c == new_ptr_34_value ? ghv_28 : _GEN_4067; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4069 = 8'h1d == new_ptr_34_value ? ghv_29 : _GEN_4068; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4070 = 8'h1e == new_ptr_34_value ? ghv_30 : _GEN_4069; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4071 = 8'h1f == new_ptr_34_value ? ghv_31 : _GEN_4070; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4072 = 8'h20 == new_ptr_34_value ? ghv_32 : _GEN_4071; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4073 = 8'h21 == new_ptr_34_value ? ghv_33 : _GEN_4072; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4074 = 8'h22 == new_ptr_34_value ? ghv_34 : _GEN_4073; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4075 = 8'h23 == new_ptr_34_value ? ghv_35 : _GEN_4074; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4076 = 8'h24 == new_ptr_34_value ? ghv_36 : _GEN_4075; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4077 = 8'h25 == new_ptr_34_value ? ghv_37 : _GEN_4076; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4078 = 8'h26 == new_ptr_34_value ? ghv_38 : _GEN_4077; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4079 = 8'h27 == new_ptr_34_value ? ghv_39 : _GEN_4078; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4080 = 8'h28 == new_ptr_34_value ? ghv_40 : _GEN_4079; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4081 = 8'h29 == new_ptr_34_value ? ghv_41 : _GEN_4080; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4082 = 8'h2a == new_ptr_34_value ? ghv_42 : _GEN_4081; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4083 = 8'h2b == new_ptr_34_value ? ghv_43 : _GEN_4082; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4084 = 8'h2c == new_ptr_34_value ? ghv_44 : _GEN_4083; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4085 = 8'h2d == new_ptr_34_value ? ghv_45 : _GEN_4084; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4086 = 8'h2e == new_ptr_34_value ? ghv_46 : _GEN_4085; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4087 = 8'h2f == new_ptr_34_value ? ghv_47 : _GEN_4086; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4088 = 8'h30 == new_ptr_34_value ? ghv_48 : _GEN_4087; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4089 = 8'h31 == new_ptr_34_value ? ghv_49 : _GEN_4088; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4090 = 8'h32 == new_ptr_34_value ? ghv_50 : _GEN_4089; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4091 = 8'h33 == new_ptr_34_value ? ghv_51 : _GEN_4090; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4092 = 8'h34 == new_ptr_34_value ? ghv_52 : _GEN_4091; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4093 = 8'h35 == new_ptr_34_value ? ghv_53 : _GEN_4092; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4094 = 8'h36 == new_ptr_34_value ? ghv_54 : _GEN_4093; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4095 = 8'h37 == new_ptr_34_value ? ghv_55 : _GEN_4094; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4096 = 8'h38 == new_ptr_34_value ? ghv_56 : _GEN_4095; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4097 = 8'h39 == new_ptr_34_value ? ghv_57 : _GEN_4096; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4098 = 8'h3a == new_ptr_34_value ? ghv_58 : _GEN_4097; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4099 = 8'h3b == new_ptr_34_value ? ghv_59 : _GEN_4098; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4100 = 8'h3c == new_ptr_34_value ? ghv_60 : _GEN_4099; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4101 = 8'h3d == new_ptr_34_value ? ghv_61 : _GEN_4100; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4102 = 8'h3e == new_ptr_34_value ? ghv_62 : _GEN_4101; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4103 = 8'h3f == new_ptr_34_value ? ghv_63 : _GEN_4102; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4104 = 8'h40 == new_ptr_34_value ? ghv_64 : _GEN_4103; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4105 = 8'h41 == new_ptr_34_value ? ghv_65 : _GEN_4104; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4106 = 8'h42 == new_ptr_34_value ? ghv_66 : _GEN_4105; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4107 = 8'h43 == new_ptr_34_value ? ghv_67 : _GEN_4106; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4108 = 8'h44 == new_ptr_34_value ? ghv_68 : _GEN_4107; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4109 = 8'h45 == new_ptr_34_value ? ghv_69 : _GEN_4108; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4110 = 8'h46 == new_ptr_34_value ? ghv_70 : _GEN_4109; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4111 = 8'h47 == new_ptr_34_value ? ghv_71 : _GEN_4110; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4112 = 8'h48 == new_ptr_34_value ? ghv_72 : _GEN_4111; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4113 = 8'h49 == new_ptr_34_value ? ghv_73 : _GEN_4112; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4114 = 8'h4a == new_ptr_34_value ? ghv_74 : _GEN_4113; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4115 = 8'h4b == new_ptr_34_value ? ghv_75 : _GEN_4114; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4116 = 8'h4c == new_ptr_34_value ? ghv_76 : _GEN_4115; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4117 = 8'h4d == new_ptr_34_value ? ghv_77 : _GEN_4116; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4118 = 8'h4e == new_ptr_34_value ? ghv_78 : _GEN_4117; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4119 = 8'h4f == new_ptr_34_value ? ghv_79 : _GEN_4118; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4120 = 8'h50 == new_ptr_34_value ? ghv_80 : _GEN_4119; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4121 = 8'h51 == new_ptr_34_value ? ghv_81 : _GEN_4120; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4122 = 8'h52 == new_ptr_34_value ? ghv_82 : _GEN_4121; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4123 = 8'h53 == new_ptr_34_value ? ghv_83 : _GEN_4122; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4124 = 8'h54 == new_ptr_34_value ? ghv_84 : _GEN_4123; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4125 = 8'h55 == new_ptr_34_value ? ghv_85 : _GEN_4124; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4126 = 8'h56 == new_ptr_34_value ? ghv_86 : _GEN_4125; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4127 = 8'h57 == new_ptr_34_value ? ghv_87 : _GEN_4126; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4128 = 8'h58 == new_ptr_34_value ? ghv_88 : _GEN_4127; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4129 = 8'h59 == new_ptr_34_value ? ghv_89 : _GEN_4128; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4130 = 8'h5a == new_ptr_34_value ? ghv_90 : _GEN_4129; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4131 = 8'h5b == new_ptr_34_value ? ghv_91 : _GEN_4130; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4132 = 8'h5c == new_ptr_34_value ? ghv_92 : _GEN_4131; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4133 = 8'h5d == new_ptr_34_value ? ghv_93 : _GEN_4132; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4134 = 8'h5e == new_ptr_34_value ? ghv_94 : _GEN_4133; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4135 = 8'h5f == new_ptr_34_value ? ghv_95 : _GEN_4134; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4136 = 8'h60 == new_ptr_34_value ? ghv_96 : _GEN_4135; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4137 = 8'h61 == new_ptr_34_value ? ghv_97 : _GEN_4136; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4138 = 8'h62 == new_ptr_34_value ? ghv_98 : _GEN_4137; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4139 = 8'h63 == new_ptr_34_value ? ghv_99 : _GEN_4138; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4140 = 8'h64 == new_ptr_34_value ? ghv_100 : _GEN_4139; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4141 = 8'h65 == new_ptr_34_value ? ghv_101 : _GEN_4140; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4142 = 8'h66 == new_ptr_34_value ? ghv_102 : _GEN_4141; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4143 = 8'h67 == new_ptr_34_value ? ghv_103 : _GEN_4142; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4144 = 8'h68 == new_ptr_34_value ? ghv_104 : _GEN_4143; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4145 = 8'h69 == new_ptr_34_value ? ghv_105 : _GEN_4144; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4146 = 8'h6a == new_ptr_34_value ? ghv_106 : _GEN_4145; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4147 = 8'h6b == new_ptr_34_value ? ghv_107 : _GEN_4146; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4148 = 8'h6c == new_ptr_34_value ? ghv_108 : _GEN_4147; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4149 = 8'h6d == new_ptr_34_value ? ghv_109 : _GEN_4148; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4150 = 8'h6e == new_ptr_34_value ? ghv_110 : _GEN_4149; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4151 = 8'h6f == new_ptr_34_value ? ghv_111 : _GEN_4150; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4152 = 8'h70 == new_ptr_34_value ? ghv_112 : _GEN_4151; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4153 = 8'h71 == new_ptr_34_value ? ghv_113 : _GEN_4152; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4154 = 8'h72 == new_ptr_34_value ? ghv_114 : _GEN_4153; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4155 = 8'h73 == new_ptr_34_value ? ghv_115 : _GEN_4154; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4156 = 8'h74 == new_ptr_34_value ? ghv_116 : _GEN_4155; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4157 = 8'h75 == new_ptr_34_value ? ghv_117 : _GEN_4156; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4158 = 8'h76 == new_ptr_34_value ? ghv_118 : _GEN_4157; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4159 = 8'h77 == new_ptr_34_value ? ghv_119 : _GEN_4158; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4160 = 8'h78 == new_ptr_34_value ? ghv_120 : _GEN_4159; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4161 = 8'h79 == new_ptr_34_value ? ghv_121 : _GEN_4160; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4162 = 8'h7a == new_ptr_34_value ? ghv_122 : _GEN_4161; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4163 = 8'h7b == new_ptr_34_value ? ghv_123 : _GEN_4162; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4164 = 8'h7c == new_ptr_34_value ? ghv_124 : _GEN_4163; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4165 = 8'h7d == new_ptr_34_value ? ghv_125 : _GEN_4164; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4166 = 8'h7e == new_ptr_34_value ? ghv_126 : _GEN_4165; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4167 = 8'h7f == new_ptr_34_value ? ghv_127 : _GEN_4166; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4168 = 8'h80 == new_ptr_34_value ? ghv_128 : _GEN_4167; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4169 = 8'h81 == new_ptr_34_value ? ghv_129 : _GEN_4168; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4170 = 8'h82 == new_ptr_34_value ? ghv_130 : _GEN_4169; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4171 = 8'h83 == new_ptr_34_value ? ghv_131 : _GEN_4170; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4172 = 8'h84 == new_ptr_34_value ? ghv_132 : _GEN_4171; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4173 = 8'h85 == new_ptr_34_value ? ghv_133 : _GEN_4172; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4174 = 8'h86 == new_ptr_34_value ? ghv_134 : _GEN_4173; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4175 = 8'h87 == new_ptr_34_value ? ghv_135 : _GEN_4174; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4176 = 8'h88 == new_ptr_34_value ? ghv_136 : _GEN_4175; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4177 = 8'h89 == new_ptr_34_value ? ghv_137 : _GEN_4176; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4178 = 8'h8a == new_ptr_34_value ? ghv_138 : _GEN_4177; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4179 = 8'h8b == new_ptr_34_value ? ghv_139 : _GEN_4178; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4180 = 8'h8c == new_ptr_34_value ? ghv_140 : _GEN_4179; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4181 = 8'h8d == new_ptr_34_value ? ghv_141 : _GEN_4180; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4182 = 8'h8e == new_ptr_34_value ? ghv_142 : _GEN_4181; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_37_value = _new_ptr_value_T_75[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_4185 = 8'h1 == new_ptr_37_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4186 = 8'h2 == new_ptr_37_value ? ghv_2 : _GEN_4185; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4187 = 8'h3 == new_ptr_37_value ? ghv_3 : _GEN_4186; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4188 = 8'h4 == new_ptr_37_value ? ghv_4 : _GEN_4187; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4189 = 8'h5 == new_ptr_37_value ? ghv_5 : _GEN_4188; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4190 = 8'h6 == new_ptr_37_value ? ghv_6 : _GEN_4189; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4191 = 8'h7 == new_ptr_37_value ? ghv_7 : _GEN_4190; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4192 = 8'h8 == new_ptr_37_value ? ghv_8 : _GEN_4191; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4193 = 8'h9 == new_ptr_37_value ? ghv_9 : _GEN_4192; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4194 = 8'ha == new_ptr_37_value ? ghv_10 : _GEN_4193; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4195 = 8'hb == new_ptr_37_value ? ghv_11 : _GEN_4194; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4196 = 8'hc == new_ptr_37_value ? ghv_12 : _GEN_4195; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4197 = 8'hd == new_ptr_37_value ? ghv_13 : _GEN_4196; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4198 = 8'he == new_ptr_37_value ? ghv_14 : _GEN_4197; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4199 = 8'hf == new_ptr_37_value ? ghv_15 : _GEN_4198; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4200 = 8'h10 == new_ptr_37_value ? ghv_16 : _GEN_4199; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4201 = 8'h11 == new_ptr_37_value ? ghv_17 : _GEN_4200; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4202 = 8'h12 == new_ptr_37_value ? ghv_18 : _GEN_4201; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4203 = 8'h13 == new_ptr_37_value ? ghv_19 : _GEN_4202; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4204 = 8'h14 == new_ptr_37_value ? ghv_20 : _GEN_4203; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4205 = 8'h15 == new_ptr_37_value ? ghv_21 : _GEN_4204; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4206 = 8'h16 == new_ptr_37_value ? ghv_22 : _GEN_4205; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4207 = 8'h17 == new_ptr_37_value ? ghv_23 : _GEN_4206; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4208 = 8'h18 == new_ptr_37_value ? ghv_24 : _GEN_4207; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4209 = 8'h19 == new_ptr_37_value ? ghv_25 : _GEN_4208; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4210 = 8'h1a == new_ptr_37_value ? ghv_26 : _GEN_4209; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4211 = 8'h1b == new_ptr_37_value ? ghv_27 : _GEN_4210; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4212 = 8'h1c == new_ptr_37_value ? ghv_28 : _GEN_4211; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4213 = 8'h1d == new_ptr_37_value ? ghv_29 : _GEN_4212; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4214 = 8'h1e == new_ptr_37_value ? ghv_30 : _GEN_4213; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4215 = 8'h1f == new_ptr_37_value ? ghv_31 : _GEN_4214; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4216 = 8'h20 == new_ptr_37_value ? ghv_32 : _GEN_4215; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4217 = 8'h21 == new_ptr_37_value ? ghv_33 : _GEN_4216; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4218 = 8'h22 == new_ptr_37_value ? ghv_34 : _GEN_4217; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4219 = 8'h23 == new_ptr_37_value ? ghv_35 : _GEN_4218; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4220 = 8'h24 == new_ptr_37_value ? ghv_36 : _GEN_4219; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4221 = 8'h25 == new_ptr_37_value ? ghv_37 : _GEN_4220; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4222 = 8'h26 == new_ptr_37_value ? ghv_38 : _GEN_4221; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4223 = 8'h27 == new_ptr_37_value ? ghv_39 : _GEN_4222; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4224 = 8'h28 == new_ptr_37_value ? ghv_40 : _GEN_4223; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4225 = 8'h29 == new_ptr_37_value ? ghv_41 : _GEN_4224; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4226 = 8'h2a == new_ptr_37_value ? ghv_42 : _GEN_4225; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4227 = 8'h2b == new_ptr_37_value ? ghv_43 : _GEN_4226; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4228 = 8'h2c == new_ptr_37_value ? ghv_44 : _GEN_4227; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4229 = 8'h2d == new_ptr_37_value ? ghv_45 : _GEN_4228; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4230 = 8'h2e == new_ptr_37_value ? ghv_46 : _GEN_4229; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4231 = 8'h2f == new_ptr_37_value ? ghv_47 : _GEN_4230; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4232 = 8'h30 == new_ptr_37_value ? ghv_48 : _GEN_4231; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4233 = 8'h31 == new_ptr_37_value ? ghv_49 : _GEN_4232; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4234 = 8'h32 == new_ptr_37_value ? ghv_50 : _GEN_4233; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4235 = 8'h33 == new_ptr_37_value ? ghv_51 : _GEN_4234; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4236 = 8'h34 == new_ptr_37_value ? ghv_52 : _GEN_4235; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4237 = 8'h35 == new_ptr_37_value ? ghv_53 : _GEN_4236; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4238 = 8'h36 == new_ptr_37_value ? ghv_54 : _GEN_4237; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4239 = 8'h37 == new_ptr_37_value ? ghv_55 : _GEN_4238; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4240 = 8'h38 == new_ptr_37_value ? ghv_56 : _GEN_4239; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4241 = 8'h39 == new_ptr_37_value ? ghv_57 : _GEN_4240; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4242 = 8'h3a == new_ptr_37_value ? ghv_58 : _GEN_4241; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4243 = 8'h3b == new_ptr_37_value ? ghv_59 : _GEN_4242; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4244 = 8'h3c == new_ptr_37_value ? ghv_60 : _GEN_4243; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4245 = 8'h3d == new_ptr_37_value ? ghv_61 : _GEN_4244; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4246 = 8'h3e == new_ptr_37_value ? ghv_62 : _GEN_4245; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4247 = 8'h3f == new_ptr_37_value ? ghv_63 : _GEN_4246; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4248 = 8'h40 == new_ptr_37_value ? ghv_64 : _GEN_4247; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4249 = 8'h41 == new_ptr_37_value ? ghv_65 : _GEN_4248; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4250 = 8'h42 == new_ptr_37_value ? ghv_66 : _GEN_4249; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4251 = 8'h43 == new_ptr_37_value ? ghv_67 : _GEN_4250; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4252 = 8'h44 == new_ptr_37_value ? ghv_68 : _GEN_4251; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4253 = 8'h45 == new_ptr_37_value ? ghv_69 : _GEN_4252; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4254 = 8'h46 == new_ptr_37_value ? ghv_70 : _GEN_4253; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4255 = 8'h47 == new_ptr_37_value ? ghv_71 : _GEN_4254; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4256 = 8'h48 == new_ptr_37_value ? ghv_72 : _GEN_4255; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4257 = 8'h49 == new_ptr_37_value ? ghv_73 : _GEN_4256; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4258 = 8'h4a == new_ptr_37_value ? ghv_74 : _GEN_4257; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4259 = 8'h4b == new_ptr_37_value ? ghv_75 : _GEN_4258; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4260 = 8'h4c == new_ptr_37_value ? ghv_76 : _GEN_4259; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4261 = 8'h4d == new_ptr_37_value ? ghv_77 : _GEN_4260; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4262 = 8'h4e == new_ptr_37_value ? ghv_78 : _GEN_4261; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4263 = 8'h4f == new_ptr_37_value ? ghv_79 : _GEN_4262; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4264 = 8'h50 == new_ptr_37_value ? ghv_80 : _GEN_4263; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4265 = 8'h51 == new_ptr_37_value ? ghv_81 : _GEN_4264; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4266 = 8'h52 == new_ptr_37_value ? ghv_82 : _GEN_4265; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4267 = 8'h53 == new_ptr_37_value ? ghv_83 : _GEN_4266; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4268 = 8'h54 == new_ptr_37_value ? ghv_84 : _GEN_4267; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4269 = 8'h55 == new_ptr_37_value ? ghv_85 : _GEN_4268; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4270 = 8'h56 == new_ptr_37_value ? ghv_86 : _GEN_4269; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4271 = 8'h57 == new_ptr_37_value ? ghv_87 : _GEN_4270; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4272 = 8'h58 == new_ptr_37_value ? ghv_88 : _GEN_4271; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4273 = 8'h59 == new_ptr_37_value ? ghv_89 : _GEN_4272; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4274 = 8'h5a == new_ptr_37_value ? ghv_90 : _GEN_4273; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4275 = 8'h5b == new_ptr_37_value ? ghv_91 : _GEN_4274; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4276 = 8'h5c == new_ptr_37_value ? ghv_92 : _GEN_4275; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4277 = 8'h5d == new_ptr_37_value ? ghv_93 : _GEN_4276; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4278 = 8'h5e == new_ptr_37_value ? ghv_94 : _GEN_4277; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4279 = 8'h5f == new_ptr_37_value ? ghv_95 : _GEN_4278; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4280 = 8'h60 == new_ptr_37_value ? ghv_96 : _GEN_4279; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4281 = 8'h61 == new_ptr_37_value ? ghv_97 : _GEN_4280; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4282 = 8'h62 == new_ptr_37_value ? ghv_98 : _GEN_4281; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4283 = 8'h63 == new_ptr_37_value ? ghv_99 : _GEN_4282; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4284 = 8'h64 == new_ptr_37_value ? ghv_100 : _GEN_4283; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4285 = 8'h65 == new_ptr_37_value ? ghv_101 : _GEN_4284; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4286 = 8'h66 == new_ptr_37_value ? ghv_102 : _GEN_4285; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4287 = 8'h67 == new_ptr_37_value ? ghv_103 : _GEN_4286; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4288 = 8'h68 == new_ptr_37_value ? ghv_104 : _GEN_4287; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4289 = 8'h69 == new_ptr_37_value ? ghv_105 : _GEN_4288; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4290 = 8'h6a == new_ptr_37_value ? ghv_106 : _GEN_4289; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4291 = 8'h6b == new_ptr_37_value ? ghv_107 : _GEN_4290; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4292 = 8'h6c == new_ptr_37_value ? ghv_108 : _GEN_4291; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4293 = 8'h6d == new_ptr_37_value ? ghv_109 : _GEN_4292; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4294 = 8'h6e == new_ptr_37_value ? ghv_110 : _GEN_4293; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4295 = 8'h6f == new_ptr_37_value ? ghv_111 : _GEN_4294; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4296 = 8'h70 == new_ptr_37_value ? ghv_112 : _GEN_4295; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4297 = 8'h71 == new_ptr_37_value ? ghv_113 : _GEN_4296; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4298 = 8'h72 == new_ptr_37_value ? ghv_114 : _GEN_4297; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4299 = 8'h73 == new_ptr_37_value ? ghv_115 : _GEN_4298; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4300 = 8'h74 == new_ptr_37_value ? ghv_116 : _GEN_4299; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4301 = 8'h75 == new_ptr_37_value ? ghv_117 : _GEN_4300; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4302 = 8'h76 == new_ptr_37_value ? ghv_118 : _GEN_4301; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4303 = 8'h77 == new_ptr_37_value ? ghv_119 : _GEN_4302; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4304 = 8'h78 == new_ptr_37_value ? ghv_120 : _GEN_4303; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4305 = 8'h79 == new_ptr_37_value ? ghv_121 : _GEN_4304; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4306 = 8'h7a == new_ptr_37_value ? ghv_122 : _GEN_4305; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4307 = 8'h7b == new_ptr_37_value ? ghv_123 : _GEN_4306; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4308 = 8'h7c == new_ptr_37_value ? ghv_124 : _GEN_4307; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4309 = 8'h7d == new_ptr_37_value ? ghv_125 : _GEN_4308; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4310 = 8'h7e == new_ptr_37_value ? ghv_126 : _GEN_4309; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4311 = 8'h7f == new_ptr_37_value ? ghv_127 : _GEN_4310; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4312 = 8'h80 == new_ptr_37_value ? ghv_128 : _GEN_4311; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4313 = 8'h81 == new_ptr_37_value ? ghv_129 : _GEN_4312; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4314 = 8'h82 == new_ptr_37_value ? ghv_130 : _GEN_4313; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4315 = 8'h83 == new_ptr_37_value ? ghv_131 : _GEN_4314; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4316 = 8'h84 == new_ptr_37_value ? ghv_132 : _GEN_4315; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4317 = 8'h85 == new_ptr_37_value ? ghv_133 : _GEN_4316; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4318 = 8'h86 == new_ptr_37_value ? ghv_134 : _GEN_4317; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4319 = 8'h87 == new_ptr_37_value ? ghv_135 : _GEN_4318; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4320 = 8'h88 == new_ptr_37_value ? ghv_136 : _GEN_4319; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4321 = 8'h89 == new_ptr_37_value ? ghv_137 : _GEN_4320; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4322 = 8'h8a == new_ptr_37_value ? ghv_138 : _GEN_4321; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4323 = 8'h8b == new_ptr_37_value ? ghv_139 : _GEN_4322; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4324 = 8'h8c == new_ptr_37_value ? ghv_140 : _GEN_4323; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4325 = 8'h8d == new_ptr_37_value ? ghv_141 : _GEN_4324; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4326 = 8'h8e == new_ptr_37_value ? ghv_142 : _GEN_4325; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_24_value = _new_ptr_value_T_49[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_4329 = 8'h1 == new_ptr_24_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4330 = 8'h2 == new_ptr_24_value ? ghv_2 : _GEN_4329; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4331 = 8'h3 == new_ptr_24_value ? ghv_3 : _GEN_4330; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4332 = 8'h4 == new_ptr_24_value ? ghv_4 : _GEN_4331; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4333 = 8'h5 == new_ptr_24_value ? ghv_5 : _GEN_4332; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4334 = 8'h6 == new_ptr_24_value ? ghv_6 : _GEN_4333; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4335 = 8'h7 == new_ptr_24_value ? ghv_7 : _GEN_4334; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4336 = 8'h8 == new_ptr_24_value ? ghv_8 : _GEN_4335; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4337 = 8'h9 == new_ptr_24_value ? ghv_9 : _GEN_4336; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4338 = 8'ha == new_ptr_24_value ? ghv_10 : _GEN_4337; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4339 = 8'hb == new_ptr_24_value ? ghv_11 : _GEN_4338; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4340 = 8'hc == new_ptr_24_value ? ghv_12 : _GEN_4339; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4341 = 8'hd == new_ptr_24_value ? ghv_13 : _GEN_4340; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4342 = 8'he == new_ptr_24_value ? ghv_14 : _GEN_4341; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4343 = 8'hf == new_ptr_24_value ? ghv_15 : _GEN_4342; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4344 = 8'h10 == new_ptr_24_value ? ghv_16 : _GEN_4343; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4345 = 8'h11 == new_ptr_24_value ? ghv_17 : _GEN_4344; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4346 = 8'h12 == new_ptr_24_value ? ghv_18 : _GEN_4345; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4347 = 8'h13 == new_ptr_24_value ? ghv_19 : _GEN_4346; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4348 = 8'h14 == new_ptr_24_value ? ghv_20 : _GEN_4347; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4349 = 8'h15 == new_ptr_24_value ? ghv_21 : _GEN_4348; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4350 = 8'h16 == new_ptr_24_value ? ghv_22 : _GEN_4349; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4351 = 8'h17 == new_ptr_24_value ? ghv_23 : _GEN_4350; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4352 = 8'h18 == new_ptr_24_value ? ghv_24 : _GEN_4351; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4353 = 8'h19 == new_ptr_24_value ? ghv_25 : _GEN_4352; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4354 = 8'h1a == new_ptr_24_value ? ghv_26 : _GEN_4353; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4355 = 8'h1b == new_ptr_24_value ? ghv_27 : _GEN_4354; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4356 = 8'h1c == new_ptr_24_value ? ghv_28 : _GEN_4355; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4357 = 8'h1d == new_ptr_24_value ? ghv_29 : _GEN_4356; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4358 = 8'h1e == new_ptr_24_value ? ghv_30 : _GEN_4357; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4359 = 8'h1f == new_ptr_24_value ? ghv_31 : _GEN_4358; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4360 = 8'h20 == new_ptr_24_value ? ghv_32 : _GEN_4359; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4361 = 8'h21 == new_ptr_24_value ? ghv_33 : _GEN_4360; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4362 = 8'h22 == new_ptr_24_value ? ghv_34 : _GEN_4361; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4363 = 8'h23 == new_ptr_24_value ? ghv_35 : _GEN_4362; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4364 = 8'h24 == new_ptr_24_value ? ghv_36 : _GEN_4363; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4365 = 8'h25 == new_ptr_24_value ? ghv_37 : _GEN_4364; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4366 = 8'h26 == new_ptr_24_value ? ghv_38 : _GEN_4365; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4367 = 8'h27 == new_ptr_24_value ? ghv_39 : _GEN_4366; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4368 = 8'h28 == new_ptr_24_value ? ghv_40 : _GEN_4367; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4369 = 8'h29 == new_ptr_24_value ? ghv_41 : _GEN_4368; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4370 = 8'h2a == new_ptr_24_value ? ghv_42 : _GEN_4369; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4371 = 8'h2b == new_ptr_24_value ? ghv_43 : _GEN_4370; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4372 = 8'h2c == new_ptr_24_value ? ghv_44 : _GEN_4371; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4373 = 8'h2d == new_ptr_24_value ? ghv_45 : _GEN_4372; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4374 = 8'h2e == new_ptr_24_value ? ghv_46 : _GEN_4373; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4375 = 8'h2f == new_ptr_24_value ? ghv_47 : _GEN_4374; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4376 = 8'h30 == new_ptr_24_value ? ghv_48 : _GEN_4375; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4377 = 8'h31 == new_ptr_24_value ? ghv_49 : _GEN_4376; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4378 = 8'h32 == new_ptr_24_value ? ghv_50 : _GEN_4377; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4379 = 8'h33 == new_ptr_24_value ? ghv_51 : _GEN_4378; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4380 = 8'h34 == new_ptr_24_value ? ghv_52 : _GEN_4379; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4381 = 8'h35 == new_ptr_24_value ? ghv_53 : _GEN_4380; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4382 = 8'h36 == new_ptr_24_value ? ghv_54 : _GEN_4381; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4383 = 8'h37 == new_ptr_24_value ? ghv_55 : _GEN_4382; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4384 = 8'h38 == new_ptr_24_value ? ghv_56 : _GEN_4383; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4385 = 8'h39 == new_ptr_24_value ? ghv_57 : _GEN_4384; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4386 = 8'h3a == new_ptr_24_value ? ghv_58 : _GEN_4385; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4387 = 8'h3b == new_ptr_24_value ? ghv_59 : _GEN_4386; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4388 = 8'h3c == new_ptr_24_value ? ghv_60 : _GEN_4387; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4389 = 8'h3d == new_ptr_24_value ? ghv_61 : _GEN_4388; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4390 = 8'h3e == new_ptr_24_value ? ghv_62 : _GEN_4389; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4391 = 8'h3f == new_ptr_24_value ? ghv_63 : _GEN_4390; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4392 = 8'h40 == new_ptr_24_value ? ghv_64 : _GEN_4391; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4393 = 8'h41 == new_ptr_24_value ? ghv_65 : _GEN_4392; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4394 = 8'h42 == new_ptr_24_value ? ghv_66 : _GEN_4393; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4395 = 8'h43 == new_ptr_24_value ? ghv_67 : _GEN_4394; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4396 = 8'h44 == new_ptr_24_value ? ghv_68 : _GEN_4395; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4397 = 8'h45 == new_ptr_24_value ? ghv_69 : _GEN_4396; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4398 = 8'h46 == new_ptr_24_value ? ghv_70 : _GEN_4397; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4399 = 8'h47 == new_ptr_24_value ? ghv_71 : _GEN_4398; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4400 = 8'h48 == new_ptr_24_value ? ghv_72 : _GEN_4399; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4401 = 8'h49 == new_ptr_24_value ? ghv_73 : _GEN_4400; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4402 = 8'h4a == new_ptr_24_value ? ghv_74 : _GEN_4401; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4403 = 8'h4b == new_ptr_24_value ? ghv_75 : _GEN_4402; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4404 = 8'h4c == new_ptr_24_value ? ghv_76 : _GEN_4403; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4405 = 8'h4d == new_ptr_24_value ? ghv_77 : _GEN_4404; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4406 = 8'h4e == new_ptr_24_value ? ghv_78 : _GEN_4405; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4407 = 8'h4f == new_ptr_24_value ? ghv_79 : _GEN_4406; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4408 = 8'h50 == new_ptr_24_value ? ghv_80 : _GEN_4407; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4409 = 8'h51 == new_ptr_24_value ? ghv_81 : _GEN_4408; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4410 = 8'h52 == new_ptr_24_value ? ghv_82 : _GEN_4409; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4411 = 8'h53 == new_ptr_24_value ? ghv_83 : _GEN_4410; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4412 = 8'h54 == new_ptr_24_value ? ghv_84 : _GEN_4411; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4413 = 8'h55 == new_ptr_24_value ? ghv_85 : _GEN_4412; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4414 = 8'h56 == new_ptr_24_value ? ghv_86 : _GEN_4413; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4415 = 8'h57 == new_ptr_24_value ? ghv_87 : _GEN_4414; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4416 = 8'h58 == new_ptr_24_value ? ghv_88 : _GEN_4415; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4417 = 8'h59 == new_ptr_24_value ? ghv_89 : _GEN_4416; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4418 = 8'h5a == new_ptr_24_value ? ghv_90 : _GEN_4417; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4419 = 8'h5b == new_ptr_24_value ? ghv_91 : _GEN_4418; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4420 = 8'h5c == new_ptr_24_value ? ghv_92 : _GEN_4419; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4421 = 8'h5d == new_ptr_24_value ? ghv_93 : _GEN_4420; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4422 = 8'h5e == new_ptr_24_value ? ghv_94 : _GEN_4421; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4423 = 8'h5f == new_ptr_24_value ? ghv_95 : _GEN_4422; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4424 = 8'h60 == new_ptr_24_value ? ghv_96 : _GEN_4423; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4425 = 8'h61 == new_ptr_24_value ? ghv_97 : _GEN_4424; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4426 = 8'h62 == new_ptr_24_value ? ghv_98 : _GEN_4425; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4427 = 8'h63 == new_ptr_24_value ? ghv_99 : _GEN_4426; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4428 = 8'h64 == new_ptr_24_value ? ghv_100 : _GEN_4427; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4429 = 8'h65 == new_ptr_24_value ? ghv_101 : _GEN_4428; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4430 = 8'h66 == new_ptr_24_value ? ghv_102 : _GEN_4429; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4431 = 8'h67 == new_ptr_24_value ? ghv_103 : _GEN_4430; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4432 = 8'h68 == new_ptr_24_value ? ghv_104 : _GEN_4431; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4433 = 8'h69 == new_ptr_24_value ? ghv_105 : _GEN_4432; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4434 = 8'h6a == new_ptr_24_value ? ghv_106 : _GEN_4433; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4435 = 8'h6b == new_ptr_24_value ? ghv_107 : _GEN_4434; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4436 = 8'h6c == new_ptr_24_value ? ghv_108 : _GEN_4435; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4437 = 8'h6d == new_ptr_24_value ? ghv_109 : _GEN_4436; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4438 = 8'h6e == new_ptr_24_value ? ghv_110 : _GEN_4437; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4439 = 8'h6f == new_ptr_24_value ? ghv_111 : _GEN_4438; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4440 = 8'h70 == new_ptr_24_value ? ghv_112 : _GEN_4439; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4441 = 8'h71 == new_ptr_24_value ? ghv_113 : _GEN_4440; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4442 = 8'h72 == new_ptr_24_value ? ghv_114 : _GEN_4441; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4443 = 8'h73 == new_ptr_24_value ? ghv_115 : _GEN_4442; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4444 = 8'h74 == new_ptr_24_value ? ghv_116 : _GEN_4443; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4445 = 8'h75 == new_ptr_24_value ? ghv_117 : _GEN_4444; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4446 = 8'h76 == new_ptr_24_value ? ghv_118 : _GEN_4445; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4447 = 8'h77 == new_ptr_24_value ? ghv_119 : _GEN_4446; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4448 = 8'h78 == new_ptr_24_value ? ghv_120 : _GEN_4447; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4449 = 8'h79 == new_ptr_24_value ? ghv_121 : _GEN_4448; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4450 = 8'h7a == new_ptr_24_value ? ghv_122 : _GEN_4449; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4451 = 8'h7b == new_ptr_24_value ? ghv_123 : _GEN_4450; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4452 = 8'h7c == new_ptr_24_value ? ghv_124 : _GEN_4451; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4453 = 8'h7d == new_ptr_24_value ? ghv_125 : _GEN_4452; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4454 = 8'h7e == new_ptr_24_value ? ghv_126 : _GEN_4453; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4455 = 8'h7f == new_ptr_24_value ? ghv_127 : _GEN_4454; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4456 = 8'h80 == new_ptr_24_value ? ghv_128 : _GEN_4455; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4457 = 8'h81 == new_ptr_24_value ? ghv_129 : _GEN_4456; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4458 = 8'h82 == new_ptr_24_value ? ghv_130 : _GEN_4457; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4459 = 8'h83 == new_ptr_24_value ? ghv_131 : _GEN_4458; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4460 = 8'h84 == new_ptr_24_value ? ghv_132 : _GEN_4459; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4461 = 8'h85 == new_ptr_24_value ? ghv_133 : _GEN_4460; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4462 = 8'h86 == new_ptr_24_value ? ghv_134 : _GEN_4461; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4463 = 8'h87 == new_ptr_24_value ? ghv_135 : _GEN_4462; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4464 = 8'h88 == new_ptr_24_value ? ghv_136 : _GEN_4463; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4465 = 8'h89 == new_ptr_24_value ? ghv_137 : _GEN_4464; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4466 = 8'h8a == new_ptr_24_value ? ghv_138 : _GEN_4465; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4467 = 8'h8b == new_ptr_24_value ? ghv_139 : _GEN_4466; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4468 = 8'h8c == new_ptr_24_value ? ghv_140 : _GEN_4467; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4469 = 8'h8d == new_ptr_24_value ? ghv_141 : _GEN_4468; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4470 = 8'h8e == new_ptr_24_value ? ghv_142 : _GEN_4469; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_28_value = _new_ptr_value_T_57[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_4473 = 8'h1 == new_ptr_28_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4474 = 8'h2 == new_ptr_28_value ? ghv_2 : _GEN_4473; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4475 = 8'h3 == new_ptr_28_value ? ghv_3 : _GEN_4474; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4476 = 8'h4 == new_ptr_28_value ? ghv_4 : _GEN_4475; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4477 = 8'h5 == new_ptr_28_value ? ghv_5 : _GEN_4476; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4478 = 8'h6 == new_ptr_28_value ? ghv_6 : _GEN_4477; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4479 = 8'h7 == new_ptr_28_value ? ghv_7 : _GEN_4478; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4480 = 8'h8 == new_ptr_28_value ? ghv_8 : _GEN_4479; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4481 = 8'h9 == new_ptr_28_value ? ghv_9 : _GEN_4480; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4482 = 8'ha == new_ptr_28_value ? ghv_10 : _GEN_4481; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4483 = 8'hb == new_ptr_28_value ? ghv_11 : _GEN_4482; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4484 = 8'hc == new_ptr_28_value ? ghv_12 : _GEN_4483; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4485 = 8'hd == new_ptr_28_value ? ghv_13 : _GEN_4484; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4486 = 8'he == new_ptr_28_value ? ghv_14 : _GEN_4485; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4487 = 8'hf == new_ptr_28_value ? ghv_15 : _GEN_4486; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4488 = 8'h10 == new_ptr_28_value ? ghv_16 : _GEN_4487; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4489 = 8'h11 == new_ptr_28_value ? ghv_17 : _GEN_4488; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4490 = 8'h12 == new_ptr_28_value ? ghv_18 : _GEN_4489; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4491 = 8'h13 == new_ptr_28_value ? ghv_19 : _GEN_4490; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4492 = 8'h14 == new_ptr_28_value ? ghv_20 : _GEN_4491; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4493 = 8'h15 == new_ptr_28_value ? ghv_21 : _GEN_4492; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4494 = 8'h16 == new_ptr_28_value ? ghv_22 : _GEN_4493; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4495 = 8'h17 == new_ptr_28_value ? ghv_23 : _GEN_4494; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4496 = 8'h18 == new_ptr_28_value ? ghv_24 : _GEN_4495; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4497 = 8'h19 == new_ptr_28_value ? ghv_25 : _GEN_4496; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4498 = 8'h1a == new_ptr_28_value ? ghv_26 : _GEN_4497; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4499 = 8'h1b == new_ptr_28_value ? ghv_27 : _GEN_4498; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4500 = 8'h1c == new_ptr_28_value ? ghv_28 : _GEN_4499; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4501 = 8'h1d == new_ptr_28_value ? ghv_29 : _GEN_4500; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4502 = 8'h1e == new_ptr_28_value ? ghv_30 : _GEN_4501; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4503 = 8'h1f == new_ptr_28_value ? ghv_31 : _GEN_4502; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4504 = 8'h20 == new_ptr_28_value ? ghv_32 : _GEN_4503; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4505 = 8'h21 == new_ptr_28_value ? ghv_33 : _GEN_4504; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4506 = 8'h22 == new_ptr_28_value ? ghv_34 : _GEN_4505; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4507 = 8'h23 == new_ptr_28_value ? ghv_35 : _GEN_4506; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4508 = 8'h24 == new_ptr_28_value ? ghv_36 : _GEN_4507; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4509 = 8'h25 == new_ptr_28_value ? ghv_37 : _GEN_4508; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4510 = 8'h26 == new_ptr_28_value ? ghv_38 : _GEN_4509; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4511 = 8'h27 == new_ptr_28_value ? ghv_39 : _GEN_4510; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4512 = 8'h28 == new_ptr_28_value ? ghv_40 : _GEN_4511; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4513 = 8'h29 == new_ptr_28_value ? ghv_41 : _GEN_4512; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4514 = 8'h2a == new_ptr_28_value ? ghv_42 : _GEN_4513; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4515 = 8'h2b == new_ptr_28_value ? ghv_43 : _GEN_4514; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4516 = 8'h2c == new_ptr_28_value ? ghv_44 : _GEN_4515; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4517 = 8'h2d == new_ptr_28_value ? ghv_45 : _GEN_4516; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4518 = 8'h2e == new_ptr_28_value ? ghv_46 : _GEN_4517; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4519 = 8'h2f == new_ptr_28_value ? ghv_47 : _GEN_4518; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4520 = 8'h30 == new_ptr_28_value ? ghv_48 : _GEN_4519; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4521 = 8'h31 == new_ptr_28_value ? ghv_49 : _GEN_4520; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4522 = 8'h32 == new_ptr_28_value ? ghv_50 : _GEN_4521; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4523 = 8'h33 == new_ptr_28_value ? ghv_51 : _GEN_4522; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4524 = 8'h34 == new_ptr_28_value ? ghv_52 : _GEN_4523; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4525 = 8'h35 == new_ptr_28_value ? ghv_53 : _GEN_4524; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4526 = 8'h36 == new_ptr_28_value ? ghv_54 : _GEN_4525; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4527 = 8'h37 == new_ptr_28_value ? ghv_55 : _GEN_4526; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4528 = 8'h38 == new_ptr_28_value ? ghv_56 : _GEN_4527; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4529 = 8'h39 == new_ptr_28_value ? ghv_57 : _GEN_4528; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4530 = 8'h3a == new_ptr_28_value ? ghv_58 : _GEN_4529; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4531 = 8'h3b == new_ptr_28_value ? ghv_59 : _GEN_4530; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4532 = 8'h3c == new_ptr_28_value ? ghv_60 : _GEN_4531; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4533 = 8'h3d == new_ptr_28_value ? ghv_61 : _GEN_4532; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4534 = 8'h3e == new_ptr_28_value ? ghv_62 : _GEN_4533; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4535 = 8'h3f == new_ptr_28_value ? ghv_63 : _GEN_4534; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4536 = 8'h40 == new_ptr_28_value ? ghv_64 : _GEN_4535; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4537 = 8'h41 == new_ptr_28_value ? ghv_65 : _GEN_4536; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4538 = 8'h42 == new_ptr_28_value ? ghv_66 : _GEN_4537; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4539 = 8'h43 == new_ptr_28_value ? ghv_67 : _GEN_4538; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4540 = 8'h44 == new_ptr_28_value ? ghv_68 : _GEN_4539; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4541 = 8'h45 == new_ptr_28_value ? ghv_69 : _GEN_4540; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4542 = 8'h46 == new_ptr_28_value ? ghv_70 : _GEN_4541; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4543 = 8'h47 == new_ptr_28_value ? ghv_71 : _GEN_4542; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4544 = 8'h48 == new_ptr_28_value ? ghv_72 : _GEN_4543; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4545 = 8'h49 == new_ptr_28_value ? ghv_73 : _GEN_4544; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4546 = 8'h4a == new_ptr_28_value ? ghv_74 : _GEN_4545; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4547 = 8'h4b == new_ptr_28_value ? ghv_75 : _GEN_4546; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4548 = 8'h4c == new_ptr_28_value ? ghv_76 : _GEN_4547; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4549 = 8'h4d == new_ptr_28_value ? ghv_77 : _GEN_4548; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4550 = 8'h4e == new_ptr_28_value ? ghv_78 : _GEN_4549; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4551 = 8'h4f == new_ptr_28_value ? ghv_79 : _GEN_4550; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4552 = 8'h50 == new_ptr_28_value ? ghv_80 : _GEN_4551; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4553 = 8'h51 == new_ptr_28_value ? ghv_81 : _GEN_4552; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4554 = 8'h52 == new_ptr_28_value ? ghv_82 : _GEN_4553; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4555 = 8'h53 == new_ptr_28_value ? ghv_83 : _GEN_4554; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4556 = 8'h54 == new_ptr_28_value ? ghv_84 : _GEN_4555; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4557 = 8'h55 == new_ptr_28_value ? ghv_85 : _GEN_4556; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4558 = 8'h56 == new_ptr_28_value ? ghv_86 : _GEN_4557; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4559 = 8'h57 == new_ptr_28_value ? ghv_87 : _GEN_4558; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4560 = 8'h58 == new_ptr_28_value ? ghv_88 : _GEN_4559; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4561 = 8'h59 == new_ptr_28_value ? ghv_89 : _GEN_4560; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4562 = 8'h5a == new_ptr_28_value ? ghv_90 : _GEN_4561; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4563 = 8'h5b == new_ptr_28_value ? ghv_91 : _GEN_4562; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4564 = 8'h5c == new_ptr_28_value ? ghv_92 : _GEN_4563; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4565 = 8'h5d == new_ptr_28_value ? ghv_93 : _GEN_4564; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4566 = 8'h5e == new_ptr_28_value ? ghv_94 : _GEN_4565; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4567 = 8'h5f == new_ptr_28_value ? ghv_95 : _GEN_4566; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4568 = 8'h60 == new_ptr_28_value ? ghv_96 : _GEN_4567; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4569 = 8'h61 == new_ptr_28_value ? ghv_97 : _GEN_4568; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4570 = 8'h62 == new_ptr_28_value ? ghv_98 : _GEN_4569; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4571 = 8'h63 == new_ptr_28_value ? ghv_99 : _GEN_4570; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4572 = 8'h64 == new_ptr_28_value ? ghv_100 : _GEN_4571; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4573 = 8'h65 == new_ptr_28_value ? ghv_101 : _GEN_4572; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4574 = 8'h66 == new_ptr_28_value ? ghv_102 : _GEN_4573; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4575 = 8'h67 == new_ptr_28_value ? ghv_103 : _GEN_4574; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4576 = 8'h68 == new_ptr_28_value ? ghv_104 : _GEN_4575; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4577 = 8'h69 == new_ptr_28_value ? ghv_105 : _GEN_4576; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4578 = 8'h6a == new_ptr_28_value ? ghv_106 : _GEN_4577; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4579 = 8'h6b == new_ptr_28_value ? ghv_107 : _GEN_4578; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4580 = 8'h6c == new_ptr_28_value ? ghv_108 : _GEN_4579; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4581 = 8'h6d == new_ptr_28_value ? ghv_109 : _GEN_4580; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4582 = 8'h6e == new_ptr_28_value ? ghv_110 : _GEN_4581; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4583 = 8'h6f == new_ptr_28_value ? ghv_111 : _GEN_4582; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4584 = 8'h70 == new_ptr_28_value ? ghv_112 : _GEN_4583; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4585 = 8'h71 == new_ptr_28_value ? ghv_113 : _GEN_4584; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4586 = 8'h72 == new_ptr_28_value ? ghv_114 : _GEN_4585; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4587 = 8'h73 == new_ptr_28_value ? ghv_115 : _GEN_4586; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4588 = 8'h74 == new_ptr_28_value ? ghv_116 : _GEN_4587; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4589 = 8'h75 == new_ptr_28_value ? ghv_117 : _GEN_4588; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4590 = 8'h76 == new_ptr_28_value ? ghv_118 : _GEN_4589; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4591 = 8'h77 == new_ptr_28_value ? ghv_119 : _GEN_4590; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4592 = 8'h78 == new_ptr_28_value ? ghv_120 : _GEN_4591; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4593 = 8'h79 == new_ptr_28_value ? ghv_121 : _GEN_4592; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4594 = 8'h7a == new_ptr_28_value ? ghv_122 : _GEN_4593; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4595 = 8'h7b == new_ptr_28_value ? ghv_123 : _GEN_4594; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4596 = 8'h7c == new_ptr_28_value ? ghv_124 : _GEN_4595; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4597 = 8'h7d == new_ptr_28_value ? ghv_125 : _GEN_4596; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4598 = 8'h7e == new_ptr_28_value ? ghv_126 : _GEN_4597; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4599 = 8'h7f == new_ptr_28_value ? ghv_127 : _GEN_4598; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4600 = 8'h80 == new_ptr_28_value ? ghv_128 : _GEN_4599; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4601 = 8'h81 == new_ptr_28_value ? ghv_129 : _GEN_4600; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4602 = 8'h82 == new_ptr_28_value ? ghv_130 : _GEN_4601; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4603 = 8'h83 == new_ptr_28_value ? ghv_131 : _GEN_4602; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4604 = 8'h84 == new_ptr_28_value ? ghv_132 : _GEN_4603; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4605 = 8'h85 == new_ptr_28_value ? ghv_133 : _GEN_4604; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4606 = 8'h86 == new_ptr_28_value ? ghv_134 : _GEN_4605; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4607 = 8'h87 == new_ptr_28_value ? ghv_135 : _GEN_4606; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4608 = 8'h88 == new_ptr_28_value ? ghv_136 : _GEN_4607; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4609 = 8'h89 == new_ptr_28_value ? ghv_137 : _GEN_4608; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4610 = 8'h8a == new_ptr_28_value ? ghv_138 : _GEN_4609; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4611 = 8'h8b == new_ptr_28_value ? ghv_139 : _GEN_4610; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4612 = 8'h8c == new_ptr_28_value ? ghv_140 : _GEN_4611; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4613 = 8'h8d == new_ptr_28_value ? ghv_141 : _GEN_4612; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4614 = 8'h8e == new_ptr_28_value ? ghv_142 : _GEN_4613; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_39_value = _new_ptr_value_T_79[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_4617 = 8'h1 == new_ptr_39_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4618 = 8'h2 == new_ptr_39_value ? ghv_2 : _GEN_4617; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4619 = 8'h3 == new_ptr_39_value ? ghv_3 : _GEN_4618; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4620 = 8'h4 == new_ptr_39_value ? ghv_4 : _GEN_4619; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4621 = 8'h5 == new_ptr_39_value ? ghv_5 : _GEN_4620; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4622 = 8'h6 == new_ptr_39_value ? ghv_6 : _GEN_4621; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4623 = 8'h7 == new_ptr_39_value ? ghv_7 : _GEN_4622; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4624 = 8'h8 == new_ptr_39_value ? ghv_8 : _GEN_4623; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4625 = 8'h9 == new_ptr_39_value ? ghv_9 : _GEN_4624; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4626 = 8'ha == new_ptr_39_value ? ghv_10 : _GEN_4625; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4627 = 8'hb == new_ptr_39_value ? ghv_11 : _GEN_4626; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4628 = 8'hc == new_ptr_39_value ? ghv_12 : _GEN_4627; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4629 = 8'hd == new_ptr_39_value ? ghv_13 : _GEN_4628; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4630 = 8'he == new_ptr_39_value ? ghv_14 : _GEN_4629; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4631 = 8'hf == new_ptr_39_value ? ghv_15 : _GEN_4630; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4632 = 8'h10 == new_ptr_39_value ? ghv_16 : _GEN_4631; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4633 = 8'h11 == new_ptr_39_value ? ghv_17 : _GEN_4632; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4634 = 8'h12 == new_ptr_39_value ? ghv_18 : _GEN_4633; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4635 = 8'h13 == new_ptr_39_value ? ghv_19 : _GEN_4634; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4636 = 8'h14 == new_ptr_39_value ? ghv_20 : _GEN_4635; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4637 = 8'h15 == new_ptr_39_value ? ghv_21 : _GEN_4636; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4638 = 8'h16 == new_ptr_39_value ? ghv_22 : _GEN_4637; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4639 = 8'h17 == new_ptr_39_value ? ghv_23 : _GEN_4638; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4640 = 8'h18 == new_ptr_39_value ? ghv_24 : _GEN_4639; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4641 = 8'h19 == new_ptr_39_value ? ghv_25 : _GEN_4640; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4642 = 8'h1a == new_ptr_39_value ? ghv_26 : _GEN_4641; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4643 = 8'h1b == new_ptr_39_value ? ghv_27 : _GEN_4642; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4644 = 8'h1c == new_ptr_39_value ? ghv_28 : _GEN_4643; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4645 = 8'h1d == new_ptr_39_value ? ghv_29 : _GEN_4644; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4646 = 8'h1e == new_ptr_39_value ? ghv_30 : _GEN_4645; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4647 = 8'h1f == new_ptr_39_value ? ghv_31 : _GEN_4646; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4648 = 8'h20 == new_ptr_39_value ? ghv_32 : _GEN_4647; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4649 = 8'h21 == new_ptr_39_value ? ghv_33 : _GEN_4648; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4650 = 8'h22 == new_ptr_39_value ? ghv_34 : _GEN_4649; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4651 = 8'h23 == new_ptr_39_value ? ghv_35 : _GEN_4650; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4652 = 8'h24 == new_ptr_39_value ? ghv_36 : _GEN_4651; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4653 = 8'h25 == new_ptr_39_value ? ghv_37 : _GEN_4652; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4654 = 8'h26 == new_ptr_39_value ? ghv_38 : _GEN_4653; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4655 = 8'h27 == new_ptr_39_value ? ghv_39 : _GEN_4654; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4656 = 8'h28 == new_ptr_39_value ? ghv_40 : _GEN_4655; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4657 = 8'h29 == new_ptr_39_value ? ghv_41 : _GEN_4656; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4658 = 8'h2a == new_ptr_39_value ? ghv_42 : _GEN_4657; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4659 = 8'h2b == new_ptr_39_value ? ghv_43 : _GEN_4658; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4660 = 8'h2c == new_ptr_39_value ? ghv_44 : _GEN_4659; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4661 = 8'h2d == new_ptr_39_value ? ghv_45 : _GEN_4660; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4662 = 8'h2e == new_ptr_39_value ? ghv_46 : _GEN_4661; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4663 = 8'h2f == new_ptr_39_value ? ghv_47 : _GEN_4662; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4664 = 8'h30 == new_ptr_39_value ? ghv_48 : _GEN_4663; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4665 = 8'h31 == new_ptr_39_value ? ghv_49 : _GEN_4664; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4666 = 8'h32 == new_ptr_39_value ? ghv_50 : _GEN_4665; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4667 = 8'h33 == new_ptr_39_value ? ghv_51 : _GEN_4666; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4668 = 8'h34 == new_ptr_39_value ? ghv_52 : _GEN_4667; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4669 = 8'h35 == new_ptr_39_value ? ghv_53 : _GEN_4668; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4670 = 8'h36 == new_ptr_39_value ? ghv_54 : _GEN_4669; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4671 = 8'h37 == new_ptr_39_value ? ghv_55 : _GEN_4670; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4672 = 8'h38 == new_ptr_39_value ? ghv_56 : _GEN_4671; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4673 = 8'h39 == new_ptr_39_value ? ghv_57 : _GEN_4672; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4674 = 8'h3a == new_ptr_39_value ? ghv_58 : _GEN_4673; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4675 = 8'h3b == new_ptr_39_value ? ghv_59 : _GEN_4674; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4676 = 8'h3c == new_ptr_39_value ? ghv_60 : _GEN_4675; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4677 = 8'h3d == new_ptr_39_value ? ghv_61 : _GEN_4676; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4678 = 8'h3e == new_ptr_39_value ? ghv_62 : _GEN_4677; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4679 = 8'h3f == new_ptr_39_value ? ghv_63 : _GEN_4678; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4680 = 8'h40 == new_ptr_39_value ? ghv_64 : _GEN_4679; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4681 = 8'h41 == new_ptr_39_value ? ghv_65 : _GEN_4680; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4682 = 8'h42 == new_ptr_39_value ? ghv_66 : _GEN_4681; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4683 = 8'h43 == new_ptr_39_value ? ghv_67 : _GEN_4682; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4684 = 8'h44 == new_ptr_39_value ? ghv_68 : _GEN_4683; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4685 = 8'h45 == new_ptr_39_value ? ghv_69 : _GEN_4684; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4686 = 8'h46 == new_ptr_39_value ? ghv_70 : _GEN_4685; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4687 = 8'h47 == new_ptr_39_value ? ghv_71 : _GEN_4686; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4688 = 8'h48 == new_ptr_39_value ? ghv_72 : _GEN_4687; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4689 = 8'h49 == new_ptr_39_value ? ghv_73 : _GEN_4688; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4690 = 8'h4a == new_ptr_39_value ? ghv_74 : _GEN_4689; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4691 = 8'h4b == new_ptr_39_value ? ghv_75 : _GEN_4690; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4692 = 8'h4c == new_ptr_39_value ? ghv_76 : _GEN_4691; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4693 = 8'h4d == new_ptr_39_value ? ghv_77 : _GEN_4692; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4694 = 8'h4e == new_ptr_39_value ? ghv_78 : _GEN_4693; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4695 = 8'h4f == new_ptr_39_value ? ghv_79 : _GEN_4694; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4696 = 8'h50 == new_ptr_39_value ? ghv_80 : _GEN_4695; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4697 = 8'h51 == new_ptr_39_value ? ghv_81 : _GEN_4696; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4698 = 8'h52 == new_ptr_39_value ? ghv_82 : _GEN_4697; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4699 = 8'h53 == new_ptr_39_value ? ghv_83 : _GEN_4698; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4700 = 8'h54 == new_ptr_39_value ? ghv_84 : _GEN_4699; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4701 = 8'h55 == new_ptr_39_value ? ghv_85 : _GEN_4700; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4702 = 8'h56 == new_ptr_39_value ? ghv_86 : _GEN_4701; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4703 = 8'h57 == new_ptr_39_value ? ghv_87 : _GEN_4702; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4704 = 8'h58 == new_ptr_39_value ? ghv_88 : _GEN_4703; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4705 = 8'h59 == new_ptr_39_value ? ghv_89 : _GEN_4704; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4706 = 8'h5a == new_ptr_39_value ? ghv_90 : _GEN_4705; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4707 = 8'h5b == new_ptr_39_value ? ghv_91 : _GEN_4706; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4708 = 8'h5c == new_ptr_39_value ? ghv_92 : _GEN_4707; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4709 = 8'h5d == new_ptr_39_value ? ghv_93 : _GEN_4708; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4710 = 8'h5e == new_ptr_39_value ? ghv_94 : _GEN_4709; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4711 = 8'h5f == new_ptr_39_value ? ghv_95 : _GEN_4710; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4712 = 8'h60 == new_ptr_39_value ? ghv_96 : _GEN_4711; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4713 = 8'h61 == new_ptr_39_value ? ghv_97 : _GEN_4712; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4714 = 8'h62 == new_ptr_39_value ? ghv_98 : _GEN_4713; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4715 = 8'h63 == new_ptr_39_value ? ghv_99 : _GEN_4714; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4716 = 8'h64 == new_ptr_39_value ? ghv_100 : _GEN_4715; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4717 = 8'h65 == new_ptr_39_value ? ghv_101 : _GEN_4716; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4718 = 8'h66 == new_ptr_39_value ? ghv_102 : _GEN_4717; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4719 = 8'h67 == new_ptr_39_value ? ghv_103 : _GEN_4718; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4720 = 8'h68 == new_ptr_39_value ? ghv_104 : _GEN_4719; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4721 = 8'h69 == new_ptr_39_value ? ghv_105 : _GEN_4720; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4722 = 8'h6a == new_ptr_39_value ? ghv_106 : _GEN_4721; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4723 = 8'h6b == new_ptr_39_value ? ghv_107 : _GEN_4722; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4724 = 8'h6c == new_ptr_39_value ? ghv_108 : _GEN_4723; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4725 = 8'h6d == new_ptr_39_value ? ghv_109 : _GEN_4724; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4726 = 8'h6e == new_ptr_39_value ? ghv_110 : _GEN_4725; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4727 = 8'h6f == new_ptr_39_value ? ghv_111 : _GEN_4726; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4728 = 8'h70 == new_ptr_39_value ? ghv_112 : _GEN_4727; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4729 = 8'h71 == new_ptr_39_value ? ghv_113 : _GEN_4728; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4730 = 8'h72 == new_ptr_39_value ? ghv_114 : _GEN_4729; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4731 = 8'h73 == new_ptr_39_value ? ghv_115 : _GEN_4730; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4732 = 8'h74 == new_ptr_39_value ? ghv_116 : _GEN_4731; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4733 = 8'h75 == new_ptr_39_value ? ghv_117 : _GEN_4732; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4734 = 8'h76 == new_ptr_39_value ? ghv_118 : _GEN_4733; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4735 = 8'h77 == new_ptr_39_value ? ghv_119 : _GEN_4734; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4736 = 8'h78 == new_ptr_39_value ? ghv_120 : _GEN_4735; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4737 = 8'h79 == new_ptr_39_value ? ghv_121 : _GEN_4736; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4738 = 8'h7a == new_ptr_39_value ? ghv_122 : _GEN_4737; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4739 = 8'h7b == new_ptr_39_value ? ghv_123 : _GEN_4738; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4740 = 8'h7c == new_ptr_39_value ? ghv_124 : _GEN_4739; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4741 = 8'h7d == new_ptr_39_value ? ghv_125 : _GEN_4740; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4742 = 8'h7e == new_ptr_39_value ? ghv_126 : _GEN_4741; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4743 = 8'h7f == new_ptr_39_value ? ghv_127 : _GEN_4742; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4744 = 8'h80 == new_ptr_39_value ? ghv_128 : _GEN_4743; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4745 = 8'h81 == new_ptr_39_value ? ghv_129 : _GEN_4744; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4746 = 8'h82 == new_ptr_39_value ? ghv_130 : _GEN_4745; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4747 = 8'h83 == new_ptr_39_value ? ghv_131 : _GEN_4746; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4748 = 8'h84 == new_ptr_39_value ? ghv_132 : _GEN_4747; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4749 = 8'h85 == new_ptr_39_value ? ghv_133 : _GEN_4748; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4750 = 8'h86 == new_ptr_39_value ? ghv_134 : _GEN_4749; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4751 = 8'h87 == new_ptr_39_value ? ghv_135 : _GEN_4750; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4752 = 8'h88 == new_ptr_39_value ? ghv_136 : _GEN_4751; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4753 = 8'h89 == new_ptr_39_value ? ghv_137 : _GEN_4752; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4754 = 8'h8a == new_ptr_39_value ? ghv_138 : _GEN_4753; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4755 = 8'h8b == new_ptr_39_value ? ghv_139 : _GEN_4754; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4756 = 8'h8c == new_ptr_39_value ? ghv_140 : _GEN_4755; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4757 = 8'h8d == new_ptr_39_value ? ghv_141 : _GEN_4756; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4758 = 8'h8e == new_ptr_39_value ? ghv_142 : _GEN_4757; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_23_value = _new_ptr_value_T_47[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_4761 = 8'h1 == new_ptr_23_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4762 = 8'h2 == new_ptr_23_value ? ghv_2 : _GEN_4761; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4763 = 8'h3 == new_ptr_23_value ? ghv_3 : _GEN_4762; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4764 = 8'h4 == new_ptr_23_value ? ghv_4 : _GEN_4763; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4765 = 8'h5 == new_ptr_23_value ? ghv_5 : _GEN_4764; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4766 = 8'h6 == new_ptr_23_value ? ghv_6 : _GEN_4765; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4767 = 8'h7 == new_ptr_23_value ? ghv_7 : _GEN_4766; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4768 = 8'h8 == new_ptr_23_value ? ghv_8 : _GEN_4767; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4769 = 8'h9 == new_ptr_23_value ? ghv_9 : _GEN_4768; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4770 = 8'ha == new_ptr_23_value ? ghv_10 : _GEN_4769; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4771 = 8'hb == new_ptr_23_value ? ghv_11 : _GEN_4770; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4772 = 8'hc == new_ptr_23_value ? ghv_12 : _GEN_4771; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4773 = 8'hd == new_ptr_23_value ? ghv_13 : _GEN_4772; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4774 = 8'he == new_ptr_23_value ? ghv_14 : _GEN_4773; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4775 = 8'hf == new_ptr_23_value ? ghv_15 : _GEN_4774; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4776 = 8'h10 == new_ptr_23_value ? ghv_16 : _GEN_4775; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4777 = 8'h11 == new_ptr_23_value ? ghv_17 : _GEN_4776; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4778 = 8'h12 == new_ptr_23_value ? ghv_18 : _GEN_4777; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4779 = 8'h13 == new_ptr_23_value ? ghv_19 : _GEN_4778; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4780 = 8'h14 == new_ptr_23_value ? ghv_20 : _GEN_4779; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4781 = 8'h15 == new_ptr_23_value ? ghv_21 : _GEN_4780; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4782 = 8'h16 == new_ptr_23_value ? ghv_22 : _GEN_4781; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4783 = 8'h17 == new_ptr_23_value ? ghv_23 : _GEN_4782; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4784 = 8'h18 == new_ptr_23_value ? ghv_24 : _GEN_4783; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4785 = 8'h19 == new_ptr_23_value ? ghv_25 : _GEN_4784; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4786 = 8'h1a == new_ptr_23_value ? ghv_26 : _GEN_4785; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4787 = 8'h1b == new_ptr_23_value ? ghv_27 : _GEN_4786; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4788 = 8'h1c == new_ptr_23_value ? ghv_28 : _GEN_4787; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4789 = 8'h1d == new_ptr_23_value ? ghv_29 : _GEN_4788; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4790 = 8'h1e == new_ptr_23_value ? ghv_30 : _GEN_4789; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4791 = 8'h1f == new_ptr_23_value ? ghv_31 : _GEN_4790; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4792 = 8'h20 == new_ptr_23_value ? ghv_32 : _GEN_4791; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4793 = 8'h21 == new_ptr_23_value ? ghv_33 : _GEN_4792; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4794 = 8'h22 == new_ptr_23_value ? ghv_34 : _GEN_4793; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4795 = 8'h23 == new_ptr_23_value ? ghv_35 : _GEN_4794; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4796 = 8'h24 == new_ptr_23_value ? ghv_36 : _GEN_4795; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4797 = 8'h25 == new_ptr_23_value ? ghv_37 : _GEN_4796; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4798 = 8'h26 == new_ptr_23_value ? ghv_38 : _GEN_4797; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4799 = 8'h27 == new_ptr_23_value ? ghv_39 : _GEN_4798; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4800 = 8'h28 == new_ptr_23_value ? ghv_40 : _GEN_4799; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4801 = 8'h29 == new_ptr_23_value ? ghv_41 : _GEN_4800; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4802 = 8'h2a == new_ptr_23_value ? ghv_42 : _GEN_4801; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4803 = 8'h2b == new_ptr_23_value ? ghv_43 : _GEN_4802; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4804 = 8'h2c == new_ptr_23_value ? ghv_44 : _GEN_4803; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4805 = 8'h2d == new_ptr_23_value ? ghv_45 : _GEN_4804; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4806 = 8'h2e == new_ptr_23_value ? ghv_46 : _GEN_4805; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4807 = 8'h2f == new_ptr_23_value ? ghv_47 : _GEN_4806; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4808 = 8'h30 == new_ptr_23_value ? ghv_48 : _GEN_4807; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4809 = 8'h31 == new_ptr_23_value ? ghv_49 : _GEN_4808; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4810 = 8'h32 == new_ptr_23_value ? ghv_50 : _GEN_4809; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4811 = 8'h33 == new_ptr_23_value ? ghv_51 : _GEN_4810; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4812 = 8'h34 == new_ptr_23_value ? ghv_52 : _GEN_4811; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4813 = 8'h35 == new_ptr_23_value ? ghv_53 : _GEN_4812; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4814 = 8'h36 == new_ptr_23_value ? ghv_54 : _GEN_4813; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4815 = 8'h37 == new_ptr_23_value ? ghv_55 : _GEN_4814; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4816 = 8'h38 == new_ptr_23_value ? ghv_56 : _GEN_4815; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4817 = 8'h39 == new_ptr_23_value ? ghv_57 : _GEN_4816; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4818 = 8'h3a == new_ptr_23_value ? ghv_58 : _GEN_4817; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4819 = 8'h3b == new_ptr_23_value ? ghv_59 : _GEN_4818; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4820 = 8'h3c == new_ptr_23_value ? ghv_60 : _GEN_4819; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4821 = 8'h3d == new_ptr_23_value ? ghv_61 : _GEN_4820; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4822 = 8'h3e == new_ptr_23_value ? ghv_62 : _GEN_4821; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4823 = 8'h3f == new_ptr_23_value ? ghv_63 : _GEN_4822; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4824 = 8'h40 == new_ptr_23_value ? ghv_64 : _GEN_4823; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4825 = 8'h41 == new_ptr_23_value ? ghv_65 : _GEN_4824; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4826 = 8'h42 == new_ptr_23_value ? ghv_66 : _GEN_4825; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4827 = 8'h43 == new_ptr_23_value ? ghv_67 : _GEN_4826; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4828 = 8'h44 == new_ptr_23_value ? ghv_68 : _GEN_4827; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4829 = 8'h45 == new_ptr_23_value ? ghv_69 : _GEN_4828; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4830 = 8'h46 == new_ptr_23_value ? ghv_70 : _GEN_4829; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4831 = 8'h47 == new_ptr_23_value ? ghv_71 : _GEN_4830; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4832 = 8'h48 == new_ptr_23_value ? ghv_72 : _GEN_4831; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4833 = 8'h49 == new_ptr_23_value ? ghv_73 : _GEN_4832; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4834 = 8'h4a == new_ptr_23_value ? ghv_74 : _GEN_4833; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4835 = 8'h4b == new_ptr_23_value ? ghv_75 : _GEN_4834; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4836 = 8'h4c == new_ptr_23_value ? ghv_76 : _GEN_4835; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4837 = 8'h4d == new_ptr_23_value ? ghv_77 : _GEN_4836; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4838 = 8'h4e == new_ptr_23_value ? ghv_78 : _GEN_4837; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4839 = 8'h4f == new_ptr_23_value ? ghv_79 : _GEN_4838; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4840 = 8'h50 == new_ptr_23_value ? ghv_80 : _GEN_4839; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4841 = 8'h51 == new_ptr_23_value ? ghv_81 : _GEN_4840; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4842 = 8'h52 == new_ptr_23_value ? ghv_82 : _GEN_4841; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4843 = 8'h53 == new_ptr_23_value ? ghv_83 : _GEN_4842; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4844 = 8'h54 == new_ptr_23_value ? ghv_84 : _GEN_4843; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4845 = 8'h55 == new_ptr_23_value ? ghv_85 : _GEN_4844; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4846 = 8'h56 == new_ptr_23_value ? ghv_86 : _GEN_4845; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4847 = 8'h57 == new_ptr_23_value ? ghv_87 : _GEN_4846; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4848 = 8'h58 == new_ptr_23_value ? ghv_88 : _GEN_4847; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4849 = 8'h59 == new_ptr_23_value ? ghv_89 : _GEN_4848; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4850 = 8'h5a == new_ptr_23_value ? ghv_90 : _GEN_4849; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4851 = 8'h5b == new_ptr_23_value ? ghv_91 : _GEN_4850; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4852 = 8'h5c == new_ptr_23_value ? ghv_92 : _GEN_4851; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4853 = 8'h5d == new_ptr_23_value ? ghv_93 : _GEN_4852; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4854 = 8'h5e == new_ptr_23_value ? ghv_94 : _GEN_4853; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4855 = 8'h5f == new_ptr_23_value ? ghv_95 : _GEN_4854; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4856 = 8'h60 == new_ptr_23_value ? ghv_96 : _GEN_4855; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4857 = 8'h61 == new_ptr_23_value ? ghv_97 : _GEN_4856; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4858 = 8'h62 == new_ptr_23_value ? ghv_98 : _GEN_4857; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4859 = 8'h63 == new_ptr_23_value ? ghv_99 : _GEN_4858; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4860 = 8'h64 == new_ptr_23_value ? ghv_100 : _GEN_4859; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4861 = 8'h65 == new_ptr_23_value ? ghv_101 : _GEN_4860; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4862 = 8'h66 == new_ptr_23_value ? ghv_102 : _GEN_4861; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4863 = 8'h67 == new_ptr_23_value ? ghv_103 : _GEN_4862; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4864 = 8'h68 == new_ptr_23_value ? ghv_104 : _GEN_4863; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4865 = 8'h69 == new_ptr_23_value ? ghv_105 : _GEN_4864; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4866 = 8'h6a == new_ptr_23_value ? ghv_106 : _GEN_4865; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4867 = 8'h6b == new_ptr_23_value ? ghv_107 : _GEN_4866; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4868 = 8'h6c == new_ptr_23_value ? ghv_108 : _GEN_4867; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4869 = 8'h6d == new_ptr_23_value ? ghv_109 : _GEN_4868; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4870 = 8'h6e == new_ptr_23_value ? ghv_110 : _GEN_4869; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4871 = 8'h6f == new_ptr_23_value ? ghv_111 : _GEN_4870; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4872 = 8'h70 == new_ptr_23_value ? ghv_112 : _GEN_4871; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4873 = 8'h71 == new_ptr_23_value ? ghv_113 : _GEN_4872; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4874 = 8'h72 == new_ptr_23_value ? ghv_114 : _GEN_4873; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4875 = 8'h73 == new_ptr_23_value ? ghv_115 : _GEN_4874; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4876 = 8'h74 == new_ptr_23_value ? ghv_116 : _GEN_4875; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4877 = 8'h75 == new_ptr_23_value ? ghv_117 : _GEN_4876; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4878 = 8'h76 == new_ptr_23_value ? ghv_118 : _GEN_4877; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4879 = 8'h77 == new_ptr_23_value ? ghv_119 : _GEN_4878; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4880 = 8'h78 == new_ptr_23_value ? ghv_120 : _GEN_4879; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4881 = 8'h79 == new_ptr_23_value ? ghv_121 : _GEN_4880; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4882 = 8'h7a == new_ptr_23_value ? ghv_122 : _GEN_4881; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4883 = 8'h7b == new_ptr_23_value ? ghv_123 : _GEN_4882; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4884 = 8'h7c == new_ptr_23_value ? ghv_124 : _GEN_4883; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4885 = 8'h7d == new_ptr_23_value ? ghv_125 : _GEN_4884; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4886 = 8'h7e == new_ptr_23_value ? ghv_126 : _GEN_4885; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4887 = 8'h7f == new_ptr_23_value ? ghv_127 : _GEN_4886; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4888 = 8'h80 == new_ptr_23_value ? ghv_128 : _GEN_4887; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4889 = 8'h81 == new_ptr_23_value ? ghv_129 : _GEN_4888; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4890 = 8'h82 == new_ptr_23_value ? ghv_130 : _GEN_4889; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4891 = 8'h83 == new_ptr_23_value ? ghv_131 : _GEN_4890; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4892 = 8'h84 == new_ptr_23_value ? ghv_132 : _GEN_4891; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4893 = 8'h85 == new_ptr_23_value ? ghv_133 : _GEN_4892; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4894 = 8'h86 == new_ptr_23_value ? ghv_134 : _GEN_4893; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4895 = 8'h87 == new_ptr_23_value ? ghv_135 : _GEN_4894; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4896 = 8'h88 == new_ptr_23_value ? ghv_136 : _GEN_4895; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4897 = 8'h89 == new_ptr_23_value ? ghv_137 : _GEN_4896; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4898 = 8'h8a == new_ptr_23_value ? ghv_138 : _GEN_4897; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4899 = 8'h8b == new_ptr_23_value ? ghv_139 : _GEN_4898; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4900 = 8'h8c == new_ptr_23_value ? ghv_140 : _GEN_4899; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4901 = 8'h8d == new_ptr_23_value ? ghv_141 : _GEN_4900; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4902 = 8'h8e == new_ptr_23_value ? ghv_142 : _GEN_4901; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_30_value = _new_ptr_value_T_61[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_4905 = 8'h1 == new_ptr_30_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4906 = 8'h2 == new_ptr_30_value ? ghv_2 : _GEN_4905; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4907 = 8'h3 == new_ptr_30_value ? ghv_3 : _GEN_4906; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4908 = 8'h4 == new_ptr_30_value ? ghv_4 : _GEN_4907; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4909 = 8'h5 == new_ptr_30_value ? ghv_5 : _GEN_4908; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4910 = 8'h6 == new_ptr_30_value ? ghv_6 : _GEN_4909; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4911 = 8'h7 == new_ptr_30_value ? ghv_7 : _GEN_4910; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4912 = 8'h8 == new_ptr_30_value ? ghv_8 : _GEN_4911; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4913 = 8'h9 == new_ptr_30_value ? ghv_9 : _GEN_4912; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4914 = 8'ha == new_ptr_30_value ? ghv_10 : _GEN_4913; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4915 = 8'hb == new_ptr_30_value ? ghv_11 : _GEN_4914; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4916 = 8'hc == new_ptr_30_value ? ghv_12 : _GEN_4915; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4917 = 8'hd == new_ptr_30_value ? ghv_13 : _GEN_4916; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4918 = 8'he == new_ptr_30_value ? ghv_14 : _GEN_4917; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4919 = 8'hf == new_ptr_30_value ? ghv_15 : _GEN_4918; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4920 = 8'h10 == new_ptr_30_value ? ghv_16 : _GEN_4919; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4921 = 8'h11 == new_ptr_30_value ? ghv_17 : _GEN_4920; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4922 = 8'h12 == new_ptr_30_value ? ghv_18 : _GEN_4921; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4923 = 8'h13 == new_ptr_30_value ? ghv_19 : _GEN_4922; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4924 = 8'h14 == new_ptr_30_value ? ghv_20 : _GEN_4923; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4925 = 8'h15 == new_ptr_30_value ? ghv_21 : _GEN_4924; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4926 = 8'h16 == new_ptr_30_value ? ghv_22 : _GEN_4925; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4927 = 8'h17 == new_ptr_30_value ? ghv_23 : _GEN_4926; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4928 = 8'h18 == new_ptr_30_value ? ghv_24 : _GEN_4927; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4929 = 8'h19 == new_ptr_30_value ? ghv_25 : _GEN_4928; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4930 = 8'h1a == new_ptr_30_value ? ghv_26 : _GEN_4929; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4931 = 8'h1b == new_ptr_30_value ? ghv_27 : _GEN_4930; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4932 = 8'h1c == new_ptr_30_value ? ghv_28 : _GEN_4931; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4933 = 8'h1d == new_ptr_30_value ? ghv_29 : _GEN_4932; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4934 = 8'h1e == new_ptr_30_value ? ghv_30 : _GEN_4933; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4935 = 8'h1f == new_ptr_30_value ? ghv_31 : _GEN_4934; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4936 = 8'h20 == new_ptr_30_value ? ghv_32 : _GEN_4935; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4937 = 8'h21 == new_ptr_30_value ? ghv_33 : _GEN_4936; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4938 = 8'h22 == new_ptr_30_value ? ghv_34 : _GEN_4937; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4939 = 8'h23 == new_ptr_30_value ? ghv_35 : _GEN_4938; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4940 = 8'h24 == new_ptr_30_value ? ghv_36 : _GEN_4939; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4941 = 8'h25 == new_ptr_30_value ? ghv_37 : _GEN_4940; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4942 = 8'h26 == new_ptr_30_value ? ghv_38 : _GEN_4941; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4943 = 8'h27 == new_ptr_30_value ? ghv_39 : _GEN_4942; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4944 = 8'h28 == new_ptr_30_value ? ghv_40 : _GEN_4943; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4945 = 8'h29 == new_ptr_30_value ? ghv_41 : _GEN_4944; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4946 = 8'h2a == new_ptr_30_value ? ghv_42 : _GEN_4945; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4947 = 8'h2b == new_ptr_30_value ? ghv_43 : _GEN_4946; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4948 = 8'h2c == new_ptr_30_value ? ghv_44 : _GEN_4947; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4949 = 8'h2d == new_ptr_30_value ? ghv_45 : _GEN_4948; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4950 = 8'h2e == new_ptr_30_value ? ghv_46 : _GEN_4949; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4951 = 8'h2f == new_ptr_30_value ? ghv_47 : _GEN_4950; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4952 = 8'h30 == new_ptr_30_value ? ghv_48 : _GEN_4951; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4953 = 8'h31 == new_ptr_30_value ? ghv_49 : _GEN_4952; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4954 = 8'h32 == new_ptr_30_value ? ghv_50 : _GEN_4953; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4955 = 8'h33 == new_ptr_30_value ? ghv_51 : _GEN_4954; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4956 = 8'h34 == new_ptr_30_value ? ghv_52 : _GEN_4955; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4957 = 8'h35 == new_ptr_30_value ? ghv_53 : _GEN_4956; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4958 = 8'h36 == new_ptr_30_value ? ghv_54 : _GEN_4957; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4959 = 8'h37 == new_ptr_30_value ? ghv_55 : _GEN_4958; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4960 = 8'h38 == new_ptr_30_value ? ghv_56 : _GEN_4959; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4961 = 8'h39 == new_ptr_30_value ? ghv_57 : _GEN_4960; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4962 = 8'h3a == new_ptr_30_value ? ghv_58 : _GEN_4961; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4963 = 8'h3b == new_ptr_30_value ? ghv_59 : _GEN_4962; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4964 = 8'h3c == new_ptr_30_value ? ghv_60 : _GEN_4963; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4965 = 8'h3d == new_ptr_30_value ? ghv_61 : _GEN_4964; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4966 = 8'h3e == new_ptr_30_value ? ghv_62 : _GEN_4965; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4967 = 8'h3f == new_ptr_30_value ? ghv_63 : _GEN_4966; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4968 = 8'h40 == new_ptr_30_value ? ghv_64 : _GEN_4967; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4969 = 8'h41 == new_ptr_30_value ? ghv_65 : _GEN_4968; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4970 = 8'h42 == new_ptr_30_value ? ghv_66 : _GEN_4969; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4971 = 8'h43 == new_ptr_30_value ? ghv_67 : _GEN_4970; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4972 = 8'h44 == new_ptr_30_value ? ghv_68 : _GEN_4971; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4973 = 8'h45 == new_ptr_30_value ? ghv_69 : _GEN_4972; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4974 = 8'h46 == new_ptr_30_value ? ghv_70 : _GEN_4973; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4975 = 8'h47 == new_ptr_30_value ? ghv_71 : _GEN_4974; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4976 = 8'h48 == new_ptr_30_value ? ghv_72 : _GEN_4975; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4977 = 8'h49 == new_ptr_30_value ? ghv_73 : _GEN_4976; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4978 = 8'h4a == new_ptr_30_value ? ghv_74 : _GEN_4977; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4979 = 8'h4b == new_ptr_30_value ? ghv_75 : _GEN_4978; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4980 = 8'h4c == new_ptr_30_value ? ghv_76 : _GEN_4979; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4981 = 8'h4d == new_ptr_30_value ? ghv_77 : _GEN_4980; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4982 = 8'h4e == new_ptr_30_value ? ghv_78 : _GEN_4981; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4983 = 8'h4f == new_ptr_30_value ? ghv_79 : _GEN_4982; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4984 = 8'h50 == new_ptr_30_value ? ghv_80 : _GEN_4983; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4985 = 8'h51 == new_ptr_30_value ? ghv_81 : _GEN_4984; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4986 = 8'h52 == new_ptr_30_value ? ghv_82 : _GEN_4985; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4987 = 8'h53 == new_ptr_30_value ? ghv_83 : _GEN_4986; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4988 = 8'h54 == new_ptr_30_value ? ghv_84 : _GEN_4987; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4989 = 8'h55 == new_ptr_30_value ? ghv_85 : _GEN_4988; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4990 = 8'h56 == new_ptr_30_value ? ghv_86 : _GEN_4989; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4991 = 8'h57 == new_ptr_30_value ? ghv_87 : _GEN_4990; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4992 = 8'h58 == new_ptr_30_value ? ghv_88 : _GEN_4991; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4993 = 8'h59 == new_ptr_30_value ? ghv_89 : _GEN_4992; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4994 = 8'h5a == new_ptr_30_value ? ghv_90 : _GEN_4993; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4995 = 8'h5b == new_ptr_30_value ? ghv_91 : _GEN_4994; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4996 = 8'h5c == new_ptr_30_value ? ghv_92 : _GEN_4995; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4997 = 8'h5d == new_ptr_30_value ? ghv_93 : _GEN_4996; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4998 = 8'h5e == new_ptr_30_value ? ghv_94 : _GEN_4997; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_4999 = 8'h5f == new_ptr_30_value ? ghv_95 : _GEN_4998; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5000 = 8'h60 == new_ptr_30_value ? ghv_96 : _GEN_4999; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5001 = 8'h61 == new_ptr_30_value ? ghv_97 : _GEN_5000; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5002 = 8'h62 == new_ptr_30_value ? ghv_98 : _GEN_5001; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5003 = 8'h63 == new_ptr_30_value ? ghv_99 : _GEN_5002; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5004 = 8'h64 == new_ptr_30_value ? ghv_100 : _GEN_5003; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5005 = 8'h65 == new_ptr_30_value ? ghv_101 : _GEN_5004; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5006 = 8'h66 == new_ptr_30_value ? ghv_102 : _GEN_5005; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5007 = 8'h67 == new_ptr_30_value ? ghv_103 : _GEN_5006; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5008 = 8'h68 == new_ptr_30_value ? ghv_104 : _GEN_5007; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5009 = 8'h69 == new_ptr_30_value ? ghv_105 : _GEN_5008; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5010 = 8'h6a == new_ptr_30_value ? ghv_106 : _GEN_5009; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5011 = 8'h6b == new_ptr_30_value ? ghv_107 : _GEN_5010; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5012 = 8'h6c == new_ptr_30_value ? ghv_108 : _GEN_5011; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5013 = 8'h6d == new_ptr_30_value ? ghv_109 : _GEN_5012; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5014 = 8'h6e == new_ptr_30_value ? ghv_110 : _GEN_5013; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5015 = 8'h6f == new_ptr_30_value ? ghv_111 : _GEN_5014; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5016 = 8'h70 == new_ptr_30_value ? ghv_112 : _GEN_5015; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5017 = 8'h71 == new_ptr_30_value ? ghv_113 : _GEN_5016; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5018 = 8'h72 == new_ptr_30_value ? ghv_114 : _GEN_5017; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5019 = 8'h73 == new_ptr_30_value ? ghv_115 : _GEN_5018; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5020 = 8'h74 == new_ptr_30_value ? ghv_116 : _GEN_5019; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5021 = 8'h75 == new_ptr_30_value ? ghv_117 : _GEN_5020; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5022 = 8'h76 == new_ptr_30_value ? ghv_118 : _GEN_5021; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5023 = 8'h77 == new_ptr_30_value ? ghv_119 : _GEN_5022; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5024 = 8'h78 == new_ptr_30_value ? ghv_120 : _GEN_5023; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5025 = 8'h79 == new_ptr_30_value ? ghv_121 : _GEN_5024; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5026 = 8'h7a == new_ptr_30_value ? ghv_122 : _GEN_5025; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5027 = 8'h7b == new_ptr_30_value ? ghv_123 : _GEN_5026; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5028 = 8'h7c == new_ptr_30_value ? ghv_124 : _GEN_5027; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5029 = 8'h7d == new_ptr_30_value ? ghv_125 : _GEN_5028; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5030 = 8'h7e == new_ptr_30_value ? ghv_126 : _GEN_5029; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5031 = 8'h7f == new_ptr_30_value ? ghv_127 : _GEN_5030; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5032 = 8'h80 == new_ptr_30_value ? ghv_128 : _GEN_5031; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5033 = 8'h81 == new_ptr_30_value ? ghv_129 : _GEN_5032; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5034 = 8'h82 == new_ptr_30_value ? ghv_130 : _GEN_5033; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5035 = 8'h83 == new_ptr_30_value ? ghv_131 : _GEN_5034; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5036 = 8'h84 == new_ptr_30_value ? ghv_132 : _GEN_5035; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5037 = 8'h85 == new_ptr_30_value ? ghv_133 : _GEN_5036; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5038 = 8'h86 == new_ptr_30_value ? ghv_134 : _GEN_5037; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5039 = 8'h87 == new_ptr_30_value ? ghv_135 : _GEN_5038; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5040 = 8'h88 == new_ptr_30_value ? ghv_136 : _GEN_5039; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5041 = 8'h89 == new_ptr_30_value ? ghv_137 : _GEN_5040; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5042 = 8'h8a == new_ptr_30_value ? ghv_138 : _GEN_5041; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5043 = 8'h8b == new_ptr_30_value ? ghv_139 : _GEN_5042; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5044 = 8'h8c == new_ptr_30_value ? ghv_140 : _GEN_5043; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5045 = 8'h8d == new_ptr_30_value ? ghv_141 : _GEN_5044; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5046 = 8'h8e == new_ptr_30_value ? ghv_142 : _GEN_5045; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_21_value = _new_ptr_value_T_43[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_5049 = 8'h1 == new_ptr_21_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5050 = 8'h2 == new_ptr_21_value ? ghv_2 : _GEN_5049; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5051 = 8'h3 == new_ptr_21_value ? ghv_3 : _GEN_5050; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5052 = 8'h4 == new_ptr_21_value ? ghv_4 : _GEN_5051; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5053 = 8'h5 == new_ptr_21_value ? ghv_5 : _GEN_5052; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5054 = 8'h6 == new_ptr_21_value ? ghv_6 : _GEN_5053; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5055 = 8'h7 == new_ptr_21_value ? ghv_7 : _GEN_5054; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5056 = 8'h8 == new_ptr_21_value ? ghv_8 : _GEN_5055; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5057 = 8'h9 == new_ptr_21_value ? ghv_9 : _GEN_5056; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5058 = 8'ha == new_ptr_21_value ? ghv_10 : _GEN_5057; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5059 = 8'hb == new_ptr_21_value ? ghv_11 : _GEN_5058; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5060 = 8'hc == new_ptr_21_value ? ghv_12 : _GEN_5059; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5061 = 8'hd == new_ptr_21_value ? ghv_13 : _GEN_5060; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5062 = 8'he == new_ptr_21_value ? ghv_14 : _GEN_5061; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5063 = 8'hf == new_ptr_21_value ? ghv_15 : _GEN_5062; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5064 = 8'h10 == new_ptr_21_value ? ghv_16 : _GEN_5063; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5065 = 8'h11 == new_ptr_21_value ? ghv_17 : _GEN_5064; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5066 = 8'h12 == new_ptr_21_value ? ghv_18 : _GEN_5065; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5067 = 8'h13 == new_ptr_21_value ? ghv_19 : _GEN_5066; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5068 = 8'h14 == new_ptr_21_value ? ghv_20 : _GEN_5067; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5069 = 8'h15 == new_ptr_21_value ? ghv_21 : _GEN_5068; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5070 = 8'h16 == new_ptr_21_value ? ghv_22 : _GEN_5069; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5071 = 8'h17 == new_ptr_21_value ? ghv_23 : _GEN_5070; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5072 = 8'h18 == new_ptr_21_value ? ghv_24 : _GEN_5071; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5073 = 8'h19 == new_ptr_21_value ? ghv_25 : _GEN_5072; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5074 = 8'h1a == new_ptr_21_value ? ghv_26 : _GEN_5073; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5075 = 8'h1b == new_ptr_21_value ? ghv_27 : _GEN_5074; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5076 = 8'h1c == new_ptr_21_value ? ghv_28 : _GEN_5075; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5077 = 8'h1d == new_ptr_21_value ? ghv_29 : _GEN_5076; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5078 = 8'h1e == new_ptr_21_value ? ghv_30 : _GEN_5077; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5079 = 8'h1f == new_ptr_21_value ? ghv_31 : _GEN_5078; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5080 = 8'h20 == new_ptr_21_value ? ghv_32 : _GEN_5079; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5081 = 8'h21 == new_ptr_21_value ? ghv_33 : _GEN_5080; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5082 = 8'h22 == new_ptr_21_value ? ghv_34 : _GEN_5081; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5083 = 8'h23 == new_ptr_21_value ? ghv_35 : _GEN_5082; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5084 = 8'h24 == new_ptr_21_value ? ghv_36 : _GEN_5083; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5085 = 8'h25 == new_ptr_21_value ? ghv_37 : _GEN_5084; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5086 = 8'h26 == new_ptr_21_value ? ghv_38 : _GEN_5085; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5087 = 8'h27 == new_ptr_21_value ? ghv_39 : _GEN_5086; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5088 = 8'h28 == new_ptr_21_value ? ghv_40 : _GEN_5087; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5089 = 8'h29 == new_ptr_21_value ? ghv_41 : _GEN_5088; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5090 = 8'h2a == new_ptr_21_value ? ghv_42 : _GEN_5089; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5091 = 8'h2b == new_ptr_21_value ? ghv_43 : _GEN_5090; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5092 = 8'h2c == new_ptr_21_value ? ghv_44 : _GEN_5091; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5093 = 8'h2d == new_ptr_21_value ? ghv_45 : _GEN_5092; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5094 = 8'h2e == new_ptr_21_value ? ghv_46 : _GEN_5093; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5095 = 8'h2f == new_ptr_21_value ? ghv_47 : _GEN_5094; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5096 = 8'h30 == new_ptr_21_value ? ghv_48 : _GEN_5095; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5097 = 8'h31 == new_ptr_21_value ? ghv_49 : _GEN_5096; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5098 = 8'h32 == new_ptr_21_value ? ghv_50 : _GEN_5097; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5099 = 8'h33 == new_ptr_21_value ? ghv_51 : _GEN_5098; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5100 = 8'h34 == new_ptr_21_value ? ghv_52 : _GEN_5099; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5101 = 8'h35 == new_ptr_21_value ? ghv_53 : _GEN_5100; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5102 = 8'h36 == new_ptr_21_value ? ghv_54 : _GEN_5101; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5103 = 8'h37 == new_ptr_21_value ? ghv_55 : _GEN_5102; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5104 = 8'h38 == new_ptr_21_value ? ghv_56 : _GEN_5103; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5105 = 8'h39 == new_ptr_21_value ? ghv_57 : _GEN_5104; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5106 = 8'h3a == new_ptr_21_value ? ghv_58 : _GEN_5105; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5107 = 8'h3b == new_ptr_21_value ? ghv_59 : _GEN_5106; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5108 = 8'h3c == new_ptr_21_value ? ghv_60 : _GEN_5107; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5109 = 8'h3d == new_ptr_21_value ? ghv_61 : _GEN_5108; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5110 = 8'h3e == new_ptr_21_value ? ghv_62 : _GEN_5109; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5111 = 8'h3f == new_ptr_21_value ? ghv_63 : _GEN_5110; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5112 = 8'h40 == new_ptr_21_value ? ghv_64 : _GEN_5111; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5113 = 8'h41 == new_ptr_21_value ? ghv_65 : _GEN_5112; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5114 = 8'h42 == new_ptr_21_value ? ghv_66 : _GEN_5113; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5115 = 8'h43 == new_ptr_21_value ? ghv_67 : _GEN_5114; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5116 = 8'h44 == new_ptr_21_value ? ghv_68 : _GEN_5115; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5117 = 8'h45 == new_ptr_21_value ? ghv_69 : _GEN_5116; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5118 = 8'h46 == new_ptr_21_value ? ghv_70 : _GEN_5117; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5119 = 8'h47 == new_ptr_21_value ? ghv_71 : _GEN_5118; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5120 = 8'h48 == new_ptr_21_value ? ghv_72 : _GEN_5119; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5121 = 8'h49 == new_ptr_21_value ? ghv_73 : _GEN_5120; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5122 = 8'h4a == new_ptr_21_value ? ghv_74 : _GEN_5121; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5123 = 8'h4b == new_ptr_21_value ? ghv_75 : _GEN_5122; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5124 = 8'h4c == new_ptr_21_value ? ghv_76 : _GEN_5123; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5125 = 8'h4d == new_ptr_21_value ? ghv_77 : _GEN_5124; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5126 = 8'h4e == new_ptr_21_value ? ghv_78 : _GEN_5125; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5127 = 8'h4f == new_ptr_21_value ? ghv_79 : _GEN_5126; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5128 = 8'h50 == new_ptr_21_value ? ghv_80 : _GEN_5127; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5129 = 8'h51 == new_ptr_21_value ? ghv_81 : _GEN_5128; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5130 = 8'h52 == new_ptr_21_value ? ghv_82 : _GEN_5129; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5131 = 8'h53 == new_ptr_21_value ? ghv_83 : _GEN_5130; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5132 = 8'h54 == new_ptr_21_value ? ghv_84 : _GEN_5131; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5133 = 8'h55 == new_ptr_21_value ? ghv_85 : _GEN_5132; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5134 = 8'h56 == new_ptr_21_value ? ghv_86 : _GEN_5133; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5135 = 8'h57 == new_ptr_21_value ? ghv_87 : _GEN_5134; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5136 = 8'h58 == new_ptr_21_value ? ghv_88 : _GEN_5135; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5137 = 8'h59 == new_ptr_21_value ? ghv_89 : _GEN_5136; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5138 = 8'h5a == new_ptr_21_value ? ghv_90 : _GEN_5137; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5139 = 8'h5b == new_ptr_21_value ? ghv_91 : _GEN_5138; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5140 = 8'h5c == new_ptr_21_value ? ghv_92 : _GEN_5139; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5141 = 8'h5d == new_ptr_21_value ? ghv_93 : _GEN_5140; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5142 = 8'h5e == new_ptr_21_value ? ghv_94 : _GEN_5141; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5143 = 8'h5f == new_ptr_21_value ? ghv_95 : _GEN_5142; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5144 = 8'h60 == new_ptr_21_value ? ghv_96 : _GEN_5143; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5145 = 8'h61 == new_ptr_21_value ? ghv_97 : _GEN_5144; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5146 = 8'h62 == new_ptr_21_value ? ghv_98 : _GEN_5145; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5147 = 8'h63 == new_ptr_21_value ? ghv_99 : _GEN_5146; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5148 = 8'h64 == new_ptr_21_value ? ghv_100 : _GEN_5147; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5149 = 8'h65 == new_ptr_21_value ? ghv_101 : _GEN_5148; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5150 = 8'h66 == new_ptr_21_value ? ghv_102 : _GEN_5149; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5151 = 8'h67 == new_ptr_21_value ? ghv_103 : _GEN_5150; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5152 = 8'h68 == new_ptr_21_value ? ghv_104 : _GEN_5151; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5153 = 8'h69 == new_ptr_21_value ? ghv_105 : _GEN_5152; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5154 = 8'h6a == new_ptr_21_value ? ghv_106 : _GEN_5153; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5155 = 8'h6b == new_ptr_21_value ? ghv_107 : _GEN_5154; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5156 = 8'h6c == new_ptr_21_value ? ghv_108 : _GEN_5155; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5157 = 8'h6d == new_ptr_21_value ? ghv_109 : _GEN_5156; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5158 = 8'h6e == new_ptr_21_value ? ghv_110 : _GEN_5157; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5159 = 8'h6f == new_ptr_21_value ? ghv_111 : _GEN_5158; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5160 = 8'h70 == new_ptr_21_value ? ghv_112 : _GEN_5159; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5161 = 8'h71 == new_ptr_21_value ? ghv_113 : _GEN_5160; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5162 = 8'h72 == new_ptr_21_value ? ghv_114 : _GEN_5161; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5163 = 8'h73 == new_ptr_21_value ? ghv_115 : _GEN_5162; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5164 = 8'h74 == new_ptr_21_value ? ghv_116 : _GEN_5163; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5165 = 8'h75 == new_ptr_21_value ? ghv_117 : _GEN_5164; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5166 = 8'h76 == new_ptr_21_value ? ghv_118 : _GEN_5165; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5167 = 8'h77 == new_ptr_21_value ? ghv_119 : _GEN_5166; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5168 = 8'h78 == new_ptr_21_value ? ghv_120 : _GEN_5167; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5169 = 8'h79 == new_ptr_21_value ? ghv_121 : _GEN_5168; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5170 = 8'h7a == new_ptr_21_value ? ghv_122 : _GEN_5169; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5171 = 8'h7b == new_ptr_21_value ? ghv_123 : _GEN_5170; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5172 = 8'h7c == new_ptr_21_value ? ghv_124 : _GEN_5171; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5173 = 8'h7d == new_ptr_21_value ? ghv_125 : _GEN_5172; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5174 = 8'h7e == new_ptr_21_value ? ghv_126 : _GEN_5173; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5175 = 8'h7f == new_ptr_21_value ? ghv_127 : _GEN_5174; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5176 = 8'h80 == new_ptr_21_value ? ghv_128 : _GEN_5175; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5177 = 8'h81 == new_ptr_21_value ? ghv_129 : _GEN_5176; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5178 = 8'h82 == new_ptr_21_value ? ghv_130 : _GEN_5177; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5179 = 8'h83 == new_ptr_21_value ? ghv_131 : _GEN_5178; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5180 = 8'h84 == new_ptr_21_value ? ghv_132 : _GEN_5179; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5181 = 8'h85 == new_ptr_21_value ? ghv_133 : _GEN_5180; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5182 = 8'h86 == new_ptr_21_value ? ghv_134 : _GEN_5181; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5183 = 8'h87 == new_ptr_21_value ? ghv_135 : _GEN_5182; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5184 = 8'h88 == new_ptr_21_value ? ghv_136 : _GEN_5183; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5185 = 8'h89 == new_ptr_21_value ? ghv_137 : _GEN_5184; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5186 = 8'h8a == new_ptr_21_value ? ghv_138 : _GEN_5185; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5187 = 8'h8b == new_ptr_21_value ? ghv_139 : _GEN_5186; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5188 = 8'h8c == new_ptr_21_value ? ghv_140 : _GEN_5187; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5189 = 8'h8d == new_ptr_21_value ? ghv_141 : _GEN_5188; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5190 = 8'h8e == new_ptr_21_value ? ghv_142 : _GEN_5189; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_38_value = _new_ptr_value_T_77[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_5193 = 8'h1 == new_ptr_38_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5194 = 8'h2 == new_ptr_38_value ? ghv_2 : _GEN_5193; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5195 = 8'h3 == new_ptr_38_value ? ghv_3 : _GEN_5194; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5196 = 8'h4 == new_ptr_38_value ? ghv_4 : _GEN_5195; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5197 = 8'h5 == new_ptr_38_value ? ghv_5 : _GEN_5196; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5198 = 8'h6 == new_ptr_38_value ? ghv_6 : _GEN_5197; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5199 = 8'h7 == new_ptr_38_value ? ghv_7 : _GEN_5198; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5200 = 8'h8 == new_ptr_38_value ? ghv_8 : _GEN_5199; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5201 = 8'h9 == new_ptr_38_value ? ghv_9 : _GEN_5200; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5202 = 8'ha == new_ptr_38_value ? ghv_10 : _GEN_5201; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5203 = 8'hb == new_ptr_38_value ? ghv_11 : _GEN_5202; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5204 = 8'hc == new_ptr_38_value ? ghv_12 : _GEN_5203; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5205 = 8'hd == new_ptr_38_value ? ghv_13 : _GEN_5204; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5206 = 8'he == new_ptr_38_value ? ghv_14 : _GEN_5205; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5207 = 8'hf == new_ptr_38_value ? ghv_15 : _GEN_5206; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5208 = 8'h10 == new_ptr_38_value ? ghv_16 : _GEN_5207; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5209 = 8'h11 == new_ptr_38_value ? ghv_17 : _GEN_5208; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5210 = 8'h12 == new_ptr_38_value ? ghv_18 : _GEN_5209; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5211 = 8'h13 == new_ptr_38_value ? ghv_19 : _GEN_5210; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5212 = 8'h14 == new_ptr_38_value ? ghv_20 : _GEN_5211; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5213 = 8'h15 == new_ptr_38_value ? ghv_21 : _GEN_5212; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5214 = 8'h16 == new_ptr_38_value ? ghv_22 : _GEN_5213; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5215 = 8'h17 == new_ptr_38_value ? ghv_23 : _GEN_5214; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5216 = 8'h18 == new_ptr_38_value ? ghv_24 : _GEN_5215; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5217 = 8'h19 == new_ptr_38_value ? ghv_25 : _GEN_5216; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5218 = 8'h1a == new_ptr_38_value ? ghv_26 : _GEN_5217; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5219 = 8'h1b == new_ptr_38_value ? ghv_27 : _GEN_5218; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5220 = 8'h1c == new_ptr_38_value ? ghv_28 : _GEN_5219; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5221 = 8'h1d == new_ptr_38_value ? ghv_29 : _GEN_5220; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5222 = 8'h1e == new_ptr_38_value ? ghv_30 : _GEN_5221; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5223 = 8'h1f == new_ptr_38_value ? ghv_31 : _GEN_5222; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5224 = 8'h20 == new_ptr_38_value ? ghv_32 : _GEN_5223; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5225 = 8'h21 == new_ptr_38_value ? ghv_33 : _GEN_5224; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5226 = 8'h22 == new_ptr_38_value ? ghv_34 : _GEN_5225; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5227 = 8'h23 == new_ptr_38_value ? ghv_35 : _GEN_5226; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5228 = 8'h24 == new_ptr_38_value ? ghv_36 : _GEN_5227; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5229 = 8'h25 == new_ptr_38_value ? ghv_37 : _GEN_5228; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5230 = 8'h26 == new_ptr_38_value ? ghv_38 : _GEN_5229; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5231 = 8'h27 == new_ptr_38_value ? ghv_39 : _GEN_5230; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5232 = 8'h28 == new_ptr_38_value ? ghv_40 : _GEN_5231; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5233 = 8'h29 == new_ptr_38_value ? ghv_41 : _GEN_5232; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5234 = 8'h2a == new_ptr_38_value ? ghv_42 : _GEN_5233; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5235 = 8'h2b == new_ptr_38_value ? ghv_43 : _GEN_5234; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5236 = 8'h2c == new_ptr_38_value ? ghv_44 : _GEN_5235; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5237 = 8'h2d == new_ptr_38_value ? ghv_45 : _GEN_5236; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5238 = 8'h2e == new_ptr_38_value ? ghv_46 : _GEN_5237; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5239 = 8'h2f == new_ptr_38_value ? ghv_47 : _GEN_5238; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5240 = 8'h30 == new_ptr_38_value ? ghv_48 : _GEN_5239; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5241 = 8'h31 == new_ptr_38_value ? ghv_49 : _GEN_5240; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5242 = 8'h32 == new_ptr_38_value ? ghv_50 : _GEN_5241; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5243 = 8'h33 == new_ptr_38_value ? ghv_51 : _GEN_5242; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5244 = 8'h34 == new_ptr_38_value ? ghv_52 : _GEN_5243; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5245 = 8'h35 == new_ptr_38_value ? ghv_53 : _GEN_5244; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5246 = 8'h36 == new_ptr_38_value ? ghv_54 : _GEN_5245; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5247 = 8'h37 == new_ptr_38_value ? ghv_55 : _GEN_5246; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5248 = 8'h38 == new_ptr_38_value ? ghv_56 : _GEN_5247; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5249 = 8'h39 == new_ptr_38_value ? ghv_57 : _GEN_5248; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5250 = 8'h3a == new_ptr_38_value ? ghv_58 : _GEN_5249; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5251 = 8'h3b == new_ptr_38_value ? ghv_59 : _GEN_5250; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5252 = 8'h3c == new_ptr_38_value ? ghv_60 : _GEN_5251; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5253 = 8'h3d == new_ptr_38_value ? ghv_61 : _GEN_5252; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5254 = 8'h3e == new_ptr_38_value ? ghv_62 : _GEN_5253; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5255 = 8'h3f == new_ptr_38_value ? ghv_63 : _GEN_5254; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5256 = 8'h40 == new_ptr_38_value ? ghv_64 : _GEN_5255; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5257 = 8'h41 == new_ptr_38_value ? ghv_65 : _GEN_5256; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5258 = 8'h42 == new_ptr_38_value ? ghv_66 : _GEN_5257; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5259 = 8'h43 == new_ptr_38_value ? ghv_67 : _GEN_5258; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5260 = 8'h44 == new_ptr_38_value ? ghv_68 : _GEN_5259; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5261 = 8'h45 == new_ptr_38_value ? ghv_69 : _GEN_5260; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5262 = 8'h46 == new_ptr_38_value ? ghv_70 : _GEN_5261; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5263 = 8'h47 == new_ptr_38_value ? ghv_71 : _GEN_5262; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5264 = 8'h48 == new_ptr_38_value ? ghv_72 : _GEN_5263; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5265 = 8'h49 == new_ptr_38_value ? ghv_73 : _GEN_5264; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5266 = 8'h4a == new_ptr_38_value ? ghv_74 : _GEN_5265; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5267 = 8'h4b == new_ptr_38_value ? ghv_75 : _GEN_5266; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5268 = 8'h4c == new_ptr_38_value ? ghv_76 : _GEN_5267; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5269 = 8'h4d == new_ptr_38_value ? ghv_77 : _GEN_5268; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5270 = 8'h4e == new_ptr_38_value ? ghv_78 : _GEN_5269; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5271 = 8'h4f == new_ptr_38_value ? ghv_79 : _GEN_5270; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5272 = 8'h50 == new_ptr_38_value ? ghv_80 : _GEN_5271; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5273 = 8'h51 == new_ptr_38_value ? ghv_81 : _GEN_5272; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5274 = 8'h52 == new_ptr_38_value ? ghv_82 : _GEN_5273; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5275 = 8'h53 == new_ptr_38_value ? ghv_83 : _GEN_5274; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5276 = 8'h54 == new_ptr_38_value ? ghv_84 : _GEN_5275; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5277 = 8'h55 == new_ptr_38_value ? ghv_85 : _GEN_5276; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5278 = 8'h56 == new_ptr_38_value ? ghv_86 : _GEN_5277; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5279 = 8'h57 == new_ptr_38_value ? ghv_87 : _GEN_5278; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5280 = 8'h58 == new_ptr_38_value ? ghv_88 : _GEN_5279; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5281 = 8'h59 == new_ptr_38_value ? ghv_89 : _GEN_5280; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5282 = 8'h5a == new_ptr_38_value ? ghv_90 : _GEN_5281; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5283 = 8'h5b == new_ptr_38_value ? ghv_91 : _GEN_5282; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5284 = 8'h5c == new_ptr_38_value ? ghv_92 : _GEN_5283; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5285 = 8'h5d == new_ptr_38_value ? ghv_93 : _GEN_5284; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5286 = 8'h5e == new_ptr_38_value ? ghv_94 : _GEN_5285; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5287 = 8'h5f == new_ptr_38_value ? ghv_95 : _GEN_5286; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5288 = 8'h60 == new_ptr_38_value ? ghv_96 : _GEN_5287; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5289 = 8'h61 == new_ptr_38_value ? ghv_97 : _GEN_5288; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5290 = 8'h62 == new_ptr_38_value ? ghv_98 : _GEN_5289; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5291 = 8'h63 == new_ptr_38_value ? ghv_99 : _GEN_5290; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5292 = 8'h64 == new_ptr_38_value ? ghv_100 : _GEN_5291; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5293 = 8'h65 == new_ptr_38_value ? ghv_101 : _GEN_5292; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5294 = 8'h66 == new_ptr_38_value ? ghv_102 : _GEN_5293; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5295 = 8'h67 == new_ptr_38_value ? ghv_103 : _GEN_5294; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5296 = 8'h68 == new_ptr_38_value ? ghv_104 : _GEN_5295; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5297 = 8'h69 == new_ptr_38_value ? ghv_105 : _GEN_5296; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5298 = 8'h6a == new_ptr_38_value ? ghv_106 : _GEN_5297; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5299 = 8'h6b == new_ptr_38_value ? ghv_107 : _GEN_5298; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5300 = 8'h6c == new_ptr_38_value ? ghv_108 : _GEN_5299; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5301 = 8'h6d == new_ptr_38_value ? ghv_109 : _GEN_5300; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5302 = 8'h6e == new_ptr_38_value ? ghv_110 : _GEN_5301; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5303 = 8'h6f == new_ptr_38_value ? ghv_111 : _GEN_5302; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5304 = 8'h70 == new_ptr_38_value ? ghv_112 : _GEN_5303; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5305 = 8'h71 == new_ptr_38_value ? ghv_113 : _GEN_5304; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5306 = 8'h72 == new_ptr_38_value ? ghv_114 : _GEN_5305; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5307 = 8'h73 == new_ptr_38_value ? ghv_115 : _GEN_5306; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5308 = 8'h74 == new_ptr_38_value ? ghv_116 : _GEN_5307; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5309 = 8'h75 == new_ptr_38_value ? ghv_117 : _GEN_5308; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5310 = 8'h76 == new_ptr_38_value ? ghv_118 : _GEN_5309; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5311 = 8'h77 == new_ptr_38_value ? ghv_119 : _GEN_5310; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5312 = 8'h78 == new_ptr_38_value ? ghv_120 : _GEN_5311; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5313 = 8'h79 == new_ptr_38_value ? ghv_121 : _GEN_5312; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5314 = 8'h7a == new_ptr_38_value ? ghv_122 : _GEN_5313; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5315 = 8'h7b == new_ptr_38_value ? ghv_123 : _GEN_5314; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5316 = 8'h7c == new_ptr_38_value ? ghv_124 : _GEN_5315; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5317 = 8'h7d == new_ptr_38_value ? ghv_125 : _GEN_5316; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5318 = 8'h7e == new_ptr_38_value ? ghv_126 : _GEN_5317; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5319 = 8'h7f == new_ptr_38_value ? ghv_127 : _GEN_5318; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5320 = 8'h80 == new_ptr_38_value ? ghv_128 : _GEN_5319; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5321 = 8'h81 == new_ptr_38_value ? ghv_129 : _GEN_5320; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5322 = 8'h82 == new_ptr_38_value ? ghv_130 : _GEN_5321; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5323 = 8'h83 == new_ptr_38_value ? ghv_131 : _GEN_5322; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5324 = 8'h84 == new_ptr_38_value ? ghv_132 : _GEN_5323; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5325 = 8'h85 == new_ptr_38_value ? ghv_133 : _GEN_5324; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5326 = 8'h86 == new_ptr_38_value ? ghv_134 : _GEN_5325; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5327 = 8'h87 == new_ptr_38_value ? ghv_135 : _GEN_5326; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5328 = 8'h88 == new_ptr_38_value ? ghv_136 : _GEN_5327; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5329 = 8'h89 == new_ptr_38_value ? ghv_137 : _GEN_5328; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5330 = 8'h8a == new_ptr_38_value ? ghv_138 : _GEN_5329; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5331 = 8'h8b == new_ptr_38_value ? ghv_139 : _GEN_5330; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5332 = 8'h8c == new_ptr_38_value ? ghv_140 : _GEN_5331; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5333 = 8'h8d == new_ptr_38_value ? ghv_141 : _GEN_5332; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5334 = 8'h8e == new_ptr_38_value ? ghv_142 : _GEN_5333; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_31_value = _new_ptr_value_T_63[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_5337 = 8'h1 == new_ptr_31_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5338 = 8'h2 == new_ptr_31_value ? ghv_2 : _GEN_5337; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5339 = 8'h3 == new_ptr_31_value ? ghv_3 : _GEN_5338; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5340 = 8'h4 == new_ptr_31_value ? ghv_4 : _GEN_5339; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5341 = 8'h5 == new_ptr_31_value ? ghv_5 : _GEN_5340; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5342 = 8'h6 == new_ptr_31_value ? ghv_6 : _GEN_5341; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5343 = 8'h7 == new_ptr_31_value ? ghv_7 : _GEN_5342; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5344 = 8'h8 == new_ptr_31_value ? ghv_8 : _GEN_5343; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5345 = 8'h9 == new_ptr_31_value ? ghv_9 : _GEN_5344; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5346 = 8'ha == new_ptr_31_value ? ghv_10 : _GEN_5345; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5347 = 8'hb == new_ptr_31_value ? ghv_11 : _GEN_5346; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5348 = 8'hc == new_ptr_31_value ? ghv_12 : _GEN_5347; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5349 = 8'hd == new_ptr_31_value ? ghv_13 : _GEN_5348; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5350 = 8'he == new_ptr_31_value ? ghv_14 : _GEN_5349; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5351 = 8'hf == new_ptr_31_value ? ghv_15 : _GEN_5350; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5352 = 8'h10 == new_ptr_31_value ? ghv_16 : _GEN_5351; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5353 = 8'h11 == new_ptr_31_value ? ghv_17 : _GEN_5352; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5354 = 8'h12 == new_ptr_31_value ? ghv_18 : _GEN_5353; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5355 = 8'h13 == new_ptr_31_value ? ghv_19 : _GEN_5354; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5356 = 8'h14 == new_ptr_31_value ? ghv_20 : _GEN_5355; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5357 = 8'h15 == new_ptr_31_value ? ghv_21 : _GEN_5356; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5358 = 8'h16 == new_ptr_31_value ? ghv_22 : _GEN_5357; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5359 = 8'h17 == new_ptr_31_value ? ghv_23 : _GEN_5358; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5360 = 8'h18 == new_ptr_31_value ? ghv_24 : _GEN_5359; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5361 = 8'h19 == new_ptr_31_value ? ghv_25 : _GEN_5360; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5362 = 8'h1a == new_ptr_31_value ? ghv_26 : _GEN_5361; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5363 = 8'h1b == new_ptr_31_value ? ghv_27 : _GEN_5362; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5364 = 8'h1c == new_ptr_31_value ? ghv_28 : _GEN_5363; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5365 = 8'h1d == new_ptr_31_value ? ghv_29 : _GEN_5364; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5366 = 8'h1e == new_ptr_31_value ? ghv_30 : _GEN_5365; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5367 = 8'h1f == new_ptr_31_value ? ghv_31 : _GEN_5366; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5368 = 8'h20 == new_ptr_31_value ? ghv_32 : _GEN_5367; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5369 = 8'h21 == new_ptr_31_value ? ghv_33 : _GEN_5368; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5370 = 8'h22 == new_ptr_31_value ? ghv_34 : _GEN_5369; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5371 = 8'h23 == new_ptr_31_value ? ghv_35 : _GEN_5370; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5372 = 8'h24 == new_ptr_31_value ? ghv_36 : _GEN_5371; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5373 = 8'h25 == new_ptr_31_value ? ghv_37 : _GEN_5372; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5374 = 8'h26 == new_ptr_31_value ? ghv_38 : _GEN_5373; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5375 = 8'h27 == new_ptr_31_value ? ghv_39 : _GEN_5374; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5376 = 8'h28 == new_ptr_31_value ? ghv_40 : _GEN_5375; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5377 = 8'h29 == new_ptr_31_value ? ghv_41 : _GEN_5376; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5378 = 8'h2a == new_ptr_31_value ? ghv_42 : _GEN_5377; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5379 = 8'h2b == new_ptr_31_value ? ghv_43 : _GEN_5378; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5380 = 8'h2c == new_ptr_31_value ? ghv_44 : _GEN_5379; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5381 = 8'h2d == new_ptr_31_value ? ghv_45 : _GEN_5380; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5382 = 8'h2e == new_ptr_31_value ? ghv_46 : _GEN_5381; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5383 = 8'h2f == new_ptr_31_value ? ghv_47 : _GEN_5382; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5384 = 8'h30 == new_ptr_31_value ? ghv_48 : _GEN_5383; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5385 = 8'h31 == new_ptr_31_value ? ghv_49 : _GEN_5384; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5386 = 8'h32 == new_ptr_31_value ? ghv_50 : _GEN_5385; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5387 = 8'h33 == new_ptr_31_value ? ghv_51 : _GEN_5386; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5388 = 8'h34 == new_ptr_31_value ? ghv_52 : _GEN_5387; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5389 = 8'h35 == new_ptr_31_value ? ghv_53 : _GEN_5388; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5390 = 8'h36 == new_ptr_31_value ? ghv_54 : _GEN_5389; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5391 = 8'h37 == new_ptr_31_value ? ghv_55 : _GEN_5390; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5392 = 8'h38 == new_ptr_31_value ? ghv_56 : _GEN_5391; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5393 = 8'h39 == new_ptr_31_value ? ghv_57 : _GEN_5392; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5394 = 8'h3a == new_ptr_31_value ? ghv_58 : _GEN_5393; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5395 = 8'h3b == new_ptr_31_value ? ghv_59 : _GEN_5394; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5396 = 8'h3c == new_ptr_31_value ? ghv_60 : _GEN_5395; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5397 = 8'h3d == new_ptr_31_value ? ghv_61 : _GEN_5396; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5398 = 8'h3e == new_ptr_31_value ? ghv_62 : _GEN_5397; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5399 = 8'h3f == new_ptr_31_value ? ghv_63 : _GEN_5398; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5400 = 8'h40 == new_ptr_31_value ? ghv_64 : _GEN_5399; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5401 = 8'h41 == new_ptr_31_value ? ghv_65 : _GEN_5400; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5402 = 8'h42 == new_ptr_31_value ? ghv_66 : _GEN_5401; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5403 = 8'h43 == new_ptr_31_value ? ghv_67 : _GEN_5402; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5404 = 8'h44 == new_ptr_31_value ? ghv_68 : _GEN_5403; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5405 = 8'h45 == new_ptr_31_value ? ghv_69 : _GEN_5404; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5406 = 8'h46 == new_ptr_31_value ? ghv_70 : _GEN_5405; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5407 = 8'h47 == new_ptr_31_value ? ghv_71 : _GEN_5406; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5408 = 8'h48 == new_ptr_31_value ? ghv_72 : _GEN_5407; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5409 = 8'h49 == new_ptr_31_value ? ghv_73 : _GEN_5408; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5410 = 8'h4a == new_ptr_31_value ? ghv_74 : _GEN_5409; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5411 = 8'h4b == new_ptr_31_value ? ghv_75 : _GEN_5410; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5412 = 8'h4c == new_ptr_31_value ? ghv_76 : _GEN_5411; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5413 = 8'h4d == new_ptr_31_value ? ghv_77 : _GEN_5412; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5414 = 8'h4e == new_ptr_31_value ? ghv_78 : _GEN_5413; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5415 = 8'h4f == new_ptr_31_value ? ghv_79 : _GEN_5414; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5416 = 8'h50 == new_ptr_31_value ? ghv_80 : _GEN_5415; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5417 = 8'h51 == new_ptr_31_value ? ghv_81 : _GEN_5416; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5418 = 8'h52 == new_ptr_31_value ? ghv_82 : _GEN_5417; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5419 = 8'h53 == new_ptr_31_value ? ghv_83 : _GEN_5418; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5420 = 8'h54 == new_ptr_31_value ? ghv_84 : _GEN_5419; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5421 = 8'h55 == new_ptr_31_value ? ghv_85 : _GEN_5420; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5422 = 8'h56 == new_ptr_31_value ? ghv_86 : _GEN_5421; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5423 = 8'h57 == new_ptr_31_value ? ghv_87 : _GEN_5422; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5424 = 8'h58 == new_ptr_31_value ? ghv_88 : _GEN_5423; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5425 = 8'h59 == new_ptr_31_value ? ghv_89 : _GEN_5424; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5426 = 8'h5a == new_ptr_31_value ? ghv_90 : _GEN_5425; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5427 = 8'h5b == new_ptr_31_value ? ghv_91 : _GEN_5426; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5428 = 8'h5c == new_ptr_31_value ? ghv_92 : _GEN_5427; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5429 = 8'h5d == new_ptr_31_value ? ghv_93 : _GEN_5428; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5430 = 8'h5e == new_ptr_31_value ? ghv_94 : _GEN_5429; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5431 = 8'h5f == new_ptr_31_value ? ghv_95 : _GEN_5430; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5432 = 8'h60 == new_ptr_31_value ? ghv_96 : _GEN_5431; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5433 = 8'h61 == new_ptr_31_value ? ghv_97 : _GEN_5432; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5434 = 8'h62 == new_ptr_31_value ? ghv_98 : _GEN_5433; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5435 = 8'h63 == new_ptr_31_value ? ghv_99 : _GEN_5434; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5436 = 8'h64 == new_ptr_31_value ? ghv_100 : _GEN_5435; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5437 = 8'h65 == new_ptr_31_value ? ghv_101 : _GEN_5436; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5438 = 8'h66 == new_ptr_31_value ? ghv_102 : _GEN_5437; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5439 = 8'h67 == new_ptr_31_value ? ghv_103 : _GEN_5438; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5440 = 8'h68 == new_ptr_31_value ? ghv_104 : _GEN_5439; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5441 = 8'h69 == new_ptr_31_value ? ghv_105 : _GEN_5440; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5442 = 8'h6a == new_ptr_31_value ? ghv_106 : _GEN_5441; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5443 = 8'h6b == new_ptr_31_value ? ghv_107 : _GEN_5442; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5444 = 8'h6c == new_ptr_31_value ? ghv_108 : _GEN_5443; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5445 = 8'h6d == new_ptr_31_value ? ghv_109 : _GEN_5444; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5446 = 8'h6e == new_ptr_31_value ? ghv_110 : _GEN_5445; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5447 = 8'h6f == new_ptr_31_value ? ghv_111 : _GEN_5446; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5448 = 8'h70 == new_ptr_31_value ? ghv_112 : _GEN_5447; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5449 = 8'h71 == new_ptr_31_value ? ghv_113 : _GEN_5448; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5450 = 8'h72 == new_ptr_31_value ? ghv_114 : _GEN_5449; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5451 = 8'h73 == new_ptr_31_value ? ghv_115 : _GEN_5450; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5452 = 8'h74 == new_ptr_31_value ? ghv_116 : _GEN_5451; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5453 = 8'h75 == new_ptr_31_value ? ghv_117 : _GEN_5452; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5454 = 8'h76 == new_ptr_31_value ? ghv_118 : _GEN_5453; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5455 = 8'h77 == new_ptr_31_value ? ghv_119 : _GEN_5454; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5456 = 8'h78 == new_ptr_31_value ? ghv_120 : _GEN_5455; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5457 = 8'h79 == new_ptr_31_value ? ghv_121 : _GEN_5456; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5458 = 8'h7a == new_ptr_31_value ? ghv_122 : _GEN_5457; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5459 = 8'h7b == new_ptr_31_value ? ghv_123 : _GEN_5458; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5460 = 8'h7c == new_ptr_31_value ? ghv_124 : _GEN_5459; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5461 = 8'h7d == new_ptr_31_value ? ghv_125 : _GEN_5460; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5462 = 8'h7e == new_ptr_31_value ? ghv_126 : _GEN_5461; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5463 = 8'h7f == new_ptr_31_value ? ghv_127 : _GEN_5462; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5464 = 8'h80 == new_ptr_31_value ? ghv_128 : _GEN_5463; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5465 = 8'h81 == new_ptr_31_value ? ghv_129 : _GEN_5464; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5466 = 8'h82 == new_ptr_31_value ? ghv_130 : _GEN_5465; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5467 = 8'h83 == new_ptr_31_value ? ghv_131 : _GEN_5466; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5468 = 8'h84 == new_ptr_31_value ? ghv_132 : _GEN_5467; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5469 = 8'h85 == new_ptr_31_value ? ghv_133 : _GEN_5468; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5470 = 8'h86 == new_ptr_31_value ? ghv_134 : _GEN_5469; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5471 = 8'h87 == new_ptr_31_value ? ghv_135 : _GEN_5470; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5472 = 8'h88 == new_ptr_31_value ? ghv_136 : _GEN_5471; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5473 = 8'h89 == new_ptr_31_value ? ghv_137 : _GEN_5472; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5474 = 8'h8a == new_ptr_31_value ? ghv_138 : _GEN_5473; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5475 = 8'h8b == new_ptr_31_value ? ghv_139 : _GEN_5474; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5476 = 8'h8c == new_ptr_31_value ? ghv_140 : _GEN_5475; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5477 = 8'h8d == new_ptr_31_value ? ghv_141 : _GEN_5476; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5478 = 8'h8e == new_ptr_31_value ? ghv_142 : _GEN_5477; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_27_value = _new_ptr_value_T_55[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_5481 = 8'h1 == new_ptr_27_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5482 = 8'h2 == new_ptr_27_value ? ghv_2 : _GEN_5481; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5483 = 8'h3 == new_ptr_27_value ? ghv_3 : _GEN_5482; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5484 = 8'h4 == new_ptr_27_value ? ghv_4 : _GEN_5483; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5485 = 8'h5 == new_ptr_27_value ? ghv_5 : _GEN_5484; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5486 = 8'h6 == new_ptr_27_value ? ghv_6 : _GEN_5485; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5487 = 8'h7 == new_ptr_27_value ? ghv_7 : _GEN_5486; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5488 = 8'h8 == new_ptr_27_value ? ghv_8 : _GEN_5487; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5489 = 8'h9 == new_ptr_27_value ? ghv_9 : _GEN_5488; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5490 = 8'ha == new_ptr_27_value ? ghv_10 : _GEN_5489; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5491 = 8'hb == new_ptr_27_value ? ghv_11 : _GEN_5490; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5492 = 8'hc == new_ptr_27_value ? ghv_12 : _GEN_5491; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5493 = 8'hd == new_ptr_27_value ? ghv_13 : _GEN_5492; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5494 = 8'he == new_ptr_27_value ? ghv_14 : _GEN_5493; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5495 = 8'hf == new_ptr_27_value ? ghv_15 : _GEN_5494; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5496 = 8'h10 == new_ptr_27_value ? ghv_16 : _GEN_5495; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5497 = 8'h11 == new_ptr_27_value ? ghv_17 : _GEN_5496; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5498 = 8'h12 == new_ptr_27_value ? ghv_18 : _GEN_5497; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5499 = 8'h13 == new_ptr_27_value ? ghv_19 : _GEN_5498; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5500 = 8'h14 == new_ptr_27_value ? ghv_20 : _GEN_5499; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5501 = 8'h15 == new_ptr_27_value ? ghv_21 : _GEN_5500; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5502 = 8'h16 == new_ptr_27_value ? ghv_22 : _GEN_5501; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5503 = 8'h17 == new_ptr_27_value ? ghv_23 : _GEN_5502; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5504 = 8'h18 == new_ptr_27_value ? ghv_24 : _GEN_5503; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5505 = 8'h19 == new_ptr_27_value ? ghv_25 : _GEN_5504; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5506 = 8'h1a == new_ptr_27_value ? ghv_26 : _GEN_5505; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5507 = 8'h1b == new_ptr_27_value ? ghv_27 : _GEN_5506; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5508 = 8'h1c == new_ptr_27_value ? ghv_28 : _GEN_5507; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5509 = 8'h1d == new_ptr_27_value ? ghv_29 : _GEN_5508; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5510 = 8'h1e == new_ptr_27_value ? ghv_30 : _GEN_5509; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5511 = 8'h1f == new_ptr_27_value ? ghv_31 : _GEN_5510; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5512 = 8'h20 == new_ptr_27_value ? ghv_32 : _GEN_5511; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5513 = 8'h21 == new_ptr_27_value ? ghv_33 : _GEN_5512; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5514 = 8'h22 == new_ptr_27_value ? ghv_34 : _GEN_5513; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5515 = 8'h23 == new_ptr_27_value ? ghv_35 : _GEN_5514; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5516 = 8'h24 == new_ptr_27_value ? ghv_36 : _GEN_5515; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5517 = 8'h25 == new_ptr_27_value ? ghv_37 : _GEN_5516; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5518 = 8'h26 == new_ptr_27_value ? ghv_38 : _GEN_5517; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5519 = 8'h27 == new_ptr_27_value ? ghv_39 : _GEN_5518; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5520 = 8'h28 == new_ptr_27_value ? ghv_40 : _GEN_5519; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5521 = 8'h29 == new_ptr_27_value ? ghv_41 : _GEN_5520; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5522 = 8'h2a == new_ptr_27_value ? ghv_42 : _GEN_5521; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5523 = 8'h2b == new_ptr_27_value ? ghv_43 : _GEN_5522; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5524 = 8'h2c == new_ptr_27_value ? ghv_44 : _GEN_5523; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5525 = 8'h2d == new_ptr_27_value ? ghv_45 : _GEN_5524; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5526 = 8'h2e == new_ptr_27_value ? ghv_46 : _GEN_5525; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5527 = 8'h2f == new_ptr_27_value ? ghv_47 : _GEN_5526; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5528 = 8'h30 == new_ptr_27_value ? ghv_48 : _GEN_5527; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5529 = 8'h31 == new_ptr_27_value ? ghv_49 : _GEN_5528; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5530 = 8'h32 == new_ptr_27_value ? ghv_50 : _GEN_5529; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5531 = 8'h33 == new_ptr_27_value ? ghv_51 : _GEN_5530; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5532 = 8'h34 == new_ptr_27_value ? ghv_52 : _GEN_5531; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5533 = 8'h35 == new_ptr_27_value ? ghv_53 : _GEN_5532; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5534 = 8'h36 == new_ptr_27_value ? ghv_54 : _GEN_5533; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5535 = 8'h37 == new_ptr_27_value ? ghv_55 : _GEN_5534; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5536 = 8'h38 == new_ptr_27_value ? ghv_56 : _GEN_5535; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5537 = 8'h39 == new_ptr_27_value ? ghv_57 : _GEN_5536; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5538 = 8'h3a == new_ptr_27_value ? ghv_58 : _GEN_5537; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5539 = 8'h3b == new_ptr_27_value ? ghv_59 : _GEN_5538; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5540 = 8'h3c == new_ptr_27_value ? ghv_60 : _GEN_5539; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5541 = 8'h3d == new_ptr_27_value ? ghv_61 : _GEN_5540; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5542 = 8'h3e == new_ptr_27_value ? ghv_62 : _GEN_5541; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5543 = 8'h3f == new_ptr_27_value ? ghv_63 : _GEN_5542; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5544 = 8'h40 == new_ptr_27_value ? ghv_64 : _GEN_5543; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5545 = 8'h41 == new_ptr_27_value ? ghv_65 : _GEN_5544; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5546 = 8'h42 == new_ptr_27_value ? ghv_66 : _GEN_5545; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5547 = 8'h43 == new_ptr_27_value ? ghv_67 : _GEN_5546; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5548 = 8'h44 == new_ptr_27_value ? ghv_68 : _GEN_5547; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5549 = 8'h45 == new_ptr_27_value ? ghv_69 : _GEN_5548; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5550 = 8'h46 == new_ptr_27_value ? ghv_70 : _GEN_5549; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5551 = 8'h47 == new_ptr_27_value ? ghv_71 : _GEN_5550; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5552 = 8'h48 == new_ptr_27_value ? ghv_72 : _GEN_5551; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5553 = 8'h49 == new_ptr_27_value ? ghv_73 : _GEN_5552; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5554 = 8'h4a == new_ptr_27_value ? ghv_74 : _GEN_5553; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5555 = 8'h4b == new_ptr_27_value ? ghv_75 : _GEN_5554; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5556 = 8'h4c == new_ptr_27_value ? ghv_76 : _GEN_5555; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5557 = 8'h4d == new_ptr_27_value ? ghv_77 : _GEN_5556; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5558 = 8'h4e == new_ptr_27_value ? ghv_78 : _GEN_5557; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5559 = 8'h4f == new_ptr_27_value ? ghv_79 : _GEN_5558; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5560 = 8'h50 == new_ptr_27_value ? ghv_80 : _GEN_5559; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5561 = 8'h51 == new_ptr_27_value ? ghv_81 : _GEN_5560; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5562 = 8'h52 == new_ptr_27_value ? ghv_82 : _GEN_5561; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5563 = 8'h53 == new_ptr_27_value ? ghv_83 : _GEN_5562; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5564 = 8'h54 == new_ptr_27_value ? ghv_84 : _GEN_5563; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5565 = 8'h55 == new_ptr_27_value ? ghv_85 : _GEN_5564; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5566 = 8'h56 == new_ptr_27_value ? ghv_86 : _GEN_5565; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5567 = 8'h57 == new_ptr_27_value ? ghv_87 : _GEN_5566; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5568 = 8'h58 == new_ptr_27_value ? ghv_88 : _GEN_5567; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5569 = 8'h59 == new_ptr_27_value ? ghv_89 : _GEN_5568; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5570 = 8'h5a == new_ptr_27_value ? ghv_90 : _GEN_5569; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5571 = 8'h5b == new_ptr_27_value ? ghv_91 : _GEN_5570; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5572 = 8'h5c == new_ptr_27_value ? ghv_92 : _GEN_5571; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5573 = 8'h5d == new_ptr_27_value ? ghv_93 : _GEN_5572; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5574 = 8'h5e == new_ptr_27_value ? ghv_94 : _GEN_5573; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5575 = 8'h5f == new_ptr_27_value ? ghv_95 : _GEN_5574; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5576 = 8'h60 == new_ptr_27_value ? ghv_96 : _GEN_5575; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5577 = 8'h61 == new_ptr_27_value ? ghv_97 : _GEN_5576; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5578 = 8'h62 == new_ptr_27_value ? ghv_98 : _GEN_5577; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5579 = 8'h63 == new_ptr_27_value ? ghv_99 : _GEN_5578; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5580 = 8'h64 == new_ptr_27_value ? ghv_100 : _GEN_5579; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5581 = 8'h65 == new_ptr_27_value ? ghv_101 : _GEN_5580; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5582 = 8'h66 == new_ptr_27_value ? ghv_102 : _GEN_5581; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5583 = 8'h67 == new_ptr_27_value ? ghv_103 : _GEN_5582; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5584 = 8'h68 == new_ptr_27_value ? ghv_104 : _GEN_5583; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5585 = 8'h69 == new_ptr_27_value ? ghv_105 : _GEN_5584; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5586 = 8'h6a == new_ptr_27_value ? ghv_106 : _GEN_5585; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5587 = 8'h6b == new_ptr_27_value ? ghv_107 : _GEN_5586; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5588 = 8'h6c == new_ptr_27_value ? ghv_108 : _GEN_5587; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5589 = 8'h6d == new_ptr_27_value ? ghv_109 : _GEN_5588; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5590 = 8'h6e == new_ptr_27_value ? ghv_110 : _GEN_5589; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5591 = 8'h6f == new_ptr_27_value ? ghv_111 : _GEN_5590; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5592 = 8'h70 == new_ptr_27_value ? ghv_112 : _GEN_5591; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5593 = 8'h71 == new_ptr_27_value ? ghv_113 : _GEN_5592; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5594 = 8'h72 == new_ptr_27_value ? ghv_114 : _GEN_5593; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5595 = 8'h73 == new_ptr_27_value ? ghv_115 : _GEN_5594; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5596 = 8'h74 == new_ptr_27_value ? ghv_116 : _GEN_5595; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5597 = 8'h75 == new_ptr_27_value ? ghv_117 : _GEN_5596; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5598 = 8'h76 == new_ptr_27_value ? ghv_118 : _GEN_5597; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5599 = 8'h77 == new_ptr_27_value ? ghv_119 : _GEN_5598; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5600 = 8'h78 == new_ptr_27_value ? ghv_120 : _GEN_5599; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5601 = 8'h79 == new_ptr_27_value ? ghv_121 : _GEN_5600; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5602 = 8'h7a == new_ptr_27_value ? ghv_122 : _GEN_5601; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5603 = 8'h7b == new_ptr_27_value ? ghv_123 : _GEN_5602; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5604 = 8'h7c == new_ptr_27_value ? ghv_124 : _GEN_5603; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5605 = 8'h7d == new_ptr_27_value ? ghv_125 : _GEN_5604; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5606 = 8'h7e == new_ptr_27_value ? ghv_126 : _GEN_5605; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5607 = 8'h7f == new_ptr_27_value ? ghv_127 : _GEN_5606; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5608 = 8'h80 == new_ptr_27_value ? ghv_128 : _GEN_5607; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5609 = 8'h81 == new_ptr_27_value ? ghv_129 : _GEN_5608; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5610 = 8'h82 == new_ptr_27_value ? ghv_130 : _GEN_5609; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5611 = 8'h83 == new_ptr_27_value ? ghv_131 : _GEN_5610; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5612 = 8'h84 == new_ptr_27_value ? ghv_132 : _GEN_5611; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5613 = 8'h85 == new_ptr_27_value ? ghv_133 : _GEN_5612; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5614 = 8'h86 == new_ptr_27_value ? ghv_134 : _GEN_5613; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5615 = 8'h87 == new_ptr_27_value ? ghv_135 : _GEN_5614; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5616 = 8'h88 == new_ptr_27_value ? ghv_136 : _GEN_5615; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5617 = 8'h89 == new_ptr_27_value ? ghv_137 : _GEN_5616; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5618 = 8'h8a == new_ptr_27_value ? ghv_138 : _GEN_5617; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5619 = 8'h8b == new_ptr_27_value ? ghv_139 : _GEN_5618; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5620 = 8'h8c == new_ptr_27_value ? ghv_140 : _GEN_5619; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5621 = 8'h8d == new_ptr_27_value ? ghv_141 : _GEN_5620; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5622 = 8'h8e == new_ptr_27_value ? ghv_142 : _GEN_5621; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_25_value = _new_ptr_value_T_51[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_5625 = 8'h1 == new_ptr_25_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5626 = 8'h2 == new_ptr_25_value ? ghv_2 : _GEN_5625; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5627 = 8'h3 == new_ptr_25_value ? ghv_3 : _GEN_5626; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5628 = 8'h4 == new_ptr_25_value ? ghv_4 : _GEN_5627; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5629 = 8'h5 == new_ptr_25_value ? ghv_5 : _GEN_5628; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5630 = 8'h6 == new_ptr_25_value ? ghv_6 : _GEN_5629; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5631 = 8'h7 == new_ptr_25_value ? ghv_7 : _GEN_5630; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5632 = 8'h8 == new_ptr_25_value ? ghv_8 : _GEN_5631; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5633 = 8'h9 == new_ptr_25_value ? ghv_9 : _GEN_5632; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5634 = 8'ha == new_ptr_25_value ? ghv_10 : _GEN_5633; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5635 = 8'hb == new_ptr_25_value ? ghv_11 : _GEN_5634; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5636 = 8'hc == new_ptr_25_value ? ghv_12 : _GEN_5635; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5637 = 8'hd == new_ptr_25_value ? ghv_13 : _GEN_5636; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5638 = 8'he == new_ptr_25_value ? ghv_14 : _GEN_5637; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5639 = 8'hf == new_ptr_25_value ? ghv_15 : _GEN_5638; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5640 = 8'h10 == new_ptr_25_value ? ghv_16 : _GEN_5639; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5641 = 8'h11 == new_ptr_25_value ? ghv_17 : _GEN_5640; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5642 = 8'h12 == new_ptr_25_value ? ghv_18 : _GEN_5641; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5643 = 8'h13 == new_ptr_25_value ? ghv_19 : _GEN_5642; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5644 = 8'h14 == new_ptr_25_value ? ghv_20 : _GEN_5643; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5645 = 8'h15 == new_ptr_25_value ? ghv_21 : _GEN_5644; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5646 = 8'h16 == new_ptr_25_value ? ghv_22 : _GEN_5645; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5647 = 8'h17 == new_ptr_25_value ? ghv_23 : _GEN_5646; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5648 = 8'h18 == new_ptr_25_value ? ghv_24 : _GEN_5647; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5649 = 8'h19 == new_ptr_25_value ? ghv_25 : _GEN_5648; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5650 = 8'h1a == new_ptr_25_value ? ghv_26 : _GEN_5649; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5651 = 8'h1b == new_ptr_25_value ? ghv_27 : _GEN_5650; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5652 = 8'h1c == new_ptr_25_value ? ghv_28 : _GEN_5651; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5653 = 8'h1d == new_ptr_25_value ? ghv_29 : _GEN_5652; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5654 = 8'h1e == new_ptr_25_value ? ghv_30 : _GEN_5653; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5655 = 8'h1f == new_ptr_25_value ? ghv_31 : _GEN_5654; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5656 = 8'h20 == new_ptr_25_value ? ghv_32 : _GEN_5655; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5657 = 8'h21 == new_ptr_25_value ? ghv_33 : _GEN_5656; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5658 = 8'h22 == new_ptr_25_value ? ghv_34 : _GEN_5657; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5659 = 8'h23 == new_ptr_25_value ? ghv_35 : _GEN_5658; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5660 = 8'h24 == new_ptr_25_value ? ghv_36 : _GEN_5659; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5661 = 8'h25 == new_ptr_25_value ? ghv_37 : _GEN_5660; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5662 = 8'h26 == new_ptr_25_value ? ghv_38 : _GEN_5661; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5663 = 8'h27 == new_ptr_25_value ? ghv_39 : _GEN_5662; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5664 = 8'h28 == new_ptr_25_value ? ghv_40 : _GEN_5663; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5665 = 8'h29 == new_ptr_25_value ? ghv_41 : _GEN_5664; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5666 = 8'h2a == new_ptr_25_value ? ghv_42 : _GEN_5665; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5667 = 8'h2b == new_ptr_25_value ? ghv_43 : _GEN_5666; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5668 = 8'h2c == new_ptr_25_value ? ghv_44 : _GEN_5667; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5669 = 8'h2d == new_ptr_25_value ? ghv_45 : _GEN_5668; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5670 = 8'h2e == new_ptr_25_value ? ghv_46 : _GEN_5669; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5671 = 8'h2f == new_ptr_25_value ? ghv_47 : _GEN_5670; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5672 = 8'h30 == new_ptr_25_value ? ghv_48 : _GEN_5671; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5673 = 8'h31 == new_ptr_25_value ? ghv_49 : _GEN_5672; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5674 = 8'h32 == new_ptr_25_value ? ghv_50 : _GEN_5673; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5675 = 8'h33 == new_ptr_25_value ? ghv_51 : _GEN_5674; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5676 = 8'h34 == new_ptr_25_value ? ghv_52 : _GEN_5675; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5677 = 8'h35 == new_ptr_25_value ? ghv_53 : _GEN_5676; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5678 = 8'h36 == new_ptr_25_value ? ghv_54 : _GEN_5677; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5679 = 8'h37 == new_ptr_25_value ? ghv_55 : _GEN_5678; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5680 = 8'h38 == new_ptr_25_value ? ghv_56 : _GEN_5679; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5681 = 8'h39 == new_ptr_25_value ? ghv_57 : _GEN_5680; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5682 = 8'h3a == new_ptr_25_value ? ghv_58 : _GEN_5681; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5683 = 8'h3b == new_ptr_25_value ? ghv_59 : _GEN_5682; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5684 = 8'h3c == new_ptr_25_value ? ghv_60 : _GEN_5683; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5685 = 8'h3d == new_ptr_25_value ? ghv_61 : _GEN_5684; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5686 = 8'h3e == new_ptr_25_value ? ghv_62 : _GEN_5685; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5687 = 8'h3f == new_ptr_25_value ? ghv_63 : _GEN_5686; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5688 = 8'h40 == new_ptr_25_value ? ghv_64 : _GEN_5687; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5689 = 8'h41 == new_ptr_25_value ? ghv_65 : _GEN_5688; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5690 = 8'h42 == new_ptr_25_value ? ghv_66 : _GEN_5689; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5691 = 8'h43 == new_ptr_25_value ? ghv_67 : _GEN_5690; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5692 = 8'h44 == new_ptr_25_value ? ghv_68 : _GEN_5691; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5693 = 8'h45 == new_ptr_25_value ? ghv_69 : _GEN_5692; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5694 = 8'h46 == new_ptr_25_value ? ghv_70 : _GEN_5693; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5695 = 8'h47 == new_ptr_25_value ? ghv_71 : _GEN_5694; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5696 = 8'h48 == new_ptr_25_value ? ghv_72 : _GEN_5695; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5697 = 8'h49 == new_ptr_25_value ? ghv_73 : _GEN_5696; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5698 = 8'h4a == new_ptr_25_value ? ghv_74 : _GEN_5697; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5699 = 8'h4b == new_ptr_25_value ? ghv_75 : _GEN_5698; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5700 = 8'h4c == new_ptr_25_value ? ghv_76 : _GEN_5699; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5701 = 8'h4d == new_ptr_25_value ? ghv_77 : _GEN_5700; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5702 = 8'h4e == new_ptr_25_value ? ghv_78 : _GEN_5701; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5703 = 8'h4f == new_ptr_25_value ? ghv_79 : _GEN_5702; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5704 = 8'h50 == new_ptr_25_value ? ghv_80 : _GEN_5703; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5705 = 8'h51 == new_ptr_25_value ? ghv_81 : _GEN_5704; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5706 = 8'h52 == new_ptr_25_value ? ghv_82 : _GEN_5705; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5707 = 8'h53 == new_ptr_25_value ? ghv_83 : _GEN_5706; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5708 = 8'h54 == new_ptr_25_value ? ghv_84 : _GEN_5707; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5709 = 8'h55 == new_ptr_25_value ? ghv_85 : _GEN_5708; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5710 = 8'h56 == new_ptr_25_value ? ghv_86 : _GEN_5709; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5711 = 8'h57 == new_ptr_25_value ? ghv_87 : _GEN_5710; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5712 = 8'h58 == new_ptr_25_value ? ghv_88 : _GEN_5711; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5713 = 8'h59 == new_ptr_25_value ? ghv_89 : _GEN_5712; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5714 = 8'h5a == new_ptr_25_value ? ghv_90 : _GEN_5713; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5715 = 8'h5b == new_ptr_25_value ? ghv_91 : _GEN_5714; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5716 = 8'h5c == new_ptr_25_value ? ghv_92 : _GEN_5715; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5717 = 8'h5d == new_ptr_25_value ? ghv_93 : _GEN_5716; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5718 = 8'h5e == new_ptr_25_value ? ghv_94 : _GEN_5717; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5719 = 8'h5f == new_ptr_25_value ? ghv_95 : _GEN_5718; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5720 = 8'h60 == new_ptr_25_value ? ghv_96 : _GEN_5719; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5721 = 8'h61 == new_ptr_25_value ? ghv_97 : _GEN_5720; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5722 = 8'h62 == new_ptr_25_value ? ghv_98 : _GEN_5721; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5723 = 8'h63 == new_ptr_25_value ? ghv_99 : _GEN_5722; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5724 = 8'h64 == new_ptr_25_value ? ghv_100 : _GEN_5723; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5725 = 8'h65 == new_ptr_25_value ? ghv_101 : _GEN_5724; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5726 = 8'h66 == new_ptr_25_value ? ghv_102 : _GEN_5725; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5727 = 8'h67 == new_ptr_25_value ? ghv_103 : _GEN_5726; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5728 = 8'h68 == new_ptr_25_value ? ghv_104 : _GEN_5727; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5729 = 8'h69 == new_ptr_25_value ? ghv_105 : _GEN_5728; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5730 = 8'h6a == new_ptr_25_value ? ghv_106 : _GEN_5729; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5731 = 8'h6b == new_ptr_25_value ? ghv_107 : _GEN_5730; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5732 = 8'h6c == new_ptr_25_value ? ghv_108 : _GEN_5731; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5733 = 8'h6d == new_ptr_25_value ? ghv_109 : _GEN_5732; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5734 = 8'h6e == new_ptr_25_value ? ghv_110 : _GEN_5733; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5735 = 8'h6f == new_ptr_25_value ? ghv_111 : _GEN_5734; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5736 = 8'h70 == new_ptr_25_value ? ghv_112 : _GEN_5735; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5737 = 8'h71 == new_ptr_25_value ? ghv_113 : _GEN_5736; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5738 = 8'h72 == new_ptr_25_value ? ghv_114 : _GEN_5737; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5739 = 8'h73 == new_ptr_25_value ? ghv_115 : _GEN_5738; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5740 = 8'h74 == new_ptr_25_value ? ghv_116 : _GEN_5739; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5741 = 8'h75 == new_ptr_25_value ? ghv_117 : _GEN_5740; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5742 = 8'h76 == new_ptr_25_value ? ghv_118 : _GEN_5741; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5743 = 8'h77 == new_ptr_25_value ? ghv_119 : _GEN_5742; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5744 = 8'h78 == new_ptr_25_value ? ghv_120 : _GEN_5743; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5745 = 8'h79 == new_ptr_25_value ? ghv_121 : _GEN_5744; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5746 = 8'h7a == new_ptr_25_value ? ghv_122 : _GEN_5745; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5747 = 8'h7b == new_ptr_25_value ? ghv_123 : _GEN_5746; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5748 = 8'h7c == new_ptr_25_value ? ghv_124 : _GEN_5747; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5749 = 8'h7d == new_ptr_25_value ? ghv_125 : _GEN_5748; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5750 = 8'h7e == new_ptr_25_value ? ghv_126 : _GEN_5749; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5751 = 8'h7f == new_ptr_25_value ? ghv_127 : _GEN_5750; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5752 = 8'h80 == new_ptr_25_value ? ghv_128 : _GEN_5751; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5753 = 8'h81 == new_ptr_25_value ? ghv_129 : _GEN_5752; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5754 = 8'h82 == new_ptr_25_value ? ghv_130 : _GEN_5753; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5755 = 8'h83 == new_ptr_25_value ? ghv_131 : _GEN_5754; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5756 = 8'h84 == new_ptr_25_value ? ghv_132 : _GEN_5755; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5757 = 8'h85 == new_ptr_25_value ? ghv_133 : _GEN_5756; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5758 = 8'h86 == new_ptr_25_value ? ghv_134 : _GEN_5757; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5759 = 8'h87 == new_ptr_25_value ? ghv_135 : _GEN_5758; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5760 = 8'h88 == new_ptr_25_value ? ghv_136 : _GEN_5759; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5761 = 8'h89 == new_ptr_25_value ? ghv_137 : _GEN_5760; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5762 = 8'h8a == new_ptr_25_value ? ghv_138 : _GEN_5761; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5763 = 8'h8b == new_ptr_25_value ? ghv_139 : _GEN_5762; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5764 = 8'h8c == new_ptr_25_value ? ghv_140 : _GEN_5763; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5765 = 8'h8d == new_ptr_25_value ? ghv_141 : _GEN_5764; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5766 = 8'h8e == new_ptr_25_value ? ghv_142 : _GEN_5765; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_20_value = _new_ptr_value_T_41[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_5769 = 8'h1 == new_ptr_20_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5770 = 8'h2 == new_ptr_20_value ? ghv_2 : _GEN_5769; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5771 = 8'h3 == new_ptr_20_value ? ghv_3 : _GEN_5770; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5772 = 8'h4 == new_ptr_20_value ? ghv_4 : _GEN_5771; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5773 = 8'h5 == new_ptr_20_value ? ghv_5 : _GEN_5772; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5774 = 8'h6 == new_ptr_20_value ? ghv_6 : _GEN_5773; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5775 = 8'h7 == new_ptr_20_value ? ghv_7 : _GEN_5774; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5776 = 8'h8 == new_ptr_20_value ? ghv_8 : _GEN_5775; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5777 = 8'h9 == new_ptr_20_value ? ghv_9 : _GEN_5776; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5778 = 8'ha == new_ptr_20_value ? ghv_10 : _GEN_5777; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5779 = 8'hb == new_ptr_20_value ? ghv_11 : _GEN_5778; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5780 = 8'hc == new_ptr_20_value ? ghv_12 : _GEN_5779; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5781 = 8'hd == new_ptr_20_value ? ghv_13 : _GEN_5780; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5782 = 8'he == new_ptr_20_value ? ghv_14 : _GEN_5781; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5783 = 8'hf == new_ptr_20_value ? ghv_15 : _GEN_5782; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5784 = 8'h10 == new_ptr_20_value ? ghv_16 : _GEN_5783; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5785 = 8'h11 == new_ptr_20_value ? ghv_17 : _GEN_5784; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5786 = 8'h12 == new_ptr_20_value ? ghv_18 : _GEN_5785; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5787 = 8'h13 == new_ptr_20_value ? ghv_19 : _GEN_5786; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5788 = 8'h14 == new_ptr_20_value ? ghv_20 : _GEN_5787; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5789 = 8'h15 == new_ptr_20_value ? ghv_21 : _GEN_5788; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5790 = 8'h16 == new_ptr_20_value ? ghv_22 : _GEN_5789; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5791 = 8'h17 == new_ptr_20_value ? ghv_23 : _GEN_5790; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5792 = 8'h18 == new_ptr_20_value ? ghv_24 : _GEN_5791; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5793 = 8'h19 == new_ptr_20_value ? ghv_25 : _GEN_5792; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5794 = 8'h1a == new_ptr_20_value ? ghv_26 : _GEN_5793; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5795 = 8'h1b == new_ptr_20_value ? ghv_27 : _GEN_5794; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5796 = 8'h1c == new_ptr_20_value ? ghv_28 : _GEN_5795; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5797 = 8'h1d == new_ptr_20_value ? ghv_29 : _GEN_5796; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5798 = 8'h1e == new_ptr_20_value ? ghv_30 : _GEN_5797; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5799 = 8'h1f == new_ptr_20_value ? ghv_31 : _GEN_5798; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5800 = 8'h20 == new_ptr_20_value ? ghv_32 : _GEN_5799; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5801 = 8'h21 == new_ptr_20_value ? ghv_33 : _GEN_5800; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5802 = 8'h22 == new_ptr_20_value ? ghv_34 : _GEN_5801; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5803 = 8'h23 == new_ptr_20_value ? ghv_35 : _GEN_5802; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5804 = 8'h24 == new_ptr_20_value ? ghv_36 : _GEN_5803; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5805 = 8'h25 == new_ptr_20_value ? ghv_37 : _GEN_5804; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5806 = 8'h26 == new_ptr_20_value ? ghv_38 : _GEN_5805; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5807 = 8'h27 == new_ptr_20_value ? ghv_39 : _GEN_5806; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5808 = 8'h28 == new_ptr_20_value ? ghv_40 : _GEN_5807; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5809 = 8'h29 == new_ptr_20_value ? ghv_41 : _GEN_5808; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5810 = 8'h2a == new_ptr_20_value ? ghv_42 : _GEN_5809; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5811 = 8'h2b == new_ptr_20_value ? ghv_43 : _GEN_5810; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5812 = 8'h2c == new_ptr_20_value ? ghv_44 : _GEN_5811; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5813 = 8'h2d == new_ptr_20_value ? ghv_45 : _GEN_5812; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5814 = 8'h2e == new_ptr_20_value ? ghv_46 : _GEN_5813; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5815 = 8'h2f == new_ptr_20_value ? ghv_47 : _GEN_5814; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5816 = 8'h30 == new_ptr_20_value ? ghv_48 : _GEN_5815; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5817 = 8'h31 == new_ptr_20_value ? ghv_49 : _GEN_5816; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5818 = 8'h32 == new_ptr_20_value ? ghv_50 : _GEN_5817; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5819 = 8'h33 == new_ptr_20_value ? ghv_51 : _GEN_5818; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5820 = 8'h34 == new_ptr_20_value ? ghv_52 : _GEN_5819; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5821 = 8'h35 == new_ptr_20_value ? ghv_53 : _GEN_5820; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5822 = 8'h36 == new_ptr_20_value ? ghv_54 : _GEN_5821; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5823 = 8'h37 == new_ptr_20_value ? ghv_55 : _GEN_5822; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5824 = 8'h38 == new_ptr_20_value ? ghv_56 : _GEN_5823; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5825 = 8'h39 == new_ptr_20_value ? ghv_57 : _GEN_5824; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5826 = 8'h3a == new_ptr_20_value ? ghv_58 : _GEN_5825; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5827 = 8'h3b == new_ptr_20_value ? ghv_59 : _GEN_5826; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5828 = 8'h3c == new_ptr_20_value ? ghv_60 : _GEN_5827; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5829 = 8'h3d == new_ptr_20_value ? ghv_61 : _GEN_5828; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5830 = 8'h3e == new_ptr_20_value ? ghv_62 : _GEN_5829; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5831 = 8'h3f == new_ptr_20_value ? ghv_63 : _GEN_5830; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5832 = 8'h40 == new_ptr_20_value ? ghv_64 : _GEN_5831; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5833 = 8'h41 == new_ptr_20_value ? ghv_65 : _GEN_5832; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5834 = 8'h42 == new_ptr_20_value ? ghv_66 : _GEN_5833; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5835 = 8'h43 == new_ptr_20_value ? ghv_67 : _GEN_5834; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5836 = 8'h44 == new_ptr_20_value ? ghv_68 : _GEN_5835; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5837 = 8'h45 == new_ptr_20_value ? ghv_69 : _GEN_5836; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5838 = 8'h46 == new_ptr_20_value ? ghv_70 : _GEN_5837; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5839 = 8'h47 == new_ptr_20_value ? ghv_71 : _GEN_5838; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5840 = 8'h48 == new_ptr_20_value ? ghv_72 : _GEN_5839; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5841 = 8'h49 == new_ptr_20_value ? ghv_73 : _GEN_5840; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5842 = 8'h4a == new_ptr_20_value ? ghv_74 : _GEN_5841; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5843 = 8'h4b == new_ptr_20_value ? ghv_75 : _GEN_5842; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5844 = 8'h4c == new_ptr_20_value ? ghv_76 : _GEN_5843; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5845 = 8'h4d == new_ptr_20_value ? ghv_77 : _GEN_5844; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5846 = 8'h4e == new_ptr_20_value ? ghv_78 : _GEN_5845; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5847 = 8'h4f == new_ptr_20_value ? ghv_79 : _GEN_5846; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5848 = 8'h50 == new_ptr_20_value ? ghv_80 : _GEN_5847; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5849 = 8'h51 == new_ptr_20_value ? ghv_81 : _GEN_5848; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5850 = 8'h52 == new_ptr_20_value ? ghv_82 : _GEN_5849; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5851 = 8'h53 == new_ptr_20_value ? ghv_83 : _GEN_5850; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5852 = 8'h54 == new_ptr_20_value ? ghv_84 : _GEN_5851; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5853 = 8'h55 == new_ptr_20_value ? ghv_85 : _GEN_5852; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5854 = 8'h56 == new_ptr_20_value ? ghv_86 : _GEN_5853; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5855 = 8'h57 == new_ptr_20_value ? ghv_87 : _GEN_5854; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5856 = 8'h58 == new_ptr_20_value ? ghv_88 : _GEN_5855; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5857 = 8'h59 == new_ptr_20_value ? ghv_89 : _GEN_5856; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5858 = 8'h5a == new_ptr_20_value ? ghv_90 : _GEN_5857; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5859 = 8'h5b == new_ptr_20_value ? ghv_91 : _GEN_5858; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5860 = 8'h5c == new_ptr_20_value ? ghv_92 : _GEN_5859; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5861 = 8'h5d == new_ptr_20_value ? ghv_93 : _GEN_5860; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5862 = 8'h5e == new_ptr_20_value ? ghv_94 : _GEN_5861; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5863 = 8'h5f == new_ptr_20_value ? ghv_95 : _GEN_5862; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5864 = 8'h60 == new_ptr_20_value ? ghv_96 : _GEN_5863; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5865 = 8'h61 == new_ptr_20_value ? ghv_97 : _GEN_5864; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5866 = 8'h62 == new_ptr_20_value ? ghv_98 : _GEN_5865; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5867 = 8'h63 == new_ptr_20_value ? ghv_99 : _GEN_5866; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5868 = 8'h64 == new_ptr_20_value ? ghv_100 : _GEN_5867; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5869 = 8'h65 == new_ptr_20_value ? ghv_101 : _GEN_5868; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5870 = 8'h66 == new_ptr_20_value ? ghv_102 : _GEN_5869; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5871 = 8'h67 == new_ptr_20_value ? ghv_103 : _GEN_5870; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5872 = 8'h68 == new_ptr_20_value ? ghv_104 : _GEN_5871; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5873 = 8'h69 == new_ptr_20_value ? ghv_105 : _GEN_5872; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5874 = 8'h6a == new_ptr_20_value ? ghv_106 : _GEN_5873; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5875 = 8'h6b == new_ptr_20_value ? ghv_107 : _GEN_5874; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5876 = 8'h6c == new_ptr_20_value ? ghv_108 : _GEN_5875; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5877 = 8'h6d == new_ptr_20_value ? ghv_109 : _GEN_5876; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5878 = 8'h6e == new_ptr_20_value ? ghv_110 : _GEN_5877; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5879 = 8'h6f == new_ptr_20_value ? ghv_111 : _GEN_5878; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5880 = 8'h70 == new_ptr_20_value ? ghv_112 : _GEN_5879; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5881 = 8'h71 == new_ptr_20_value ? ghv_113 : _GEN_5880; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5882 = 8'h72 == new_ptr_20_value ? ghv_114 : _GEN_5881; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5883 = 8'h73 == new_ptr_20_value ? ghv_115 : _GEN_5882; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5884 = 8'h74 == new_ptr_20_value ? ghv_116 : _GEN_5883; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5885 = 8'h75 == new_ptr_20_value ? ghv_117 : _GEN_5884; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5886 = 8'h76 == new_ptr_20_value ? ghv_118 : _GEN_5885; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5887 = 8'h77 == new_ptr_20_value ? ghv_119 : _GEN_5886; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5888 = 8'h78 == new_ptr_20_value ? ghv_120 : _GEN_5887; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5889 = 8'h79 == new_ptr_20_value ? ghv_121 : _GEN_5888; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5890 = 8'h7a == new_ptr_20_value ? ghv_122 : _GEN_5889; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5891 = 8'h7b == new_ptr_20_value ? ghv_123 : _GEN_5890; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5892 = 8'h7c == new_ptr_20_value ? ghv_124 : _GEN_5891; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5893 = 8'h7d == new_ptr_20_value ? ghv_125 : _GEN_5892; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5894 = 8'h7e == new_ptr_20_value ? ghv_126 : _GEN_5893; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5895 = 8'h7f == new_ptr_20_value ? ghv_127 : _GEN_5894; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5896 = 8'h80 == new_ptr_20_value ? ghv_128 : _GEN_5895; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5897 = 8'h81 == new_ptr_20_value ? ghv_129 : _GEN_5896; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5898 = 8'h82 == new_ptr_20_value ? ghv_130 : _GEN_5897; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5899 = 8'h83 == new_ptr_20_value ? ghv_131 : _GEN_5898; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5900 = 8'h84 == new_ptr_20_value ? ghv_132 : _GEN_5899; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5901 = 8'h85 == new_ptr_20_value ? ghv_133 : _GEN_5900; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5902 = 8'h86 == new_ptr_20_value ? ghv_134 : _GEN_5901; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5903 = 8'h87 == new_ptr_20_value ? ghv_135 : _GEN_5902; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5904 = 8'h88 == new_ptr_20_value ? ghv_136 : _GEN_5903; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5905 = 8'h89 == new_ptr_20_value ? ghv_137 : _GEN_5904; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5906 = 8'h8a == new_ptr_20_value ? ghv_138 : _GEN_5905; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5907 = 8'h8b == new_ptr_20_value ? ghv_139 : _GEN_5906; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5908 = 8'h8c == new_ptr_20_value ? ghv_140 : _GEN_5907; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5909 = 8'h8d == new_ptr_20_value ? ghv_141 : _GEN_5908; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5910 = 8'h8e == new_ptr_20_value ? ghv_142 : _GEN_5909; // @[FrontendBundle.scala 329:{20,20}]
  wire  _s2_ghv_wens_T_26 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_0_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_53 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_1_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_0_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_1_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_80 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_1_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_1_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_1_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_107 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_3_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_1_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_3_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_134 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_3_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_2_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_3_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_161 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_5_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_2_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_5_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_188 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_5_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_3_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_5_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_215 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_7_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_3_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_7_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_242 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_7_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_4_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_7_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_269 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_9_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_4_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_9_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_296 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_9_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_5_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_9_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_323 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_11_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_5_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_11_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_350 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_11_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
    ; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_6_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_11_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_377 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_13_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_6_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_13_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_404 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_13_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
    ; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_7_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_13_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_431 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_15_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_7_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_15_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_458 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_15_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
    ; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_8_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_15_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_485 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_17_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_8_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_17_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_512 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_17_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
    ; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_9_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_17_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_539 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_19_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_9_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_19_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_566 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_19_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
    ; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_10_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_19_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_593 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_21_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_10_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_21_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_620 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_21_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
    ; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_11_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_21_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_647 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_23_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_11_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_23_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_674 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_23_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
    ; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_12_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_23_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_701 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_25_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_12_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_25_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_728 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_25_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
    ; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_13_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_25_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_755 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_27_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_13_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_27_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_782 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_27_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
    ; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_14_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_27_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_809 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_29_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_14_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_29_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_836 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_29_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
    ; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_15_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_29_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_863 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_31_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_15_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_31_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_890 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_31_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
    ; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_16_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_31_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_917 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_33_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_16_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_33_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_944 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_33_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
    ; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_17_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_33_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_971 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_35_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_17_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_35_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_998 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_35_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
    ; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_18_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_35_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_1025 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_37_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_18_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_37_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_1052 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_37_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_19_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_37_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_1079 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_39_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_19_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_39_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_1106 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_39_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_20_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_39_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_1133 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_41_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_20_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_41_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_1160 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_41_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_21_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_41_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_1187 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_43_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_21_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_43_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_1214 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_43_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_22_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_43_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_1241 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_45_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_22_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_45_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_1268 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_45_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_23_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_45_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_1295 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_47_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_23_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_47_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_1322 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_47_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_24_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_47_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_1349 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_49_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_24_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_49_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_1376 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_49_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_25_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_49_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_1403 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_51_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_25_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_51_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_1430 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_51_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_26_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_51_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_1457 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_53_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_26_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_53_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_1484 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_53_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_27_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_53_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_1511 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_55_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_27_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_55_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_1538 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_55_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_28_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_55_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_1565 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_57_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_28_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_57_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_1592 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_57_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_29_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_57_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_1619 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_59_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_29_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_59_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_1646 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_59_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_30_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_59_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_1673 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_61_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_30_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_61_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_1700 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_61_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_31_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_61_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_1727 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_63_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_31_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_63_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_1754 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_63_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_32_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_63_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_1781 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_65_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_32_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_65_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_1808 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_65_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_33_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_65_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_1835 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_67_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_33_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_67_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_1862 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_67_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_34_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_67_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_1889 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_69_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_34_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_69_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_1916 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_69_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_35_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_69_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_1943 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_71_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_35_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_71_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_1970 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_71_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_36_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_71_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_1997 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_73_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_36_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_73_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_2024 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_73_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_37_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_73_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_2051 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_75_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_37_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_75_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_2078 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_75_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_38_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_75_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_2105 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_77_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_38_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_77_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_2132 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_77_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_39_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_77_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_2159 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_79_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_39_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_79_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_2186 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_79_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_40_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_79_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_2213 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_81_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_40_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_81_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_2240 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_81_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_41_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_81_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_2267 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_83_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_41_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_83_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_2294 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_83_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_42_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_83_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_2321 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_85_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_42_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_85_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_2348 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_85_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_43_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_85_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_2375 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_87_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_43_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_87_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_2402 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_87_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_44_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_87_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_2429 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_89_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_44_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_89_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_2456 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_89_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_45_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_89_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_2483 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_91_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_45_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_91_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_2510 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_91_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_46_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_91_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_2537 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_93_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_46_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_93_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_2564 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_93_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_47_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_93_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_2591 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_95_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_47_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_95_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_2618 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_95_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_48_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_95_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_2645 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_97_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_48_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_97_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_2672 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_97_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_49_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_97_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_2699 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_99_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_49_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_99_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_2726 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_99_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_50_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_99_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_2753 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_101_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_50_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_101_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_2780 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_101_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_51_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_101_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_2807 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_103_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_51_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_103_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_2834 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_103_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_52_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_103_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_2861 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_105_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_52_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_105_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_2888 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_105_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_53_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_105_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_2915 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_107_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_53_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_107_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_2942 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_107_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_54_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_107_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_2969 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_109_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_54_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_109_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_2996 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_109_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_55_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_109_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_3023 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_111_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_55_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_111_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_3050 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_111_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_56_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_111_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_3077 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_113_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_56_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_113_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_3104 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_113_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_57_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_113_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_3131 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_115_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_57_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_115_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_3158 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_115_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_58_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_115_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_3185 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_117_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_58_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_117_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_3212 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_117_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_59_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_117_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_3239 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_119_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_59_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_119_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_3266 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_119_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_60_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_119_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_3293 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_121_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_60_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_121_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_3320 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_121_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_61_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_121_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_3347 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_123_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_61_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_123_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_3374 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_123_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_62_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_123_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_3401 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_125_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_62_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_125_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_3428 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_125_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_63_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_125_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_3455 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_127_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_63_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_127_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_3482 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_127_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_64_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_127_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_3509 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_129_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_64_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_129_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_3536 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_129_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_65_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_129_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_3563 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_131_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_65_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_131_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_3590 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_131_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_66_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_131_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_3617 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_133_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_66_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_133_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_3644 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_133_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_67_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_133_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_3671 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_135_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_67_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_135_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_3698 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_135_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_68_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_135_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_3725 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_137_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_68_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_137_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_3752 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_137_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_69_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_137_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_3779 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_139_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_69_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_139_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_3806 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_139_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_70_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_139_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_3833 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_141_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_70_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_141_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_3860 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_141_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_71_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_141_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_3887 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_143_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_71_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_143_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_3914 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_143_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_72_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_143_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_3941 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_145_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_72_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_145_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_3968 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_145_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_73_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_145_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_3995 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_147_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_73_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_147_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_4022 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_147_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_74_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_147_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_4049 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_149_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_74_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_149_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_4076 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_149_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_75_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_149_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_4103 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_151_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_75_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_151_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_4130 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_151_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_76_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_151_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_4157 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_153_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_76_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_153_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_4184 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_153_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_77_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_153_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_4211 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_155_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_77_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_155_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_4238 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_155_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_78_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_155_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_4265 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_157_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_78_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_157_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_4292 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_157_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_79_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_157_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_4319 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_159_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_79_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_159_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_4346 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_159_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_80_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_159_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_4373 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_161_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_80_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_161_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_4400 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_161_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_81_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_161_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_4427 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_163_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_81_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_163_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_4454 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_163_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_82_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_163_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_4481 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_165_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_82_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_165_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_4508 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_165_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_83_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_165_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_4535 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_167_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_83_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_167_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_4562 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_167_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_84_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_167_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_4589 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_169_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_84_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_169_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_4616 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_169_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_85_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_169_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_4643 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_171_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_85_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_171_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_4670 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_171_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_86_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_171_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_4697 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_173_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_86_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_173_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_4724 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_173_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_87_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_173_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_4751 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_175_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_87_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_175_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_4778 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_175_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_88_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_175_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_4805 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_177_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_88_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_177_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_4832 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_177_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_89_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_177_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_4859 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_179_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_89_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_179_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_4886 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_179_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_90_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_179_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_4913 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_181_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_90_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_181_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_4940 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_181_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_91_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_181_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_4967 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_183_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_91_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_183_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_4994 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_183_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_92_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_183_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_5021 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_185_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_92_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_185_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_5048 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_185_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_93_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_185_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_5075 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_187_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_93_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_187_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_5102 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_187_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_94_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_187_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_5129 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_189_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_94_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_189_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_5156 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_189_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_95_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_189_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_5183 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_191_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_95_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_191_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_5210 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_191_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_96_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_191_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_5237 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_193_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_96_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_193_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_5264 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_193_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_97_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_193_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_5291 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_195_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_97_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_195_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_5318 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_195_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_98_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_195_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_5345 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_197_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_98_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_197_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_5372 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_197_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_99_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_197_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_5399 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_199_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_99_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_199_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_5426 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_199_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_100_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_199_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_5453 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_201_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_100_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_201_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_5480 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_201_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_101_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_201_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_5507 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_203_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_101_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_203_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_5534 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_203_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_102_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_203_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_5561 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_205_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_102_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_205_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_5588 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_205_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_103_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_205_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_5615 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_207_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_103_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_207_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_5642 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_207_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_104_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_207_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_5669 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_209_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_104_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_209_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_5696 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_209_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_105_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_209_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_5723 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_211_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_105_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_211_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_5750 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_211_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_106_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_211_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_5777 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_213_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_106_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_213_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_5804 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_213_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_107_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_213_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_5831 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_215_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_107_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_215_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_5858 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_215_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_108_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_215_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_5885 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_217_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_108_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_217_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_5912 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_217_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_109_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_217_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_5939 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_219_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_109_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_219_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_5966 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_219_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_110_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_219_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_5993 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_221_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_110_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_221_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_6020 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_221_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_111_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_221_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_6047 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_223_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_111_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_223_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_6074 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_223_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_112_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_223_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_6101 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_225_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_112_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_225_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_6128 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_225_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_113_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_225_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_6155 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_227_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_113_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_227_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_6182 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_227_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_114_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_227_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_6209 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_229_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_114_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_229_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_6236 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_229_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_115_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_229_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_6263 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_231_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_115_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_231_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_6290 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_231_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_116_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_231_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_6317 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_233_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_116_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_233_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_6344 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_233_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_117_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_233_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_6371 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_235_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_117_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_235_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_6398 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_235_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_118_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_235_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_6425 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_237_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_118_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_237_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_6452 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_237_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_119_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_237_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_6479 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_239_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_119_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_239_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_6506 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_239_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_120_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_239_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_6533 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_241_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_120_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_241_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_6560 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_241_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_121_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_241_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_6587 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_243_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_121_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_243_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_6614 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_243_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_122_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_243_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_6641 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_245_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_122_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_245_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_6668 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_245_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_123_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_245_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_6695 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_247_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_123_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_247_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_6722 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_247_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_124_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_247_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_6749 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_249_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_124_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_249_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_6776 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_249_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_125_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_249_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_6803 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_251_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_125_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_251_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_6830 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_251_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_126_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_251_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_6857 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_253_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_126_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_253_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_6884 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_253_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_127_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_253_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_6911 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_255_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_127_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_255_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_6938 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_255_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_128_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_255_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_6965 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_257_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_128_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_257_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_6992 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_257_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_129_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_257_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_7019 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_259_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_129_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_259_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_7046 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_259_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_130_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_259_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_7073 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_261_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_130_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_261_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_7100 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_261_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_131_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_261_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_7127 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_263_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_131_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_263_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_7154 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_263_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_132_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_263_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_7181 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_265_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_132_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_265_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_7208 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_265_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_133_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_265_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_7235 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_267_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_133_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_267_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_7262 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_267_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_134_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_267_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_7289 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_269_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_134_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_269_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_7316 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_269_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_135_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_269_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_7343 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_271_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_135_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_271_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_7370 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_271_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_136_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_271_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_7397 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_273_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_136_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_273_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_7424 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_273_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_137_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_273_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_7451 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_275_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_137_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_275_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_7478 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_275_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_138_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_275_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_7505 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_277_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_138_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_277_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_7532 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_277_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_139_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_277_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_7559 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_279_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_139_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_279_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_7586 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_279_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_140_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_279_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_7613 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_281_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_140_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_281_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_7640 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_281_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_141_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_281_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_7667 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_283_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_141_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_283_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_7694 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_283_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_142_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_283_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_7721 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_285_value & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_142_1 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_285_value & _s2_redirect_s1_last_pred_vec_T_53 &
    s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_7748 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_285_value &
    _s2_redirect_s1_last_pred_vec_WIRE_2_0; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_143_0 = s2_ghist_ptr_value == s1_ghv_wens_new_ptr_285_value & _s2_redirect_s1_last_pred_vec_WIRE_2_0
     & s2_redirect; // @[BPU.scala 483:119]
  wire  _s2_ghv_wens_T_7775 = s2_ghist_ptr_value == 8'h0 & _s2_redirect_s1_last_pred_vec_T_53; // @[BPU.scala 483:90]
  wire  s2_ghv_wens_143_1 = s2_ghist_ptr_value == 8'h0 & _s2_redirect_s1_last_pred_vec_T_53 & s2_redirect; // @[BPU.scala 483:119]
  wire [1:0] _s1_pred_info_taken_cfiIndex_valid_T_7 = {_s1_predicted_ghist_ptr_T_12,_s1_predicted_ghist_ptr_T_11}; // @[FrontendBundle.scala 492:46]
  wire  cfiIndex_valid = |_s1_pred_info_taken_cfiIndex_valid_T_7; // @[FrontendBundle.scala 492:53]
  wire [2:0] _s1_pred_info_taken_cfiIndex_bits_T_8 = _s1_predicted_ghist_ptr_T_11 ?
    predictors_io_out_s1_full_pred_offsets_0 : predictors_io_out_s1_full_pred_offsets_1; // @[ParallelMux.scala 90:77]
  wire  _s1_pred_info_taken_cfiIndex_bits_T_18 = ~cfiIndex_valid; // @[FrontendBundle.scala 496:37]
  wire [2:0] _s1_pred_info_taken_cfiIndex_bits_T_20 = _s1_pred_info_taken_cfiIndex_bits_T_18 ? 3'h7 : 3'h0; // @[Bitwise.scala 74:12]
  wire [2:0] cfiIndex_bits = _s1_pred_info_taken_cfiIndex_bits_T_8 | _s1_pred_info_taken_cfiIndex_bits_T_20; // @[FrontendBundle.scala 495:60]
  wire  _T_385 = s2_ghv_wens_0_0 | s2_ghv_wens_0_1; // @[BPU.scala 511:26]
  wire  _T_386 = s2_ghv_wens_1_0 | s2_ghv_wens_1_1; // @[BPU.scala 511:26]
  wire  _T_387 = s2_ghv_wens_2_0 | s2_ghv_wens_2_1; // @[BPU.scala 511:26]
  wire  _T_388 = s2_ghv_wens_3_0 | s2_ghv_wens_3_1; // @[BPU.scala 511:26]
  wire  _T_389 = s2_ghv_wens_4_0 | s2_ghv_wens_4_1; // @[BPU.scala 511:26]
  wire  _T_390 = s2_ghv_wens_5_0 | s2_ghv_wens_5_1; // @[BPU.scala 511:26]
  wire  _T_391 = s2_ghv_wens_6_0 | s2_ghv_wens_6_1; // @[BPU.scala 511:26]
  wire  _T_392 = s2_ghv_wens_7_0 | s2_ghv_wens_7_1; // @[BPU.scala 511:26]
  wire  _T_393 = s2_ghv_wens_8_0 | s2_ghv_wens_8_1; // @[BPU.scala 511:26]
  wire  _T_394 = s2_ghv_wens_9_0 | s2_ghv_wens_9_1; // @[BPU.scala 511:26]
  wire  _T_395 = s2_ghv_wens_10_0 | s2_ghv_wens_10_1; // @[BPU.scala 511:26]
  wire  _T_396 = s2_ghv_wens_11_0 | s2_ghv_wens_11_1; // @[BPU.scala 511:26]
  wire  _T_397 = s2_ghv_wens_12_0 | s2_ghv_wens_12_1; // @[BPU.scala 511:26]
  wire  _T_398 = s2_ghv_wens_13_0 | s2_ghv_wens_13_1; // @[BPU.scala 511:26]
  wire  _T_399 = s2_ghv_wens_14_0 | s2_ghv_wens_14_1; // @[BPU.scala 511:26]
  wire  _T_400 = s2_ghv_wens_15_0 | s2_ghv_wens_15_1; // @[BPU.scala 511:26]
  wire  _T_401 = s2_ghv_wens_16_0 | s2_ghv_wens_16_1; // @[BPU.scala 511:26]
  wire  _T_402 = s2_ghv_wens_17_0 | s2_ghv_wens_17_1; // @[BPU.scala 511:26]
  wire  _T_403 = s2_ghv_wens_18_0 | s2_ghv_wens_18_1; // @[BPU.scala 511:26]
  wire  _T_404 = s2_ghv_wens_19_0 | s2_ghv_wens_19_1; // @[BPU.scala 511:26]
  wire  _T_405 = s2_ghv_wens_20_0 | s2_ghv_wens_20_1; // @[BPU.scala 511:26]
  wire  _T_406 = s2_ghv_wens_21_0 | s2_ghv_wens_21_1; // @[BPU.scala 511:26]
  wire  _T_407 = s2_ghv_wens_22_0 | s2_ghv_wens_22_1; // @[BPU.scala 511:26]
  wire  _T_408 = s2_ghv_wens_23_0 | s2_ghv_wens_23_1; // @[BPU.scala 511:26]
  wire  _T_409 = s2_ghv_wens_24_0 | s2_ghv_wens_24_1; // @[BPU.scala 511:26]
  wire  _T_410 = s2_ghv_wens_25_0 | s2_ghv_wens_25_1; // @[BPU.scala 511:26]
  wire  _T_411 = s2_ghv_wens_26_0 | s2_ghv_wens_26_1; // @[BPU.scala 511:26]
  wire  _T_412 = s2_ghv_wens_27_0 | s2_ghv_wens_27_1; // @[BPU.scala 511:26]
  wire  _T_413 = s2_ghv_wens_28_0 | s2_ghv_wens_28_1; // @[BPU.scala 511:26]
  wire  _T_414 = s2_ghv_wens_29_0 | s2_ghv_wens_29_1; // @[BPU.scala 511:26]
  wire  _T_415 = s2_ghv_wens_30_0 | s2_ghv_wens_30_1; // @[BPU.scala 511:26]
  wire  _T_416 = s2_ghv_wens_31_0 | s2_ghv_wens_31_1; // @[BPU.scala 511:26]
  wire  _T_417 = s2_ghv_wens_32_0 | s2_ghv_wens_32_1; // @[BPU.scala 511:26]
  wire  _T_418 = s2_ghv_wens_33_0 | s2_ghv_wens_33_1; // @[BPU.scala 511:26]
  wire  _T_419 = s2_ghv_wens_34_0 | s2_ghv_wens_34_1; // @[BPU.scala 511:26]
  wire  _T_420 = s2_ghv_wens_35_0 | s2_ghv_wens_35_1; // @[BPU.scala 511:26]
  wire  _T_421 = s2_ghv_wens_36_0 | s2_ghv_wens_36_1; // @[BPU.scala 511:26]
  wire  _T_422 = s2_ghv_wens_37_0 | s2_ghv_wens_37_1; // @[BPU.scala 511:26]
  wire  _T_423 = s2_ghv_wens_38_0 | s2_ghv_wens_38_1; // @[BPU.scala 511:26]
  wire  _T_424 = s2_ghv_wens_39_0 | s2_ghv_wens_39_1; // @[BPU.scala 511:26]
  wire  _T_425 = s2_ghv_wens_40_0 | s2_ghv_wens_40_1; // @[BPU.scala 511:26]
  wire  _T_426 = s2_ghv_wens_41_0 | s2_ghv_wens_41_1; // @[BPU.scala 511:26]
  wire  _T_427 = s2_ghv_wens_42_0 | s2_ghv_wens_42_1; // @[BPU.scala 511:26]
  wire  _T_428 = s2_ghv_wens_43_0 | s2_ghv_wens_43_1; // @[BPU.scala 511:26]
  wire  _T_429 = s2_ghv_wens_44_0 | s2_ghv_wens_44_1; // @[BPU.scala 511:26]
  wire  _T_430 = s2_ghv_wens_45_0 | s2_ghv_wens_45_1; // @[BPU.scala 511:26]
  wire  _T_431 = s2_ghv_wens_46_0 | s2_ghv_wens_46_1; // @[BPU.scala 511:26]
  wire  _T_432 = s2_ghv_wens_47_0 | s2_ghv_wens_47_1; // @[BPU.scala 511:26]
  wire  _T_433 = s2_ghv_wens_48_0 | s2_ghv_wens_48_1; // @[BPU.scala 511:26]
  wire  _T_434 = s2_ghv_wens_49_0 | s2_ghv_wens_49_1; // @[BPU.scala 511:26]
  wire  _T_435 = s2_ghv_wens_50_0 | s2_ghv_wens_50_1; // @[BPU.scala 511:26]
  wire  _T_436 = s2_ghv_wens_51_0 | s2_ghv_wens_51_1; // @[BPU.scala 511:26]
  wire  _T_437 = s2_ghv_wens_52_0 | s2_ghv_wens_52_1; // @[BPU.scala 511:26]
  wire  _T_438 = s2_ghv_wens_53_0 | s2_ghv_wens_53_1; // @[BPU.scala 511:26]
  wire  _T_439 = s2_ghv_wens_54_0 | s2_ghv_wens_54_1; // @[BPU.scala 511:26]
  wire  _T_440 = s2_ghv_wens_55_0 | s2_ghv_wens_55_1; // @[BPU.scala 511:26]
  wire  _T_441 = s2_ghv_wens_56_0 | s2_ghv_wens_56_1; // @[BPU.scala 511:26]
  wire  _T_442 = s2_ghv_wens_57_0 | s2_ghv_wens_57_1; // @[BPU.scala 511:26]
  wire  _T_443 = s2_ghv_wens_58_0 | s2_ghv_wens_58_1; // @[BPU.scala 511:26]
  wire  _T_444 = s2_ghv_wens_59_0 | s2_ghv_wens_59_1; // @[BPU.scala 511:26]
  wire  _T_445 = s2_ghv_wens_60_0 | s2_ghv_wens_60_1; // @[BPU.scala 511:26]
  wire  _T_446 = s2_ghv_wens_61_0 | s2_ghv_wens_61_1; // @[BPU.scala 511:26]
  wire  _T_447 = s2_ghv_wens_62_0 | s2_ghv_wens_62_1; // @[BPU.scala 511:26]
  wire  _T_448 = s2_ghv_wens_63_0 | s2_ghv_wens_63_1; // @[BPU.scala 511:26]
  wire  _T_449 = s2_ghv_wens_64_0 | s2_ghv_wens_64_1; // @[BPU.scala 511:26]
  wire  _T_450 = s2_ghv_wens_65_0 | s2_ghv_wens_65_1; // @[BPU.scala 511:26]
  wire  _T_451 = s2_ghv_wens_66_0 | s2_ghv_wens_66_1; // @[BPU.scala 511:26]
  wire  _T_452 = s2_ghv_wens_67_0 | s2_ghv_wens_67_1; // @[BPU.scala 511:26]
  wire  _T_453 = s2_ghv_wens_68_0 | s2_ghv_wens_68_1; // @[BPU.scala 511:26]
  wire  _T_454 = s2_ghv_wens_69_0 | s2_ghv_wens_69_1; // @[BPU.scala 511:26]
  wire  _T_455 = s2_ghv_wens_70_0 | s2_ghv_wens_70_1; // @[BPU.scala 511:26]
  wire  _T_456 = s2_ghv_wens_71_0 | s2_ghv_wens_71_1; // @[BPU.scala 511:26]
  wire  _T_457 = s2_ghv_wens_72_0 | s2_ghv_wens_72_1; // @[BPU.scala 511:26]
  wire  _T_458 = s2_ghv_wens_73_0 | s2_ghv_wens_73_1; // @[BPU.scala 511:26]
  wire  _T_459 = s2_ghv_wens_74_0 | s2_ghv_wens_74_1; // @[BPU.scala 511:26]
  wire  _T_460 = s2_ghv_wens_75_0 | s2_ghv_wens_75_1; // @[BPU.scala 511:26]
  wire  _T_461 = s2_ghv_wens_76_0 | s2_ghv_wens_76_1; // @[BPU.scala 511:26]
  wire  _T_462 = s2_ghv_wens_77_0 | s2_ghv_wens_77_1; // @[BPU.scala 511:26]
  wire  _T_463 = s2_ghv_wens_78_0 | s2_ghv_wens_78_1; // @[BPU.scala 511:26]
  wire  _T_464 = s2_ghv_wens_79_0 | s2_ghv_wens_79_1; // @[BPU.scala 511:26]
  wire  _T_465 = s2_ghv_wens_80_0 | s2_ghv_wens_80_1; // @[BPU.scala 511:26]
  wire  _T_466 = s2_ghv_wens_81_0 | s2_ghv_wens_81_1; // @[BPU.scala 511:26]
  wire  _T_467 = s2_ghv_wens_82_0 | s2_ghv_wens_82_1; // @[BPU.scala 511:26]
  wire  _T_468 = s2_ghv_wens_83_0 | s2_ghv_wens_83_1; // @[BPU.scala 511:26]
  wire  _T_469 = s2_ghv_wens_84_0 | s2_ghv_wens_84_1; // @[BPU.scala 511:26]
  wire  _T_470 = s2_ghv_wens_85_0 | s2_ghv_wens_85_1; // @[BPU.scala 511:26]
  wire  _T_471 = s2_ghv_wens_86_0 | s2_ghv_wens_86_1; // @[BPU.scala 511:26]
  wire  _T_472 = s2_ghv_wens_87_0 | s2_ghv_wens_87_1; // @[BPU.scala 511:26]
  wire  _T_473 = s2_ghv_wens_88_0 | s2_ghv_wens_88_1; // @[BPU.scala 511:26]
  wire  _T_474 = s2_ghv_wens_89_0 | s2_ghv_wens_89_1; // @[BPU.scala 511:26]
  wire  _T_475 = s2_ghv_wens_90_0 | s2_ghv_wens_90_1; // @[BPU.scala 511:26]
  wire  _T_476 = s2_ghv_wens_91_0 | s2_ghv_wens_91_1; // @[BPU.scala 511:26]
  wire  _T_477 = s2_ghv_wens_92_0 | s2_ghv_wens_92_1; // @[BPU.scala 511:26]
  wire  _T_478 = s2_ghv_wens_93_0 | s2_ghv_wens_93_1; // @[BPU.scala 511:26]
  wire  _T_479 = s2_ghv_wens_94_0 | s2_ghv_wens_94_1; // @[BPU.scala 511:26]
  wire  _T_480 = s2_ghv_wens_95_0 | s2_ghv_wens_95_1; // @[BPU.scala 511:26]
  wire  _T_481 = s2_ghv_wens_96_0 | s2_ghv_wens_96_1; // @[BPU.scala 511:26]
  wire  _T_482 = s2_ghv_wens_97_0 | s2_ghv_wens_97_1; // @[BPU.scala 511:26]
  wire  _T_483 = s2_ghv_wens_98_0 | s2_ghv_wens_98_1; // @[BPU.scala 511:26]
  wire  _T_484 = s2_ghv_wens_99_0 | s2_ghv_wens_99_1; // @[BPU.scala 511:26]
  wire  _T_485 = s2_ghv_wens_100_0 | s2_ghv_wens_100_1; // @[BPU.scala 511:26]
  wire  _T_486 = s2_ghv_wens_101_0 | s2_ghv_wens_101_1; // @[BPU.scala 511:26]
  wire  _T_487 = s2_ghv_wens_102_0 | s2_ghv_wens_102_1; // @[BPU.scala 511:26]
  wire  _T_488 = s2_ghv_wens_103_0 | s2_ghv_wens_103_1; // @[BPU.scala 511:26]
  wire  _T_489 = s2_ghv_wens_104_0 | s2_ghv_wens_104_1; // @[BPU.scala 511:26]
  wire  _T_490 = s2_ghv_wens_105_0 | s2_ghv_wens_105_1; // @[BPU.scala 511:26]
  wire  _T_491 = s2_ghv_wens_106_0 | s2_ghv_wens_106_1; // @[BPU.scala 511:26]
  wire  _T_492 = s2_ghv_wens_107_0 | s2_ghv_wens_107_1; // @[BPU.scala 511:26]
  wire  _T_493 = s2_ghv_wens_108_0 | s2_ghv_wens_108_1; // @[BPU.scala 511:26]
  wire  _T_494 = s2_ghv_wens_109_0 | s2_ghv_wens_109_1; // @[BPU.scala 511:26]
  wire  _T_495 = s2_ghv_wens_110_0 | s2_ghv_wens_110_1; // @[BPU.scala 511:26]
  wire  _T_496 = s2_ghv_wens_111_0 | s2_ghv_wens_111_1; // @[BPU.scala 511:26]
  wire  _T_497 = s2_ghv_wens_112_0 | s2_ghv_wens_112_1; // @[BPU.scala 511:26]
  wire  _T_498 = s2_ghv_wens_113_0 | s2_ghv_wens_113_1; // @[BPU.scala 511:26]
  wire  _T_499 = s2_ghv_wens_114_0 | s2_ghv_wens_114_1; // @[BPU.scala 511:26]
  wire  _T_500 = s2_ghv_wens_115_0 | s2_ghv_wens_115_1; // @[BPU.scala 511:26]
  wire  _T_501 = s2_ghv_wens_116_0 | s2_ghv_wens_116_1; // @[BPU.scala 511:26]
  wire  _T_502 = s2_ghv_wens_117_0 | s2_ghv_wens_117_1; // @[BPU.scala 511:26]
  wire  _T_503 = s2_ghv_wens_118_0 | s2_ghv_wens_118_1; // @[BPU.scala 511:26]
  wire  _T_504 = s2_ghv_wens_119_0 | s2_ghv_wens_119_1; // @[BPU.scala 511:26]
  wire  _T_505 = s2_ghv_wens_120_0 | s2_ghv_wens_120_1; // @[BPU.scala 511:26]
  wire  _T_506 = s2_ghv_wens_121_0 | s2_ghv_wens_121_1; // @[BPU.scala 511:26]
  wire  _T_507 = s2_ghv_wens_122_0 | s2_ghv_wens_122_1; // @[BPU.scala 511:26]
  wire  _T_508 = s2_ghv_wens_123_0 | s2_ghv_wens_123_1; // @[BPU.scala 511:26]
  wire  _T_509 = s2_ghv_wens_124_0 | s2_ghv_wens_124_1; // @[BPU.scala 511:26]
  wire  _T_510 = s2_ghv_wens_125_0 | s2_ghv_wens_125_1; // @[BPU.scala 511:26]
  wire  _T_511 = s2_ghv_wens_126_0 | s2_ghv_wens_126_1; // @[BPU.scala 511:26]
  wire  _T_512 = s2_ghv_wens_127_0 | s2_ghv_wens_127_1; // @[BPU.scala 511:26]
  wire  _T_513 = s2_ghv_wens_128_0 | s2_ghv_wens_128_1; // @[BPU.scala 511:26]
  wire  _T_514 = s2_ghv_wens_129_0 | s2_ghv_wens_129_1; // @[BPU.scala 511:26]
  wire  _T_515 = s2_ghv_wens_130_0 | s2_ghv_wens_130_1; // @[BPU.scala 511:26]
  wire  _T_516 = s2_ghv_wens_131_0 | s2_ghv_wens_131_1; // @[BPU.scala 511:26]
  wire  _T_517 = s2_ghv_wens_132_0 | s2_ghv_wens_132_1; // @[BPU.scala 511:26]
  wire  _T_518 = s2_ghv_wens_133_0 | s2_ghv_wens_133_1; // @[BPU.scala 511:26]
  wire  _T_519 = s2_ghv_wens_134_0 | s2_ghv_wens_134_1; // @[BPU.scala 511:26]
  wire  _T_520 = s2_ghv_wens_135_0 | s2_ghv_wens_135_1; // @[BPU.scala 511:26]
  wire  _T_521 = s2_ghv_wens_136_0 | s2_ghv_wens_136_1; // @[BPU.scala 511:26]
  wire  _T_522 = s2_ghv_wens_137_0 | s2_ghv_wens_137_1; // @[BPU.scala 511:26]
  wire  _T_523 = s2_ghv_wens_138_0 | s2_ghv_wens_138_1; // @[BPU.scala 511:26]
  wire  _T_524 = s2_ghv_wens_139_0 | s2_ghv_wens_139_1; // @[BPU.scala 511:26]
  wire  _T_525 = s2_ghv_wens_140_0 | s2_ghv_wens_140_1; // @[BPU.scala 511:26]
  wire  _T_526 = s2_ghv_wens_141_0 | s2_ghv_wens_141_1; // @[BPU.scala 511:26]
  wire  _T_527 = s2_ghv_wens_142_0 | s2_ghv_wens_142_1; // @[BPU.scala 511:26]
  wire  _T_528 = s2_ghv_wens_143_0 | s2_ghv_wens_143_1; // @[BPU.scala 511:26]
  wire [8:0] s3_possible_predicted_ghist_ptrs_flipped_new_ptr_new_value = s3_ghist_ptr_value +
    _s1_possible_predicted_ghist_ptrs_flipped_new_ptr_T_1; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _s3_possible_predicted_ghist_ptrs_flipped_new_ptr_diff_T_1 = {1'h0,
    s3_possible_predicted_ghist_ptrs_flipped_new_ptr_new_value}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] s3_possible_predicted_ghist_ptrs_flipped_new_ptr_diff = $signed(
    _s3_possible_predicted_ghist_ptrs_flipped_new_ptr_diff_T_1) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s3_possible_predicted_ghist_ptrs_flipped_new_ptr_reverse_flag = $signed(
    s3_possible_predicted_ghist_ptrs_flipped_new_ptr_diff) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire  s3_possible_predicted_ghist_ptrs_flipped_new_ptr_flag =
    s3_possible_predicted_ghist_ptrs_flipped_new_ptr_reverse_flag ? ~s3_ghist_ptr_flag : s3_ghist_ptr_flag; // @[CircularQueuePtr.scala 44:26]
  wire [9:0] _s3_possible_predicted_ghist_ptrs_flipped_new_ptr_new_ptr_value_T = $signed(
    _s3_possible_predicted_ghist_ptrs_flipped_new_ptr_diff_T_1) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s3_possible_predicted_ghist_ptrs_flipped_new_ptr_new_ptr_value_T_1 =
    s3_possible_predicted_ghist_ptrs_flipped_new_ptr_reverse_flag ?
    _s3_possible_predicted_ghist_ptrs_flipped_new_ptr_new_ptr_value_T : {{1'd0},
    s3_possible_predicted_ghist_ptrs_flipped_new_ptr_new_value}; // @[CircularQueuePtr.scala 45:27]
  wire  s3_possible_predicted_ghist_ptrs_0_flag = ~s3_possible_predicted_ghist_ptrs_flipped_new_ptr_flag; // @[CircularQueuePtr.scala 56:21]
  wire [8:0] s3_possible_predicted_ghist_ptrs_flipped_new_ptr_new_value_1 = s3_ghist_ptr_value +
    _s1_possible_predicted_ghist_ptrs_flipped_new_ptr_T_3; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _s3_possible_predicted_ghist_ptrs_flipped_new_ptr_diff_T_7 = {1'h0,
    s3_possible_predicted_ghist_ptrs_flipped_new_ptr_new_value_1}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] s3_possible_predicted_ghist_ptrs_flipped_new_ptr_diff_1 = $signed(
    _s3_possible_predicted_ghist_ptrs_flipped_new_ptr_diff_T_7) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s3_possible_predicted_ghist_ptrs_flipped_new_ptr_reverse_flag_1 = $signed(
    s3_possible_predicted_ghist_ptrs_flipped_new_ptr_diff_1) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire  s3_possible_predicted_ghist_ptrs_flipped_new_ptr_1_flag =
    s3_possible_predicted_ghist_ptrs_flipped_new_ptr_reverse_flag_1 ? ~s3_ghist_ptr_flag : s3_ghist_ptr_flag; // @[CircularQueuePtr.scala 44:26]
  wire [9:0] _s3_possible_predicted_ghist_ptrs_flipped_new_ptr_new_ptr_value_T_2 = $signed(
    _s3_possible_predicted_ghist_ptrs_flipped_new_ptr_diff_T_7) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s3_possible_predicted_ghist_ptrs_flipped_new_ptr_new_ptr_value_T_3 =
    s3_possible_predicted_ghist_ptrs_flipped_new_ptr_reverse_flag_1 ?
    _s3_possible_predicted_ghist_ptrs_flipped_new_ptr_new_ptr_value_T_2 : {{1'd0},
    s3_possible_predicted_ghist_ptrs_flipped_new_ptr_new_value_1}; // @[CircularQueuePtr.scala 45:27]
  wire  s3_possible_predicted_ghist_ptrs_1_flag = ~s3_possible_predicted_ghist_ptrs_flipped_new_ptr_1_flag; // @[CircularQueuePtr.scala 56:21]
  wire [8:0] s3_possible_predicted_ghist_ptrs_flipped_new_ptr_new_value_2 = s3_ghist_ptr_value +
    _s1_possible_predicted_ghist_ptrs_flipped_new_ptr_T_5; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _s3_possible_predicted_ghist_ptrs_flipped_new_ptr_diff_T_13 = {1'h0,
    s3_possible_predicted_ghist_ptrs_flipped_new_ptr_new_value_2}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] s3_possible_predicted_ghist_ptrs_flipped_new_ptr_diff_2 = $signed(
    _s3_possible_predicted_ghist_ptrs_flipped_new_ptr_diff_T_13) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  s3_possible_predicted_ghist_ptrs_flipped_new_ptr_reverse_flag_2 = $signed(
    s3_possible_predicted_ghist_ptrs_flipped_new_ptr_diff_2) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire  s3_possible_predicted_ghist_ptrs_flipped_new_ptr_2_flag =
    s3_possible_predicted_ghist_ptrs_flipped_new_ptr_reverse_flag_2 ? ~s3_ghist_ptr_flag : s3_ghist_ptr_flag; // @[CircularQueuePtr.scala 44:26]
  wire [9:0] _s3_possible_predicted_ghist_ptrs_flipped_new_ptr_new_ptr_value_T_4 = $signed(
    _s3_possible_predicted_ghist_ptrs_flipped_new_ptr_diff_T_13) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _s3_possible_predicted_ghist_ptrs_flipped_new_ptr_new_ptr_value_T_5 =
    s3_possible_predicted_ghist_ptrs_flipped_new_ptr_reverse_flag_2 ?
    _s3_possible_predicted_ghist_ptrs_flipped_new_ptr_new_ptr_value_T_4 : {{1'd0},
    s3_possible_predicted_ghist_ptrs_flipped_new_ptr_new_value_2}; // @[CircularQueuePtr.scala 45:27]
  wire  s3_possible_predicted_ghist_ptrs_2_flag = ~s3_possible_predicted_ghist_ptrs_flipped_new_ptr_2_flag; // @[CircularQueuePtr.scala 56:21]
  wire  _s3_predicted_ghist_ptr_T_1 = predictors_io_out_s3_full_pred_slot_valids_1 &
    predictors_io_out_s3_full_pred_is_br_sharing; // @[FrontendBundle.scala 430:48]
  wire  _s3_predicted_ghist_ptr_WIRE__0 = predictors_io_out_s3_full_pred_slot_valids_0; // @[FrontendBundle.scala 430:{12,12}]
  wire  _s3_predicted_ghist_ptr_T_4 = selVecOH_3_3 | ~(_s3_predicted_ghist_ptr_WIRE__0 | _s3_predicted_ghist_ptr_T_1); // @[FrontendBundle.scala 461:19]
  wire  _s3_predicted_ghist_ptr_T_30 = _s3_redirect_on_br_taken_T_5 | ~_s3_predicted_ghist_ptr_T_1; // @[FrontendBundle.scala 465:34]
  wire  _s3_predicted_ghist_ptr_T_31 = _s3_predicted_ghist_ptr_WIRE__0 & _s3_predicted_ghist_ptr_T_30; // @[FrontendBundle.scala 464:75]
  wire  _s3_predicted_ghist_ptr_T_32 = _s3_predicted_ghist_ptr_T_31 & predictors_io_out_s3_full_pred_hit; // @[FrontendBundle.scala 465:97]
  wire  _s3_predicted_ghist_ptr_T_44 = ~_s3_redirect_on_br_taken_T_5; // @[FrontendBundle.scala 464:9]
  wire  _s3_predicted_ghist_ptr_T_45 = _s3_predicted_ghist_ptr_T_1 & _s3_predicted_ghist_ptr_T_44; // @[FrontendBundle.scala 463:22]
  wire  _s3_predicted_ghist_ptr_T_60 = _s3_predicted_ghist_ptr_T_45 & predictors_io_out_s3_full_pred_hit; // @[FrontendBundle.scala 465:97]
  wire [7:0] s3_possible_predicted_ghist_ptrs_flipped_new_ptr_value =
    _s3_possible_predicted_ghist_ptrs_flipped_new_ptr_new_ptr_value_T_1[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire [7:0] _s3_predicted_ghist_ptr_T_61 = _s3_predicted_ghist_ptr_T_4 ?
    s3_possible_predicted_ghist_ptrs_flipped_new_ptr_value : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] s3_possible_predicted_ghist_ptrs_flipped_new_ptr_1_value =
    _s3_possible_predicted_ghist_ptrs_flipped_new_ptr_new_ptr_value_T_3[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire [7:0] _s3_predicted_ghist_ptr_T_62 = _s3_predicted_ghist_ptr_T_32 ?
    s3_possible_predicted_ghist_ptrs_flipped_new_ptr_1_value : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] s3_possible_predicted_ghist_ptrs_flipped_new_ptr_2_value =
    _s3_possible_predicted_ghist_ptrs_flipped_new_ptr_new_ptr_value_T_5[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire [7:0] _s3_predicted_ghist_ptr_T_63 = _s3_predicted_ghist_ptr_T_60 ?
    s3_possible_predicted_ghist_ptrs_flipped_new_ptr_2_value : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _s3_predicted_ghist_ptr_T_64 = _s3_predicted_ghist_ptr_T_61 | _s3_predicted_ghist_ptr_T_62; // @[Mux.scala 27:73]
  wire  s3_possible_predicted_fhs_ob__0 = s3_last_br_num_oh[0] & s3_ahead_fh_oldest_bits_afhob_3_bits_0 |
    s3_last_br_num_oh[1] & s3_ahead_fh_oldest_bits_afhob_3_bits_1 | s3_last_br_num_oh[2] &
    s3_ahead_fh_oldest_bits_afhob_3_bits_2; // @[Mux.scala 27:73]
  wire  s3_possible_predicted_fhs_ob__1 = s3_last_br_num_oh[0] & s3_ahead_fh_oldest_bits_afhob_3_bits_1 |
    s3_last_br_num_oh[1] & s3_ahead_fh_oldest_bits_afhob_3_bits_2 | s3_last_br_num_oh[2] &
    s3_ahead_fh_oldest_bits_afhob_3_bits_3; // @[Mux.scala 27:73]
  wire  s3_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__0 = s3_folded_gh_hist_0_folded_hist[0
    ]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__1 = s3_folded_gh_hist_0_folded_hist[1
    ]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__2 = s3_folded_gh_hist_0_folded_hist[2
    ]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__3 = s3_folded_gh_hist_0_folded_hist[3
    ]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__4 = s3_folded_gh_hist_0_folded_hist[4
    ]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__5 = s3_folded_gh_hist_0_folded_hist[5
    ]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__6 = s3_folded_gh_hist_0_folded_hist[6
    ]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__7 = s3_folded_gh_hist_0_folded_hist[7
    ]; // @[FrontendBundle.scala 280:54]
  wire [7:0] s3_possible_predicted_fhs_res_hist_0_new_folded_hist_xored = {
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__7,
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__6,
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__5,
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__4,
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__3,
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__1,
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [15:0] s3_possible_predicted_fhs_res_hist_0_new_folded_hist_src_doubled = {
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__7,
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__6,
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__5,
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__4,
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__3,
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__1,
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__0,
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_xored}; // @[Cat.scala 31:58]
  wire [7:0] s3_possible_predicted_fhs_res_hist_0_new_folded_hist =
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_src_doubled[15:8]; // @[FrontendBundle.scala 221:30]
  wire  s3_possible_predicted_fhs_ob_1_0 = s3_last_br_num_oh[0] & s3_ahead_fh_oldest_bits_afhob_2_bits_0 |
    s3_last_br_num_oh[1] & s3_ahead_fh_oldest_bits_afhob_2_bits_1 | s3_last_br_num_oh[2] &
    s3_ahead_fh_oldest_bits_afhob_2_bits_2; // @[Mux.scala 27:73]
  wire  s3_possible_predicted_fhs_ob_1_1 = s3_last_br_num_oh[0] & s3_ahead_fh_oldest_bits_afhob_2_bits_1 |
    s3_last_br_num_oh[1] & s3_ahead_fh_oldest_bits_afhob_2_bits_2 | s3_last_br_num_oh[2] &
    s3_ahead_fh_oldest_bits_afhob_2_bits_3; // @[Mux.scala 27:73]
  wire  s3_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__0 = s3_folded_gh_hist_1_folded_hist[0
    ]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__1 = s3_folded_gh_hist_1_folded_hist[1
    ]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__2 = s3_folded_gh_hist_1_folded_hist[2
    ]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__3 = s3_folded_gh_hist_1_folded_hist[3
    ]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__4 = s3_folded_gh_hist_1_folded_hist[4
    ]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__5 = s3_folded_gh_hist_1_folded_hist[5
    ]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__6 = s3_folded_gh_hist_1_folded_hist[6
    ]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__7 = s3_folded_gh_hist_1_folded_hist[7
    ]; // @[FrontendBundle.scala 280:54]
  wire [7:0] s3_possible_predicted_fhs_res_hist_1_new_folded_hist_xored = {
    s3_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__7,
    s3_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__6,
    s3_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__5,
    s3_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__4,
    s3_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__3,
    s3_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__1,
    s3_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [15:0] s3_possible_predicted_fhs_res_hist_1_new_folded_hist_src_doubled = {
    s3_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__7,
    s3_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__6,
    s3_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__5,
    s3_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__4,
    s3_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__3,
    s3_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__1,
    s3_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__0,
    s3_possible_predicted_fhs_res_hist_1_new_folded_hist_xored}; // @[Cat.scala 31:58]
  wire [7:0] s3_possible_predicted_fhs_res_hist_1_new_folded_hist =
    s3_possible_predicted_fhs_res_hist_1_new_folded_hist_src_doubled[15:8]; // @[FrontendBundle.scala 221:30]
  wire  s3_possible_predicted_fhs_ob_2_0 = s3_last_br_num_oh[0] & s3_ahead_fh_oldest_bits_afhob_5_bits_0 |
    s3_last_br_num_oh[1] & s3_ahead_fh_oldest_bits_afhob_5_bits_1 | s3_last_br_num_oh[2] &
    s3_ahead_fh_oldest_bits_afhob_5_bits_2; // @[Mux.scala 27:73]
  wire  s3_possible_predicted_fhs_ob_2_1 = s3_last_br_num_oh[0] & s3_ahead_fh_oldest_bits_afhob_5_bits_1 |
    s3_last_br_num_oh[1] & s3_ahead_fh_oldest_bits_afhob_5_bits_2 | s3_last_br_num_oh[2] &
    s3_ahead_fh_oldest_bits_afhob_5_bits_3; // @[Mux.scala 27:73]
  wire  s3_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__0 = s3_folded_gh_hist_2_folded_hist[0
    ]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__1 = s3_folded_gh_hist_2_folded_hist[1
    ]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__2 = s3_folded_gh_hist_2_folded_hist[2
    ]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__3 = s3_folded_gh_hist_2_folded_hist[3
    ]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__4 = s3_folded_gh_hist_2_folded_hist[4
    ]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__5 = s3_folded_gh_hist_2_folded_hist[5
    ]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__6 = s3_folded_gh_hist_2_folded_hist[6
    ]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__7 = s3_folded_gh_hist_2_folded_hist[7
    ]; // @[FrontendBundle.scala 280:54]
  wire [7:0] s3_possible_predicted_fhs_res_hist_2_new_folded_hist_xored = {
    s3_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__7,
    s3_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__6,
    s3_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__5,
    s3_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__4,
    s3_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__3,
    s3_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__1,
    s3_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [15:0] s3_possible_predicted_fhs_res_hist_2_new_folded_hist_src_doubled = {
    s3_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__7,
    s3_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__6,
    s3_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__5,
    s3_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__4,
    s3_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__3,
    s3_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__1,
    s3_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__0,
    s3_possible_predicted_fhs_res_hist_2_new_folded_hist_xored}; // @[Cat.scala 31:58]
  wire [7:0] s3_possible_predicted_fhs_res_hist_2_new_folded_hist =
    s3_possible_predicted_fhs_res_hist_2_new_folded_hist_src_doubled[15:8]; // @[FrontendBundle.scala 221:30]
  wire  s3_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__0 = s3_folded_gh_hist_3_folded_hist[0
    ]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__1 = s3_folded_gh_hist_3_folded_hist[1
    ]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__2 = s3_folded_gh_hist_3_folded_hist[2
    ]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__3 = s3_folded_gh_hist_3_folded_hist[3
    ]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__4 = s3_folded_gh_hist_3_folded_hist[4
    ]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__5 = s3_folded_gh_hist_3_folded_hist[5
    ]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__6 = s3_folded_gh_hist_3_folded_hist[6
    ]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__7 = s3_folded_gh_hist_3_folded_hist[7
    ]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__8 = s3_folded_gh_hist_3_folded_hist[8
    ]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__9 = s3_folded_gh_hist_3_folded_hist[9
    ]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__10 = s3_folded_gh_hist_3_folded_hist[
    10]; // @[FrontendBundle.scala 280:54]
  wire [4:0] s3_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_lo = {
    s3_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__4,
    s3_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__3,
    s3_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__1,
    s3_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [10:0] s3_possible_predicted_fhs_res_hist_3_new_folded_hist_xored = {
    s3_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__10,
    s3_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__9,
    s3_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__8,
    s3_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__7,
    s3_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__6,
    s3_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__5,
    s3_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_lo}; // @[FrontendBundle.scala 258:11]
  wire [21:0] s3_possible_predicted_fhs_res_hist_3_new_folded_hist_src_doubled = {
    s3_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__10,
    s3_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__9,
    s3_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__8,
    s3_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__7,
    s3_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__6,
    s3_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__5,
    s3_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_lo,
    s3_possible_predicted_fhs_res_hist_3_new_folded_hist_xored}; // @[Cat.scala 31:58]
  wire [10:0] s3_possible_predicted_fhs_res_hist_3_new_folded_hist =
    s3_possible_predicted_fhs_res_hist_3_new_folded_hist_src_doubled[21:11]; // @[FrontendBundle.scala 221:30]
  wire  s3_possible_predicted_fhs_ob_4_0 = s3_last_br_num_oh[0] & s3_ahead_fh_oldest_bits_afhob_1_bits_0 |
    s3_last_br_num_oh[1] & s3_ahead_fh_oldest_bits_afhob_1_bits_1 | s3_last_br_num_oh[2] &
    s3_ahead_fh_oldest_bits_afhob_1_bits_2; // @[Mux.scala 27:73]
  wire  s3_possible_predicted_fhs_ob_4_1 = s3_last_br_num_oh[0] & s3_ahead_fh_oldest_bits_afhob_1_bits_1 |
    s3_last_br_num_oh[1] & s3_ahead_fh_oldest_bits_afhob_1_bits_2 | s3_last_br_num_oh[2] &
    s3_ahead_fh_oldest_bits_afhob_1_bits_3; // @[Mux.scala 27:73]
  wire  s3_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__0 = s3_folded_gh_hist_5_folded_hist[0
    ]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__1 = s3_folded_gh_hist_5_folded_hist[1
    ]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__2 = s3_folded_gh_hist_5_folded_hist[2
    ]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__3 = s3_folded_gh_hist_5_folded_hist[3
    ]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__4 = s3_folded_gh_hist_5_folded_hist[4
    ]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__5 = s3_folded_gh_hist_5_folded_hist[5
    ]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__6 = s3_folded_gh_hist_5_folded_hist[6
    ]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__7 = s3_folded_gh_hist_5_folded_hist[7
    ]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__8 = s3_folded_gh_hist_5_folded_hist[8
    ]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__9 = s3_folded_gh_hist_5_folded_hist[9
    ]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__10 = s3_folded_gh_hist_5_folded_hist[
    10]; // @[FrontendBundle.scala 280:54]
  wire [4:0] s3_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_lo = {
    s3_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__4,
    s3_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__3,
    s3_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__1,
    s3_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [10:0] s3_possible_predicted_fhs_res_hist_5_new_folded_hist_xored = {
    s3_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__10,
    s3_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__9,
    s3_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__8,
    s3_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__7,
    s3_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__6,
    s3_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__5,
    s3_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_lo}; // @[FrontendBundle.scala 258:11]
  wire [21:0] s3_possible_predicted_fhs_res_hist_5_new_folded_hist_src_doubled = {
    s3_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__10,
    s3_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__9,
    s3_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__8,
    s3_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__7,
    s3_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__6,
    s3_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__5,
    s3_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_lo,
    s3_possible_predicted_fhs_res_hist_5_new_folded_hist_xored}; // @[Cat.scala 31:58]
  wire [10:0] s3_possible_predicted_fhs_res_hist_5_new_folded_hist =
    s3_possible_predicted_fhs_res_hist_5_new_folded_hist_src_doubled[21:11]; // @[FrontendBundle.scala 221:30]
  wire  s3_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__0 = s3_folded_gh_hist_6_folded_hist[0
    ]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__1 = s3_folded_gh_hist_6_folded_hist[1
    ]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__2 = s3_folded_gh_hist_6_folded_hist[2
    ]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__3 = s3_folded_gh_hist_6_folded_hist[3
    ]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__4 = s3_folded_gh_hist_6_folded_hist[4
    ]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__5 = s3_folded_gh_hist_6_folded_hist[5
    ]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__6 = s3_folded_gh_hist_6_folded_hist[6
    ]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__7 = s3_folded_gh_hist_6_folded_hist[7
    ]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__8 = s3_folded_gh_hist_6_folded_hist[8
    ]; // @[FrontendBundle.scala 280:54]
  wire [8:0] s3_possible_predicted_fhs_res_hist_6_new_folded_hist_xored = {
    s3_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__8,
    s3_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__7,
    s3_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__6,
    s3_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__5,
    s3_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__4,
    s3_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__3,
    s3_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__1,
    s3_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [17:0] s3_possible_predicted_fhs_res_hist_6_new_folded_hist_src_doubled = {
    s3_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__8,
    s3_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__7,
    s3_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__6,
    s3_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__5,
    s3_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__4,
    s3_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__3,
    s3_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__1,
    s3_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__0,
    s3_possible_predicted_fhs_res_hist_6_new_folded_hist_xored}; // @[Cat.scala 31:58]
  wire [8:0] s3_possible_predicted_fhs_res_hist_6_new_folded_hist =
    s3_possible_predicted_fhs_res_hist_6_new_folded_hist_src_doubled[17:9]; // @[FrontendBundle.scala 221:30]
  wire  s3_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__0 = s3_folded_gh_hist_7_folded_hist[0
    ]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__1 = s3_folded_gh_hist_7_folded_hist[1
    ]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__2 = s3_folded_gh_hist_7_folded_hist[2
    ]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__3 = s3_folded_gh_hist_7_folded_hist[3
    ]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__4 = s3_folded_gh_hist_7_folded_hist[4
    ]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__5 = s3_folded_gh_hist_7_folded_hist[5
    ]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__6 = s3_folded_gh_hist_7_folded_hist[6
    ]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__7 = s3_folded_gh_hist_7_folded_hist[7
    ]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__8 = s3_folded_gh_hist_7_folded_hist[8
    ]; // @[FrontendBundle.scala 280:54]
  wire [8:0] s3_possible_predicted_fhs_res_hist_7_new_folded_hist_xored = {
    s3_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__8,
    s3_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__7,
    s3_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__6,
    s3_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__5,
    s3_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__4,
    s3_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__3,
    s3_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__1,
    s3_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [17:0] s3_possible_predicted_fhs_res_hist_7_new_folded_hist_src_doubled = {
    s3_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__8,
    s3_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__7,
    s3_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__6,
    s3_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__5,
    s3_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__4,
    s3_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__3,
    s3_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__1,
    s3_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__0,
    s3_possible_predicted_fhs_res_hist_7_new_folded_hist_xored}; // @[Cat.scala 31:58]
  wire [8:0] s3_possible_predicted_fhs_res_hist_7_new_folded_hist =
    s3_possible_predicted_fhs_res_hist_7_new_folded_hist_src_doubled[17:9]; // @[FrontendBundle.scala 221:30]
  wire  s3_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__0 = s3_folded_gh_hist_9_folded_hist[0
    ]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__1 = s3_folded_gh_hist_9_folded_hist[1
    ]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__2 = s3_folded_gh_hist_9_folded_hist[2
    ]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__3 = s3_folded_gh_hist_9_folded_hist[3
    ]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__4 = s3_folded_gh_hist_9_folded_hist[4
    ]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__5 = s3_folded_gh_hist_9_folded_hist[5
    ]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__6 = s3_folded_gh_hist_9_folded_hist[6
    ]; // @[FrontendBundle.scala 280:54]
  wire [6:0] s3_possible_predicted_fhs_res_hist_9_new_folded_hist_xored = {
    s3_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__6,
    s3_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__5,
    s3_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__4,
    s3_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__3,
    s3_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__1,
    s3_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [13:0] s3_possible_predicted_fhs_res_hist_9_new_folded_hist_src_doubled = {
    s3_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__6,
    s3_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__5,
    s3_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__4,
    s3_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__3,
    s3_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__1,
    s3_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__0,
    s3_possible_predicted_fhs_res_hist_9_new_folded_hist_xored}; // @[Cat.scala 31:58]
  wire [6:0] s3_possible_predicted_fhs_res_hist_9_new_folded_hist =
    s3_possible_predicted_fhs_res_hist_9_new_folded_hist_src_doubled[13:7]; // @[FrontendBundle.scala 221:30]
  wire  s3_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__0 = s3_folded_gh_hist_10_folded_hist
    [0]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__1 = s3_folded_gh_hist_10_folded_hist
    [1]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__2 = s3_folded_gh_hist_10_folded_hist
    [2]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__3 = s3_folded_gh_hist_10_folded_hist
    [3]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__4 = s3_folded_gh_hist_10_folded_hist
    [4]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__5 = s3_folded_gh_hist_10_folded_hist
    [5]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__6 = s3_folded_gh_hist_10_folded_hist
    [6]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__7 = s3_folded_gh_hist_10_folded_hist
    [7]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__8 = s3_folded_gh_hist_10_folded_hist
    [8]; // @[FrontendBundle.scala 280:54]
  wire [8:0] s3_possible_predicted_fhs_res_hist_10_new_folded_hist_xored = {
    s3_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__8,
    s3_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__7,
    s3_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__6,
    s3_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__5,
    s3_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__4,
    s3_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__3,
    s3_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__1,
    s3_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [17:0] s3_possible_predicted_fhs_res_hist_10_new_folded_hist_src_doubled = {
    s3_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__8,
    s3_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__7,
    s3_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__6,
    s3_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__5,
    s3_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__4,
    s3_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__3,
    s3_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__1,
    s3_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__0,
    s3_possible_predicted_fhs_res_hist_10_new_folded_hist_xored}; // @[Cat.scala 31:58]
  wire [8:0] s3_possible_predicted_fhs_res_hist_10_new_folded_hist =
    s3_possible_predicted_fhs_res_hist_10_new_folded_hist_src_doubled[17:9]; // @[FrontendBundle.scala 221:30]
  wire  s3_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__0 = s3_folded_gh_hist_12_folded_hist
    [0]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__1 = s3_folded_gh_hist_12_folded_hist
    [1]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__2 = s3_folded_gh_hist_12_folded_hist
    [2]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__3 = s3_folded_gh_hist_12_folded_hist
    [3]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__4 = s3_folded_gh_hist_12_folded_hist
    [4]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__5 = s3_folded_gh_hist_12_folded_hist
    [5]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__6 = s3_folded_gh_hist_12_folded_hist
    [6]; // @[FrontendBundle.scala 280:54]
  wire [6:0] s3_possible_predicted_fhs_res_hist_12_new_folded_hist_xored = {
    s3_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__6,
    s3_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__5,
    s3_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__4,
    s3_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__3,
    s3_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__1,
    s3_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [13:0] s3_possible_predicted_fhs_res_hist_12_new_folded_hist_src_doubled = {
    s3_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__6,
    s3_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__5,
    s3_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__4,
    s3_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__3,
    s3_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__1,
    s3_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__0,
    s3_possible_predicted_fhs_res_hist_12_new_folded_hist_xored}; // @[Cat.scala 31:58]
  wire [6:0] s3_possible_predicted_fhs_res_hist_12_new_folded_hist =
    s3_possible_predicted_fhs_res_hist_12_new_folded_hist_src_doubled[13:7]; // @[FrontendBundle.scala 221:30]
  wire  s3_possible_predicted_fhs_ob_10_0 = s3_last_br_num_oh[0] & s3_ahead_fh_oldest_bits_afhob_4_bits_0 |
    s3_last_br_num_oh[1] & s3_ahead_fh_oldest_bits_afhob_4_bits_1 | s3_last_br_num_oh[2] &
    s3_ahead_fh_oldest_bits_afhob_4_bits_2; // @[Mux.scala 27:73]
  wire  s3_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__0 = s3_folded_gh_hist_13_folded_hist
    [0]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__1 = s3_folded_gh_hist_13_folded_hist
    [1]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__2 = s3_folded_gh_hist_13_folded_hist
    [2]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__3 = s3_folded_gh_hist_13_folded_hist
    [3]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__4 = s3_folded_gh_hist_13_folded_hist
    [4]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__5 = s3_folded_gh_hist_13_folded_hist
    [5]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__6 = s3_folded_gh_hist_13_folded_hist
    [6]; // @[FrontendBundle.scala 280:54]
  wire [6:0] s3_possible_predicted_fhs_res_hist_13_new_folded_hist_xored = {
    s3_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__6,
    s3_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__5,
    s3_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__4,
    s3_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__3,
    s3_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__1,
    s3_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [13:0] s3_possible_predicted_fhs_res_hist_13_new_folded_hist_src_doubled = {
    s3_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__6,
    s3_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__5,
    s3_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__4,
    s3_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__3,
    s3_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__1,
    s3_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__0,
    s3_possible_predicted_fhs_res_hist_13_new_folded_hist_xored}; // @[Cat.scala 31:58]
  wire [6:0] s3_possible_predicted_fhs_res_hist_13_new_folded_hist =
    s3_possible_predicted_fhs_res_hist_13_new_folded_hist_src_doubled[13:7]; // @[FrontendBundle.scala 221:30]
  wire  s3_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__0 = s3_folded_gh_hist_14_folded_hist
    [0]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__1 = s3_folded_gh_hist_14_folded_hist
    [1]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__2 = s3_folded_gh_hist_14_folded_hist
    [2]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__3 = s3_folded_gh_hist_14_folded_hist
    [3]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__4 = s3_folded_gh_hist_14_folded_hist
    [4]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__5 = s3_folded_gh_hist_14_folded_hist
    [5]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__6 = s3_folded_gh_hist_14_folded_hist
    [6]; // @[FrontendBundle.scala 280:54]
  wire [6:0] s3_possible_predicted_fhs_res_hist_14_new_folded_hist_xored = {
    s3_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__6,
    s3_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__5,
    s3_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__4,
    s3_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__3,
    s3_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__1,
    s3_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [13:0] s3_possible_predicted_fhs_res_hist_14_new_folded_hist_src_doubled = {
    s3_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__6,
    s3_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__5,
    s3_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__4,
    s3_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__3,
    s3_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__1,
    s3_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__0,
    s3_possible_predicted_fhs_res_hist_14_new_folded_hist_xored}; // @[Cat.scala 31:58]
  wire [6:0] s3_possible_predicted_fhs_res_hist_14_new_folded_hist =
    s3_possible_predicted_fhs_res_hist_14_new_folded_hist_src_doubled[13:7]; // @[FrontendBundle.scala 221:30]
  wire  s3_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__0 = s3_folded_gh_hist_15_folded_hist
    [0]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__1 = s3_folded_gh_hist_15_folded_hist
    [1]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__2 = s3_folded_gh_hist_15_folded_hist
    [2]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__3 = s3_folded_gh_hist_15_folded_hist
    [3]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__4 = s3_folded_gh_hist_15_folded_hist
    [4]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__5 = s3_folded_gh_hist_15_folded_hist
    [5]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__6 = s3_folded_gh_hist_15_folded_hist
    [6]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__7 = s3_folded_gh_hist_15_folded_hist
    [7]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__8 = s3_folded_gh_hist_15_folded_hist
    [8]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__9 = s3_folded_gh_hist_15_folded_hist
    [9]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__10 =
    s3_folded_gh_hist_15_folded_hist[10]; // @[FrontendBundle.scala 280:54]
  wire [4:0] s3_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_lo = {
    s3_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__4,
    s3_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__3,
    s3_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__1,
    s3_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [10:0] s3_possible_predicted_fhs_res_hist_15_new_folded_hist_xored = {
    s3_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__10,
    s3_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__9,
    s3_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__8,
    s3_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__7,
    s3_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__6,
    s3_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__5,
    s3_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_lo}; // @[FrontendBundle.scala 258:11]
  wire [21:0] s3_possible_predicted_fhs_res_hist_15_new_folded_hist_src_doubled = {
    s3_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__10,
    s3_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__9,
    s3_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__8,
    s3_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__7,
    s3_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__6,
    s3_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__5,
    s3_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_lo,
    s3_possible_predicted_fhs_res_hist_15_new_folded_hist_xored}; // @[Cat.scala 31:58]
  wire [10:0] s3_possible_predicted_fhs_res_hist_15_new_folded_hist =
    s3_possible_predicted_fhs_res_hist_15_new_folded_hist_src_doubled[21:11]; // @[FrontendBundle.scala 221:30]
  wire  s3_possible_predicted_fhs_ob_13_0 = s3_last_br_num_oh[0] & s3_ahead_fh_oldest_bits_afhob_0_bits_0 |
    s3_last_br_num_oh[1] & s3_ahead_fh_oldest_bits_afhob_0_bits_1 | s3_last_br_num_oh[2] &
    s3_ahead_fh_oldest_bits_afhob_0_bits_2; // @[Mux.scala 27:73]
  wire  s3_possible_predicted_fhs_ob_13_1 = s3_last_br_num_oh[0] & s3_ahead_fh_oldest_bits_afhob_0_bits_1 |
    s3_last_br_num_oh[1] & s3_ahead_fh_oldest_bits_afhob_0_bits_2 | s3_last_br_num_oh[2] &
    s3_ahead_fh_oldest_bits_afhob_0_bits_3; // @[Mux.scala 27:73]
  wire  s3_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__0 = s3_folded_gh_hist_16_folded_hist
    [0]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__1 = s3_folded_gh_hist_16_folded_hist
    [1]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__2 = s3_folded_gh_hist_16_folded_hist
    [2]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__3 = s3_folded_gh_hist_16_folded_hist
    [3]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__4 = s3_folded_gh_hist_16_folded_hist
    [4]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__5 = s3_folded_gh_hist_16_folded_hist
    [5]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__6 = s3_folded_gh_hist_16_folded_hist
    [6]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__7 = s3_folded_gh_hist_16_folded_hist
    [7]; // @[FrontendBundle.scala 280:54]
  wire [7:0] s3_possible_predicted_fhs_res_hist_16_new_folded_hist_xored = {
    s3_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__7,
    s3_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__6,
    s3_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__5,
    s3_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__4,
    s3_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__3,
    s3_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__1,
    s3_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [15:0] s3_possible_predicted_fhs_res_hist_16_new_folded_hist_src_doubled = {
    s3_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__7,
    s3_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__6,
    s3_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__5,
    s3_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__4,
    s3_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__3,
    s3_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__1,
    s3_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__0,
    s3_possible_predicted_fhs_res_hist_16_new_folded_hist_xored}; // @[Cat.scala 31:58]
  wire [7:0] s3_possible_predicted_fhs_res_hist_16_new_folded_hist =
    s3_possible_predicted_fhs_res_hist_16_new_folded_hist_src_doubled[15:8]; // @[FrontendBundle.scala 221:30]
  wire  s3_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__0 = s3_folded_gh_hist_17_folded_hist
    [0]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__1 = s3_folded_gh_hist_17_folded_hist
    [1]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__2 = s3_folded_gh_hist_17_folded_hist
    [2]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__3 = s3_folded_gh_hist_17_folded_hist
    [3]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__4 = s3_folded_gh_hist_17_folded_hist
    [4]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__5 = s3_folded_gh_hist_17_folded_hist
    [5]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__6 = s3_folded_gh_hist_17_folded_hist
    [6]; // @[FrontendBundle.scala 280:54]
  wire  s3_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__7 = s3_folded_gh_hist_17_folded_hist
    [7]; // @[FrontendBundle.scala 280:54]
  wire [7:0] s3_possible_predicted_fhs_res_hist_17_new_folded_hist_xored = {
    s3_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__7,
    s3_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__6,
    s3_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__5,
    s3_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__4,
    s3_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__3,
    s3_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__1,
    s3_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [15:0] s3_possible_predicted_fhs_res_hist_17_new_folded_hist_src_doubled = {
    s3_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__7,
    s3_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__6,
    s3_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__5,
    s3_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__4,
    s3_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__3,
    s3_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__1,
    s3_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__0,
    s3_possible_predicted_fhs_res_hist_17_new_folded_hist_xored}; // @[Cat.scala 31:58]
  wire [7:0] s3_possible_predicted_fhs_res_hist_17_new_folded_hist =
    s3_possible_predicted_fhs_res_hist_17_new_folded_hist_src_doubled[15:8]; // @[FrontendBundle.scala 221:30]
  wire  _s3_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_T_2 =
    predictors_io_out_s3_full_pred_br_taken_mask_0; // @[FrontendBundle.scala 274:80]
  wire [1:0] s3_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1 = {1'h0,
    _s3_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_T_2}; // @[FrontendBundle.scala 274:102]
  wire  s3_possible_predicted_fhs_res_hist_0_new_folded_hist_xored_res_1_6 =
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[1] ^
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__6; // @[FrontendBundle.scala 256:48]
  wire  s3_possible_predicted_fhs_res_hist_0_new_folded_hist_xored_res_1_7 =
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[0] ^ s3_possible_predicted_fhs_ob__0 ^
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__7; // @[FrontendBundle.scala 256:48]
  wire [7:0] s3_possible_predicted_fhs_res_hist_0_new_folded_hist_xored_1 = {
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_xored_res_1_7,
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_xored_res_1_6,
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__5,
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__4,
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__3,
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__1,
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [15:0] s3_possible_predicted_fhs_res_hist_0_new_folded_hist_src_doubled_1 = {
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_xored_res_1_7,
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_xored_res_1_6,
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__5,
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__4,
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__3,
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__1,
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__0,
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_xored_1}; // @[Cat.scala 31:58]
  wire [7:0] s3_possible_predicted_fhs_res_hist_0_new_folded_hist_1 =
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_src_doubled_1[14:7]; // @[FrontendBundle.scala 221:30]
  wire  s3_possible_predicted_fhs_res_hist_1_new_folded_hist_xored_res_1_6 =
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[1] ^
    s3_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__6; // @[FrontendBundle.scala 256:48]
  wire  s3_possible_predicted_fhs_res_hist_1_new_folded_hist_xored_res_1_7 =
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[0] ^ s3_possible_predicted_fhs_ob_1_0 ^
    s3_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__7; // @[FrontendBundle.scala 256:48]
  wire [7:0] s3_possible_predicted_fhs_res_hist_1_new_folded_hist_xored_1 = {
    s3_possible_predicted_fhs_res_hist_1_new_folded_hist_xored_res_1_7,
    s3_possible_predicted_fhs_res_hist_1_new_folded_hist_xored_res_1_6,
    s3_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__5,
    s3_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__4,
    s3_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__3,
    s3_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__1,
    s3_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [15:0] s3_possible_predicted_fhs_res_hist_1_new_folded_hist_src_doubled_1 = {
    s3_possible_predicted_fhs_res_hist_1_new_folded_hist_xored_res_1_7,
    s3_possible_predicted_fhs_res_hist_1_new_folded_hist_xored_res_1_6,
    s3_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__5,
    s3_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__4,
    s3_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__3,
    s3_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__1,
    s3_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__0,
    s3_possible_predicted_fhs_res_hist_1_new_folded_hist_xored_1}; // @[Cat.scala 31:58]
  wire [7:0] s3_possible_predicted_fhs_res_hist_1_new_folded_hist_1 =
    s3_possible_predicted_fhs_res_hist_1_new_folded_hist_src_doubled_1[14:7]; // @[FrontendBundle.scala 221:30]
  wire  s3_possible_predicted_fhs_res_hist_2_new_folded_hist_xored_res_1_6 =
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[1] ^ s3_possible_predicted_fhs_ob_2_0 ^
    s3_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__6; // @[FrontendBundle.scala 256:48]
  wire  s3_possible_predicted_fhs_res_hist_2_new_folded_hist_xored_res_1_7 =
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[0] ^
    s3_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__7; // @[FrontendBundle.scala 256:48]
  wire [7:0] s3_possible_predicted_fhs_res_hist_2_new_folded_hist_xored_1 = {
    s3_possible_predicted_fhs_res_hist_2_new_folded_hist_xored_res_1_7,
    s3_possible_predicted_fhs_res_hist_2_new_folded_hist_xored_res_1_6,
    s3_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__5,
    s3_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__4,
    s3_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__3,
    s3_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__1,
    s3_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [15:0] s3_possible_predicted_fhs_res_hist_2_new_folded_hist_src_doubled_1 = {
    s3_possible_predicted_fhs_res_hist_2_new_folded_hist_xored_res_1_7,
    s3_possible_predicted_fhs_res_hist_2_new_folded_hist_xored_res_1_6,
    s3_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__5,
    s3_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__4,
    s3_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__3,
    s3_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__1,
    s3_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__0,
    s3_possible_predicted_fhs_res_hist_2_new_folded_hist_xored_1}; // @[Cat.scala 31:58]
  wire [7:0] s3_possible_predicted_fhs_res_hist_2_new_folded_hist_1 =
    s3_possible_predicted_fhs_res_hist_2_new_folded_hist_src_doubled_1[14:7]; // @[FrontendBundle.scala 221:30]
  wire  s3_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_res_1_9 =
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[1] ^ s3_possible_predicted_fhs_ob_1_0 ^
    s3_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__9; // @[FrontendBundle.scala 256:48]
  wire  s3_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_res_1_10 =
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[0] ^
    s3_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__10; // @[FrontendBundle.scala 256:48]
  wire [10:0] s3_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_1 = {
    s3_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_res_1_10,
    s3_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_res_1_9,
    s3_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__8,
    s3_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__7,
    s3_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__6,
    s3_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__5,
    s3_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_lo}; // @[FrontendBundle.scala 258:11]
  wire [21:0] s3_possible_predicted_fhs_res_hist_3_new_folded_hist_src_doubled_1 = {
    s3_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_res_1_10,
    s3_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_res_1_9,
    s3_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__8,
    s3_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__7,
    s3_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__6,
    s3_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__5,
    s3_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_lo,
    s3_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_1}; // @[Cat.scala 31:58]
  wire [10:0] s3_possible_predicted_fhs_res_hist_3_new_folded_hist_1 =
    s3_possible_predicted_fhs_res_hist_3_new_folded_hist_src_doubled_1[20:10]; // @[FrontendBundle.scala 221:30]
  wire [4:0] _s3_possible_predicted_fhs_res_hist_4_new_folded_hist_T_2 = {s3_folded_gh_hist_4_folded_hist, 1'h0}; // @[FrontendBundle.scala 290:21]
  wire [4:0] _GEN_11925 = {{4'd0}, predictors_io_out_s3_full_pred_br_taken_mask_0}; // @[FrontendBundle.scala 290:29]
  wire [4:0] _s3_possible_predicted_fhs_res_hist_4_new_folded_hist_T_3 =
    _s3_possible_predicted_fhs_res_hist_4_new_folded_hist_T_2 | _GEN_11925; // @[FrontendBundle.scala 290:29]
  wire [3:0] s3_possible_predicted_fhs_res_hist_4_new_folded_hist_1 =
    _s3_possible_predicted_fhs_res_hist_4_new_folded_hist_T_3[3:0]; // @[FrontendBundle.scala 290:37]
  wire  s3_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_res_1_1 = s3_possible_predicted_fhs_ob_4_0 ^
    s3_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__1; // @[FrontendBundle.scala 256:48]
  wire  s3_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_res_1_9 =
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[1] ^
    s3_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__9; // @[FrontendBundle.scala 256:48]
  wire  s3_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_res_1_10 =
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[0] ^
    s3_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__10; // @[FrontendBundle.scala 256:48]
  wire [4:0] s3_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_lo_1 = {
    s3_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__4,
    s3_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__3,
    s3_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_res_1_1,
    s3_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [10:0] s3_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_1 = {
    s3_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_res_1_10,
    s3_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_res_1_9,
    s3_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__8,
    s3_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__7,
    s3_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__6,
    s3_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__5,
    s3_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_lo_1}; // @[FrontendBundle.scala 258:11]
  wire [21:0] s3_possible_predicted_fhs_res_hist_5_new_folded_hist_src_doubled_1 = {
    s3_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_res_1_10,
    s3_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_res_1_9,
    s3_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__8,
    s3_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__7,
    s3_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__6,
    s3_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__5,
    s3_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_lo_1,
    s3_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_1}; // @[Cat.scala 31:58]
  wire [10:0] s3_possible_predicted_fhs_res_hist_5_new_folded_hist_1 =
    s3_possible_predicted_fhs_res_hist_5_new_folded_hist_src_doubled_1[20:10]; // @[FrontendBundle.scala 221:30]
  wire  s3_possible_predicted_fhs_res_hist_6_new_folded_hist_xored_res_1_3 = s3_possible_predicted_fhs_ob_4_0 ^
    s3_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__3; // @[FrontendBundle.scala 256:48]
  wire  s3_possible_predicted_fhs_res_hist_6_new_folded_hist_xored_res_1_7 =
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[1] ^
    s3_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__7; // @[FrontendBundle.scala 256:48]
  wire  s3_possible_predicted_fhs_res_hist_6_new_folded_hist_xored_res_1_8 =
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[0] ^
    s3_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__8; // @[FrontendBundle.scala 256:48]
  wire [8:0] s3_possible_predicted_fhs_res_hist_6_new_folded_hist_xored_1 = {
    s3_possible_predicted_fhs_res_hist_6_new_folded_hist_xored_res_1_8,
    s3_possible_predicted_fhs_res_hist_6_new_folded_hist_xored_res_1_7,
    s3_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__6,
    s3_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__5,
    s3_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__4,
    s3_possible_predicted_fhs_res_hist_6_new_folded_hist_xored_res_1_3,
    s3_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__1,
    s3_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [17:0] s3_possible_predicted_fhs_res_hist_6_new_folded_hist_src_doubled_1 = {
    s3_possible_predicted_fhs_res_hist_6_new_folded_hist_xored_res_1_8,
    s3_possible_predicted_fhs_res_hist_6_new_folded_hist_xored_res_1_7,
    s3_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__6,
    s3_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__5,
    s3_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__4,
    s3_possible_predicted_fhs_res_hist_6_new_folded_hist_xored_res_1_3,
    s3_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__1,
    s3_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__0,
    s3_possible_predicted_fhs_res_hist_6_new_folded_hist_xored_1}; // @[Cat.scala 31:58]
  wire [8:0] s3_possible_predicted_fhs_res_hist_6_new_folded_hist_1 =
    s3_possible_predicted_fhs_res_hist_6_new_folded_hist_src_doubled_1[16:8]; // @[FrontendBundle.scala 221:30]
  wire  s3_possible_predicted_fhs_res_hist_7_new_folded_hist_xored_res_1_6 = s3_possible_predicted_fhs_ob__0 ^
    s3_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__6; // @[FrontendBundle.scala 256:48]
  wire  s3_possible_predicted_fhs_res_hist_7_new_folded_hist_xored_res_1_7 =
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[1] ^
    s3_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__7; // @[FrontendBundle.scala 256:48]
  wire  s3_possible_predicted_fhs_res_hist_7_new_folded_hist_xored_res_1_8 =
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[0] ^
    s3_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__8; // @[FrontendBundle.scala 256:48]
  wire [8:0] s3_possible_predicted_fhs_res_hist_7_new_folded_hist_xored_1 = {
    s3_possible_predicted_fhs_res_hist_7_new_folded_hist_xored_res_1_8,
    s3_possible_predicted_fhs_res_hist_7_new_folded_hist_xored_res_1_7,
    s3_possible_predicted_fhs_res_hist_7_new_folded_hist_xored_res_1_6,
    s3_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__5,
    s3_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__4,
    s3_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__3,
    s3_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__1,
    s3_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [17:0] s3_possible_predicted_fhs_res_hist_7_new_folded_hist_src_doubled_1 = {
    s3_possible_predicted_fhs_res_hist_7_new_folded_hist_xored_res_1_8,
    s3_possible_predicted_fhs_res_hist_7_new_folded_hist_xored_res_1_7,
    s3_possible_predicted_fhs_res_hist_7_new_folded_hist_xored_res_1_6,
    s3_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__5,
    s3_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__4,
    s3_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__3,
    s3_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__1,
    s3_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__0,
    s3_possible_predicted_fhs_res_hist_7_new_folded_hist_xored_1}; // @[Cat.scala 31:58]
  wire [8:0] s3_possible_predicted_fhs_res_hist_7_new_folded_hist_1 =
    s3_possible_predicted_fhs_res_hist_7_new_folded_hist_src_doubled_1[16:8]; // @[FrontendBundle.scala 221:30]
  wire [8:0] _s3_possible_predicted_fhs_res_hist_8_new_folded_hist_T_2 = {s3_folded_gh_hist_8_folded_hist, 1'h0}; // @[FrontendBundle.scala 290:21]
  wire [8:0] _GEN_11926 = {{8'd0}, predictors_io_out_s3_full_pred_br_taken_mask_0}; // @[FrontendBundle.scala 290:29]
  wire [8:0] _s3_possible_predicted_fhs_res_hist_8_new_folded_hist_T_3 =
    _s3_possible_predicted_fhs_res_hist_8_new_folded_hist_T_2 | _GEN_11926; // @[FrontendBundle.scala 290:29]
  wire [7:0] s3_possible_predicted_fhs_res_hist_8_new_folded_hist_1 =
    _s3_possible_predicted_fhs_res_hist_8_new_folded_hist_T_3[7:0]; // @[FrontendBundle.scala 290:37]
  wire  s3_possible_predicted_fhs_res_hist_9_new_folded_hist_xored_res_1_3 = s3_possible_predicted_fhs_ob_1_0 ^
    s3_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__3; // @[FrontendBundle.scala 256:48]
  wire  s3_possible_predicted_fhs_res_hist_9_new_folded_hist_xored_res_1_5 =
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[1] ^
    s3_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__5; // @[FrontendBundle.scala 256:48]
  wire  s3_possible_predicted_fhs_res_hist_9_new_folded_hist_xored_res_1_6 =
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[0] ^
    s3_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__6; // @[FrontendBundle.scala 256:48]
  wire [6:0] s3_possible_predicted_fhs_res_hist_9_new_folded_hist_xored_1 = {
    s3_possible_predicted_fhs_res_hist_9_new_folded_hist_xored_res_1_6,
    s3_possible_predicted_fhs_res_hist_9_new_folded_hist_xored_res_1_5,
    s3_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__4,
    s3_possible_predicted_fhs_res_hist_9_new_folded_hist_xored_res_1_3,
    s3_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__1,
    s3_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [13:0] s3_possible_predicted_fhs_res_hist_9_new_folded_hist_src_doubled_1 = {
    s3_possible_predicted_fhs_res_hist_9_new_folded_hist_xored_res_1_6,
    s3_possible_predicted_fhs_res_hist_9_new_folded_hist_xored_res_1_5,
    s3_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__4,
    s3_possible_predicted_fhs_res_hist_9_new_folded_hist_xored_res_1_3,
    s3_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__1,
    s3_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__0,
    s3_possible_predicted_fhs_res_hist_9_new_folded_hist_xored_1}; // @[Cat.scala 31:58]
  wire [6:0] s3_possible_predicted_fhs_res_hist_9_new_folded_hist_1 =
    s3_possible_predicted_fhs_res_hist_9_new_folded_hist_src_doubled_1[12:6]; // @[FrontendBundle.scala 221:30]
  wire  s3_possible_predicted_fhs_res_hist_10_new_folded_hist_xored_res_1_4 = s3_possible_predicted_fhs_ob_1_0 ^
    s3_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__4; // @[FrontendBundle.scala 256:48]
  wire  s3_possible_predicted_fhs_res_hist_10_new_folded_hist_xored_res_1_7 =
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[1] ^
    s3_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__7; // @[FrontendBundle.scala 256:48]
  wire  s3_possible_predicted_fhs_res_hist_10_new_folded_hist_xored_res_1_8 =
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[0] ^
    s3_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__8; // @[FrontendBundle.scala 256:48]
  wire [8:0] s3_possible_predicted_fhs_res_hist_10_new_folded_hist_xored_1 = {
    s3_possible_predicted_fhs_res_hist_10_new_folded_hist_xored_res_1_8,
    s3_possible_predicted_fhs_res_hist_10_new_folded_hist_xored_res_1_7,
    s3_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__6,
    s3_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__5,
    s3_possible_predicted_fhs_res_hist_10_new_folded_hist_xored_res_1_4,
    s3_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__3,
    s3_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__1,
    s3_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [17:0] s3_possible_predicted_fhs_res_hist_10_new_folded_hist_src_doubled_1 = {
    s3_possible_predicted_fhs_res_hist_10_new_folded_hist_xored_res_1_8,
    s3_possible_predicted_fhs_res_hist_10_new_folded_hist_xored_res_1_7,
    s3_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__6,
    s3_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__5,
    s3_possible_predicted_fhs_res_hist_10_new_folded_hist_xored_res_1_4,
    s3_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__3,
    s3_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__1,
    s3_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__0,
    s3_possible_predicted_fhs_res_hist_10_new_folded_hist_xored_1}; // @[Cat.scala 31:58]
  wire [8:0] s3_possible_predicted_fhs_res_hist_10_new_folded_hist_1 =
    s3_possible_predicted_fhs_res_hist_10_new_folded_hist_src_doubled_1[16:8]; // @[FrontendBundle.scala 221:30]
  wire [8:0] _s3_possible_predicted_fhs_res_hist_11_new_folded_hist_T_2 = {s3_folded_gh_hist_11_folded_hist, 1'h0}; // @[FrontendBundle.scala 290:21]
  wire [8:0] _s3_possible_predicted_fhs_res_hist_11_new_folded_hist_T_3 =
    _s3_possible_predicted_fhs_res_hist_11_new_folded_hist_T_2 | _GEN_11926; // @[FrontendBundle.scala 290:29]
  wire [7:0] s3_possible_predicted_fhs_res_hist_11_new_folded_hist_1 =
    _s3_possible_predicted_fhs_res_hist_11_new_folded_hist_T_3[7:0]; // @[FrontendBundle.scala 290:37]
  wire  s3_possible_predicted_fhs_res_hist_12_new_folded_hist_xored_res_1_5 =
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[1] ^ s3_possible_predicted_fhs_ob_4_0 ^
    s3_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__5; // @[FrontendBundle.scala 256:48]
  wire  s3_possible_predicted_fhs_res_hist_12_new_folded_hist_xored_res_1_6 =
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[0] ^
    s3_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__6; // @[FrontendBundle.scala 256:48]
  wire [6:0] s3_possible_predicted_fhs_res_hist_12_new_folded_hist_xored_1 = {
    s3_possible_predicted_fhs_res_hist_12_new_folded_hist_xored_res_1_6,
    s3_possible_predicted_fhs_res_hist_12_new_folded_hist_xored_res_1_5,
    s3_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__4,
    s3_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__3,
    s3_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__1,
    s3_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [13:0] s3_possible_predicted_fhs_res_hist_12_new_folded_hist_src_doubled_1 = {
    s3_possible_predicted_fhs_res_hist_12_new_folded_hist_xored_res_1_6,
    s3_possible_predicted_fhs_res_hist_12_new_folded_hist_xored_res_1_5,
    s3_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__4,
    s3_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__3,
    s3_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__1,
    s3_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__0,
    s3_possible_predicted_fhs_res_hist_12_new_folded_hist_xored_1}; // @[Cat.scala 31:58]
  wire [6:0] s3_possible_predicted_fhs_res_hist_12_new_folded_hist_1 =
    s3_possible_predicted_fhs_res_hist_12_new_folded_hist_src_doubled_1[12:6]; // @[FrontendBundle.scala 221:30]
  wire  s3_possible_predicted_fhs_res_hist_13_new_folded_hist_xored_res_1_0 = s3_possible_predicted_fhs_ob_10_0 ^
    s3_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__0; // @[FrontendBundle.scala 256:48]
  wire  s3_possible_predicted_fhs_res_hist_13_new_folded_hist_xored_res_1_5 =
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[1] ^
    s3_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__5; // @[FrontendBundle.scala 256:48]
  wire  s3_possible_predicted_fhs_res_hist_13_new_folded_hist_xored_res_1_6 =
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[0] ^
    s3_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__6; // @[FrontendBundle.scala 256:48]
  wire [6:0] s3_possible_predicted_fhs_res_hist_13_new_folded_hist_xored_1 = {
    s3_possible_predicted_fhs_res_hist_13_new_folded_hist_xored_res_1_6,
    s3_possible_predicted_fhs_res_hist_13_new_folded_hist_xored_res_1_5,
    s3_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__4,
    s3_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__3,
    s3_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__1,
    s3_possible_predicted_fhs_res_hist_13_new_folded_hist_xored_res_1_0}; // @[FrontendBundle.scala 258:11]
  wire [13:0] s3_possible_predicted_fhs_res_hist_13_new_folded_hist_src_doubled_1 = {
    s3_possible_predicted_fhs_res_hist_13_new_folded_hist_xored_res_1_6,
    s3_possible_predicted_fhs_res_hist_13_new_folded_hist_xored_res_1_5,
    s3_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__4,
    s3_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__3,
    s3_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__1,
    s3_possible_predicted_fhs_res_hist_13_new_folded_hist_xored_res_1_0,
    s3_possible_predicted_fhs_res_hist_13_new_folded_hist_xored_1}; // @[Cat.scala 31:58]
  wire [6:0] s3_possible_predicted_fhs_res_hist_13_new_folded_hist_1 =
    s3_possible_predicted_fhs_res_hist_13_new_folded_hist_src_doubled_1[12:6]; // @[FrontendBundle.scala 221:30]
  wire  s3_possible_predicted_fhs_res_hist_14_new_folded_hist_xored_res_1_5 =
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[1] ^
    s3_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__5; // @[FrontendBundle.scala 256:48]
  wire  s3_possible_predicted_fhs_res_hist_14_new_folded_hist_xored_res_1_6 =
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[0] ^ s3_possible_predicted_fhs_ob_2_0 ^
    s3_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__6; // @[FrontendBundle.scala 256:48]
  wire [6:0] s3_possible_predicted_fhs_res_hist_14_new_folded_hist_xored_1 = {
    s3_possible_predicted_fhs_res_hist_14_new_folded_hist_xored_res_1_6,
    s3_possible_predicted_fhs_res_hist_14_new_folded_hist_xored_res_1_5,
    s3_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__4,
    s3_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__3,
    s3_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__1,
    s3_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [13:0] s3_possible_predicted_fhs_res_hist_14_new_folded_hist_src_doubled_1 = {
    s3_possible_predicted_fhs_res_hist_14_new_folded_hist_xored_res_1_6,
    s3_possible_predicted_fhs_res_hist_14_new_folded_hist_xored_res_1_5,
    s3_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__4,
    s3_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__3,
    s3_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__1,
    s3_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__0,
    s3_possible_predicted_fhs_res_hist_14_new_folded_hist_xored_1}; // @[Cat.scala 31:58]
  wire [6:0] s3_possible_predicted_fhs_res_hist_14_new_folded_hist_1 =
    s3_possible_predicted_fhs_res_hist_14_new_folded_hist_src_doubled_1[12:6]; // @[FrontendBundle.scala 221:30]
  wire  s3_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_res_1_8 = s3_possible_predicted_fhs_ob_2_0 ^
    s3_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__8; // @[FrontendBundle.scala 256:48]
  wire  s3_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_res_1_9 =
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[1] ^
    s3_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__9; // @[FrontendBundle.scala 256:48]
  wire  s3_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_res_1_10 =
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[0] ^
    s3_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__10; // @[FrontendBundle.scala 256:48]
  wire [10:0] s3_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_1 = {
    s3_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_res_1_10,
    s3_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_res_1_9,
    s3_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_res_1_8,
    s3_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__7,
    s3_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__6,
    s3_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__5,
    s3_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_lo}; // @[FrontendBundle.scala 258:11]
  wire [21:0] s3_possible_predicted_fhs_res_hist_15_new_folded_hist_src_doubled_1 = {
    s3_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_res_1_10,
    s3_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_res_1_9,
    s3_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_res_1_8,
    s3_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__7,
    s3_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__6,
    s3_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__5,
    s3_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_lo,
    s3_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_1}; // @[Cat.scala 31:58]
  wire [10:0] s3_possible_predicted_fhs_res_hist_15_new_folded_hist_1 =
    s3_possible_predicted_fhs_res_hist_15_new_folded_hist_src_doubled_1[20:10]; // @[FrontendBundle.scala 221:30]
  wire  s3_possible_predicted_fhs_res_hist_16_new_folded_hist_xored_res_1_1 = s3_possible_predicted_fhs_ob_13_0 ^
    s3_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__1; // @[FrontendBundle.scala 256:48]
  wire  s3_possible_predicted_fhs_res_hist_16_new_folded_hist_xored_res_1_6 =
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[1] ^
    s3_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__6; // @[FrontendBundle.scala 256:48]
  wire  s3_possible_predicted_fhs_res_hist_16_new_folded_hist_xored_res_1_7 =
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[0] ^
    s3_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__7; // @[FrontendBundle.scala 256:48]
  wire [7:0] s3_possible_predicted_fhs_res_hist_16_new_folded_hist_xored_1 = {
    s3_possible_predicted_fhs_res_hist_16_new_folded_hist_xored_res_1_7,
    s3_possible_predicted_fhs_res_hist_16_new_folded_hist_xored_res_1_6,
    s3_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__5,
    s3_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__4,
    s3_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__3,
    s3_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_16_new_folded_hist_xored_res_1_1,
    s3_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [15:0] s3_possible_predicted_fhs_res_hist_16_new_folded_hist_src_doubled_1 = {
    s3_possible_predicted_fhs_res_hist_16_new_folded_hist_xored_res_1_7,
    s3_possible_predicted_fhs_res_hist_16_new_folded_hist_xored_res_1_6,
    s3_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__5,
    s3_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__4,
    s3_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__3,
    s3_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_16_new_folded_hist_xored_res_1_1,
    s3_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__0,
    s3_possible_predicted_fhs_res_hist_16_new_folded_hist_xored_1}; // @[Cat.scala 31:58]
  wire [7:0] s3_possible_predicted_fhs_res_hist_16_new_folded_hist_1 =
    s3_possible_predicted_fhs_res_hist_16_new_folded_hist_src_doubled_1[14:7]; // @[FrontendBundle.scala 221:30]
  wire  s3_possible_predicted_fhs_res_hist_17_new_folded_hist_xored_res_1_4 = s3_possible_predicted_fhs_ob_4_0 ^
    s3_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__4; // @[FrontendBundle.scala 256:48]
  wire  s3_possible_predicted_fhs_res_hist_17_new_folded_hist_xored_res_1_6 =
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[1] ^
    s3_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__6; // @[FrontendBundle.scala 256:48]
  wire  s3_possible_predicted_fhs_res_hist_17_new_folded_hist_xored_res_1_7 =
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_1[0] ^
    s3_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__7; // @[FrontendBundle.scala 256:48]
  wire [7:0] s3_possible_predicted_fhs_res_hist_17_new_folded_hist_xored_1 = {
    s3_possible_predicted_fhs_res_hist_17_new_folded_hist_xored_res_1_7,
    s3_possible_predicted_fhs_res_hist_17_new_folded_hist_xored_res_1_6,
    s3_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__5,
    s3_possible_predicted_fhs_res_hist_17_new_folded_hist_xored_res_1_4,
    s3_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__3,
    s3_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__1,
    s3_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [15:0] s3_possible_predicted_fhs_res_hist_17_new_folded_hist_src_doubled_1 = {
    s3_possible_predicted_fhs_res_hist_17_new_folded_hist_xored_res_1_7,
    s3_possible_predicted_fhs_res_hist_17_new_folded_hist_xored_res_1_6,
    s3_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__5,
    s3_possible_predicted_fhs_res_hist_17_new_folded_hist_xored_res_1_4,
    s3_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__3,
    s3_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__1,
    s3_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__0,
    s3_possible_predicted_fhs_res_hist_17_new_folded_hist_xored_1}; // @[Cat.scala 31:58]
  wire [7:0] s3_possible_predicted_fhs_res_hist_17_new_folded_hist_1 =
    s3_possible_predicted_fhs_res_hist_17_new_folded_hist_src_doubled_1[14:7]; // @[FrontendBundle.scala 221:30]
  wire  _s3_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_T_5 =
    predictors_io_out_s3_full_pred_br_taken_mask_1; // @[FrontendBundle.scala 274:80]
  wire [1:0] s3_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2 = {
    _s3_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_T_5,1'h0}; // @[FrontendBundle.scala 274:102]
  wire  s3_possible_predicted_fhs_res_hist_0_new_folded_hist_xored_res_2_6 =
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[1] ^ s3_possible_predicted_fhs_ob__1 ^
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__6; // @[FrontendBundle.scala 256:48]
  wire  s3_possible_predicted_fhs_res_hist_0_new_folded_hist_xored_res_2_7 =
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[0] ^ s3_possible_predicted_fhs_ob__0 ^
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__7; // @[FrontendBundle.scala 256:48]
  wire [7:0] s3_possible_predicted_fhs_res_hist_0_new_folded_hist_xored_2 = {
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_xored_res_2_7,
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_xored_res_2_6,
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__5,
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__4,
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__3,
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__1,
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [15:0] s3_possible_predicted_fhs_res_hist_0_new_folded_hist_src_doubled_2 = {
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_xored_res_2_7,
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_xored_res_2_6,
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__5,
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__4,
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__3,
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__1,
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_original_bits_masked__0,
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_xored_2}; // @[Cat.scala 31:58]
  wire [7:0] s3_possible_predicted_fhs_res_hist_0_new_folded_hist_2 =
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_src_doubled_2[13:6]; // @[FrontendBundle.scala 221:30]
  wire  s3_possible_predicted_fhs_res_hist_1_new_folded_hist_xored_res_2_6 =
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[1] ^ s3_possible_predicted_fhs_ob_1_1 ^
    s3_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__6; // @[FrontendBundle.scala 256:48]
  wire  s3_possible_predicted_fhs_res_hist_1_new_folded_hist_xored_res_2_7 =
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[0] ^ s3_possible_predicted_fhs_ob_1_0 ^
    s3_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__7; // @[FrontendBundle.scala 256:48]
  wire [7:0] s3_possible_predicted_fhs_res_hist_1_new_folded_hist_xored_2 = {
    s3_possible_predicted_fhs_res_hist_1_new_folded_hist_xored_res_2_7,
    s3_possible_predicted_fhs_res_hist_1_new_folded_hist_xored_res_2_6,
    s3_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__5,
    s3_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__4,
    s3_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__3,
    s3_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__1,
    s3_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [15:0] s3_possible_predicted_fhs_res_hist_1_new_folded_hist_src_doubled_2 = {
    s3_possible_predicted_fhs_res_hist_1_new_folded_hist_xored_res_2_7,
    s3_possible_predicted_fhs_res_hist_1_new_folded_hist_xored_res_2_6,
    s3_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__5,
    s3_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__4,
    s3_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__3,
    s3_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__1,
    s3_possible_predicted_fhs_res_hist_1_new_folded_hist_original_bits_masked__0,
    s3_possible_predicted_fhs_res_hist_1_new_folded_hist_xored_2}; // @[Cat.scala 31:58]
  wire [7:0] s3_possible_predicted_fhs_res_hist_1_new_folded_hist_2 =
    s3_possible_predicted_fhs_res_hist_1_new_folded_hist_src_doubled_2[13:6]; // @[FrontendBundle.scala 221:30]
  wire  s3_possible_predicted_fhs_res_hist_2_new_folded_hist_xored_res_2_5 = s3_possible_predicted_fhs_ob_2_1 ^
    s3_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__5; // @[FrontendBundle.scala 256:48]
  wire  s3_possible_predicted_fhs_res_hist_2_new_folded_hist_xored_res_2_6 =
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[1] ^ s3_possible_predicted_fhs_ob_2_0 ^
    s3_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__6; // @[FrontendBundle.scala 256:48]
  wire  s3_possible_predicted_fhs_res_hist_2_new_folded_hist_xored_res_2_7 =
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[0] ^
    s3_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__7; // @[FrontendBundle.scala 256:48]
  wire [7:0] s3_possible_predicted_fhs_res_hist_2_new_folded_hist_xored_2 = {
    s3_possible_predicted_fhs_res_hist_2_new_folded_hist_xored_res_2_7,
    s3_possible_predicted_fhs_res_hist_2_new_folded_hist_xored_res_2_6,
    s3_possible_predicted_fhs_res_hist_2_new_folded_hist_xored_res_2_5,
    s3_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__4,
    s3_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__3,
    s3_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__1,
    s3_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [15:0] s3_possible_predicted_fhs_res_hist_2_new_folded_hist_src_doubled_2 = {
    s3_possible_predicted_fhs_res_hist_2_new_folded_hist_xored_res_2_7,
    s3_possible_predicted_fhs_res_hist_2_new_folded_hist_xored_res_2_6,
    s3_possible_predicted_fhs_res_hist_2_new_folded_hist_xored_res_2_5,
    s3_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__4,
    s3_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__3,
    s3_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__1,
    s3_possible_predicted_fhs_res_hist_2_new_folded_hist_original_bits_masked__0,
    s3_possible_predicted_fhs_res_hist_2_new_folded_hist_xored_2}; // @[Cat.scala 31:58]
  wire [7:0] s3_possible_predicted_fhs_res_hist_2_new_folded_hist_2 =
    s3_possible_predicted_fhs_res_hist_2_new_folded_hist_src_doubled_2[13:6]; // @[FrontendBundle.scala 221:30]
  wire  s3_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_res_2_8 = s3_possible_predicted_fhs_ob_1_1 ^
    s3_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__8; // @[FrontendBundle.scala 256:48]
  wire  s3_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_res_2_9 =
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[1] ^ s3_possible_predicted_fhs_ob_1_0 ^
    s3_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__9; // @[FrontendBundle.scala 256:48]
  wire  s3_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_res_2_10 =
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[0] ^
    s3_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__10; // @[FrontendBundle.scala 256:48]
  wire [10:0] s3_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_2 = {
    s3_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_res_2_10,
    s3_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_res_2_9,
    s3_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_res_2_8,
    s3_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__7,
    s3_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__6,
    s3_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__5,
    s3_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_lo}; // @[FrontendBundle.scala 258:11]
  wire [21:0] s3_possible_predicted_fhs_res_hist_3_new_folded_hist_src_doubled_2 = {
    s3_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_res_2_10,
    s3_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_res_2_9,
    s3_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_res_2_8,
    s3_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__7,
    s3_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__6,
    s3_possible_predicted_fhs_res_hist_3_new_folded_hist_original_bits_masked__5,
    s3_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_lo,
    s3_possible_predicted_fhs_res_hist_3_new_folded_hist_xored_2}; // @[Cat.scala 31:58]
  wire [10:0] s3_possible_predicted_fhs_res_hist_3_new_folded_hist_2 =
    s3_possible_predicted_fhs_res_hist_3_new_folded_hist_src_doubled_2[19:9]; // @[FrontendBundle.scala 221:30]
  wire [5:0] _s3_possible_predicted_fhs_res_hist_4_new_folded_hist_T_4 = {s3_folded_gh_hist_4_folded_hist, 2'h0}; // @[FrontendBundle.scala 290:21]
  wire [5:0] _GEN_11928 = {{5'd0}, predictors_io_out_s3_full_pred_br_taken_mask_1}; // @[FrontendBundle.scala 290:29]
  wire [5:0] _s3_possible_predicted_fhs_res_hist_4_new_folded_hist_T_5 =
    _s3_possible_predicted_fhs_res_hist_4_new_folded_hist_T_4 | _GEN_11928; // @[FrontendBundle.scala 290:29]
  wire [3:0] s3_possible_predicted_fhs_res_hist_4_new_folded_hist_2 =
    _s3_possible_predicted_fhs_res_hist_4_new_folded_hist_T_5[3:0]; // @[FrontendBundle.scala 290:37]
  wire  s3_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_res_2_0 = s3_possible_predicted_fhs_ob_4_1 ^
    s3_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__0; // @[FrontendBundle.scala 256:48]
  wire  s3_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_res_2_9 =
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[1] ^
    s3_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__9; // @[FrontendBundle.scala 256:48]
  wire  s3_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_res_2_10 =
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[0] ^
    s3_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__10; // @[FrontendBundle.scala 256:48]
  wire [4:0] s3_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_lo_2 = {
    s3_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__4,
    s3_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__3,
    s3_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_res_1_1,
    s3_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_res_2_0}; // @[FrontendBundle.scala 258:11]
  wire [10:0] s3_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_2 = {
    s3_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_res_2_10,
    s3_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_res_2_9,
    s3_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__8,
    s3_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__7,
    s3_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__6,
    s3_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__5,
    s3_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_lo_2}; // @[FrontendBundle.scala 258:11]
  wire [21:0] s3_possible_predicted_fhs_res_hist_5_new_folded_hist_src_doubled_2 = {
    s3_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_res_2_10,
    s3_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_res_2_9,
    s3_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__8,
    s3_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__7,
    s3_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__6,
    s3_possible_predicted_fhs_res_hist_5_new_folded_hist_original_bits_masked__5,
    s3_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_lo_2,
    s3_possible_predicted_fhs_res_hist_5_new_folded_hist_xored_2}; // @[Cat.scala 31:58]
  wire [10:0] s3_possible_predicted_fhs_res_hist_5_new_folded_hist_2 =
    s3_possible_predicted_fhs_res_hist_5_new_folded_hist_src_doubled_2[19:9]; // @[FrontendBundle.scala 221:30]
  wire  s3_possible_predicted_fhs_res_hist_6_new_folded_hist_xored_res_2_2 = s3_possible_predicted_fhs_ob_4_1 ^
    s3_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__2; // @[FrontendBundle.scala 256:48]
  wire  s3_possible_predicted_fhs_res_hist_6_new_folded_hist_xored_res_2_7 =
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[1] ^
    s3_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__7; // @[FrontendBundle.scala 256:48]
  wire  s3_possible_predicted_fhs_res_hist_6_new_folded_hist_xored_res_2_8 =
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[0] ^
    s3_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__8; // @[FrontendBundle.scala 256:48]
  wire [8:0] s3_possible_predicted_fhs_res_hist_6_new_folded_hist_xored_2 = {
    s3_possible_predicted_fhs_res_hist_6_new_folded_hist_xored_res_2_8,
    s3_possible_predicted_fhs_res_hist_6_new_folded_hist_xored_res_2_7,
    s3_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__6,
    s3_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__5,
    s3_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__4,
    s3_possible_predicted_fhs_res_hist_6_new_folded_hist_xored_res_1_3,
    s3_possible_predicted_fhs_res_hist_6_new_folded_hist_xored_res_2_2,
    s3_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__1,
    s3_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [17:0] s3_possible_predicted_fhs_res_hist_6_new_folded_hist_src_doubled_2 = {
    s3_possible_predicted_fhs_res_hist_6_new_folded_hist_xored_res_2_8,
    s3_possible_predicted_fhs_res_hist_6_new_folded_hist_xored_res_2_7,
    s3_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__6,
    s3_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__5,
    s3_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__4,
    s3_possible_predicted_fhs_res_hist_6_new_folded_hist_xored_res_1_3,
    s3_possible_predicted_fhs_res_hist_6_new_folded_hist_xored_res_2_2,
    s3_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__1,
    s3_possible_predicted_fhs_res_hist_6_new_folded_hist_original_bits_masked__0,
    s3_possible_predicted_fhs_res_hist_6_new_folded_hist_xored_2}; // @[Cat.scala 31:58]
  wire [8:0] s3_possible_predicted_fhs_res_hist_6_new_folded_hist_2 =
    s3_possible_predicted_fhs_res_hist_6_new_folded_hist_src_doubled_2[15:7]; // @[FrontendBundle.scala 221:30]
  wire  s3_possible_predicted_fhs_res_hist_7_new_folded_hist_xored_res_2_5 = s3_possible_predicted_fhs_ob__1 ^
    s3_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__5; // @[FrontendBundle.scala 256:48]
  wire  s3_possible_predicted_fhs_res_hist_7_new_folded_hist_xored_res_2_7 =
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[1] ^
    s3_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__7; // @[FrontendBundle.scala 256:48]
  wire  s3_possible_predicted_fhs_res_hist_7_new_folded_hist_xored_res_2_8 =
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[0] ^
    s3_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__8; // @[FrontendBundle.scala 256:48]
  wire [8:0] s3_possible_predicted_fhs_res_hist_7_new_folded_hist_xored_2 = {
    s3_possible_predicted_fhs_res_hist_7_new_folded_hist_xored_res_2_8,
    s3_possible_predicted_fhs_res_hist_7_new_folded_hist_xored_res_2_7,
    s3_possible_predicted_fhs_res_hist_7_new_folded_hist_xored_res_1_6,
    s3_possible_predicted_fhs_res_hist_7_new_folded_hist_xored_res_2_5,
    s3_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__4,
    s3_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__3,
    s3_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__1,
    s3_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [17:0] s3_possible_predicted_fhs_res_hist_7_new_folded_hist_src_doubled_2 = {
    s3_possible_predicted_fhs_res_hist_7_new_folded_hist_xored_res_2_8,
    s3_possible_predicted_fhs_res_hist_7_new_folded_hist_xored_res_2_7,
    s3_possible_predicted_fhs_res_hist_7_new_folded_hist_xored_res_1_6,
    s3_possible_predicted_fhs_res_hist_7_new_folded_hist_xored_res_2_5,
    s3_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__4,
    s3_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__3,
    s3_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__1,
    s3_possible_predicted_fhs_res_hist_7_new_folded_hist_original_bits_masked__0,
    s3_possible_predicted_fhs_res_hist_7_new_folded_hist_xored_2}; // @[Cat.scala 31:58]
  wire [8:0] s3_possible_predicted_fhs_res_hist_7_new_folded_hist_2 =
    s3_possible_predicted_fhs_res_hist_7_new_folded_hist_src_doubled_2[15:7]; // @[FrontendBundle.scala 221:30]
  wire [9:0] _s3_possible_predicted_fhs_res_hist_8_new_folded_hist_T_4 = {s3_folded_gh_hist_8_folded_hist, 2'h0}; // @[FrontendBundle.scala 290:21]
  wire [9:0] _GEN_11929 = {{9'd0}, predictors_io_out_s3_full_pred_br_taken_mask_1}; // @[FrontendBundle.scala 290:29]
  wire [9:0] _s3_possible_predicted_fhs_res_hist_8_new_folded_hist_T_5 =
    _s3_possible_predicted_fhs_res_hist_8_new_folded_hist_T_4 | _GEN_11929; // @[FrontendBundle.scala 290:29]
  wire [7:0] s3_possible_predicted_fhs_res_hist_8_new_folded_hist_2 =
    _s3_possible_predicted_fhs_res_hist_8_new_folded_hist_T_5[7:0]; // @[FrontendBundle.scala 290:37]
  wire  s3_possible_predicted_fhs_res_hist_9_new_folded_hist_xored_res_2_2 = s3_possible_predicted_fhs_ob_1_1 ^
    s3_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__2; // @[FrontendBundle.scala 256:48]
  wire  s3_possible_predicted_fhs_res_hist_9_new_folded_hist_xored_res_2_5 =
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[1] ^
    s3_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__5; // @[FrontendBundle.scala 256:48]
  wire  s3_possible_predicted_fhs_res_hist_9_new_folded_hist_xored_res_2_6 =
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[0] ^
    s3_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__6; // @[FrontendBundle.scala 256:48]
  wire [6:0] s3_possible_predicted_fhs_res_hist_9_new_folded_hist_xored_2 = {
    s3_possible_predicted_fhs_res_hist_9_new_folded_hist_xored_res_2_6,
    s3_possible_predicted_fhs_res_hist_9_new_folded_hist_xored_res_2_5,
    s3_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__4,
    s3_possible_predicted_fhs_res_hist_9_new_folded_hist_xored_res_1_3,
    s3_possible_predicted_fhs_res_hist_9_new_folded_hist_xored_res_2_2,
    s3_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__1,
    s3_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [13:0] s3_possible_predicted_fhs_res_hist_9_new_folded_hist_src_doubled_2 = {
    s3_possible_predicted_fhs_res_hist_9_new_folded_hist_xored_res_2_6,
    s3_possible_predicted_fhs_res_hist_9_new_folded_hist_xored_res_2_5,
    s3_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__4,
    s3_possible_predicted_fhs_res_hist_9_new_folded_hist_xored_res_1_3,
    s3_possible_predicted_fhs_res_hist_9_new_folded_hist_xored_res_2_2,
    s3_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__1,
    s3_possible_predicted_fhs_res_hist_9_new_folded_hist_original_bits_masked__0,
    s3_possible_predicted_fhs_res_hist_9_new_folded_hist_xored_2}; // @[Cat.scala 31:58]
  wire [6:0] s3_possible_predicted_fhs_res_hist_9_new_folded_hist_2 =
    s3_possible_predicted_fhs_res_hist_9_new_folded_hist_src_doubled_2[11:5]; // @[FrontendBundle.scala 221:30]
  wire  s3_possible_predicted_fhs_res_hist_10_new_folded_hist_xored_res_2_3 = s3_possible_predicted_fhs_ob_1_1 ^
    s3_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__3; // @[FrontendBundle.scala 256:48]
  wire  s3_possible_predicted_fhs_res_hist_10_new_folded_hist_xored_res_2_7 =
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[1] ^
    s3_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__7; // @[FrontendBundle.scala 256:48]
  wire  s3_possible_predicted_fhs_res_hist_10_new_folded_hist_xored_res_2_8 =
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[0] ^
    s3_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__8; // @[FrontendBundle.scala 256:48]
  wire [8:0] s3_possible_predicted_fhs_res_hist_10_new_folded_hist_xored_2 = {
    s3_possible_predicted_fhs_res_hist_10_new_folded_hist_xored_res_2_8,
    s3_possible_predicted_fhs_res_hist_10_new_folded_hist_xored_res_2_7,
    s3_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__6,
    s3_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__5,
    s3_possible_predicted_fhs_res_hist_10_new_folded_hist_xored_res_1_4,
    s3_possible_predicted_fhs_res_hist_10_new_folded_hist_xored_res_2_3,
    s3_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__1,
    s3_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [17:0] s3_possible_predicted_fhs_res_hist_10_new_folded_hist_src_doubled_2 = {
    s3_possible_predicted_fhs_res_hist_10_new_folded_hist_xored_res_2_8,
    s3_possible_predicted_fhs_res_hist_10_new_folded_hist_xored_res_2_7,
    s3_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__6,
    s3_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__5,
    s3_possible_predicted_fhs_res_hist_10_new_folded_hist_xored_res_1_4,
    s3_possible_predicted_fhs_res_hist_10_new_folded_hist_xored_res_2_3,
    s3_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__1,
    s3_possible_predicted_fhs_res_hist_10_new_folded_hist_original_bits_masked__0,
    s3_possible_predicted_fhs_res_hist_10_new_folded_hist_xored_2}; // @[Cat.scala 31:58]
  wire [8:0] s3_possible_predicted_fhs_res_hist_10_new_folded_hist_2 =
    s3_possible_predicted_fhs_res_hist_10_new_folded_hist_src_doubled_2[15:7]; // @[FrontendBundle.scala 221:30]
  wire [9:0] _s3_possible_predicted_fhs_res_hist_11_new_folded_hist_T_4 = {s3_folded_gh_hist_11_folded_hist, 2'h0}; // @[FrontendBundle.scala 290:21]
  wire [9:0] _s3_possible_predicted_fhs_res_hist_11_new_folded_hist_T_5 =
    _s3_possible_predicted_fhs_res_hist_11_new_folded_hist_T_4 | _GEN_11929; // @[FrontendBundle.scala 290:29]
  wire [7:0] s3_possible_predicted_fhs_res_hist_11_new_folded_hist_2 =
    _s3_possible_predicted_fhs_res_hist_11_new_folded_hist_T_5[7:0]; // @[FrontendBundle.scala 290:37]
  wire  s3_possible_predicted_fhs_res_hist_12_new_folded_hist_xored_res_2_4 = s3_possible_predicted_fhs_ob_4_1 ^
    s3_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__4; // @[FrontendBundle.scala 256:48]
  wire  s3_possible_predicted_fhs_res_hist_12_new_folded_hist_xored_res_2_5 =
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[1] ^ s3_possible_predicted_fhs_ob_4_0 ^
    s3_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__5; // @[FrontendBundle.scala 256:48]
  wire  s3_possible_predicted_fhs_res_hist_12_new_folded_hist_xored_res_2_6 =
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[0] ^
    s3_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__6; // @[FrontendBundle.scala 256:48]
  wire [6:0] s3_possible_predicted_fhs_res_hist_12_new_folded_hist_xored_2 = {
    s3_possible_predicted_fhs_res_hist_12_new_folded_hist_xored_res_2_6,
    s3_possible_predicted_fhs_res_hist_12_new_folded_hist_xored_res_2_5,
    s3_possible_predicted_fhs_res_hist_12_new_folded_hist_xored_res_2_4,
    s3_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__3,
    s3_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__1,
    s3_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [13:0] s3_possible_predicted_fhs_res_hist_12_new_folded_hist_src_doubled_2 = {
    s3_possible_predicted_fhs_res_hist_12_new_folded_hist_xored_res_2_6,
    s3_possible_predicted_fhs_res_hist_12_new_folded_hist_xored_res_2_5,
    s3_possible_predicted_fhs_res_hist_12_new_folded_hist_xored_res_2_4,
    s3_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__3,
    s3_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__1,
    s3_possible_predicted_fhs_res_hist_12_new_folded_hist_original_bits_masked__0,
    s3_possible_predicted_fhs_res_hist_12_new_folded_hist_xored_2}; // @[Cat.scala 31:58]
  wire [6:0] s3_possible_predicted_fhs_res_hist_12_new_folded_hist_2 =
    s3_possible_predicted_fhs_res_hist_12_new_folded_hist_src_doubled_2[11:5]; // @[FrontendBundle.scala 221:30]
  wire  s3_possible_predicted_fhs_res_hist_13_new_folded_hist_xored_res_2_5 =
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[1] ^
    s3_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__5; // @[FrontendBundle.scala 256:48]
  wire [6:0] s3_possible_predicted_fhs_res_hist_13_new_folded_hist_xored_2 = {
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[0],
    s3_possible_predicted_fhs_res_hist_13_new_folded_hist_xored_res_2_5,
    s3_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__4,
    s3_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__3,
    s3_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__1,
    s3_possible_predicted_fhs_res_hist_13_new_folded_hist_xored_res_1_0}; // @[FrontendBundle.scala 258:11]
  wire [13:0] s3_possible_predicted_fhs_res_hist_13_new_folded_hist_src_doubled_2 = {
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[0],
    s3_possible_predicted_fhs_res_hist_13_new_folded_hist_xored_res_2_5,
    s3_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__4,
    s3_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__3,
    s3_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_13_new_folded_hist_original_bits_masked__1,
    s3_possible_predicted_fhs_res_hist_13_new_folded_hist_xored_res_1_0,
    s3_possible_predicted_fhs_res_hist_13_new_folded_hist_xored_2}; // @[Cat.scala 31:58]
  wire [6:0] s3_possible_predicted_fhs_res_hist_13_new_folded_hist_2 =
    s3_possible_predicted_fhs_res_hist_13_new_folded_hist_src_doubled_2[11:5]; // @[FrontendBundle.scala 221:30]
  wire  s3_possible_predicted_fhs_res_hist_14_new_folded_hist_xored_res_2_5 =
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[1] ^ s3_possible_predicted_fhs_ob_2_1 ^
    s3_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__5; // @[FrontendBundle.scala 256:48]
  wire  s3_possible_predicted_fhs_res_hist_14_new_folded_hist_xored_res_2_6 =
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[0] ^ s3_possible_predicted_fhs_ob_2_0 ^
    s3_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__6; // @[FrontendBundle.scala 256:48]
  wire [6:0] s3_possible_predicted_fhs_res_hist_14_new_folded_hist_xored_2 = {
    s3_possible_predicted_fhs_res_hist_14_new_folded_hist_xored_res_2_6,
    s3_possible_predicted_fhs_res_hist_14_new_folded_hist_xored_res_2_5,
    s3_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__4,
    s3_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__3,
    s3_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__1,
    s3_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [13:0] s3_possible_predicted_fhs_res_hist_14_new_folded_hist_src_doubled_2 = {
    s3_possible_predicted_fhs_res_hist_14_new_folded_hist_xored_res_2_6,
    s3_possible_predicted_fhs_res_hist_14_new_folded_hist_xored_res_2_5,
    s3_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__4,
    s3_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__3,
    s3_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__1,
    s3_possible_predicted_fhs_res_hist_14_new_folded_hist_original_bits_masked__0,
    s3_possible_predicted_fhs_res_hist_14_new_folded_hist_xored_2}; // @[Cat.scala 31:58]
  wire [6:0] s3_possible_predicted_fhs_res_hist_14_new_folded_hist_2 =
    s3_possible_predicted_fhs_res_hist_14_new_folded_hist_src_doubled_2[11:5]; // @[FrontendBundle.scala 221:30]
  wire  s3_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_res_2_7 = s3_possible_predicted_fhs_ob_2_1 ^
    s3_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__7; // @[FrontendBundle.scala 256:48]
  wire  s3_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_res_2_9 =
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[1] ^
    s3_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__9; // @[FrontendBundle.scala 256:48]
  wire  s3_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_res_2_10 =
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[0] ^
    s3_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__10; // @[FrontendBundle.scala 256:48]
  wire [10:0] s3_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_2 = {
    s3_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_res_2_10,
    s3_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_res_2_9,
    s3_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_res_1_8,
    s3_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_res_2_7,
    s3_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__6,
    s3_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__5,
    s3_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_lo}; // @[FrontendBundle.scala 258:11]
  wire [21:0] s3_possible_predicted_fhs_res_hist_15_new_folded_hist_src_doubled_2 = {
    s3_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_res_2_10,
    s3_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_res_2_9,
    s3_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_res_1_8,
    s3_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_res_2_7,
    s3_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__6,
    s3_possible_predicted_fhs_res_hist_15_new_folded_hist_original_bits_masked__5,
    s3_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_lo,
    s3_possible_predicted_fhs_res_hist_15_new_folded_hist_xored_2}; // @[Cat.scala 31:58]
  wire [10:0] s3_possible_predicted_fhs_res_hist_15_new_folded_hist_2 =
    s3_possible_predicted_fhs_res_hist_15_new_folded_hist_src_doubled_2[19:9]; // @[FrontendBundle.scala 221:30]
  wire  s3_possible_predicted_fhs_res_hist_16_new_folded_hist_xored_res_2_0 = s3_possible_predicted_fhs_ob_13_1 ^
    s3_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__0; // @[FrontendBundle.scala 256:48]
  wire  s3_possible_predicted_fhs_res_hist_16_new_folded_hist_xored_res_2_6 =
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[1] ^
    s3_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__6; // @[FrontendBundle.scala 256:48]
  wire  s3_possible_predicted_fhs_res_hist_16_new_folded_hist_xored_res_2_7 =
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[0] ^
    s3_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__7; // @[FrontendBundle.scala 256:48]
  wire [7:0] s3_possible_predicted_fhs_res_hist_16_new_folded_hist_xored_2 = {
    s3_possible_predicted_fhs_res_hist_16_new_folded_hist_xored_res_2_7,
    s3_possible_predicted_fhs_res_hist_16_new_folded_hist_xored_res_2_6,
    s3_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__5,
    s3_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__4,
    s3_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__3,
    s3_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_16_new_folded_hist_xored_res_1_1,
    s3_possible_predicted_fhs_res_hist_16_new_folded_hist_xored_res_2_0}; // @[FrontendBundle.scala 258:11]
  wire [15:0] s3_possible_predicted_fhs_res_hist_16_new_folded_hist_src_doubled_2 = {
    s3_possible_predicted_fhs_res_hist_16_new_folded_hist_xored_res_2_7,
    s3_possible_predicted_fhs_res_hist_16_new_folded_hist_xored_res_2_6,
    s3_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__5,
    s3_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__4,
    s3_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__3,
    s3_possible_predicted_fhs_res_hist_16_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_16_new_folded_hist_xored_res_1_1,
    s3_possible_predicted_fhs_res_hist_16_new_folded_hist_xored_res_2_0,
    s3_possible_predicted_fhs_res_hist_16_new_folded_hist_xored_2}; // @[Cat.scala 31:58]
  wire [7:0] s3_possible_predicted_fhs_res_hist_16_new_folded_hist_2 =
    s3_possible_predicted_fhs_res_hist_16_new_folded_hist_src_doubled_2[13:6]; // @[FrontendBundle.scala 221:30]
  wire  s3_possible_predicted_fhs_res_hist_17_new_folded_hist_xored_res_2_3 = s3_possible_predicted_fhs_ob_4_1 ^
    s3_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__3; // @[FrontendBundle.scala 256:48]
  wire  s3_possible_predicted_fhs_res_hist_17_new_folded_hist_xored_res_2_6 =
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[1] ^
    s3_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__6; // @[FrontendBundle.scala 256:48]
  wire  s3_possible_predicted_fhs_res_hist_17_new_folded_hist_xored_res_2_7 =
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_newest_bits_masked_2[0] ^
    s3_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__7; // @[FrontendBundle.scala 256:48]
  wire [7:0] s3_possible_predicted_fhs_res_hist_17_new_folded_hist_xored_2 = {
    s3_possible_predicted_fhs_res_hist_17_new_folded_hist_xored_res_2_7,
    s3_possible_predicted_fhs_res_hist_17_new_folded_hist_xored_res_2_6,
    s3_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__5,
    s3_possible_predicted_fhs_res_hist_17_new_folded_hist_xored_res_1_4,
    s3_possible_predicted_fhs_res_hist_17_new_folded_hist_xored_res_2_3,
    s3_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__1,
    s3_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [15:0] s3_possible_predicted_fhs_res_hist_17_new_folded_hist_src_doubled_2 = {
    s3_possible_predicted_fhs_res_hist_17_new_folded_hist_xored_res_2_7,
    s3_possible_predicted_fhs_res_hist_17_new_folded_hist_xored_res_2_6,
    s3_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__5,
    s3_possible_predicted_fhs_res_hist_17_new_folded_hist_xored_res_1_4,
    s3_possible_predicted_fhs_res_hist_17_new_folded_hist_xored_res_2_3,
    s3_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__2,
    s3_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__1,
    s3_possible_predicted_fhs_res_hist_17_new_folded_hist_original_bits_masked__0,
    s3_possible_predicted_fhs_res_hist_17_new_folded_hist_xored_2}; // @[Cat.scala 31:58]
  wire [7:0] s3_possible_predicted_fhs_res_hist_17_new_folded_hist_2 =
    s3_possible_predicted_fhs_res_hist_17_new_folded_hist_src_doubled_2[13:6]; // @[FrontendBundle.scala 221:30]
  wire [7:0] _s3_predicted_fh_T_61 = _s3_predicted_ghist_ptr_T_4 ? s3_possible_predicted_fhs_res_hist_0_new_folded_hist
     : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _s3_predicted_fh_T_62 = _s3_predicted_ghist_ptr_T_32 ?
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _s3_predicted_fh_T_63 = _s3_predicted_ghist_ptr_T_60 ?
    s3_possible_predicted_fhs_res_hist_0_new_folded_hist_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _s3_predicted_fh_T_64 = _s3_predicted_fh_T_61 | _s3_predicted_fh_T_62; // @[Mux.scala 27:73]
  wire [7:0] _s3_predicted_fh_T_66 = _s3_predicted_ghist_ptr_T_4 ? s3_possible_predicted_fhs_res_hist_1_new_folded_hist
     : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _s3_predicted_fh_T_67 = _s3_predicted_ghist_ptr_T_32 ?
    s3_possible_predicted_fhs_res_hist_1_new_folded_hist_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _s3_predicted_fh_T_68 = _s3_predicted_ghist_ptr_T_60 ?
    s3_possible_predicted_fhs_res_hist_1_new_folded_hist_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _s3_predicted_fh_T_69 = _s3_predicted_fh_T_66 | _s3_predicted_fh_T_67; // @[Mux.scala 27:73]
  wire [7:0] _s3_predicted_fh_T_71 = _s3_predicted_ghist_ptr_T_4 ? s3_possible_predicted_fhs_res_hist_2_new_folded_hist
     : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _s3_predicted_fh_T_72 = _s3_predicted_ghist_ptr_T_32 ?
    s3_possible_predicted_fhs_res_hist_2_new_folded_hist_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _s3_predicted_fh_T_73 = _s3_predicted_ghist_ptr_T_60 ?
    s3_possible_predicted_fhs_res_hist_2_new_folded_hist_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _s3_predicted_fh_T_74 = _s3_predicted_fh_T_71 | _s3_predicted_fh_T_72; // @[Mux.scala 27:73]
  wire [10:0] _s3_predicted_fh_T_76 = _s3_predicted_ghist_ptr_T_4 ? s3_possible_predicted_fhs_res_hist_3_new_folded_hist
     : 11'h0; // @[Mux.scala 27:73]
  wire [10:0] _s3_predicted_fh_T_77 = _s3_predicted_ghist_ptr_T_32 ?
    s3_possible_predicted_fhs_res_hist_3_new_folded_hist_1 : 11'h0; // @[Mux.scala 27:73]
  wire [10:0] _s3_predicted_fh_T_78 = _s3_predicted_ghist_ptr_T_60 ?
    s3_possible_predicted_fhs_res_hist_3_new_folded_hist_2 : 11'h0; // @[Mux.scala 27:73]
  wire [10:0] _s3_predicted_fh_T_79 = _s3_predicted_fh_T_76 | _s3_predicted_fh_T_77; // @[Mux.scala 27:73]
  wire [3:0] _s3_predicted_fh_T_81 = _s3_predicted_ghist_ptr_T_4 ? s3_folded_gh_hist_4_folded_hist : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _s3_predicted_fh_T_82 = _s3_predicted_ghist_ptr_T_32 ?
    s3_possible_predicted_fhs_res_hist_4_new_folded_hist_1 : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _s3_predicted_fh_T_83 = _s3_predicted_ghist_ptr_T_60 ?
    s3_possible_predicted_fhs_res_hist_4_new_folded_hist_2 : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _s3_predicted_fh_T_84 = _s3_predicted_fh_T_81 | _s3_predicted_fh_T_82; // @[Mux.scala 27:73]
  wire [10:0] _s3_predicted_fh_T_86 = _s3_predicted_ghist_ptr_T_4 ? s3_possible_predicted_fhs_res_hist_5_new_folded_hist
     : 11'h0; // @[Mux.scala 27:73]
  wire [10:0] _s3_predicted_fh_T_87 = _s3_predicted_ghist_ptr_T_32 ?
    s3_possible_predicted_fhs_res_hist_5_new_folded_hist_1 : 11'h0; // @[Mux.scala 27:73]
  wire [10:0] _s3_predicted_fh_T_88 = _s3_predicted_ghist_ptr_T_60 ?
    s3_possible_predicted_fhs_res_hist_5_new_folded_hist_2 : 11'h0; // @[Mux.scala 27:73]
  wire [10:0] _s3_predicted_fh_T_89 = _s3_predicted_fh_T_86 | _s3_predicted_fh_T_87; // @[Mux.scala 27:73]
  wire [8:0] _s3_predicted_fh_T_91 = _s3_predicted_ghist_ptr_T_4 ? s3_possible_predicted_fhs_res_hist_6_new_folded_hist
     : 9'h0; // @[Mux.scala 27:73]
  wire [8:0] _s3_predicted_fh_T_92 = _s3_predicted_ghist_ptr_T_32 ?
    s3_possible_predicted_fhs_res_hist_6_new_folded_hist_1 : 9'h0; // @[Mux.scala 27:73]
  wire [8:0] _s3_predicted_fh_T_93 = _s3_predicted_ghist_ptr_T_60 ?
    s3_possible_predicted_fhs_res_hist_6_new_folded_hist_2 : 9'h0; // @[Mux.scala 27:73]
  wire [8:0] _s3_predicted_fh_T_94 = _s3_predicted_fh_T_91 | _s3_predicted_fh_T_92; // @[Mux.scala 27:73]
  wire [8:0] _s3_predicted_fh_T_96 = _s3_predicted_ghist_ptr_T_4 ? s3_possible_predicted_fhs_res_hist_7_new_folded_hist
     : 9'h0; // @[Mux.scala 27:73]
  wire [8:0] _s3_predicted_fh_T_97 = _s3_predicted_ghist_ptr_T_32 ?
    s3_possible_predicted_fhs_res_hist_7_new_folded_hist_1 : 9'h0; // @[Mux.scala 27:73]
  wire [8:0] _s3_predicted_fh_T_98 = _s3_predicted_ghist_ptr_T_60 ?
    s3_possible_predicted_fhs_res_hist_7_new_folded_hist_2 : 9'h0; // @[Mux.scala 27:73]
  wire [8:0] _s3_predicted_fh_T_99 = _s3_predicted_fh_T_96 | _s3_predicted_fh_T_97; // @[Mux.scala 27:73]
  wire [7:0] _s3_predicted_fh_T_101 = _s3_predicted_ghist_ptr_T_4 ? s3_folded_gh_hist_8_folded_hist : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _s3_predicted_fh_T_102 = _s3_predicted_ghist_ptr_T_32 ?
    s3_possible_predicted_fhs_res_hist_8_new_folded_hist_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _s3_predicted_fh_T_103 = _s3_predicted_ghist_ptr_T_60 ?
    s3_possible_predicted_fhs_res_hist_8_new_folded_hist_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _s3_predicted_fh_T_104 = _s3_predicted_fh_T_101 | _s3_predicted_fh_T_102; // @[Mux.scala 27:73]
  wire [6:0] _s3_predicted_fh_T_106 = _s3_predicted_ghist_ptr_T_4 ? s3_possible_predicted_fhs_res_hist_9_new_folded_hist
     : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _s3_predicted_fh_T_107 = _s3_predicted_ghist_ptr_T_32 ?
    s3_possible_predicted_fhs_res_hist_9_new_folded_hist_1 : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _s3_predicted_fh_T_108 = _s3_predicted_ghist_ptr_T_60 ?
    s3_possible_predicted_fhs_res_hist_9_new_folded_hist_2 : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _s3_predicted_fh_T_109 = _s3_predicted_fh_T_106 | _s3_predicted_fh_T_107; // @[Mux.scala 27:73]
  wire [8:0] _s3_predicted_fh_T_111 = _s3_predicted_ghist_ptr_T_4 ?
    s3_possible_predicted_fhs_res_hist_10_new_folded_hist : 9'h0; // @[Mux.scala 27:73]
  wire [8:0] _s3_predicted_fh_T_112 = _s3_predicted_ghist_ptr_T_32 ?
    s3_possible_predicted_fhs_res_hist_10_new_folded_hist_1 : 9'h0; // @[Mux.scala 27:73]
  wire [8:0] _s3_predicted_fh_T_113 = _s3_predicted_ghist_ptr_T_60 ?
    s3_possible_predicted_fhs_res_hist_10_new_folded_hist_2 : 9'h0; // @[Mux.scala 27:73]
  wire [8:0] _s3_predicted_fh_T_114 = _s3_predicted_fh_T_111 | _s3_predicted_fh_T_112; // @[Mux.scala 27:73]
  wire [7:0] _s3_predicted_fh_T_116 = _s3_predicted_ghist_ptr_T_4 ? s3_folded_gh_hist_11_folded_hist : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _s3_predicted_fh_T_117 = _s3_predicted_ghist_ptr_T_32 ?
    s3_possible_predicted_fhs_res_hist_11_new_folded_hist_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _s3_predicted_fh_T_118 = _s3_predicted_ghist_ptr_T_60 ?
    s3_possible_predicted_fhs_res_hist_11_new_folded_hist_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _s3_predicted_fh_T_119 = _s3_predicted_fh_T_116 | _s3_predicted_fh_T_117; // @[Mux.scala 27:73]
  wire [6:0] _s3_predicted_fh_T_121 = _s3_predicted_ghist_ptr_T_4 ?
    s3_possible_predicted_fhs_res_hist_12_new_folded_hist : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _s3_predicted_fh_T_122 = _s3_predicted_ghist_ptr_T_32 ?
    s3_possible_predicted_fhs_res_hist_12_new_folded_hist_1 : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _s3_predicted_fh_T_123 = _s3_predicted_ghist_ptr_T_60 ?
    s3_possible_predicted_fhs_res_hist_12_new_folded_hist_2 : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _s3_predicted_fh_T_124 = _s3_predicted_fh_T_121 | _s3_predicted_fh_T_122; // @[Mux.scala 27:73]
  wire [6:0] _s3_predicted_fh_T_126 = _s3_predicted_ghist_ptr_T_4 ?
    s3_possible_predicted_fhs_res_hist_13_new_folded_hist : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _s3_predicted_fh_T_127 = _s3_predicted_ghist_ptr_T_32 ?
    s3_possible_predicted_fhs_res_hist_13_new_folded_hist_1 : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _s3_predicted_fh_T_128 = _s3_predicted_ghist_ptr_T_60 ?
    s3_possible_predicted_fhs_res_hist_13_new_folded_hist_2 : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _s3_predicted_fh_T_129 = _s3_predicted_fh_T_126 | _s3_predicted_fh_T_127; // @[Mux.scala 27:73]
  wire [6:0] _s3_predicted_fh_T_131 = _s3_predicted_ghist_ptr_T_4 ?
    s3_possible_predicted_fhs_res_hist_14_new_folded_hist : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _s3_predicted_fh_T_132 = _s3_predicted_ghist_ptr_T_32 ?
    s3_possible_predicted_fhs_res_hist_14_new_folded_hist_1 : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _s3_predicted_fh_T_133 = _s3_predicted_ghist_ptr_T_60 ?
    s3_possible_predicted_fhs_res_hist_14_new_folded_hist_2 : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _s3_predicted_fh_T_134 = _s3_predicted_fh_T_131 | _s3_predicted_fh_T_132; // @[Mux.scala 27:73]
  wire [10:0] _s3_predicted_fh_T_136 = _s3_predicted_ghist_ptr_T_4 ?
    s3_possible_predicted_fhs_res_hist_15_new_folded_hist : 11'h0; // @[Mux.scala 27:73]
  wire [10:0] _s3_predicted_fh_T_137 = _s3_predicted_ghist_ptr_T_32 ?
    s3_possible_predicted_fhs_res_hist_15_new_folded_hist_1 : 11'h0; // @[Mux.scala 27:73]
  wire [10:0] _s3_predicted_fh_T_138 = _s3_predicted_ghist_ptr_T_60 ?
    s3_possible_predicted_fhs_res_hist_15_new_folded_hist_2 : 11'h0; // @[Mux.scala 27:73]
  wire [10:0] _s3_predicted_fh_T_139 = _s3_predicted_fh_T_136 | _s3_predicted_fh_T_137; // @[Mux.scala 27:73]
  wire [7:0] _s3_predicted_fh_T_141 = _s3_predicted_ghist_ptr_T_4 ?
    s3_possible_predicted_fhs_res_hist_16_new_folded_hist : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _s3_predicted_fh_T_142 = _s3_predicted_ghist_ptr_T_32 ?
    s3_possible_predicted_fhs_res_hist_16_new_folded_hist_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _s3_predicted_fh_T_143 = _s3_predicted_ghist_ptr_T_60 ?
    s3_possible_predicted_fhs_res_hist_16_new_folded_hist_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _s3_predicted_fh_T_144 = _s3_predicted_fh_T_141 | _s3_predicted_fh_T_142; // @[Mux.scala 27:73]
  wire [7:0] _s3_predicted_fh_T_146 = _s3_predicted_ghist_ptr_T_4 ?
    s3_possible_predicted_fhs_res_hist_17_new_folded_hist : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _s3_predicted_fh_T_147 = _s3_predicted_ghist_ptr_T_32 ?
    s3_possible_predicted_fhs_res_hist_17_new_folded_hist_1 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _s3_predicted_fh_T_148 = _s3_predicted_ghist_ptr_T_60 ?
    s3_possible_predicted_fhs_res_hist_17_new_folded_hist_2 : 8'h0; // @[Mux.scala 27:73]
  wire [7:0] _s3_predicted_fh_T_149 = _s3_predicted_fh_T_146 | _s3_predicted_fh_T_147; // @[Mux.scala 27:73]
  wire [8:0] new_value_40 = s3_ghist_ptr_value + 8'h74; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_241 = {1'h0,new_value_40}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_40 = $signed(_diff_T_241) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_40 = $signed(diff_40) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_80 = $signed(_diff_T_241) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_81 = reverse_flag_40 ? _new_ptr_value_T_80 : {{1'd0}, new_value_40}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_41 = s3_ghist_ptr_value + 8'h6; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_247 = {1'h0,new_value_41}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_41 = $signed(_diff_T_247) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_41 = $signed(diff_41) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_82 = $signed(_diff_T_247) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_83 = reverse_flag_41 ? _new_ptr_value_T_82 : {{1'd0}, new_value_41}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_42 = s3_ghist_ptr_value + 8'hb; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_253 = {1'h0,new_value_42}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_42 = $signed(_diff_T_253) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_42 = $signed(diff_42) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_84 = $signed(_diff_T_253) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_85 = reverse_flag_42 ? _new_ptr_value_T_84 : {{1'd0}, new_value_42}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_43 = s3_ghist_ptr_value + 8'hf; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_259 = {1'h0,new_value_43}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_43 = $signed(_diff_T_259) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_43 = $signed(diff_43) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_86 = $signed(_diff_T_259) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_87 = reverse_flag_43 ? _new_ptr_value_T_86 : {{1'd0}, new_value_43}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_44 = s3_ghist_ptr_value + 8'h1e; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_265 = {1'h0,new_value_44}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_44 = $signed(_diff_T_265) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_44 = $signed(diff_44) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_88 = $signed(_diff_T_265) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_89 = reverse_flag_44 ? _new_ptr_value_T_88 : {{1'd0}, new_value_44}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_45 = s3_ghist_ptr_value + 8'h75; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_271 = {1'h0,new_value_45}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_45 = $signed(_diff_T_271) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_45 = $signed(diff_45) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_90 = $signed(_diff_T_271) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_91 = reverse_flag_45 ? _new_ptr_value_T_90 : {{1'd0}, new_value_45}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_46 = s3_ghist_ptr_value + 8'h7; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_277 = {1'h0,new_value_46}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_46 = $signed(_diff_T_277) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_46 = $signed(diff_46) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_92 = $signed(_diff_T_277) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_93 = reverse_flag_46 ? _new_ptr_value_T_92 : {{1'd0}, new_value_46}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_47 = s3_ghist_ptr_value + 8'h76; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_283 = {1'h0,new_value_47}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_47 = $signed(_diff_T_283) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_47 = $signed(diff_47) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_94 = $signed(_diff_T_283) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_95 = reverse_flag_47 ? _new_ptr_value_T_94 : {{1'd0}, new_value_47}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_48 = s3_ghist_ptr_value + 8'h1d; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_289 = {1'h0,new_value_48}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_48 = $signed(_diff_T_289) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_48 = $signed(diff_48) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_96 = $signed(_diff_T_289) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_97 = reverse_flag_48 ? _new_ptr_value_T_96 : {{1'd0}, new_value_48}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_49 = s3_ghist_ptr_value + 8'ha; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_295 = {1'h0,new_value_49}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_49 = $signed(_diff_T_295) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_49 = $signed(diff_49) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_98 = $signed(_diff_T_295) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_99 = reverse_flag_49 ? _new_ptr_value_T_98 : {{1'd0}, new_value_49}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_50 = s3_ghist_ptr_value + 8'he; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_301 = {1'h0,new_value_50}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_50 = $signed(_diff_T_301) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_50 = $signed(diff_50) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_100 = $signed(_diff_T_301) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_101 = reverse_flag_50 ? _new_ptr_value_T_100 : {{1'd0}, new_value_50}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_51 = s3_ghist_ptr_value + 8'h77; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_307 = {1'h0,new_value_51}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_51 = $signed(_diff_T_307) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_51 = $signed(diff_51) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_102 = $signed(_diff_T_307) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_103 = reverse_flag_51 ? _new_ptr_value_T_102 : {{1'd0}, new_value_51}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_52 = s3_ghist_ptr_value + 8'hd; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_313 = {1'h0,new_value_52}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_52 = $signed(_diff_T_313) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_52 = $signed(diff_52) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_104 = $signed(_diff_T_313) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_105 = reverse_flag_52 ? _new_ptr_value_T_104 : {{1'd0}, new_value_52}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_53 = s3_ghist_ptr_value + 8'h8; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_319 = {1'h0,new_value_53}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_53 = $signed(_diff_T_319) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_53 = $signed(diff_53) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_106 = $signed(_diff_T_319) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_107 = reverse_flag_53 ? _new_ptr_value_T_106 : {{1'd0}, new_value_53}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_54 = s3_ghist_ptr_value + 8'h20; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_325 = {1'h0,new_value_54}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_54 = $signed(_diff_T_325) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_54 = $signed(diff_54) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_108 = $signed(_diff_T_325) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_109 = reverse_flag_54 ? _new_ptr_value_T_108 : {{1'd0}, new_value_54}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_55 = s3_ghist_ptr_value + 8'hc; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_331 = {1'h0,new_value_55}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_55 = $signed(_diff_T_331) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_55 = $signed(diff_55) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_110 = $signed(_diff_T_331) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_111 = reverse_flag_55 ? _new_ptr_value_T_110 : {{1'd0}, new_value_55}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_56 = s3_ghist_ptr_value + 8'h9; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_337 = {1'h0,new_value_56}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_56 = $signed(_diff_T_337) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_56 = $signed(diff_56) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_112 = $signed(_diff_T_337) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_113 = reverse_flag_56 ? _new_ptr_value_T_112 : {{1'd0}, new_value_56}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_57 = s3_ghist_ptr_value + 8'h1f; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_343 = {1'h0,new_value_57}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_57 = $signed(_diff_T_343) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_57 = $signed(diff_57) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_114 = $signed(_diff_T_343) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_115 = reverse_flag_57 ? _new_ptr_value_T_114 : {{1'd0}, new_value_57}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_58 = s3_ghist_ptr_value + 8'h5; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_349 = {1'h0,new_value_58}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_58 = $signed(_diff_T_349) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_58 = $signed(diff_58) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_116 = $signed(_diff_T_349) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_117 = reverse_flag_58 ? _new_ptr_value_T_116 : {{1'd0}, new_value_58}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_59 = s3_ghist_ptr_value + 8'h10; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_355 = {1'h0,new_value_59}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_59 = $signed(_diff_T_355) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_59 = $signed(diff_59) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_118 = $signed(_diff_T_355) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_119 = reverse_flag_59 ? _new_ptr_value_T_118 : {{1'd0}, new_value_59}; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] new_ptr_49_value = _new_ptr_value_T_99[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_5920 = 8'h1 == new_ptr_49_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5921 = 8'h2 == new_ptr_49_value ? ghv_2 : _GEN_5920; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5922 = 8'h3 == new_ptr_49_value ? ghv_3 : _GEN_5921; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5923 = 8'h4 == new_ptr_49_value ? ghv_4 : _GEN_5922; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5924 = 8'h5 == new_ptr_49_value ? ghv_5 : _GEN_5923; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5925 = 8'h6 == new_ptr_49_value ? ghv_6 : _GEN_5924; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5926 = 8'h7 == new_ptr_49_value ? ghv_7 : _GEN_5925; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5927 = 8'h8 == new_ptr_49_value ? ghv_8 : _GEN_5926; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5928 = 8'h9 == new_ptr_49_value ? ghv_9 : _GEN_5927; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5929 = 8'ha == new_ptr_49_value ? ghv_10 : _GEN_5928; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5930 = 8'hb == new_ptr_49_value ? ghv_11 : _GEN_5929; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5931 = 8'hc == new_ptr_49_value ? ghv_12 : _GEN_5930; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5932 = 8'hd == new_ptr_49_value ? ghv_13 : _GEN_5931; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5933 = 8'he == new_ptr_49_value ? ghv_14 : _GEN_5932; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5934 = 8'hf == new_ptr_49_value ? ghv_15 : _GEN_5933; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5935 = 8'h10 == new_ptr_49_value ? ghv_16 : _GEN_5934; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5936 = 8'h11 == new_ptr_49_value ? ghv_17 : _GEN_5935; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5937 = 8'h12 == new_ptr_49_value ? ghv_18 : _GEN_5936; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5938 = 8'h13 == new_ptr_49_value ? ghv_19 : _GEN_5937; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5939 = 8'h14 == new_ptr_49_value ? ghv_20 : _GEN_5938; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5940 = 8'h15 == new_ptr_49_value ? ghv_21 : _GEN_5939; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5941 = 8'h16 == new_ptr_49_value ? ghv_22 : _GEN_5940; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5942 = 8'h17 == new_ptr_49_value ? ghv_23 : _GEN_5941; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5943 = 8'h18 == new_ptr_49_value ? ghv_24 : _GEN_5942; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5944 = 8'h19 == new_ptr_49_value ? ghv_25 : _GEN_5943; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5945 = 8'h1a == new_ptr_49_value ? ghv_26 : _GEN_5944; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5946 = 8'h1b == new_ptr_49_value ? ghv_27 : _GEN_5945; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5947 = 8'h1c == new_ptr_49_value ? ghv_28 : _GEN_5946; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5948 = 8'h1d == new_ptr_49_value ? ghv_29 : _GEN_5947; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5949 = 8'h1e == new_ptr_49_value ? ghv_30 : _GEN_5948; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5950 = 8'h1f == new_ptr_49_value ? ghv_31 : _GEN_5949; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5951 = 8'h20 == new_ptr_49_value ? ghv_32 : _GEN_5950; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5952 = 8'h21 == new_ptr_49_value ? ghv_33 : _GEN_5951; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5953 = 8'h22 == new_ptr_49_value ? ghv_34 : _GEN_5952; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5954 = 8'h23 == new_ptr_49_value ? ghv_35 : _GEN_5953; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5955 = 8'h24 == new_ptr_49_value ? ghv_36 : _GEN_5954; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5956 = 8'h25 == new_ptr_49_value ? ghv_37 : _GEN_5955; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5957 = 8'h26 == new_ptr_49_value ? ghv_38 : _GEN_5956; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5958 = 8'h27 == new_ptr_49_value ? ghv_39 : _GEN_5957; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5959 = 8'h28 == new_ptr_49_value ? ghv_40 : _GEN_5958; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5960 = 8'h29 == new_ptr_49_value ? ghv_41 : _GEN_5959; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5961 = 8'h2a == new_ptr_49_value ? ghv_42 : _GEN_5960; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5962 = 8'h2b == new_ptr_49_value ? ghv_43 : _GEN_5961; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5963 = 8'h2c == new_ptr_49_value ? ghv_44 : _GEN_5962; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5964 = 8'h2d == new_ptr_49_value ? ghv_45 : _GEN_5963; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5965 = 8'h2e == new_ptr_49_value ? ghv_46 : _GEN_5964; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5966 = 8'h2f == new_ptr_49_value ? ghv_47 : _GEN_5965; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5967 = 8'h30 == new_ptr_49_value ? ghv_48 : _GEN_5966; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5968 = 8'h31 == new_ptr_49_value ? ghv_49 : _GEN_5967; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5969 = 8'h32 == new_ptr_49_value ? ghv_50 : _GEN_5968; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5970 = 8'h33 == new_ptr_49_value ? ghv_51 : _GEN_5969; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5971 = 8'h34 == new_ptr_49_value ? ghv_52 : _GEN_5970; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5972 = 8'h35 == new_ptr_49_value ? ghv_53 : _GEN_5971; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5973 = 8'h36 == new_ptr_49_value ? ghv_54 : _GEN_5972; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5974 = 8'h37 == new_ptr_49_value ? ghv_55 : _GEN_5973; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5975 = 8'h38 == new_ptr_49_value ? ghv_56 : _GEN_5974; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5976 = 8'h39 == new_ptr_49_value ? ghv_57 : _GEN_5975; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5977 = 8'h3a == new_ptr_49_value ? ghv_58 : _GEN_5976; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5978 = 8'h3b == new_ptr_49_value ? ghv_59 : _GEN_5977; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5979 = 8'h3c == new_ptr_49_value ? ghv_60 : _GEN_5978; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5980 = 8'h3d == new_ptr_49_value ? ghv_61 : _GEN_5979; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5981 = 8'h3e == new_ptr_49_value ? ghv_62 : _GEN_5980; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5982 = 8'h3f == new_ptr_49_value ? ghv_63 : _GEN_5981; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5983 = 8'h40 == new_ptr_49_value ? ghv_64 : _GEN_5982; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5984 = 8'h41 == new_ptr_49_value ? ghv_65 : _GEN_5983; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5985 = 8'h42 == new_ptr_49_value ? ghv_66 : _GEN_5984; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5986 = 8'h43 == new_ptr_49_value ? ghv_67 : _GEN_5985; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5987 = 8'h44 == new_ptr_49_value ? ghv_68 : _GEN_5986; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5988 = 8'h45 == new_ptr_49_value ? ghv_69 : _GEN_5987; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5989 = 8'h46 == new_ptr_49_value ? ghv_70 : _GEN_5988; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5990 = 8'h47 == new_ptr_49_value ? ghv_71 : _GEN_5989; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5991 = 8'h48 == new_ptr_49_value ? ghv_72 : _GEN_5990; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5992 = 8'h49 == new_ptr_49_value ? ghv_73 : _GEN_5991; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5993 = 8'h4a == new_ptr_49_value ? ghv_74 : _GEN_5992; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5994 = 8'h4b == new_ptr_49_value ? ghv_75 : _GEN_5993; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5995 = 8'h4c == new_ptr_49_value ? ghv_76 : _GEN_5994; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5996 = 8'h4d == new_ptr_49_value ? ghv_77 : _GEN_5995; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5997 = 8'h4e == new_ptr_49_value ? ghv_78 : _GEN_5996; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5998 = 8'h4f == new_ptr_49_value ? ghv_79 : _GEN_5997; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_5999 = 8'h50 == new_ptr_49_value ? ghv_80 : _GEN_5998; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6000 = 8'h51 == new_ptr_49_value ? ghv_81 : _GEN_5999; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6001 = 8'h52 == new_ptr_49_value ? ghv_82 : _GEN_6000; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6002 = 8'h53 == new_ptr_49_value ? ghv_83 : _GEN_6001; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6003 = 8'h54 == new_ptr_49_value ? ghv_84 : _GEN_6002; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6004 = 8'h55 == new_ptr_49_value ? ghv_85 : _GEN_6003; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6005 = 8'h56 == new_ptr_49_value ? ghv_86 : _GEN_6004; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6006 = 8'h57 == new_ptr_49_value ? ghv_87 : _GEN_6005; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6007 = 8'h58 == new_ptr_49_value ? ghv_88 : _GEN_6006; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6008 = 8'h59 == new_ptr_49_value ? ghv_89 : _GEN_6007; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6009 = 8'h5a == new_ptr_49_value ? ghv_90 : _GEN_6008; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6010 = 8'h5b == new_ptr_49_value ? ghv_91 : _GEN_6009; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6011 = 8'h5c == new_ptr_49_value ? ghv_92 : _GEN_6010; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6012 = 8'h5d == new_ptr_49_value ? ghv_93 : _GEN_6011; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6013 = 8'h5e == new_ptr_49_value ? ghv_94 : _GEN_6012; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6014 = 8'h5f == new_ptr_49_value ? ghv_95 : _GEN_6013; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6015 = 8'h60 == new_ptr_49_value ? ghv_96 : _GEN_6014; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6016 = 8'h61 == new_ptr_49_value ? ghv_97 : _GEN_6015; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6017 = 8'h62 == new_ptr_49_value ? ghv_98 : _GEN_6016; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6018 = 8'h63 == new_ptr_49_value ? ghv_99 : _GEN_6017; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6019 = 8'h64 == new_ptr_49_value ? ghv_100 : _GEN_6018; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6020 = 8'h65 == new_ptr_49_value ? ghv_101 : _GEN_6019; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6021 = 8'h66 == new_ptr_49_value ? ghv_102 : _GEN_6020; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6022 = 8'h67 == new_ptr_49_value ? ghv_103 : _GEN_6021; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6023 = 8'h68 == new_ptr_49_value ? ghv_104 : _GEN_6022; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6024 = 8'h69 == new_ptr_49_value ? ghv_105 : _GEN_6023; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6025 = 8'h6a == new_ptr_49_value ? ghv_106 : _GEN_6024; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6026 = 8'h6b == new_ptr_49_value ? ghv_107 : _GEN_6025; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6027 = 8'h6c == new_ptr_49_value ? ghv_108 : _GEN_6026; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6028 = 8'h6d == new_ptr_49_value ? ghv_109 : _GEN_6027; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6029 = 8'h6e == new_ptr_49_value ? ghv_110 : _GEN_6028; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6030 = 8'h6f == new_ptr_49_value ? ghv_111 : _GEN_6029; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6031 = 8'h70 == new_ptr_49_value ? ghv_112 : _GEN_6030; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6032 = 8'h71 == new_ptr_49_value ? ghv_113 : _GEN_6031; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6033 = 8'h72 == new_ptr_49_value ? ghv_114 : _GEN_6032; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6034 = 8'h73 == new_ptr_49_value ? ghv_115 : _GEN_6033; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6035 = 8'h74 == new_ptr_49_value ? ghv_116 : _GEN_6034; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6036 = 8'h75 == new_ptr_49_value ? ghv_117 : _GEN_6035; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6037 = 8'h76 == new_ptr_49_value ? ghv_118 : _GEN_6036; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6038 = 8'h77 == new_ptr_49_value ? ghv_119 : _GEN_6037; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6039 = 8'h78 == new_ptr_49_value ? ghv_120 : _GEN_6038; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6040 = 8'h79 == new_ptr_49_value ? ghv_121 : _GEN_6039; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6041 = 8'h7a == new_ptr_49_value ? ghv_122 : _GEN_6040; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6042 = 8'h7b == new_ptr_49_value ? ghv_123 : _GEN_6041; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6043 = 8'h7c == new_ptr_49_value ? ghv_124 : _GEN_6042; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6044 = 8'h7d == new_ptr_49_value ? ghv_125 : _GEN_6043; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6045 = 8'h7e == new_ptr_49_value ? ghv_126 : _GEN_6044; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6046 = 8'h7f == new_ptr_49_value ? ghv_127 : _GEN_6045; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6047 = 8'h80 == new_ptr_49_value ? ghv_128 : _GEN_6046; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6048 = 8'h81 == new_ptr_49_value ? ghv_129 : _GEN_6047; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6049 = 8'h82 == new_ptr_49_value ? ghv_130 : _GEN_6048; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6050 = 8'h83 == new_ptr_49_value ? ghv_131 : _GEN_6049; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6051 = 8'h84 == new_ptr_49_value ? ghv_132 : _GEN_6050; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6052 = 8'h85 == new_ptr_49_value ? ghv_133 : _GEN_6051; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6053 = 8'h86 == new_ptr_49_value ? ghv_134 : _GEN_6052; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6054 = 8'h87 == new_ptr_49_value ? ghv_135 : _GEN_6053; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6055 = 8'h88 == new_ptr_49_value ? ghv_136 : _GEN_6054; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6056 = 8'h89 == new_ptr_49_value ? ghv_137 : _GEN_6055; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6057 = 8'h8a == new_ptr_49_value ? ghv_138 : _GEN_6056; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6058 = 8'h8b == new_ptr_49_value ? ghv_139 : _GEN_6057; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6059 = 8'h8c == new_ptr_49_value ? ghv_140 : _GEN_6058; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6060 = 8'h8d == new_ptr_49_value ? ghv_141 : _GEN_6059; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6061 = 8'h8e == new_ptr_49_value ? ghv_142 : _GEN_6060; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_56_value = _new_ptr_value_T_113[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_6064 = 8'h1 == new_ptr_56_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6065 = 8'h2 == new_ptr_56_value ? ghv_2 : _GEN_6064; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6066 = 8'h3 == new_ptr_56_value ? ghv_3 : _GEN_6065; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6067 = 8'h4 == new_ptr_56_value ? ghv_4 : _GEN_6066; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6068 = 8'h5 == new_ptr_56_value ? ghv_5 : _GEN_6067; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6069 = 8'h6 == new_ptr_56_value ? ghv_6 : _GEN_6068; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6070 = 8'h7 == new_ptr_56_value ? ghv_7 : _GEN_6069; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6071 = 8'h8 == new_ptr_56_value ? ghv_8 : _GEN_6070; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6072 = 8'h9 == new_ptr_56_value ? ghv_9 : _GEN_6071; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6073 = 8'ha == new_ptr_56_value ? ghv_10 : _GEN_6072; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6074 = 8'hb == new_ptr_56_value ? ghv_11 : _GEN_6073; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6075 = 8'hc == new_ptr_56_value ? ghv_12 : _GEN_6074; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6076 = 8'hd == new_ptr_56_value ? ghv_13 : _GEN_6075; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6077 = 8'he == new_ptr_56_value ? ghv_14 : _GEN_6076; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6078 = 8'hf == new_ptr_56_value ? ghv_15 : _GEN_6077; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6079 = 8'h10 == new_ptr_56_value ? ghv_16 : _GEN_6078; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6080 = 8'h11 == new_ptr_56_value ? ghv_17 : _GEN_6079; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6081 = 8'h12 == new_ptr_56_value ? ghv_18 : _GEN_6080; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6082 = 8'h13 == new_ptr_56_value ? ghv_19 : _GEN_6081; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6083 = 8'h14 == new_ptr_56_value ? ghv_20 : _GEN_6082; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6084 = 8'h15 == new_ptr_56_value ? ghv_21 : _GEN_6083; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6085 = 8'h16 == new_ptr_56_value ? ghv_22 : _GEN_6084; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6086 = 8'h17 == new_ptr_56_value ? ghv_23 : _GEN_6085; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6087 = 8'h18 == new_ptr_56_value ? ghv_24 : _GEN_6086; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6088 = 8'h19 == new_ptr_56_value ? ghv_25 : _GEN_6087; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6089 = 8'h1a == new_ptr_56_value ? ghv_26 : _GEN_6088; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6090 = 8'h1b == new_ptr_56_value ? ghv_27 : _GEN_6089; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6091 = 8'h1c == new_ptr_56_value ? ghv_28 : _GEN_6090; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6092 = 8'h1d == new_ptr_56_value ? ghv_29 : _GEN_6091; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6093 = 8'h1e == new_ptr_56_value ? ghv_30 : _GEN_6092; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6094 = 8'h1f == new_ptr_56_value ? ghv_31 : _GEN_6093; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6095 = 8'h20 == new_ptr_56_value ? ghv_32 : _GEN_6094; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6096 = 8'h21 == new_ptr_56_value ? ghv_33 : _GEN_6095; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6097 = 8'h22 == new_ptr_56_value ? ghv_34 : _GEN_6096; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6098 = 8'h23 == new_ptr_56_value ? ghv_35 : _GEN_6097; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6099 = 8'h24 == new_ptr_56_value ? ghv_36 : _GEN_6098; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6100 = 8'h25 == new_ptr_56_value ? ghv_37 : _GEN_6099; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6101 = 8'h26 == new_ptr_56_value ? ghv_38 : _GEN_6100; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6102 = 8'h27 == new_ptr_56_value ? ghv_39 : _GEN_6101; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6103 = 8'h28 == new_ptr_56_value ? ghv_40 : _GEN_6102; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6104 = 8'h29 == new_ptr_56_value ? ghv_41 : _GEN_6103; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6105 = 8'h2a == new_ptr_56_value ? ghv_42 : _GEN_6104; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6106 = 8'h2b == new_ptr_56_value ? ghv_43 : _GEN_6105; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6107 = 8'h2c == new_ptr_56_value ? ghv_44 : _GEN_6106; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6108 = 8'h2d == new_ptr_56_value ? ghv_45 : _GEN_6107; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6109 = 8'h2e == new_ptr_56_value ? ghv_46 : _GEN_6108; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6110 = 8'h2f == new_ptr_56_value ? ghv_47 : _GEN_6109; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6111 = 8'h30 == new_ptr_56_value ? ghv_48 : _GEN_6110; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6112 = 8'h31 == new_ptr_56_value ? ghv_49 : _GEN_6111; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6113 = 8'h32 == new_ptr_56_value ? ghv_50 : _GEN_6112; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6114 = 8'h33 == new_ptr_56_value ? ghv_51 : _GEN_6113; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6115 = 8'h34 == new_ptr_56_value ? ghv_52 : _GEN_6114; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6116 = 8'h35 == new_ptr_56_value ? ghv_53 : _GEN_6115; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6117 = 8'h36 == new_ptr_56_value ? ghv_54 : _GEN_6116; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6118 = 8'h37 == new_ptr_56_value ? ghv_55 : _GEN_6117; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6119 = 8'h38 == new_ptr_56_value ? ghv_56 : _GEN_6118; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6120 = 8'h39 == new_ptr_56_value ? ghv_57 : _GEN_6119; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6121 = 8'h3a == new_ptr_56_value ? ghv_58 : _GEN_6120; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6122 = 8'h3b == new_ptr_56_value ? ghv_59 : _GEN_6121; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6123 = 8'h3c == new_ptr_56_value ? ghv_60 : _GEN_6122; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6124 = 8'h3d == new_ptr_56_value ? ghv_61 : _GEN_6123; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6125 = 8'h3e == new_ptr_56_value ? ghv_62 : _GEN_6124; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6126 = 8'h3f == new_ptr_56_value ? ghv_63 : _GEN_6125; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6127 = 8'h40 == new_ptr_56_value ? ghv_64 : _GEN_6126; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6128 = 8'h41 == new_ptr_56_value ? ghv_65 : _GEN_6127; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6129 = 8'h42 == new_ptr_56_value ? ghv_66 : _GEN_6128; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6130 = 8'h43 == new_ptr_56_value ? ghv_67 : _GEN_6129; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6131 = 8'h44 == new_ptr_56_value ? ghv_68 : _GEN_6130; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6132 = 8'h45 == new_ptr_56_value ? ghv_69 : _GEN_6131; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6133 = 8'h46 == new_ptr_56_value ? ghv_70 : _GEN_6132; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6134 = 8'h47 == new_ptr_56_value ? ghv_71 : _GEN_6133; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6135 = 8'h48 == new_ptr_56_value ? ghv_72 : _GEN_6134; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6136 = 8'h49 == new_ptr_56_value ? ghv_73 : _GEN_6135; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6137 = 8'h4a == new_ptr_56_value ? ghv_74 : _GEN_6136; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6138 = 8'h4b == new_ptr_56_value ? ghv_75 : _GEN_6137; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6139 = 8'h4c == new_ptr_56_value ? ghv_76 : _GEN_6138; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6140 = 8'h4d == new_ptr_56_value ? ghv_77 : _GEN_6139; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6141 = 8'h4e == new_ptr_56_value ? ghv_78 : _GEN_6140; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6142 = 8'h4f == new_ptr_56_value ? ghv_79 : _GEN_6141; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6143 = 8'h50 == new_ptr_56_value ? ghv_80 : _GEN_6142; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6144 = 8'h51 == new_ptr_56_value ? ghv_81 : _GEN_6143; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6145 = 8'h52 == new_ptr_56_value ? ghv_82 : _GEN_6144; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6146 = 8'h53 == new_ptr_56_value ? ghv_83 : _GEN_6145; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6147 = 8'h54 == new_ptr_56_value ? ghv_84 : _GEN_6146; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6148 = 8'h55 == new_ptr_56_value ? ghv_85 : _GEN_6147; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6149 = 8'h56 == new_ptr_56_value ? ghv_86 : _GEN_6148; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6150 = 8'h57 == new_ptr_56_value ? ghv_87 : _GEN_6149; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6151 = 8'h58 == new_ptr_56_value ? ghv_88 : _GEN_6150; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6152 = 8'h59 == new_ptr_56_value ? ghv_89 : _GEN_6151; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6153 = 8'h5a == new_ptr_56_value ? ghv_90 : _GEN_6152; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6154 = 8'h5b == new_ptr_56_value ? ghv_91 : _GEN_6153; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6155 = 8'h5c == new_ptr_56_value ? ghv_92 : _GEN_6154; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6156 = 8'h5d == new_ptr_56_value ? ghv_93 : _GEN_6155; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6157 = 8'h5e == new_ptr_56_value ? ghv_94 : _GEN_6156; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6158 = 8'h5f == new_ptr_56_value ? ghv_95 : _GEN_6157; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6159 = 8'h60 == new_ptr_56_value ? ghv_96 : _GEN_6158; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6160 = 8'h61 == new_ptr_56_value ? ghv_97 : _GEN_6159; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6161 = 8'h62 == new_ptr_56_value ? ghv_98 : _GEN_6160; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6162 = 8'h63 == new_ptr_56_value ? ghv_99 : _GEN_6161; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6163 = 8'h64 == new_ptr_56_value ? ghv_100 : _GEN_6162; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6164 = 8'h65 == new_ptr_56_value ? ghv_101 : _GEN_6163; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6165 = 8'h66 == new_ptr_56_value ? ghv_102 : _GEN_6164; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6166 = 8'h67 == new_ptr_56_value ? ghv_103 : _GEN_6165; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6167 = 8'h68 == new_ptr_56_value ? ghv_104 : _GEN_6166; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6168 = 8'h69 == new_ptr_56_value ? ghv_105 : _GEN_6167; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6169 = 8'h6a == new_ptr_56_value ? ghv_106 : _GEN_6168; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6170 = 8'h6b == new_ptr_56_value ? ghv_107 : _GEN_6169; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6171 = 8'h6c == new_ptr_56_value ? ghv_108 : _GEN_6170; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6172 = 8'h6d == new_ptr_56_value ? ghv_109 : _GEN_6171; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6173 = 8'h6e == new_ptr_56_value ? ghv_110 : _GEN_6172; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6174 = 8'h6f == new_ptr_56_value ? ghv_111 : _GEN_6173; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6175 = 8'h70 == new_ptr_56_value ? ghv_112 : _GEN_6174; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6176 = 8'h71 == new_ptr_56_value ? ghv_113 : _GEN_6175; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6177 = 8'h72 == new_ptr_56_value ? ghv_114 : _GEN_6176; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6178 = 8'h73 == new_ptr_56_value ? ghv_115 : _GEN_6177; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6179 = 8'h74 == new_ptr_56_value ? ghv_116 : _GEN_6178; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6180 = 8'h75 == new_ptr_56_value ? ghv_117 : _GEN_6179; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6181 = 8'h76 == new_ptr_56_value ? ghv_118 : _GEN_6180; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6182 = 8'h77 == new_ptr_56_value ? ghv_119 : _GEN_6181; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6183 = 8'h78 == new_ptr_56_value ? ghv_120 : _GEN_6182; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6184 = 8'h79 == new_ptr_56_value ? ghv_121 : _GEN_6183; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6185 = 8'h7a == new_ptr_56_value ? ghv_122 : _GEN_6184; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6186 = 8'h7b == new_ptr_56_value ? ghv_123 : _GEN_6185; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6187 = 8'h7c == new_ptr_56_value ? ghv_124 : _GEN_6186; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6188 = 8'h7d == new_ptr_56_value ? ghv_125 : _GEN_6187; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6189 = 8'h7e == new_ptr_56_value ? ghv_126 : _GEN_6188; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6190 = 8'h7f == new_ptr_56_value ? ghv_127 : _GEN_6189; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6191 = 8'h80 == new_ptr_56_value ? ghv_128 : _GEN_6190; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6192 = 8'h81 == new_ptr_56_value ? ghv_129 : _GEN_6191; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6193 = 8'h82 == new_ptr_56_value ? ghv_130 : _GEN_6192; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6194 = 8'h83 == new_ptr_56_value ? ghv_131 : _GEN_6193; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6195 = 8'h84 == new_ptr_56_value ? ghv_132 : _GEN_6194; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6196 = 8'h85 == new_ptr_56_value ? ghv_133 : _GEN_6195; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6197 = 8'h86 == new_ptr_56_value ? ghv_134 : _GEN_6196; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6198 = 8'h87 == new_ptr_56_value ? ghv_135 : _GEN_6197; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6199 = 8'h88 == new_ptr_56_value ? ghv_136 : _GEN_6198; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6200 = 8'h89 == new_ptr_56_value ? ghv_137 : _GEN_6199; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6201 = 8'h8a == new_ptr_56_value ? ghv_138 : _GEN_6200; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6202 = 8'h8b == new_ptr_56_value ? ghv_139 : _GEN_6201; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6203 = 8'h8c == new_ptr_56_value ? ghv_140 : _GEN_6202; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6204 = 8'h8d == new_ptr_56_value ? ghv_141 : _GEN_6203; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6205 = 8'h8e == new_ptr_56_value ? ghv_142 : _GEN_6204; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_53_value = _new_ptr_value_T_107[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_6208 = 8'h1 == new_ptr_53_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6209 = 8'h2 == new_ptr_53_value ? ghv_2 : _GEN_6208; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6210 = 8'h3 == new_ptr_53_value ? ghv_3 : _GEN_6209; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6211 = 8'h4 == new_ptr_53_value ? ghv_4 : _GEN_6210; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6212 = 8'h5 == new_ptr_53_value ? ghv_5 : _GEN_6211; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6213 = 8'h6 == new_ptr_53_value ? ghv_6 : _GEN_6212; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6214 = 8'h7 == new_ptr_53_value ? ghv_7 : _GEN_6213; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6215 = 8'h8 == new_ptr_53_value ? ghv_8 : _GEN_6214; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6216 = 8'h9 == new_ptr_53_value ? ghv_9 : _GEN_6215; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6217 = 8'ha == new_ptr_53_value ? ghv_10 : _GEN_6216; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6218 = 8'hb == new_ptr_53_value ? ghv_11 : _GEN_6217; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6219 = 8'hc == new_ptr_53_value ? ghv_12 : _GEN_6218; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6220 = 8'hd == new_ptr_53_value ? ghv_13 : _GEN_6219; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6221 = 8'he == new_ptr_53_value ? ghv_14 : _GEN_6220; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6222 = 8'hf == new_ptr_53_value ? ghv_15 : _GEN_6221; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6223 = 8'h10 == new_ptr_53_value ? ghv_16 : _GEN_6222; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6224 = 8'h11 == new_ptr_53_value ? ghv_17 : _GEN_6223; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6225 = 8'h12 == new_ptr_53_value ? ghv_18 : _GEN_6224; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6226 = 8'h13 == new_ptr_53_value ? ghv_19 : _GEN_6225; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6227 = 8'h14 == new_ptr_53_value ? ghv_20 : _GEN_6226; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6228 = 8'h15 == new_ptr_53_value ? ghv_21 : _GEN_6227; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6229 = 8'h16 == new_ptr_53_value ? ghv_22 : _GEN_6228; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6230 = 8'h17 == new_ptr_53_value ? ghv_23 : _GEN_6229; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6231 = 8'h18 == new_ptr_53_value ? ghv_24 : _GEN_6230; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6232 = 8'h19 == new_ptr_53_value ? ghv_25 : _GEN_6231; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6233 = 8'h1a == new_ptr_53_value ? ghv_26 : _GEN_6232; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6234 = 8'h1b == new_ptr_53_value ? ghv_27 : _GEN_6233; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6235 = 8'h1c == new_ptr_53_value ? ghv_28 : _GEN_6234; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6236 = 8'h1d == new_ptr_53_value ? ghv_29 : _GEN_6235; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6237 = 8'h1e == new_ptr_53_value ? ghv_30 : _GEN_6236; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6238 = 8'h1f == new_ptr_53_value ? ghv_31 : _GEN_6237; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6239 = 8'h20 == new_ptr_53_value ? ghv_32 : _GEN_6238; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6240 = 8'h21 == new_ptr_53_value ? ghv_33 : _GEN_6239; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6241 = 8'h22 == new_ptr_53_value ? ghv_34 : _GEN_6240; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6242 = 8'h23 == new_ptr_53_value ? ghv_35 : _GEN_6241; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6243 = 8'h24 == new_ptr_53_value ? ghv_36 : _GEN_6242; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6244 = 8'h25 == new_ptr_53_value ? ghv_37 : _GEN_6243; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6245 = 8'h26 == new_ptr_53_value ? ghv_38 : _GEN_6244; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6246 = 8'h27 == new_ptr_53_value ? ghv_39 : _GEN_6245; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6247 = 8'h28 == new_ptr_53_value ? ghv_40 : _GEN_6246; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6248 = 8'h29 == new_ptr_53_value ? ghv_41 : _GEN_6247; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6249 = 8'h2a == new_ptr_53_value ? ghv_42 : _GEN_6248; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6250 = 8'h2b == new_ptr_53_value ? ghv_43 : _GEN_6249; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6251 = 8'h2c == new_ptr_53_value ? ghv_44 : _GEN_6250; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6252 = 8'h2d == new_ptr_53_value ? ghv_45 : _GEN_6251; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6253 = 8'h2e == new_ptr_53_value ? ghv_46 : _GEN_6252; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6254 = 8'h2f == new_ptr_53_value ? ghv_47 : _GEN_6253; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6255 = 8'h30 == new_ptr_53_value ? ghv_48 : _GEN_6254; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6256 = 8'h31 == new_ptr_53_value ? ghv_49 : _GEN_6255; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6257 = 8'h32 == new_ptr_53_value ? ghv_50 : _GEN_6256; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6258 = 8'h33 == new_ptr_53_value ? ghv_51 : _GEN_6257; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6259 = 8'h34 == new_ptr_53_value ? ghv_52 : _GEN_6258; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6260 = 8'h35 == new_ptr_53_value ? ghv_53 : _GEN_6259; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6261 = 8'h36 == new_ptr_53_value ? ghv_54 : _GEN_6260; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6262 = 8'h37 == new_ptr_53_value ? ghv_55 : _GEN_6261; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6263 = 8'h38 == new_ptr_53_value ? ghv_56 : _GEN_6262; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6264 = 8'h39 == new_ptr_53_value ? ghv_57 : _GEN_6263; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6265 = 8'h3a == new_ptr_53_value ? ghv_58 : _GEN_6264; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6266 = 8'h3b == new_ptr_53_value ? ghv_59 : _GEN_6265; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6267 = 8'h3c == new_ptr_53_value ? ghv_60 : _GEN_6266; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6268 = 8'h3d == new_ptr_53_value ? ghv_61 : _GEN_6267; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6269 = 8'h3e == new_ptr_53_value ? ghv_62 : _GEN_6268; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6270 = 8'h3f == new_ptr_53_value ? ghv_63 : _GEN_6269; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6271 = 8'h40 == new_ptr_53_value ? ghv_64 : _GEN_6270; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6272 = 8'h41 == new_ptr_53_value ? ghv_65 : _GEN_6271; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6273 = 8'h42 == new_ptr_53_value ? ghv_66 : _GEN_6272; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6274 = 8'h43 == new_ptr_53_value ? ghv_67 : _GEN_6273; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6275 = 8'h44 == new_ptr_53_value ? ghv_68 : _GEN_6274; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6276 = 8'h45 == new_ptr_53_value ? ghv_69 : _GEN_6275; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6277 = 8'h46 == new_ptr_53_value ? ghv_70 : _GEN_6276; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6278 = 8'h47 == new_ptr_53_value ? ghv_71 : _GEN_6277; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6279 = 8'h48 == new_ptr_53_value ? ghv_72 : _GEN_6278; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6280 = 8'h49 == new_ptr_53_value ? ghv_73 : _GEN_6279; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6281 = 8'h4a == new_ptr_53_value ? ghv_74 : _GEN_6280; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6282 = 8'h4b == new_ptr_53_value ? ghv_75 : _GEN_6281; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6283 = 8'h4c == new_ptr_53_value ? ghv_76 : _GEN_6282; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6284 = 8'h4d == new_ptr_53_value ? ghv_77 : _GEN_6283; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6285 = 8'h4e == new_ptr_53_value ? ghv_78 : _GEN_6284; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6286 = 8'h4f == new_ptr_53_value ? ghv_79 : _GEN_6285; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6287 = 8'h50 == new_ptr_53_value ? ghv_80 : _GEN_6286; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6288 = 8'h51 == new_ptr_53_value ? ghv_81 : _GEN_6287; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6289 = 8'h52 == new_ptr_53_value ? ghv_82 : _GEN_6288; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6290 = 8'h53 == new_ptr_53_value ? ghv_83 : _GEN_6289; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6291 = 8'h54 == new_ptr_53_value ? ghv_84 : _GEN_6290; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6292 = 8'h55 == new_ptr_53_value ? ghv_85 : _GEN_6291; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6293 = 8'h56 == new_ptr_53_value ? ghv_86 : _GEN_6292; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6294 = 8'h57 == new_ptr_53_value ? ghv_87 : _GEN_6293; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6295 = 8'h58 == new_ptr_53_value ? ghv_88 : _GEN_6294; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6296 = 8'h59 == new_ptr_53_value ? ghv_89 : _GEN_6295; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6297 = 8'h5a == new_ptr_53_value ? ghv_90 : _GEN_6296; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6298 = 8'h5b == new_ptr_53_value ? ghv_91 : _GEN_6297; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6299 = 8'h5c == new_ptr_53_value ? ghv_92 : _GEN_6298; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6300 = 8'h5d == new_ptr_53_value ? ghv_93 : _GEN_6299; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6301 = 8'h5e == new_ptr_53_value ? ghv_94 : _GEN_6300; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6302 = 8'h5f == new_ptr_53_value ? ghv_95 : _GEN_6301; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6303 = 8'h60 == new_ptr_53_value ? ghv_96 : _GEN_6302; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6304 = 8'h61 == new_ptr_53_value ? ghv_97 : _GEN_6303; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6305 = 8'h62 == new_ptr_53_value ? ghv_98 : _GEN_6304; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6306 = 8'h63 == new_ptr_53_value ? ghv_99 : _GEN_6305; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6307 = 8'h64 == new_ptr_53_value ? ghv_100 : _GEN_6306; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6308 = 8'h65 == new_ptr_53_value ? ghv_101 : _GEN_6307; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6309 = 8'h66 == new_ptr_53_value ? ghv_102 : _GEN_6308; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6310 = 8'h67 == new_ptr_53_value ? ghv_103 : _GEN_6309; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6311 = 8'h68 == new_ptr_53_value ? ghv_104 : _GEN_6310; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6312 = 8'h69 == new_ptr_53_value ? ghv_105 : _GEN_6311; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6313 = 8'h6a == new_ptr_53_value ? ghv_106 : _GEN_6312; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6314 = 8'h6b == new_ptr_53_value ? ghv_107 : _GEN_6313; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6315 = 8'h6c == new_ptr_53_value ? ghv_108 : _GEN_6314; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6316 = 8'h6d == new_ptr_53_value ? ghv_109 : _GEN_6315; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6317 = 8'h6e == new_ptr_53_value ? ghv_110 : _GEN_6316; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6318 = 8'h6f == new_ptr_53_value ? ghv_111 : _GEN_6317; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6319 = 8'h70 == new_ptr_53_value ? ghv_112 : _GEN_6318; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6320 = 8'h71 == new_ptr_53_value ? ghv_113 : _GEN_6319; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6321 = 8'h72 == new_ptr_53_value ? ghv_114 : _GEN_6320; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6322 = 8'h73 == new_ptr_53_value ? ghv_115 : _GEN_6321; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6323 = 8'h74 == new_ptr_53_value ? ghv_116 : _GEN_6322; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6324 = 8'h75 == new_ptr_53_value ? ghv_117 : _GEN_6323; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6325 = 8'h76 == new_ptr_53_value ? ghv_118 : _GEN_6324; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6326 = 8'h77 == new_ptr_53_value ? ghv_119 : _GEN_6325; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6327 = 8'h78 == new_ptr_53_value ? ghv_120 : _GEN_6326; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6328 = 8'h79 == new_ptr_53_value ? ghv_121 : _GEN_6327; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6329 = 8'h7a == new_ptr_53_value ? ghv_122 : _GEN_6328; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6330 = 8'h7b == new_ptr_53_value ? ghv_123 : _GEN_6329; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6331 = 8'h7c == new_ptr_53_value ? ghv_124 : _GEN_6330; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6332 = 8'h7d == new_ptr_53_value ? ghv_125 : _GEN_6331; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6333 = 8'h7e == new_ptr_53_value ? ghv_126 : _GEN_6332; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6334 = 8'h7f == new_ptr_53_value ? ghv_127 : _GEN_6333; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6335 = 8'h80 == new_ptr_53_value ? ghv_128 : _GEN_6334; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6336 = 8'h81 == new_ptr_53_value ? ghv_129 : _GEN_6335; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6337 = 8'h82 == new_ptr_53_value ? ghv_130 : _GEN_6336; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6338 = 8'h83 == new_ptr_53_value ? ghv_131 : _GEN_6337; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6339 = 8'h84 == new_ptr_53_value ? ghv_132 : _GEN_6338; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6340 = 8'h85 == new_ptr_53_value ? ghv_133 : _GEN_6339; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6341 = 8'h86 == new_ptr_53_value ? ghv_134 : _GEN_6340; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6342 = 8'h87 == new_ptr_53_value ? ghv_135 : _GEN_6341; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6343 = 8'h88 == new_ptr_53_value ? ghv_136 : _GEN_6342; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6344 = 8'h89 == new_ptr_53_value ? ghv_137 : _GEN_6343; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6345 = 8'h8a == new_ptr_53_value ? ghv_138 : _GEN_6344; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6346 = 8'h8b == new_ptr_53_value ? ghv_139 : _GEN_6345; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6347 = 8'h8c == new_ptr_53_value ? ghv_140 : _GEN_6346; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6348 = 8'h8d == new_ptr_53_value ? ghv_141 : _GEN_6347; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6349 = 8'h8e == new_ptr_53_value ? ghv_142 : _GEN_6348; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_46_value = _new_ptr_value_T_93[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_6352 = 8'h1 == new_ptr_46_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6353 = 8'h2 == new_ptr_46_value ? ghv_2 : _GEN_6352; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6354 = 8'h3 == new_ptr_46_value ? ghv_3 : _GEN_6353; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6355 = 8'h4 == new_ptr_46_value ? ghv_4 : _GEN_6354; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6356 = 8'h5 == new_ptr_46_value ? ghv_5 : _GEN_6355; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6357 = 8'h6 == new_ptr_46_value ? ghv_6 : _GEN_6356; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6358 = 8'h7 == new_ptr_46_value ? ghv_7 : _GEN_6357; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6359 = 8'h8 == new_ptr_46_value ? ghv_8 : _GEN_6358; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6360 = 8'h9 == new_ptr_46_value ? ghv_9 : _GEN_6359; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6361 = 8'ha == new_ptr_46_value ? ghv_10 : _GEN_6360; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6362 = 8'hb == new_ptr_46_value ? ghv_11 : _GEN_6361; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6363 = 8'hc == new_ptr_46_value ? ghv_12 : _GEN_6362; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6364 = 8'hd == new_ptr_46_value ? ghv_13 : _GEN_6363; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6365 = 8'he == new_ptr_46_value ? ghv_14 : _GEN_6364; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6366 = 8'hf == new_ptr_46_value ? ghv_15 : _GEN_6365; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6367 = 8'h10 == new_ptr_46_value ? ghv_16 : _GEN_6366; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6368 = 8'h11 == new_ptr_46_value ? ghv_17 : _GEN_6367; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6369 = 8'h12 == new_ptr_46_value ? ghv_18 : _GEN_6368; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6370 = 8'h13 == new_ptr_46_value ? ghv_19 : _GEN_6369; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6371 = 8'h14 == new_ptr_46_value ? ghv_20 : _GEN_6370; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6372 = 8'h15 == new_ptr_46_value ? ghv_21 : _GEN_6371; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6373 = 8'h16 == new_ptr_46_value ? ghv_22 : _GEN_6372; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6374 = 8'h17 == new_ptr_46_value ? ghv_23 : _GEN_6373; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6375 = 8'h18 == new_ptr_46_value ? ghv_24 : _GEN_6374; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6376 = 8'h19 == new_ptr_46_value ? ghv_25 : _GEN_6375; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6377 = 8'h1a == new_ptr_46_value ? ghv_26 : _GEN_6376; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6378 = 8'h1b == new_ptr_46_value ? ghv_27 : _GEN_6377; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6379 = 8'h1c == new_ptr_46_value ? ghv_28 : _GEN_6378; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6380 = 8'h1d == new_ptr_46_value ? ghv_29 : _GEN_6379; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6381 = 8'h1e == new_ptr_46_value ? ghv_30 : _GEN_6380; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6382 = 8'h1f == new_ptr_46_value ? ghv_31 : _GEN_6381; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6383 = 8'h20 == new_ptr_46_value ? ghv_32 : _GEN_6382; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6384 = 8'h21 == new_ptr_46_value ? ghv_33 : _GEN_6383; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6385 = 8'h22 == new_ptr_46_value ? ghv_34 : _GEN_6384; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6386 = 8'h23 == new_ptr_46_value ? ghv_35 : _GEN_6385; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6387 = 8'h24 == new_ptr_46_value ? ghv_36 : _GEN_6386; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6388 = 8'h25 == new_ptr_46_value ? ghv_37 : _GEN_6387; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6389 = 8'h26 == new_ptr_46_value ? ghv_38 : _GEN_6388; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6390 = 8'h27 == new_ptr_46_value ? ghv_39 : _GEN_6389; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6391 = 8'h28 == new_ptr_46_value ? ghv_40 : _GEN_6390; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6392 = 8'h29 == new_ptr_46_value ? ghv_41 : _GEN_6391; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6393 = 8'h2a == new_ptr_46_value ? ghv_42 : _GEN_6392; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6394 = 8'h2b == new_ptr_46_value ? ghv_43 : _GEN_6393; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6395 = 8'h2c == new_ptr_46_value ? ghv_44 : _GEN_6394; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6396 = 8'h2d == new_ptr_46_value ? ghv_45 : _GEN_6395; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6397 = 8'h2e == new_ptr_46_value ? ghv_46 : _GEN_6396; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6398 = 8'h2f == new_ptr_46_value ? ghv_47 : _GEN_6397; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6399 = 8'h30 == new_ptr_46_value ? ghv_48 : _GEN_6398; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6400 = 8'h31 == new_ptr_46_value ? ghv_49 : _GEN_6399; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6401 = 8'h32 == new_ptr_46_value ? ghv_50 : _GEN_6400; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6402 = 8'h33 == new_ptr_46_value ? ghv_51 : _GEN_6401; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6403 = 8'h34 == new_ptr_46_value ? ghv_52 : _GEN_6402; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6404 = 8'h35 == new_ptr_46_value ? ghv_53 : _GEN_6403; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6405 = 8'h36 == new_ptr_46_value ? ghv_54 : _GEN_6404; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6406 = 8'h37 == new_ptr_46_value ? ghv_55 : _GEN_6405; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6407 = 8'h38 == new_ptr_46_value ? ghv_56 : _GEN_6406; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6408 = 8'h39 == new_ptr_46_value ? ghv_57 : _GEN_6407; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6409 = 8'h3a == new_ptr_46_value ? ghv_58 : _GEN_6408; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6410 = 8'h3b == new_ptr_46_value ? ghv_59 : _GEN_6409; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6411 = 8'h3c == new_ptr_46_value ? ghv_60 : _GEN_6410; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6412 = 8'h3d == new_ptr_46_value ? ghv_61 : _GEN_6411; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6413 = 8'h3e == new_ptr_46_value ? ghv_62 : _GEN_6412; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6414 = 8'h3f == new_ptr_46_value ? ghv_63 : _GEN_6413; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6415 = 8'h40 == new_ptr_46_value ? ghv_64 : _GEN_6414; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6416 = 8'h41 == new_ptr_46_value ? ghv_65 : _GEN_6415; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6417 = 8'h42 == new_ptr_46_value ? ghv_66 : _GEN_6416; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6418 = 8'h43 == new_ptr_46_value ? ghv_67 : _GEN_6417; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6419 = 8'h44 == new_ptr_46_value ? ghv_68 : _GEN_6418; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6420 = 8'h45 == new_ptr_46_value ? ghv_69 : _GEN_6419; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6421 = 8'h46 == new_ptr_46_value ? ghv_70 : _GEN_6420; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6422 = 8'h47 == new_ptr_46_value ? ghv_71 : _GEN_6421; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6423 = 8'h48 == new_ptr_46_value ? ghv_72 : _GEN_6422; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6424 = 8'h49 == new_ptr_46_value ? ghv_73 : _GEN_6423; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6425 = 8'h4a == new_ptr_46_value ? ghv_74 : _GEN_6424; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6426 = 8'h4b == new_ptr_46_value ? ghv_75 : _GEN_6425; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6427 = 8'h4c == new_ptr_46_value ? ghv_76 : _GEN_6426; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6428 = 8'h4d == new_ptr_46_value ? ghv_77 : _GEN_6427; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6429 = 8'h4e == new_ptr_46_value ? ghv_78 : _GEN_6428; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6430 = 8'h4f == new_ptr_46_value ? ghv_79 : _GEN_6429; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6431 = 8'h50 == new_ptr_46_value ? ghv_80 : _GEN_6430; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6432 = 8'h51 == new_ptr_46_value ? ghv_81 : _GEN_6431; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6433 = 8'h52 == new_ptr_46_value ? ghv_82 : _GEN_6432; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6434 = 8'h53 == new_ptr_46_value ? ghv_83 : _GEN_6433; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6435 = 8'h54 == new_ptr_46_value ? ghv_84 : _GEN_6434; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6436 = 8'h55 == new_ptr_46_value ? ghv_85 : _GEN_6435; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6437 = 8'h56 == new_ptr_46_value ? ghv_86 : _GEN_6436; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6438 = 8'h57 == new_ptr_46_value ? ghv_87 : _GEN_6437; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6439 = 8'h58 == new_ptr_46_value ? ghv_88 : _GEN_6438; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6440 = 8'h59 == new_ptr_46_value ? ghv_89 : _GEN_6439; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6441 = 8'h5a == new_ptr_46_value ? ghv_90 : _GEN_6440; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6442 = 8'h5b == new_ptr_46_value ? ghv_91 : _GEN_6441; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6443 = 8'h5c == new_ptr_46_value ? ghv_92 : _GEN_6442; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6444 = 8'h5d == new_ptr_46_value ? ghv_93 : _GEN_6443; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6445 = 8'h5e == new_ptr_46_value ? ghv_94 : _GEN_6444; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6446 = 8'h5f == new_ptr_46_value ? ghv_95 : _GEN_6445; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6447 = 8'h60 == new_ptr_46_value ? ghv_96 : _GEN_6446; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6448 = 8'h61 == new_ptr_46_value ? ghv_97 : _GEN_6447; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6449 = 8'h62 == new_ptr_46_value ? ghv_98 : _GEN_6448; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6450 = 8'h63 == new_ptr_46_value ? ghv_99 : _GEN_6449; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6451 = 8'h64 == new_ptr_46_value ? ghv_100 : _GEN_6450; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6452 = 8'h65 == new_ptr_46_value ? ghv_101 : _GEN_6451; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6453 = 8'h66 == new_ptr_46_value ? ghv_102 : _GEN_6452; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6454 = 8'h67 == new_ptr_46_value ? ghv_103 : _GEN_6453; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6455 = 8'h68 == new_ptr_46_value ? ghv_104 : _GEN_6454; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6456 = 8'h69 == new_ptr_46_value ? ghv_105 : _GEN_6455; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6457 = 8'h6a == new_ptr_46_value ? ghv_106 : _GEN_6456; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6458 = 8'h6b == new_ptr_46_value ? ghv_107 : _GEN_6457; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6459 = 8'h6c == new_ptr_46_value ? ghv_108 : _GEN_6458; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6460 = 8'h6d == new_ptr_46_value ? ghv_109 : _GEN_6459; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6461 = 8'h6e == new_ptr_46_value ? ghv_110 : _GEN_6460; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6462 = 8'h6f == new_ptr_46_value ? ghv_111 : _GEN_6461; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6463 = 8'h70 == new_ptr_46_value ? ghv_112 : _GEN_6462; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6464 = 8'h71 == new_ptr_46_value ? ghv_113 : _GEN_6463; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6465 = 8'h72 == new_ptr_46_value ? ghv_114 : _GEN_6464; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6466 = 8'h73 == new_ptr_46_value ? ghv_115 : _GEN_6465; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6467 = 8'h74 == new_ptr_46_value ? ghv_116 : _GEN_6466; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6468 = 8'h75 == new_ptr_46_value ? ghv_117 : _GEN_6467; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6469 = 8'h76 == new_ptr_46_value ? ghv_118 : _GEN_6468; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6470 = 8'h77 == new_ptr_46_value ? ghv_119 : _GEN_6469; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6471 = 8'h78 == new_ptr_46_value ? ghv_120 : _GEN_6470; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6472 = 8'h79 == new_ptr_46_value ? ghv_121 : _GEN_6471; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6473 = 8'h7a == new_ptr_46_value ? ghv_122 : _GEN_6472; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6474 = 8'h7b == new_ptr_46_value ? ghv_123 : _GEN_6473; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6475 = 8'h7c == new_ptr_46_value ? ghv_124 : _GEN_6474; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6476 = 8'h7d == new_ptr_46_value ? ghv_125 : _GEN_6475; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6477 = 8'h7e == new_ptr_46_value ? ghv_126 : _GEN_6476; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6478 = 8'h7f == new_ptr_46_value ? ghv_127 : _GEN_6477; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6479 = 8'h80 == new_ptr_46_value ? ghv_128 : _GEN_6478; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6480 = 8'h81 == new_ptr_46_value ? ghv_129 : _GEN_6479; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6481 = 8'h82 == new_ptr_46_value ? ghv_130 : _GEN_6480; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6482 = 8'h83 == new_ptr_46_value ? ghv_131 : _GEN_6481; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6483 = 8'h84 == new_ptr_46_value ? ghv_132 : _GEN_6482; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6484 = 8'h85 == new_ptr_46_value ? ghv_133 : _GEN_6483; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6485 = 8'h86 == new_ptr_46_value ? ghv_134 : _GEN_6484; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6486 = 8'h87 == new_ptr_46_value ? ghv_135 : _GEN_6485; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6487 = 8'h88 == new_ptr_46_value ? ghv_136 : _GEN_6486; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6488 = 8'h89 == new_ptr_46_value ? ghv_137 : _GEN_6487; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6489 = 8'h8a == new_ptr_46_value ? ghv_138 : _GEN_6488; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6490 = 8'h8b == new_ptr_46_value ? ghv_139 : _GEN_6489; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6491 = 8'h8c == new_ptr_46_value ? ghv_140 : _GEN_6490; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6492 = 8'h8d == new_ptr_46_value ? ghv_141 : _GEN_6491; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6493 = 8'h8e == new_ptr_46_value ? ghv_142 : _GEN_6492; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_52_value = _new_ptr_value_T_105[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_6496 = 8'h1 == new_ptr_52_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6497 = 8'h2 == new_ptr_52_value ? ghv_2 : _GEN_6496; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6498 = 8'h3 == new_ptr_52_value ? ghv_3 : _GEN_6497; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6499 = 8'h4 == new_ptr_52_value ? ghv_4 : _GEN_6498; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6500 = 8'h5 == new_ptr_52_value ? ghv_5 : _GEN_6499; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6501 = 8'h6 == new_ptr_52_value ? ghv_6 : _GEN_6500; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6502 = 8'h7 == new_ptr_52_value ? ghv_7 : _GEN_6501; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6503 = 8'h8 == new_ptr_52_value ? ghv_8 : _GEN_6502; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6504 = 8'h9 == new_ptr_52_value ? ghv_9 : _GEN_6503; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6505 = 8'ha == new_ptr_52_value ? ghv_10 : _GEN_6504; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6506 = 8'hb == new_ptr_52_value ? ghv_11 : _GEN_6505; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6507 = 8'hc == new_ptr_52_value ? ghv_12 : _GEN_6506; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6508 = 8'hd == new_ptr_52_value ? ghv_13 : _GEN_6507; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6509 = 8'he == new_ptr_52_value ? ghv_14 : _GEN_6508; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6510 = 8'hf == new_ptr_52_value ? ghv_15 : _GEN_6509; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6511 = 8'h10 == new_ptr_52_value ? ghv_16 : _GEN_6510; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6512 = 8'h11 == new_ptr_52_value ? ghv_17 : _GEN_6511; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6513 = 8'h12 == new_ptr_52_value ? ghv_18 : _GEN_6512; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6514 = 8'h13 == new_ptr_52_value ? ghv_19 : _GEN_6513; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6515 = 8'h14 == new_ptr_52_value ? ghv_20 : _GEN_6514; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6516 = 8'h15 == new_ptr_52_value ? ghv_21 : _GEN_6515; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6517 = 8'h16 == new_ptr_52_value ? ghv_22 : _GEN_6516; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6518 = 8'h17 == new_ptr_52_value ? ghv_23 : _GEN_6517; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6519 = 8'h18 == new_ptr_52_value ? ghv_24 : _GEN_6518; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6520 = 8'h19 == new_ptr_52_value ? ghv_25 : _GEN_6519; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6521 = 8'h1a == new_ptr_52_value ? ghv_26 : _GEN_6520; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6522 = 8'h1b == new_ptr_52_value ? ghv_27 : _GEN_6521; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6523 = 8'h1c == new_ptr_52_value ? ghv_28 : _GEN_6522; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6524 = 8'h1d == new_ptr_52_value ? ghv_29 : _GEN_6523; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6525 = 8'h1e == new_ptr_52_value ? ghv_30 : _GEN_6524; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6526 = 8'h1f == new_ptr_52_value ? ghv_31 : _GEN_6525; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6527 = 8'h20 == new_ptr_52_value ? ghv_32 : _GEN_6526; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6528 = 8'h21 == new_ptr_52_value ? ghv_33 : _GEN_6527; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6529 = 8'h22 == new_ptr_52_value ? ghv_34 : _GEN_6528; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6530 = 8'h23 == new_ptr_52_value ? ghv_35 : _GEN_6529; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6531 = 8'h24 == new_ptr_52_value ? ghv_36 : _GEN_6530; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6532 = 8'h25 == new_ptr_52_value ? ghv_37 : _GEN_6531; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6533 = 8'h26 == new_ptr_52_value ? ghv_38 : _GEN_6532; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6534 = 8'h27 == new_ptr_52_value ? ghv_39 : _GEN_6533; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6535 = 8'h28 == new_ptr_52_value ? ghv_40 : _GEN_6534; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6536 = 8'h29 == new_ptr_52_value ? ghv_41 : _GEN_6535; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6537 = 8'h2a == new_ptr_52_value ? ghv_42 : _GEN_6536; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6538 = 8'h2b == new_ptr_52_value ? ghv_43 : _GEN_6537; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6539 = 8'h2c == new_ptr_52_value ? ghv_44 : _GEN_6538; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6540 = 8'h2d == new_ptr_52_value ? ghv_45 : _GEN_6539; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6541 = 8'h2e == new_ptr_52_value ? ghv_46 : _GEN_6540; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6542 = 8'h2f == new_ptr_52_value ? ghv_47 : _GEN_6541; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6543 = 8'h30 == new_ptr_52_value ? ghv_48 : _GEN_6542; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6544 = 8'h31 == new_ptr_52_value ? ghv_49 : _GEN_6543; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6545 = 8'h32 == new_ptr_52_value ? ghv_50 : _GEN_6544; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6546 = 8'h33 == new_ptr_52_value ? ghv_51 : _GEN_6545; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6547 = 8'h34 == new_ptr_52_value ? ghv_52 : _GEN_6546; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6548 = 8'h35 == new_ptr_52_value ? ghv_53 : _GEN_6547; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6549 = 8'h36 == new_ptr_52_value ? ghv_54 : _GEN_6548; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6550 = 8'h37 == new_ptr_52_value ? ghv_55 : _GEN_6549; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6551 = 8'h38 == new_ptr_52_value ? ghv_56 : _GEN_6550; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6552 = 8'h39 == new_ptr_52_value ? ghv_57 : _GEN_6551; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6553 = 8'h3a == new_ptr_52_value ? ghv_58 : _GEN_6552; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6554 = 8'h3b == new_ptr_52_value ? ghv_59 : _GEN_6553; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6555 = 8'h3c == new_ptr_52_value ? ghv_60 : _GEN_6554; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6556 = 8'h3d == new_ptr_52_value ? ghv_61 : _GEN_6555; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6557 = 8'h3e == new_ptr_52_value ? ghv_62 : _GEN_6556; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6558 = 8'h3f == new_ptr_52_value ? ghv_63 : _GEN_6557; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6559 = 8'h40 == new_ptr_52_value ? ghv_64 : _GEN_6558; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6560 = 8'h41 == new_ptr_52_value ? ghv_65 : _GEN_6559; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6561 = 8'h42 == new_ptr_52_value ? ghv_66 : _GEN_6560; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6562 = 8'h43 == new_ptr_52_value ? ghv_67 : _GEN_6561; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6563 = 8'h44 == new_ptr_52_value ? ghv_68 : _GEN_6562; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6564 = 8'h45 == new_ptr_52_value ? ghv_69 : _GEN_6563; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6565 = 8'h46 == new_ptr_52_value ? ghv_70 : _GEN_6564; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6566 = 8'h47 == new_ptr_52_value ? ghv_71 : _GEN_6565; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6567 = 8'h48 == new_ptr_52_value ? ghv_72 : _GEN_6566; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6568 = 8'h49 == new_ptr_52_value ? ghv_73 : _GEN_6567; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6569 = 8'h4a == new_ptr_52_value ? ghv_74 : _GEN_6568; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6570 = 8'h4b == new_ptr_52_value ? ghv_75 : _GEN_6569; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6571 = 8'h4c == new_ptr_52_value ? ghv_76 : _GEN_6570; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6572 = 8'h4d == new_ptr_52_value ? ghv_77 : _GEN_6571; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6573 = 8'h4e == new_ptr_52_value ? ghv_78 : _GEN_6572; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6574 = 8'h4f == new_ptr_52_value ? ghv_79 : _GEN_6573; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6575 = 8'h50 == new_ptr_52_value ? ghv_80 : _GEN_6574; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6576 = 8'h51 == new_ptr_52_value ? ghv_81 : _GEN_6575; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6577 = 8'h52 == new_ptr_52_value ? ghv_82 : _GEN_6576; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6578 = 8'h53 == new_ptr_52_value ? ghv_83 : _GEN_6577; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6579 = 8'h54 == new_ptr_52_value ? ghv_84 : _GEN_6578; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6580 = 8'h55 == new_ptr_52_value ? ghv_85 : _GEN_6579; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6581 = 8'h56 == new_ptr_52_value ? ghv_86 : _GEN_6580; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6582 = 8'h57 == new_ptr_52_value ? ghv_87 : _GEN_6581; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6583 = 8'h58 == new_ptr_52_value ? ghv_88 : _GEN_6582; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6584 = 8'h59 == new_ptr_52_value ? ghv_89 : _GEN_6583; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6585 = 8'h5a == new_ptr_52_value ? ghv_90 : _GEN_6584; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6586 = 8'h5b == new_ptr_52_value ? ghv_91 : _GEN_6585; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6587 = 8'h5c == new_ptr_52_value ? ghv_92 : _GEN_6586; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6588 = 8'h5d == new_ptr_52_value ? ghv_93 : _GEN_6587; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6589 = 8'h5e == new_ptr_52_value ? ghv_94 : _GEN_6588; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6590 = 8'h5f == new_ptr_52_value ? ghv_95 : _GEN_6589; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6591 = 8'h60 == new_ptr_52_value ? ghv_96 : _GEN_6590; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6592 = 8'h61 == new_ptr_52_value ? ghv_97 : _GEN_6591; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6593 = 8'h62 == new_ptr_52_value ? ghv_98 : _GEN_6592; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6594 = 8'h63 == new_ptr_52_value ? ghv_99 : _GEN_6593; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6595 = 8'h64 == new_ptr_52_value ? ghv_100 : _GEN_6594; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6596 = 8'h65 == new_ptr_52_value ? ghv_101 : _GEN_6595; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6597 = 8'h66 == new_ptr_52_value ? ghv_102 : _GEN_6596; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6598 = 8'h67 == new_ptr_52_value ? ghv_103 : _GEN_6597; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6599 = 8'h68 == new_ptr_52_value ? ghv_104 : _GEN_6598; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6600 = 8'h69 == new_ptr_52_value ? ghv_105 : _GEN_6599; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6601 = 8'h6a == new_ptr_52_value ? ghv_106 : _GEN_6600; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6602 = 8'h6b == new_ptr_52_value ? ghv_107 : _GEN_6601; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6603 = 8'h6c == new_ptr_52_value ? ghv_108 : _GEN_6602; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6604 = 8'h6d == new_ptr_52_value ? ghv_109 : _GEN_6603; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6605 = 8'h6e == new_ptr_52_value ? ghv_110 : _GEN_6604; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6606 = 8'h6f == new_ptr_52_value ? ghv_111 : _GEN_6605; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6607 = 8'h70 == new_ptr_52_value ? ghv_112 : _GEN_6606; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6608 = 8'h71 == new_ptr_52_value ? ghv_113 : _GEN_6607; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6609 = 8'h72 == new_ptr_52_value ? ghv_114 : _GEN_6608; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6610 = 8'h73 == new_ptr_52_value ? ghv_115 : _GEN_6609; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6611 = 8'h74 == new_ptr_52_value ? ghv_116 : _GEN_6610; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6612 = 8'h75 == new_ptr_52_value ? ghv_117 : _GEN_6611; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6613 = 8'h76 == new_ptr_52_value ? ghv_118 : _GEN_6612; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6614 = 8'h77 == new_ptr_52_value ? ghv_119 : _GEN_6613; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6615 = 8'h78 == new_ptr_52_value ? ghv_120 : _GEN_6614; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6616 = 8'h79 == new_ptr_52_value ? ghv_121 : _GEN_6615; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6617 = 8'h7a == new_ptr_52_value ? ghv_122 : _GEN_6616; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6618 = 8'h7b == new_ptr_52_value ? ghv_123 : _GEN_6617; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6619 = 8'h7c == new_ptr_52_value ? ghv_124 : _GEN_6618; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6620 = 8'h7d == new_ptr_52_value ? ghv_125 : _GEN_6619; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6621 = 8'h7e == new_ptr_52_value ? ghv_126 : _GEN_6620; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6622 = 8'h7f == new_ptr_52_value ? ghv_127 : _GEN_6621; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6623 = 8'h80 == new_ptr_52_value ? ghv_128 : _GEN_6622; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6624 = 8'h81 == new_ptr_52_value ? ghv_129 : _GEN_6623; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6625 = 8'h82 == new_ptr_52_value ? ghv_130 : _GEN_6624; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6626 = 8'h83 == new_ptr_52_value ? ghv_131 : _GEN_6625; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6627 = 8'h84 == new_ptr_52_value ? ghv_132 : _GEN_6626; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6628 = 8'h85 == new_ptr_52_value ? ghv_133 : _GEN_6627; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6629 = 8'h86 == new_ptr_52_value ? ghv_134 : _GEN_6628; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6630 = 8'h87 == new_ptr_52_value ? ghv_135 : _GEN_6629; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6631 = 8'h88 == new_ptr_52_value ? ghv_136 : _GEN_6630; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6632 = 8'h89 == new_ptr_52_value ? ghv_137 : _GEN_6631; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6633 = 8'h8a == new_ptr_52_value ? ghv_138 : _GEN_6632; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6634 = 8'h8b == new_ptr_52_value ? ghv_139 : _GEN_6633; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6635 = 8'h8c == new_ptr_52_value ? ghv_140 : _GEN_6634; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6636 = 8'h8d == new_ptr_52_value ? ghv_141 : _GEN_6635; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6637 = 8'h8e == new_ptr_52_value ? ghv_142 : _GEN_6636; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_55_value = _new_ptr_value_T_111[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_6640 = 8'h1 == new_ptr_55_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6641 = 8'h2 == new_ptr_55_value ? ghv_2 : _GEN_6640; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6642 = 8'h3 == new_ptr_55_value ? ghv_3 : _GEN_6641; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6643 = 8'h4 == new_ptr_55_value ? ghv_4 : _GEN_6642; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6644 = 8'h5 == new_ptr_55_value ? ghv_5 : _GEN_6643; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6645 = 8'h6 == new_ptr_55_value ? ghv_6 : _GEN_6644; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6646 = 8'h7 == new_ptr_55_value ? ghv_7 : _GEN_6645; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6647 = 8'h8 == new_ptr_55_value ? ghv_8 : _GEN_6646; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6648 = 8'h9 == new_ptr_55_value ? ghv_9 : _GEN_6647; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6649 = 8'ha == new_ptr_55_value ? ghv_10 : _GEN_6648; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6650 = 8'hb == new_ptr_55_value ? ghv_11 : _GEN_6649; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6651 = 8'hc == new_ptr_55_value ? ghv_12 : _GEN_6650; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6652 = 8'hd == new_ptr_55_value ? ghv_13 : _GEN_6651; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6653 = 8'he == new_ptr_55_value ? ghv_14 : _GEN_6652; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6654 = 8'hf == new_ptr_55_value ? ghv_15 : _GEN_6653; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6655 = 8'h10 == new_ptr_55_value ? ghv_16 : _GEN_6654; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6656 = 8'h11 == new_ptr_55_value ? ghv_17 : _GEN_6655; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6657 = 8'h12 == new_ptr_55_value ? ghv_18 : _GEN_6656; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6658 = 8'h13 == new_ptr_55_value ? ghv_19 : _GEN_6657; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6659 = 8'h14 == new_ptr_55_value ? ghv_20 : _GEN_6658; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6660 = 8'h15 == new_ptr_55_value ? ghv_21 : _GEN_6659; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6661 = 8'h16 == new_ptr_55_value ? ghv_22 : _GEN_6660; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6662 = 8'h17 == new_ptr_55_value ? ghv_23 : _GEN_6661; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6663 = 8'h18 == new_ptr_55_value ? ghv_24 : _GEN_6662; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6664 = 8'h19 == new_ptr_55_value ? ghv_25 : _GEN_6663; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6665 = 8'h1a == new_ptr_55_value ? ghv_26 : _GEN_6664; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6666 = 8'h1b == new_ptr_55_value ? ghv_27 : _GEN_6665; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6667 = 8'h1c == new_ptr_55_value ? ghv_28 : _GEN_6666; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6668 = 8'h1d == new_ptr_55_value ? ghv_29 : _GEN_6667; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6669 = 8'h1e == new_ptr_55_value ? ghv_30 : _GEN_6668; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6670 = 8'h1f == new_ptr_55_value ? ghv_31 : _GEN_6669; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6671 = 8'h20 == new_ptr_55_value ? ghv_32 : _GEN_6670; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6672 = 8'h21 == new_ptr_55_value ? ghv_33 : _GEN_6671; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6673 = 8'h22 == new_ptr_55_value ? ghv_34 : _GEN_6672; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6674 = 8'h23 == new_ptr_55_value ? ghv_35 : _GEN_6673; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6675 = 8'h24 == new_ptr_55_value ? ghv_36 : _GEN_6674; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6676 = 8'h25 == new_ptr_55_value ? ghv_37 : _GEN_6675; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6677 = 8'h26 == new_ptr_55_value ? ghv_38 : _GEN_6676; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6678 = 8'h27 == new_ptr_55_value ? ghv_39 : _GEN_6677; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6679 = 8'h28 == new_ptr_55_value ? ghv_40 : _GEN_6678; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6680 = 8'h29 == new_ptr_55_value ? ghv_41 : _GEN_6679; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6681 = 8'h2a == new_ptr_55_value ? ghv_42 : _GEN_6680; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6682 = 8'h2b == new_ptr_55_value ? ghv_43 : _GEN_6681; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6683 = 8'h2c == new_ptr_55_value ? ghv_44 : _GEN_6682; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6684 = 8'h2d == new_ptr_55_value ? ghv_45 : _GEN_6683; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6685 = 8'h2e == new_ptr_55_value ? ghv_46 : _GEN_6684; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6686 = 8'h2f == new_ptr_55_value ? ghv_47 : _GEN_6685; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6687 = 8'h30 == new_ptr_55_value ? ghv_48 : _GEN_6686; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6688 = 8'h31 == new_ptr_55_value ? ghv_49 : _GEN_6687; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6689 = 8'h32 == new_ptr_55_value ? ghv_50 : _GEN_6688; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6690 = 8'h33 == new_ptr_55_value ? ghv_51 : _GEN_6689; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6691 = 8'h34 == new_ptr_55_value ? ghv_52 : _GEN_6690; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6692 = 8'h35 == new_ptr_55_value ? ghv_53 : _GEN_6691; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6693 = 8'h36 == new_ptr_55_value ? ghv_54 : _GEN_6692; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6694 = 8'h37 == new_ptr_55_value ? ghv_55 : _GEN_6693; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6695 = 8'h38 == new_ptr_55_value ? ghv_56 : _GEN_6694; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6696 = 8'h39 == new_ptr_55_value ? ghv_57 : _GEN_6695; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6697 = 8'h3a == new_ptr_55_value ? ghv_58 : _GEN_6696; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6698 = 8'h3b == new_ptr_55_value ? ghv_59 : _GEN_6697; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6699 = 8'h3c == new_ptr_55_value ? ghv_60 : _GEN_6698; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6700 = 8'h3d == new_ptr_55_value ? ghv_61 : _GEN_6699; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6701 = 8'h3e == new_ptr_55_value ? ghv_62 : _GEN_6700; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6702 = 8'h3f == new_ptr_55_value ? ghv_63 : _GEN_6701; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6703 = 8'h40 == new_ptr_55_value ? ghv_64 : _GEN_6702; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6704 = 8'h41 == new_ptr_55_value ? ghv_65 : _GEN_6703; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6705 = 8'h42 == new_ptr_55_value ? ghv_66 : _GEN_6704; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6706 = 8'h43 == new_ptr_55_value ? ghv_67 : _GEN_6705; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6707 = 8'h44 == new_ptr_55_value ? ghv_68 : _GEN_6706; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6708 = 8'h45 == new_ptr_55_value ? ghv_69 : _GEN_6707; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6709 = 8'h46 == new_ptr_55_value ? ghv_70 : _GEN_6708; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6710 = 8'h47 == new_ptr_55_value ? ghv_71 : _GEN_6709; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6711 = 8'h48 == new_ptr_55_value ? ghv_72 : _GEN_6710; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6712 = 8'h49 == new_ptr_55_value ? ghv_73 : _GEN_6711; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6713 = 8'h4a == new_ptr_55_value ? ghv_74 : _GEN_6712; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6714 = 8'h4b == new_ptr_55_value ? ghv_75 : _GEN_6713; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6715 = 8'h4c == new_ptr_55_value ? ghv_76 : _GEN_6714; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6716 = 8'h4d == new_ptr_55_value ? ghv_77 : _GEN_6715; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6717 = 8'h4e == new_ptr_55_value ? ghv_78 : _GEN_6716; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6718 = 8'h4f == new_ptr_55_value ? ghv_79 : _GEN_6717; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6719 = 8'h50 == new_ptr_55_value ? ghv_80 : _GEN_6718; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6720 = 8'h51 == new_ptr_55_value ? ghv_81 : _GEN_6719; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6721 = 8'h52 == new_ptr_55_value ? ghv_82 : _GEN_6720; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6722 = 8'h53 == new_ptr_55_value ? ghv_83 : _GEN_6721; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6723 = 8'h54 == new_ptr_55_value ? ghv_84 : _GEN_6722; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6724 = 8'h55 == new_ptr_55_value ? ghv_85 : _GEN_6723; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6725 = 8'h56 == new_ptr_55_value ? ghv_86 : _GEN_6724; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6726 = 8'h57 == new_ptr_55_value ? ghv_87 : _GEN_6725; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6727 = 8'h58 == new_ptr_55_value ? ghv_88 : _GEN_6726; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6728 = 8'h59 == new_ptr_55_value ? ghv_89 : _GEN_6727; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6729 = 8'h5a == new_ptr_55_value ? ghv_90 : _GEN_6728; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6730 = 8'h5b == new_ptr_55_value ? ghv_91 : _GEN_6729; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6731 = 8'h5c == new_ptr_55_value ? ghv_92 : _GEN_6730; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6732 = 8'h5d == new_ptr_55_value ? ghv_93 : _GEN_6731; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6733 = 8'h5e == new_ptr_55_value ? ghv_94 : _GEN_6732; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6734 = 8'h5f == new_ptr_55_value ? ghv_95 : _GEN_6733; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6735 = 8'h60 == new_ptr_55_value ? ghv_96 : _GEN_6734; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6736 = 8'h61 == new_ptr_55_value ? ghv_97 : _GEN_6735; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6737 = 8'h62 == new_ptr_55_value ? ghv_98 : _GEN_6736; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6738 = 8'h63 == new_ptr_55_value ? ghv_99 : _GEN_6737; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6739 = 8'h64 == new_ptr_55_value ? ghv_100 : _GEN_6738; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6740 = 8'h65 == new_ptr_55_value ? ghv_101 : _GEN_6739; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6741 = 8'h66 == new_ptr_55_value ? ghv_102 : _GEN_6740; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6742 = 8'h67 == new_ptr_55_value ? ghv_103 : _GEN_6741; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6743 = 8'h68 == new_ptr_55_value ? ghv_104 : _GEN_6742; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6744 = 8'h69 == new_ptr_55_value ? ghv_105 : _GEN_6743; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6745 = 8'h6a == new_ptr_55_value ? ghv_106 : _GEN_6744; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6746 = 8'h6b == new_ptr_55_value ? ghv_107 : _GEN_6745; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6747 = 8'h6c == new_ptr_55_value ? ghv_108 : _GEN_6746; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6748 = 8'h6d == new_ptr_55_value ? ghv_109 : _GEN_6747; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6749 = 8'h6e == new_ptr_55_value ? ghv_110 : _GEN_6748; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6750 = 8'h6f == new_ptr_55_value ? ghv_111 : _GEN_6749; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6751 = 8'h70 == new_ptr_55_value ? ghv_112 : _GEN_6750; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6752 = 8'h71 == new_ptr_55_value ? ghv_113 : _GEN_6751; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6753 = 8'h72 == new_ptr_55_value ? ghv_114 : _GEN_6752; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6754 = 8'h73 == new_ptr_55_value ? ghv_115 : _GEN_6753; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6755 = 8'h74 == new_ptr_55_value ? ghv_116 : _GEN_6754; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6756 = 8'h75 == new_ptr_55_value ? ghv_117 : _GEN_6755; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6757 = 8'h76 == new_ptr_55_value ? ghv_118 : _GEN_6756; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6758 = 8'h77 == new_ptr_55_value ? ghv_119 : _GEN_6757; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6759 = 8'h78 == new_ptr_55_value ? ghv_120 : _GEN_6758; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6760 = 8'h79 == new_ptr_55_value ? ghv_121 : _GEN_6759; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6761 = 8'h7a == new_ptr_55_value ? ghv_122 : _GEN_6760; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6762 = 8'h7b == new_ptr_55_value ? ghv_123 : _GEN_6761; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6763 = 8'h7c == new_ptr_55_value ? ghv_124 : _GEN_6762; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6764 = 8'h7d == new_ptr_55_value ? ghv_125 : _GEN_6763; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6765 = 8'h7e == new_ptr_55_value ? ghv_126 : _GEN_6764; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6766 = 8'h7f == new_ptr_55_value ? ghv_127 : _GEN_6765; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6767 = 8'h80 == new_ptr_55_value ? ghv_128 : _GEN_6766; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6768 = 8'h81 == new_ptr_55_value ? ghv_129 : _GEN_6767; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6769 = 8'h82 == new_ptr_55_value ? ghv_130 : _GEN_6768; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6770 = 8'h83 == new_ptr_55_value ? ghv_131 : _GEN_6769; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6771 = 8'h84 == new_ptr_55_value ? ghv_132 : _GEN_6770; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6772 = 8'h85 == new_ptr_55_value ? ghv_133 : _GEN_6771; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6773 = 8'h86 == new_ptr_55_value ? ghv_134 : _GEN_6772; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6774 = 8'h87 == new_ptr_55_value ? ghv_135 : _GEN_6773; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6775 = 8'h88 == new_ptr_55_value ? ghv_136 : _GEN_6774; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6776 = 8'h89 == new_ptr_55_value ? ghv_137 : _GEN_6775; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6777 = 8'h8a == new_ptr_55_value ? ghv_138 : _GEN_6776; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6778 = 8'h8b == new_ptr_55_value ? ghv_139 : _GEN_6777; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6779 = 8'h8c == new_ptr_55_value ? ghv_140 : _GEN_6778; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6780 = 8'h8d == new_ptr_55_value ? ghv_141 : _GEN_6779; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6781 = 8'h8e == new_ptr_55_value ? ghv_142 : _GEN_6780; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_42_value = _new_ptr_value_T_85[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_6784 = 8'h1 == new_ptr_42_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6785 = 8'h2 == new_ptr_42_value ? ghv_2 : _GEN_6784; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6786 = 8'h3 == new_ptr_42_value ? ghv_3 : _GEN_6785; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6787 = 8'h4 == new_ptr_42_value ? ghv_4 : _GEN_6786; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6788 = 8'h5 == new_ptr_42_value ? ghv_5 : _GEN_6787; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6789 = 8'h6 == new_ptr_42_value ? ghv_6 : _GEN_6788; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6790 = 8'h7 == new_ptr_42_value ? ghv_7 : _GEN_6789; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6791 = 8'h8 == new_ptr_42_value ? ghv_8 : _GEN_6790; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6792 = 8'h9 == new_ptr_42_value ? ghv_9 : _GEN_6791; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6793 = 8'ha == new_ptr_42_value ? ghv_10 : _GEN_6792; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6794 = 8'hb == new_ptr_42_value ? ghv_11 : _GEN_6793; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6795 = 8'hc == new_ptr_42_value ? ghv_12 : _GEN_6794; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6796 = 8'hd == new_ptr_42_value ? ghv_13 : _GEN_6795; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6797 = 8'he == new_ptr_42_value ? ghv_14 : _GEN_6796; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6798 = 8'hf == new_ptr_42_value ? ghv_15 : _GEN_6797; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6799 = 8'h10 == new_ptr_42_value ? ghv_16 : _GEN_6798; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6800 = 8'h11 == new_ptr_42_value ? ghv_17 : _GEN_6799; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6801 = 8'h12 == new_ptr_42_value ? ghv_18 : _GEN_6800; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6802 = 8'h13 == new_ptr_42_value ? ghv_19 : _GEN_6801; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6803 = 8'h14 == new_ptr_42_value ? ghv_20 : _GEN_6802; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6804 = 8'h15 == new_ptr_42_value ? ghv_21 : _GEN_6803; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6805 = 8'h16 == new_ptr_42_value ? ghv_22 : _GEN_6804; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6806 = 8'h17 == new_ptr_42_value ? ghv_23 : _GEN_6805; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6807 = 8'h18 == new_ptr_42_value ? ghv_24 : _GEN_6806; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6808 = 8'h19 == new_ptr_42_value ? ghv_25 : _GEN_6807; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6809 = 8'h1a == new_ptr_42_value ? ghv_26 : _GEN_6808; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6810 = 8'h1b == new_ptr_42_value ? ghv_27 : _GEN_6809; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6811 = 8'h1c == new_ptr_42_value ? ghv_28 : _GEN_6810; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6812 = 8'h1d == new_ptr_42_value ? ghv_29 : _GEN_6811; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6813 = 8'h1e == new_ptr_42_value ? ghv_30 : _GEN_6812; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6814 = 8'h1f == new_ptr_42_value ? ghv_31 : _GEN_6813; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6815 = 8'h20 == new_ptr_42_value ? ghv_32 : _GEN_6814; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6816 = 8'h21 == new_ptr_42_value ? ghv_33 : _GEN_6815; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6817 = 8'h22 == new_ptr_42_value ? ghv_34 : _GEN_6816; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6818 = 8'h23 == new_ptr_42_value ? ghv_35 : _GEN_6817; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6819 = 8'h24 == new_ptr_42_value ? ghv_36 : _GEN_6818; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6820 = 8'h25 == new_ptr_42_value ? ghv_37 : _GEN_6819; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6821 = 8'h26 == new_ptr_42_value ? ghv_38 : _GEN_6820; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6822 = 8'h27 == new_ptr_42_value ? ghv_39 : _GEN_6821; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6823 = 8'h28 == new_ptr_42_value ? ghv_40 : _GEN_6822; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6824 = 8'h29 == new_ptr_42_value ? ghv_41 : _GEN_6823; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6825 = 8'h2a == new_ptr_42_value ? ghv_42 : _GEN_6824; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6826 = 8'h2b == new_ptr_42_value ? ghv_43 : _GEN_6825; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6827 = 8'h2c == new_ptr_42_value ? ghv_44 : _GEN_6826; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6828 = 8'h2d == new_ptr_42_value ? ghv_45 : _GEN_6827; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6829 = 8'h2e == new_ptr_42_value ? ghv_46 : _GEN_6828; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6830 = 8'h2f == new_ptr_42_value ? ghv_47 : _GEN_6829; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6831 = 8'h30 == new_ptr_42_value ? ghv_48 : _GEN_6830; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6832 = 8'h31 == new_ptr_42_value ? ghv_49 : _GEN_6831; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6833 = 8'h32 == new_ptr_42_value ? ghv_50 : _GEN_6832; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6834 = 8'h33 == new_ptr_42_value ? ghv_51 : _GEN_6833; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6835 = 8'h34 == new_ptr_42_value ? ghv_52 : _GEN_6834; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6836 = 8'h35 == new_ptr_42_value ? ghv_53 : _GEN_6835; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6837 = 8'h36 == new_ptr_42_value ? ghv_54 : _GEN_6836; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6838 = 8'h37 == new_ptr_42_value ? ghv_55 : _GEN_6837; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6839 = 8'h38 == new_ptr_42_value ? ghv_56 : _GEN_6838; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6840 = 8'h39 == new_ptr_42_value ? ghv_57 : _GEN_6839; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6841 = 8'h3a == new_ptr_42_value ? ghv_58 : _GEN_6840; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6842 = 8'h3b == new_ptr_42_value ? ghv_59 : _GEN_6841; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6843 = 8'h3c == new_ptr_42_value ? ghv_60 : _GEN_6842; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6844 = 8'h3d == new_ptr_42_value ? ghv_61 : _GEN_6843; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6845 = 8'h3e == new_ptr_42_value ? ghv_62 : _GEN_6844; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6846 = 8'h3f == new_ptr_42_value ? ghv_63 : _GEN_6845; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6847 = 8'h40 == new_ptr_42_value ? ghv_64 : _GEN_6846; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6848 = 8'h41 == new_ptr_42_value ? ghv_65 : _GEN_6847; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6849 = 8'h42 == new_ptr_42_value ? ghv_66 : _GEN_6848; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6850 = 8'h43 == new_ptr_42_value ? ghv_67 : _GEN_6849; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6851 = 8'h44 == new_ptr_42_value ? ghv_68 : _GEN_6850; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6852 = 8'h45 == new_ptr_42_value ? ghv_69 : _GEN_6851; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6853 = 8'h46 == new_ptr_42_value ? ghv_70 : _GEN_6852; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6854 = 8'h47 == new_ptr_42_value ? ghv_71 : _GEN_6853; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6855 = 8'h48 == new_ptr_42_value ? ghv_72 : _GEN_6854; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6856 = 8'h49 == new_ptr_42_value ? ghv_73 : _GEN_6855; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6857 = 8'h4a == new_ptr_42_value ? ghv_74 : _GEN_6856; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6858 = 8'h4b == new_ptr_42_value ? ghv_75 : _GEN_6857; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6859 = 8'h4c == new_ptr_42_value ? ghv_76 : _GEN_6858; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6860 = 8'h4d == new_ptr_42_value ? ghv_77 : _GEN_6859; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6861 = 8'h4e == new_ptr_42_value ? ghv_78 : _GEN_6860; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6862 = 8'h4f == new_ptr_42_value ? ghv_79 : _GEN_6861; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6863 = 8'h50 == new_ptr_42_value ? ghv_80 : _GEN_6862; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6864 = 8'h51 == new_ptr_42_value ? ghv_81 : _GEN_6863; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6865 = 8'h52 == new_ptr_42_value ? ghv_82 : _GEN_6864; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6866 = 8'h53 == new_ptr_42_value ? ghv_83 : _GEN_6865; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6867 = 8'h54 == new_ptr_42_value ? ghv_84 : _GEN_6866; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6868 = 8'h55 == new_ptr_42_value ? ghv_85 : _GEN_6867; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6869 = 8'h56 == new_ptr_42_value ? ghv_86 : _GEN_6868; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6870 = 8'h57 == new_ptr_42_value ? ghv_87 : _GEN_6869; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6871 = 8'h58 == new_ptr_42_value ? ghv_88 : _GEN_6870; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6872 = 8'h59 == new_ptr_42_value ? ghv_89 : _GEN_6871; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6873 = 8'h5a == new_ptr_42_value ? ghv_90 : _GEN_6872; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6874 = 8'h5b == new_ptr_42_value ? ghv_91 : _GEN_6873; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6875 = 8'h5c == new_ptr_42_value ? ghv_92 : _GEN_6874; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6876 = 8'h5d == new_ptr_42_value ? ghv_93 : _GEN_6875; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6877 = 8'h5e == new_ptr_42_value ? ghv_94 : _GEN_6876; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6878 = 8'h5f == new_ptr_42_value ? ghv_95 : _GEN_6877; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6879 = 8'h60 == new_ptr_42_value ? ghv_96 : _GEN_6878; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6880 = 8'h61 == new_ptr_42_value ? ghv_97 : _GEN_6879; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6881 = 8'h62 == new_ptr_42_value ? ghv_98 : _GEN_6880; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6882 = 8'h63 == new_ptr_42_value ? ghv_99 : _GEN_6881; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6883 = 8'h64 == new_ptr_42_value ? ghv_100 : _GEN_6882; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6884 = 8'h65 == new_ptr_42_value ? ghv_101 : _GEN_6883; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6885 = 8'h66 == new_ptr_42_value ? ghv_102 : _GEN_6884; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6886 = 8'h67 == new_ptr_42_value ? ghv_103 : _GEN_6885; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6887 = 8'h68 == new_ptr_42_value ? ghv_104 : _GEN_6886; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6888 = 8'h69 == new_ptr_42_value ? ghv_105 : _GEN_6887; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6889 = 8'h6a == new_ptr_42_value ? ghv_106 : _GEN_6888; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6890 = 8'h6b == new_ptr_42_value ? ghv_107 : _GEN_6889; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6891 = 8'h6c == new_ptr_42_value ? ghv_108 : _GEN_6890; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6892 = 8'h6d == new_ptr_42_value ? ghv_109 : _GEN_6891; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6893 = 8'h6e == new_ptr_42_value ? ghv_110 : _GEN_6892; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6894 = 8'h6f == new_ptr_42_value ? ghv_111 : _GEN_6893; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6895 = 8'h70 == new_ptr_42_value ? ghv_112 : _GEN_6894; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6896 = 8'h71 == new_ptr_42_value ? ghv_113 : _GEN_6895; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6897 = 8'h72 == new_ptr_42_value ? ghv_114 : _GEN_6896; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6898 = 8'h73 == new_ptr_42_value ? ghv_115 : _GEN_6897; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6899 = 8'h74 == new_ptr_42_value ? ghv_116 : _GEN_6898; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6900 = 8'h75 == new_ptr_42_value ? ghv_117 : _GEN_6899; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6901 = 8'h76 == new_ptr_42_value ? ghv_118 : _GEN_6900; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6902 = 8'h77 == new_ptr_42_value ? ghv_119 : _GEN_6901; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6903 = 8'h78 == new_ptr_42_value ? ghv_120 : _GEN_6902; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6904 = 8'h79 == new_ptr_42_value ? ghv_121 : _GEN_6903; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6905 = 8'h7a == new_ptr_42_value ? ghv_122 : _GEN_6904; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6906 = 8'h7b == new_ptr_42_value ? ghv_123 : _GEN_6905; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6907 = 8'h7c == new_ptr_42_value ? ghv_124 : _GEN_6906; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6908 = 8'h7d == new_ptr_42_value ? ghv_125 : _GEN_6907; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6909 = 8'h7e == new_ptr_42_value ? ghv_126 : _GEN_6908; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6910 = 8'h7f == new_ptr_42_value ? ghv_127 : _GEN_6909; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6911 = 8'h80 == new_ptr_42_value ? ghv_128 : _GEN_6910; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6912 = 8'h81 == new_ptr_42_value ? ghv_129 : _GEN_6911; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6913 = 8'h82 == new_ptr_42_value ? ghv_130 : _GEN_6912; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6914 = 8'h83 == new_ptr_42_value ? ghv_131 : _GEN_6913; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6915 = 8'h84 == new_ptr_42_value ? ghv_132 : _GEN_6914; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6916 = 8'h85 == new_ptr_42_value ? ghv_133 : _GEN_6915; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6917 = 8'h86 == new_ptr_42_value ? ghv_134 : _GEN_6916; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6918 = 8'h87 == new_ptr_42_value ? ghv_135 : _GEN_6917; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6919 = 8'h88 == new_ptr_42_value ? ghv_136 : _GEN_6918; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6920 = 8'h89 == new_ptr_42_value ? ghv_137 : _GEN_6919; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6921 = 8'h8a == new_ptr_42_value ? ghv_138 : _GEN_6920; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6922 = 8'h8b == new_ptr_42_value ? ghv_139 : _GEN_6921; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6923 = 8'h8c == new_ptr_42_value ? ghv_140 : _GEN_6922; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6924 = 8'h8d == new_ptr_42_value ? ghv_141 : _GEN_6923; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6925 = 8'h8e == new_ptr_42_value ? ghv_142 : _GEN_6924; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_54_value = _new_ptr_value_T_109[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_6928 = 8'h1 == new_ptr_54_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6929 = 8'h2 == new_ptr_54_value ? ghv_2 : _GEN_6928; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6930 = 8'h3 == new_ptr_54_value ? ghv_3 : _GEN_6929; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6931 = 8'h4 == new_ptr_54_value ? ghv_4 : _GEN_6930; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6932 = 8'h5 == new_ptr_54_value ? ghv_5 : _GEN_6931; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6933 = 8'h6 == new_ptr_54_value ? ghv_6 : _GEN_6932; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6934 = 8'h7 == new_ptr_54_value ? ghv_7 : _GEN_6933; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6935 = 8'h8 == new_ptr_54_value ? ghv_8 : _GEN_6934; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6936 = 8'h9 == new_ptr_54_value ? ghv_9 : _GEN_6935; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6937 = 8'ha == new_ptr_54_value ? ghv_10 : _GEN_6936; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6938 = 8'hb == new_ptr_54_value ? ghv_11 : _GEN_6937; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6939 = 8'hc == new_ptr_54_value ? ghv_12 : _GEN_6938; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6940 = 8'hd == new_ptr_54_value ? ghv_13 : _GEN_6939; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6941 = 8'he == new_ptr_54_value ? ghv_14 : _GEN_6940; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6942 = 8'hf == new_ptr_54_value ? ghv_15 : _GEN_6941; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6943 = 8'h10 == new_ptr_54_value ? ghv_16 : _GEN_6942; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6944 = 8'h11 == new_ptr_54_value ? ghv_17 : _GEN_6943; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6945 = 8'h12 == new_ptr_54_value ? ghv_18 : _GEN_6944; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6946 = 8'h13 == new_ptr_54_value ? ghv_19 : _GEN_6945; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6947 = 8'h14 == new_ptr_54_value ? ghv_20 : _GEN_6946; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6948 = 8'h15 == new_ptr_54_value ? ghv_21 : _GEN_6947; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6949 = 8'h16 == new_ptr_54_value ? ghv_22 : _GEN_6948; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6950 = 8'h17 == new_ptr_54_value ? ghv_23 : _GEN_6949; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6951 = 8'h18 == new_ptr_54_value ? ghv_24 : _GEN_6950; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6952 = 8'h19 == new_ptr_54_value ? ghv_25 : _GEN_6951; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6953 = 8'h1a == new_ptr_54_value ? ghv_26 : _GEN_6952; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6954 = 8'h1b == new_ptr_54_value ? ghv_27 : _GEN_6953; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6955 = 8'h1c == new_ptr_54_value ? ghv_28 : _GEN_6954; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6956 = 8'h1d == new_ptr_54_value ? ghv_29 : _GEN_6955; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6957 = 8'h1e == new_ptr_54_value ? ghv_30 : _GEN_6956; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6958 = 8'h1f == new_ptr_54_value ? ghv_31 : _GEN_6957; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6959 = 8'h20 == new_ptr_54_value ? ghv_32 : _GEN_6958; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6960 = 8'h21 == new_ptr_54_value ? ghv_33 : _GEN_6959; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6961 = 8'h22 == new_ptr_54_value ? ghv_34 : _GEN_6960; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6962 = 8'h23 == new_ptr_54_value ? ghv_35 : _GEN_6961; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6963 = 8'h24 == new_ptr_54_value ? ghv_36 : _GEN_6962; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6964 = 8'h25 == new_ptr_54_value ? ghv_37 : _GEN_6963; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6965 = 8'h26 == new_ptr_54_value ? ghv_38 : _GEN_6964; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6966 = 8'h27 == new_ptr_54_value ? ghv_39 : _GEN_6965; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6967 = 8'h28 == new_ptr_54_value ? ghv_40 : _GEN_6966; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6968 = 8'h29 == new_ptr_54_value ? ghv_41 : _GEN_6967; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6969 = 8'h2a == new_ptr_54_value ? ghv_42 : _GEN_6968; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6970 = 8'h2b == new_ptr_54_value ? ghv_43 : _GEN_6969; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6971 = 8'h2c == new_ptr_54_value ? ghv_44 : _GEN_6970; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6972 = 8'h2d == new_ptr_54_value ? ghv_45 : _GEN_6971; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6973 = 8'h2e == new_ptr_54_value ? ghv_46 : _GEN_6972; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6974 = 8'h2f == new_ptr_54_value ? ghv_47 : _GEN_6973; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6975 = 8'h30 == new_ptr_54_value ? ghv_48 : _GEN_6974; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6976 = 8'h31 == new_ptr_54_value ? ghv_49 : _GEN_6975; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6977 = 8'h32 == new_ptr_54_value ? ghv_50 : _GEN_6976; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6978 = 8'h33 == new_ptr_54_value ? ghv_51 : _GEN_6977; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6979 = 8'h34 == new_ptr_54_value ? ghv_52 : _GEN_6978; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6980 = 8'h35 == new_ptr_54_value ? ghv_53 : _GEN_6979; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6981 = 8'h36 == new_ptr_54_value ? ghv_54 : _GEN_6980; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6982 = 8'h37 == new_ptr_54_value ? ghv_55 : _GEN_6981; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6983 = 8'h38 == new_ptr_54_value ? ghv_56 : _GEN_6982; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6984 = 8'h39 == new_ptr_54_value ? ghv_57 : _GEN_6983; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6985 = 8'h3a == new_ptr_54_value ? ghv_58 : _GEN_6984; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6986 = 8'h3b == new_ptr_54_value ? ghv_59 : _GEN_6985; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6987 = 8'h3c == new_ptr_54_value ? ghv_60 : _GEN_6986; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6988 = 8'h3d == new_ptr_54_value ? ghv_61 : _GEN_6987; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6989 = 8'h3e == new_ptr_54_value ? ghv_62 : _GEN_6988; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6990 = 8'h3f == new_ptr_54_value ? ghv_63 : _GEN_6989; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6991 = 8'h40 == new_ptr_54_value ? ghv_64 : _GEN_6990; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6992 = 8'h41 == new_ptr_54_value ? ghv_65 : _GEN_6991; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6993 = 8'h42 == new_ptr_54_value ? ghv_66 : _GEN_6992; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6994 = 8'h43 == new_ptr_54_value ? ghv_67 : _GEN_6993; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6995 = 8'h44 == new_ptr_54_value ? ghv_68 : _GEN_6994; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6996 = 8'h45 == new_ptr_54_value ? ghv_69 : _GEN_6995; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6997 = 8'h46 == new_ptr_54_value ? ghv_70 : _GEN_6996; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6998 = 8'h47 == new_ptr_54_value ? ghv_71 : _GEN_6997; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_6999 = 8'h48 == new_ptr_54_value ? ghv_72 : _GEN_6998; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7000 = 8'h49 == new_ptr_54_value ? ghv_73 : _GEN_6999; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7001 = 8'h4a == new_ptr_54_value ? ghv_74 : _GEN_7000; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7002 = 8'h4b == new_ptr_54_value ? ghv_75 : _GEN_7001; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7003 = 8'h4c == new_ptr_54_value ? ghv_76 : _GEN_7002; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7004 = 8'h4d == new_ptr_54_value ? ghv_77 : _GEN_7003; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7005 = 8'h4e == new_ptr_54_value ? ghv_78 : _GEN_7004; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7006 = 8'h4f == new_ptr_54_value ? ghv_79 : _GEN_7005; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7007 = 8'h50 == new_ptr_54_value ? ghv_80 : _GEN_7006; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7008 = 8'h51 == new_ptr_54_value ? ghv_81 : _GEN_7007; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7009 = 8'h52 == new_ptr_54_value ? ghv_82 : _GEN_7008; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7010 = 8'h53 == new_ptr_54_value ? ghv_83 : _GEN_7009; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7011 = 8'h54 == new_ptr_54_value ? ghv_84 : _GEN_7010; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7012 = 8'h55 == new_ptr_54_value ? ghv_85 : _GEN_7011; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7013 = 8'h56 == new_ptr_54_value ? ghv_86 : _GEN_7012; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7014 = 8'h57 == new_ptr_54_value ? ghv_87 : _GEN_7013; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7015 = 8'h58 == new_ptr_54_value ? ghv_88 : _GEN_7014; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7016 = 8'h59 == new_ptr_54_value ? ghv_89 : _GEN_7015; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7017 = 8'h5a == new_ptr_54_value ? ghv_90 : _GEN_7016; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7018 = 8'h5b == new_ptr_54_value ? ghv_91 : _GEN_7017; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7019 = 8'h5c == new_ptr_54_value ? ghv_92 : _GEN_7018; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7020 = 8'h5d == new_ptr_54_value ? ghv_93 : _GEN_7019; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7021 = 8'h5e == new_ptr_54_value ? ghv_94 : _GEN_7020; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7022 = 8'h5f == new_ptr_54_value ? ghv_95 : _GEN_7021; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7023 = 8'h60 == new_ptr_54_value ? ghv_96 : _GEN_7022; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7024 = 8'h61 == new_ptr_54_value ? ghv_97 : _GEN_7023; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7025 = 8'h62 == new_ptr_54_value ? ghv_98 : _GEN_7024; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7026 = 8'h63 == new_ptr_54_value ? ghv_99 : _GEN_7025; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7027 = 8'h64 == new_ptr_54_value ? ghv_100 : _GEN_7026; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7028 = 8'h65 == new_ptr_54_value ? ghv_101 : _GEN_7027; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7029 = 8'h66 == new_ptr_54_value ? ghv_102 : _GEN_7028; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7030 = 8'h67 == new_ptr_54_value ? ghv_103 : _GEN_7029; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7031 = 8'h68 == new_ptr_54_value ? ghv_104 : _GEN_7030; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7032 = 8'h69 == new_ptr_54_value ? ghv_105 : _GEN_7031; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7033 = 8'h6a == new_ptr_54_value ? ghv_106 : _GEN_7032; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7034 = 8'h6b == new_ptr_54_value ? ghv_107 : _GEN_7033; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7035 = 8'h6c == new_ptr_54_value ? ghv_108 : _GEN_7034; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7036 = 8'h6d == new_ptr_54_value ? ghv_109 : _GEN_7035; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7037 = 8'h6e == new_ptr_54_value ? ghv_110 : _GEN_7036; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7038 = 8'h6f == new_ptr_54_value ? ghv_111 : _GEN_7037; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7039 = 8'h70 == new_ptr_54_value ? ghv_112 : _GEN_7038; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7040 = 8'h71 == new_ptr_54_value ? ghv_113 : _GEN_7039; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7041 = 8'h72 == new_ptr_54_value ? ghv_114 : _GEN_7040; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7042 = 8'h73 == new_ptr_54_value ? ghv_115 : _GEN_7041; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7043 = 8'h74 == new_ptr_54_value ? ghv_116 : _GEN_7042; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7044 = 8'h75 == new_ptr_54_value ? ghv_117 : _GEN_7043; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7045 = 8'h76 == new_ptr_54_value ? ghv_118 : _GEN_7044; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7046 = 8'h77 == new_ptr_54_value ? ghv_119 : _GEN_7045; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7047 = 8'h78 == new_ptr_54_value ? ghv_120 : _GEN_7046; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7048 = 8'h79 == new_ptr_54_value ? ghv_121 : _GEN_7047; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7049 = 8'h7a == new_ptr_54_value ? ghv_122 : _GEN_7048; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7050 = 8'h7b == new_ptr_54_value ? ghv_123 : _GEN_7049; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7051 = 8'h7c == new_ptr_54_value ? ghv_124 : _GEN_7050; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7052 = 8'h7d == new_ptr_54_value ? ghv_125 : _GEN_7051; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7053 = 8'h7e == new_ptr_54_value ? ghv_126 : _GEN_7052; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7054 = 8'h7f == new_ptr_54_value ? ghv_127 : _GEN_7053; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7055 = 8'h80 == new_ptr_54_value ? ghv_128 : _GEN_7054; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7056 = 8'h81 == new_ptr_54_value ? ghv_129 : _GEN_7055; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7057 = 8'h82 == new_ptr_54_value ? ghv_130 : _GEN_7056; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7058 = 8'h83 == new_ptr_54_value ? ghv_131 : _GEN_7057; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7059 = 8'h84 == new_ptr_54_value ? ghv_132 : _GEN_7058; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7060 = 8'h85 == new_ptr_54_value ? ghv_133 : _GEN_7059; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7061 = 8'h86 == new_ptr_54_value ? ghv_134 : _GEN_7060; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7062 = 8'h87 == new_ptr_54_value ? ghv_135 : _GEN_7061; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7063 = 8'h88 == new_ptr_54_value ? ghv_136 : _GEN_7062; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7064 = 8'h89 == new_ptr_54_value ? ghv_137 : _GEN_7063; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7065 = 8'h8a == new_ptr_54_value ? ghv_138 : _GEN_7064; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7066 = 8'h8b == new_ptr_54_value ? ghv_139 : _GEN_7065; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7067 = 8'h8c == new_ptr_54_value ? ghv_140 : _GEN_7066; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7068 = 8'h8d == new_ptr_54_value ? ghv_141 : _GEN_7067; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7069 = 8'h8e == new_ptr_54_value ? ghv_142 : _GEN_7068; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_57_value = _new_ptr_value_T_115[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_7072 = 8'h1 == new_ptr_57_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7073 = 8'h2 == new_ptr_57_value ? ghv_2 : _GEN_7072; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7074 = 8'h3 == new_ptr_57_value ? ghv_3 : _GEN_7073; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7075 = 8'h4 == new_ptr_57_value ? ghv_4 : _GEN_7074; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7076 = 8'h5 == new_ptr_57_value ? ghv_5 : _GEN_7075; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7077 = 8'h6 == new_ptr_57_value ? ghv_6 : _GEN_7076; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7078 = 8'h7 == new_ptr_57_value ? ghv_7 : _GEN_7077; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7079 = 8'h8 == new_ptr_57_value ? ghv_8 : _GEN_7078; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7080 = 8'h9 == new_ptr_57_value ? ghv_9 : _GEN_7079; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7081 = 8'ha == new_ptr_57_value ? ghv_10 : _GEN_7080; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7082 = 8'hb == new_ptr_57_value ? ghv_11 : _GEN_7081; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7083 = 8'hc == new_ptr_57_value ? ghv_12 : _GEN_7082; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7084 = 8'hd == new_ptr_57_value ? ghv_13 : _GEN_7083; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7085 = 8'he == new_ptr_57_value ? ghv_14 : _GEN_7084; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7086 = 8'hf == new_ptr_57_value ? ghv_15 : _GEN_7085; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7087 = 8'h10 == new_ptr_57_value ? ghv_16 : _GEN_7086; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7088 = 8'h11 == new_ptr_57_value ? ghv_17 : _GEN_7087; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7089 = 8'h12 == new_ptr_57_value ? ghv_18 : _GEN_7088; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7090 = 8'h13 == new_ptr_57_value ? ghv_19 : _GEN_7089; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7091 = 8'h14 == new_ptr_57_value ? ghv_20 : _GEN_7090; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7092 = 8'h15 == new_ptr_57_value ? ghv_21 : _GEN_7091; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7093 = 8'h16 == new_ptr_57_value ? ghv_22 : _GEN_7092; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7094 = 8'h17 == new_ptr_57_value ? ghv_23 : _GEN_7093; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7095 = 8'h18 == new_ptr_57_value ? ghv_24 : _GEN_7094; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7096 = 8'h19 == new_ptr_57_value ? ghv_25 : _GEN_7095; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7097 = 8'h1a == new_ptr_57_value ? ghv_26 : _GEN_7096; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7098 = 8'h1b == new_ptr_57_value ? ghv_27 : _GEN_7097; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7099 = 8'h1c == new_ptr_57_value ? ghv_28 : _GEN_7098; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7100 = 8'h1d == new_ptr_57_value ? ghv_29 : _GEN_7099; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7101 = 8'h1e == new_ptr_57_value ? ghv_30 : _GEN_7100; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7102 = 8'h1f == new_ptr_57_value ? ghv_31 : _GEN_7101; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7103 = 8'h20 == new_ptr_57_value ? ghv_32 : _GEN_7102; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7104 = 8'h21 == new_ptr_57_value ? ghv_33 : _GEN_7103; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7105 = 8'h22 == new_ptr_57_value ? ghv_34 : _GEN_7104; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7106 = 8'h23 == new_ptr_57_value ? ghv_35 : _GEN_7105; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7107 = 8'h24 == new_ptr_57_value ? ghv_36 : _GEN_7106; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7108 = 8'h25 == new_ptr_57_value ? ghv_37 : _GEN_7107; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7109 = 8'h26 == new_ptr_57_value ? ghv_38 : _GEN_7108; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7110 = 8'h27 == new_ptr_57_value ? ghv_39 : _GEN_7109; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7111 = 8'h28 == new_ptr_57_value ? ghv_40 : _GEN_7110; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7112 = 8'h29 == new_ptr_57_value ? ghv_41 : _GEN_7111; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7113 = 8'h2a == new_ptr_57_value ? ghv_42 : _GEN_7112; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7114 = 8'h2b == new_ptr_57_value ? ghv_43 : _GEN_7113; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7115 = 8'h2c == new_ptr_57_value ? ghv_44 : _GEN_7114; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7116 = 8'h2d == new_ptr_57_value ? ghv_45 : _GEN_7115; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7117 = 8'h2e == new_ptr_57_value ? ghv_46 : _GEN_7116; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7118 = 8'h2f == new_ptr_57_value ? ghv_47 : _GEN_7117; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7119 = 8'h30 == new_ptr_57_value ? ghv_48 : _GEN_7118; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7120 = 8'h31 == new_ptr_57_value ? ghv_49 : _GEN_7119; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7121 = 8'h32 == new_ptr_57_value ? ghv_50 : _GEN_7120; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7122 = 8'h33 == new_ptr_57_value ? ghv_51 : _GEN_7121; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7123 = 8'h34 == new_ptr_57_value ? ghv_52 : _GEN_7122; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7124 = 8'h35 == new_ptr_57_value ? ghv_53 : _GEN_7123; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7125 = 8'h36 == new_ptr_57_value ? ghv_54 : _GEN_7124; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7126 = 8'h37 == new_ptr_57_value ? ghv_55 : _GEN_7125; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7127 = 8'h38 == new_ptr_57_value ? ghv_56 : _GEN_7126; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7128 = 8'h39 == new_ptr_57_value ? ghv_57 : _GEN_7127; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7129 = 8'h3a == new_ptr_57_value ? ghv_58 : _GEN_7128; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7130 = 8'h3b == new_ptr_57_value ? ghv_59 : _GEN_7129; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7131 = 8'h3c == new_ptr_57_value ? ghv_60 : _GEN_7130; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7132 = 8'h3d == new_ptr_57_value ? ghv_61 : _GEN_7131; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7133 = 8'h3e == new_ptr_57_value ? ghv_62 : _GEN_7132; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7134 = 8'h3f == new_ptr_57_value ? ghv_63 : _GEN_7133; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7135 = 8'h40 == new_ptr_57_value ? ghv_64 : _GEN_7134; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7136 = 8'h41 == new_ptr_57_value ? ghv_65 : _GEN_7135; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7137 = 8'h42 == new_ptr_57_value ? ghv_66 : _GEN_7136; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7138 = 8'h43 == new_ptr_57_value ? ghv_67 : _GEN_7137; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7139 = 8'h44 == new_ptr_57_value ? ghv_68 : _GEN_7138; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7140 = 8'h45 == new_ptr_57_value ? ghv_69 : _GEN_7139; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7141 = 8'h46 == new_ptr_57_value ? ghv_70 : _GEN_7140; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7142 = 8'h47 == new_ptr_57_value ? ghv_71 : _GEN_7141; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7143 = 8'h48 == new_ptr_57_value ? ghv_72 : _GEN_7142; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7144 = 8'h49 == new_ptr_57_value ? ghv_73 : _GEN_7143; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7145 = 8'h4a == new_ptr_57_value ? ghv_74 : _GEN_7144; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7146 = 8'h4b == new_ptr_57_value ? ghv_75 : _GEN_7145; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7147 = 8'h4c == new_ptr_57_value ? ghv_76 : _GEN_7146; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7148 = 8'h4d == new_ptr_57_value ? ghv_77 : _GEN_7147; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7149 = 8'h4e == new_ptr_57_value ? ghv_78 : _GEN_7148; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7150 = 8'h4f == new_ptr_57_value ? ghv_79 : _GEN_7149; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7151 = 8'h50 == new_ptr_57_value ? ghv_80 : _GEN_7150; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7152 = 8'h51 == new_ptr_57_value ? ghv_81 : _GEN_7151; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7153 = 8'h52 == new_ptr_57_value ? ghv_82 : _GEN_7152; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7154 = 8'h53 == new_ptr_57_value ? ghv_83 : _GEN_7153; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7155 = 8'h54 == new_ptr_57_value ? ghv_84 : _GEN_7154; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7156 = 8'h55 == new_ptr_57_value ? ghv_85 : _GEN_7155; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7157 = 8'h56 == new_ptr_57_value ? ghv_86 : _GEN_7156; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7158 = 8'h57 == new_ptr_57_value ? ghv_87 : _GEN_7157; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7159 = 8'h58 == new_ptr_57_value ? ghv_88 : _GEN_7158; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7160 = 8'h59 == new_ptr_57_value ? ghv_89 : _GEN_7159; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7161 = 8'h5a == new_ptr_57_value ? ghv_90 : _GEN_7160; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7162 = 8'h5b == new_ptr_57_value ? ghv_91 : _GEN_7161; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7163 = 8'h5c == new_ptr_57_value ? ghv_92 : _GEN_7162; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7164 = 8'h5d == new_ptr_57_value ? ghv_93 : _GEN_7163; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7165 = 8'h5e == new_ptr_57_value ? ghv_94 : _GEN_7164; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7166 = 8'h5f == new_ptr_57_value ? ghv_95 : _GEN_7165; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7167 = 8'h60 == new_ptr_57_value ? ghv_96 : _GEN_7166; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7168 = 8'h61 == new_ptr_57_value ? ghv_97 : _GEN_7167; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7169 = 8'h62 == new_ptr_57_value ? ghv_98 : _GEN_7168; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7170 = 8'h63 == new_ptr_57_value ? ghv_99 : _GEN_7169; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7171 = 8'h64 == new_ptr_57_value ? ghv_100 : _GEN_7170; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7172 = 8'h65 == new_ptr_57_value ? ghv_101 : _GEN_7171; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7173 = 8'h66 == new_ptr_57_value ? ghv_102 : _GEN_7172; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7174 = 8'h67 == new_ptr_57_value ? ghv_103 : _GEN_7173; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7175 = 8'h68 == new_ptr_57_value ? ghv_104 : _GEN_7174; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7176 = 8'h69 == new_ptr_57_value ? ghv_105 : _GEN_7175; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7177 = 8'h6a == new_ptr_57_value ? ghv_106 : _GEN_7176; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7178 = 8'h6b == new_ptr_57_value ? ghv_107 : _GEN_7177; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7179 = 8'h6c == new_ptr_57_value ? ghv_108 : _GEN_7178; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7180 = 8'h6d == new_ptr_57_value ? ghv_109 : _GEN_7179; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7181 = 8'h6e == new_ptr_57_value ? ghv_110 : _GEN_7180; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7182 = 8'h6f == new_ptr_57_value ? ghv_111 : _GEN_7181; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7183 = 8'h70 == new_ptr_57_value ? ghv_112 : _GEN_7182; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7184 = 8'h71 == new_ptr_57_value ? ghv_113 : _GEN_7183; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7185 = 8'h72 == new_ptr_57_value ? ghv_114 : _GEN_7184; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7186 = 8'h73 == new_ptr_57_value ? ghv_115 : _GEN_7185; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7187 = 8'h74 == new_ptr_57_value ? ghv_116 : _GEN_7186; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7188 = 8'h75 == new_ptr_57_value ? ghv_117 : _GEN_7187; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7189 = 8'h76 == new_ptr_57_value ? ghv_118 : _GEN_7188; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7190 = 8'h77 == new_ptr_57_value ? ghv_119 : _GEN_7189; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7191 = 8'h78 == new_ptr_57_value ? ghv_120 : _GEN_7190; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7192 = 8'h79 == new_ptr_57_value ? ghv_121 : _GEN_7191; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7193 = 8'h7a == new_ptr_57_value ? ghv_122 : _GEN_7192; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7194 = 8'h7b == new_ptr_57_value ? ghv_123 : _GEN_7193; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7195 = 8'h7c == new_ptr_57_value ? ghv_124 : _GEN_7194; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7196 = 8'h7d == new_ptr_57_value ? ghv_125 : _GEN_7195; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7197 = 8'h7e == new_ptr_57_value ? ghv_126 : _GEN_7196; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7198 = 8'h7f == new_ptr_57_value ? ghv_127 : _GEN_7197; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7199 = 8'h80 == new_ptr_57_value ? ghv_128 : _GEN_7198; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7200 = 8'h81 == new_ptr_57_value ? ghv_129 : _GEN_7199; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7201 = 8'h82 == new_ptr_57_value ? ghv_130 : _GEN_7200; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7202 = 8'h83 == new_ptr_57_value ? ghv_131 : _GEN_7201; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7203 = 8'h84 == new_ptr_57_value ? ghv_132 : _GEN_7202; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7204 = 8'h85 == new_ptr_57_value ? ghv_133 : _GEN_7203; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7205 = 8'h86 == new_ptr_57_value ? ghv_134 : _GEN_7204; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7206 = 8'h87 == new_ptr_57_value ? ghv_135 : _GEN_7205; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7207 = 8'h88 == new_ptr_57_value ? ghv_136 : _GEN_7206; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7208 = 8'h89 == new_ptr_57_value ? ghv_137 : _GEN_7207; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7209 = 8'h8a == new_ptr_57_value ? ghv_138 : _GEN_7208; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7210 = 8'h8b == new_ptr_57_value ? ghv_139 : _GEN_7209; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7211 = 8'h8c == new_ptr_57_value ? ghv_140 : _GEN_7210; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7212 = 8'h8d == new_ptr_57_value ? ghv_141 : _GEN_7211; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7213 = 8'h8e == new_ptr_57_value ? ghv_142 : _GEN_7212; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_44_value = _new_ptr_value_T_89[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_7216 = 8'h1 == new_ptr_44_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7217 = 8'h2 == new_ptr_44_value ? ghv_2 : _GEN_7216; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7218 = 8'h3 == new_ptr_44_value ? ghv_3 : _GEN_7217; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7219 = 8'h4 == new_ptr_44_value ? ghv_4 : _GEN_7218; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7220 = 8'h5 == new_ptr_44_value ? ghv_5 : _GEN_7219; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7221 = 8'h6 == new_ptr_44_value ? ghv_6 : _GEN_7220; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7222 = 8'h7 == new_ptr_44_value ? ghv_7 : _GEN_7221; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7223 = 8'h8 == new_ptr_44_value ? ghv_8 : _GEN_7222; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7224 = 8'h9 == new_ptr_44_value ? ghv_9 : _GEN_7223; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7225 = 8'ha == new_ptr_44_value ? ghv_10 : _GEN_7224; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7226 = 8'hb == new_ptr_44_value ? ghv_11 : _GEN_7225; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7227 = 8'hc == new_ptr_44_value ? ghv_12 : _GEN_7226; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7228 = 8'hd == new_ptr_44_value ? ghv_13 : _GEN_7227; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7229 = 8'he == new_ptr_44_value ? ghv_14 : _GEN_7228; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7230 = 8'hf == new_ptr_44_value ? ghv_15 : _GEN_7229; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7231 = 8'h10 == new_ptr_44_value ? ghv_16 : _GEN_7230; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7232 = 8'h11 == new_ptr_44_value ? ghv_17 : _GEN_7231; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7233 = 8'h12 == new_ptr_44_value ? ghv_18 : _GEN_7232; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7234 = 8'h13 == new_ptr_44_value ? ghv_19 : _GEN_7233; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7235 = 8'h14 == new_ptr_44_value ? ghv_20 : _GEN_7234; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7236 = 8'h15 == new_ptr_44_value ? ghv_21 : _GEN_7235; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7237 = 8'h16 == new_ptr_44_value ? ghv_22 : _GEN_7236; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7238 = 8'h17 == new_ptr_44_value ? ghv_23 : _GEN_7237; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7239 = 8'h18 == new_ptr_44_value ? ghv_24 : _GEN_7238; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7240 = 8'h19 == new_ptr_44_value ? ghv_25 : _GEN_7239; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7241 = 8'h1a == new_ptr_44_value ? ghv_26 : _GEN_7240; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7242 = 8'h1b == new_ptr_44_value ? ghv_27 : _GEN_7241; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7243 = 8'h1c == new_ptr_44_value ? ghv_28 : _GEN_7242; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7244 = 8'h1d == new_ptr_44_value ? ghv_29 : _GEN_7243; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7245 = 8'h1e == new_ptr_44_value ? ghv_30 : _GEN_7244; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7246 = 8'h1f == new_ptr_44_value ? ghv_31 : _GEN_7245; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7247 = 8'h20 == new_ptr_44_value ? ghv_32 : _GEN_7246; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7248 = 8'h21 == new_ptr_44_value ? ghv_33 : _GEN_7247; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7249 = 8'h22 == new_ptr_44_value ? ghv_34 : _GEN_7248; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7250 = 8'h23 == new_ptr_44_value ? ghv_35 : _GEN_7249; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7251 = 8'h24 == new_ptr_44_value ? ghv_36 : _GEN_7250; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7252 = 8'h25 == new_ptr_44_value ? ghv_37 : _GEN_7251; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7253 = 8'h26 == new_ptr_44_value ? ghv_38 : _GEN_7252; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7254 = 8'h27 == new_ptr_44_value ? ghv_39 : _GEN_7253; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7255 = 8'h28 == new_ptr_44_value ? ghv_40 : _GEN_7254; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7256 = 8'h29 == new_ptr_44_value ? ghv_41 : _GEN_7255; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7257 = 8'h2a == new_ptr_44_value ? ghv_42 : _GEN_7256; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7258 = 8'h2b == new_ptr_44_value ? ghv_43 : _GEN_7257; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7259 = 8'h2c == new_ptr_44_value ? ghv_44 : _GEN_7258; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7260 = 8'h2d == new_ptr_44_value ? ghv_45 : _GEN_7259; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7261 = 8'h2e == new_ptr_44_value ? ghv_46 : _GEN_7260; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7262 = 8'h2f == new_ptr_44_value ? ghv_47 : _GEN_7261; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7263 = 8'h30 == new_ptr_44_value ? ghv_48 : _GEN_7262; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7264 = 8'h31 == new_ptr_44_value ? ghv_49 : _GEN_7263; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7265 = 8'h32 == new_ptr_44_value ? ghv_50 : _GEN_7264; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7266 = 8'h33 == new_ptr_44_value ? ghv_51 : _GEN_7265; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7267 = 8'h34 == new_ptr_44_value ? ghv_52 : _GEN_7266; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7268 = 8'h35 == new_ptr_44_value ? ghv_53 : _GEN_7267; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7269 = 8'h36 == new_ptr_44_value ? ghv_54 : _GEN_7268; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7270 = 8'h37 == new_ptr_44_value ? ghv_55 : _GEN_7269; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7271 = 8'h38 == new_ptr_44_value ? ghv_56 : _GEN_7270; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7272 = 8'h39 == new_ptr_44_value ? ghv_57 : _GEN_7271; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7273 = 8'h3a == new_ptr_44_value ? ghv_58 : _GEN_7272; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7274 = 8'h3b == new_ptr_44_value ? ghv_59 : _GEN_7273; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7275 = 8'h3c == new_ptr_44_value ? ghv_60 : _GEN_7274; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7276 = 8'h3d == new_ptr_44_value ? ghv_61 : _GEN_7275; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7277 = 8'h3e == new_ptr_44_value ? ghv_62 : _GEN_7276; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7278 = 8'h3f == new_ptr_44_value ? ghv_63 : _GEN_7277; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7279 = 8'h40 == new_ptr_44_value ? ghv_64 : _GEN_7278; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7280 = 8'h41 == new_ptr_44_value ? ghv_65 : _GEN_7279; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7281 = 8'h42 == new_ptr_44_value ? ghv_66 : _GEN_7280; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7282 = 8'h43 == new_ptr_44_value ? ghv_67 : _GEN_7281; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7283 = 8'h44 == new_ptr_44_value ? ghv_68 : _GEN_7282; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7284 = 8'h45 == new_ptr_44_value ? ghv_69 : _GEN_7283; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7285 = 8'h46 == new_ptr_44_value ? ghv_70 : _GEN_7284; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7286 = 8'h47 == new_ptr_44_value ? ghv_71 : _GEN_7285; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7287 = 8'h48 == new_ptr_44_value ? ghv_72 : _GEN_7286; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7288 = 8'h49 == new_ptr_44_value ? ghv_73 : _GEN_7287; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7289 = 8'h4a == new_ptr_44_value ? ghv_74 : _GEN_7288; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7290 = 8'h4b == new_ptr_44_value ? ghv_75 : _GEN_7289; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7291 = 8'h4c == new_ptr_44_value ? ghv_76 : _GEN_7290; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7292 = 8'h4d == new_ptr_44_value ? ghv_77 : _GEN_7291; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7293 = 8'h4e == new_ptr_44_value ? ghv_78 : _GEN_7292; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7294 = 8'h4f == new_ptr_44_value ? ghv_79 : _GEN_7293; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7295 = 8'h50 == new_ptr_44_value ? ghv_80 : _GEN_7294; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7296 = 8'h51 == new_ptr_44_value ? ghv_81 : _GEN_7295; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7297 = 8'h52 == new_ptr_44_value ? ghv_82 : _GEN_7296; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7298 = 8'h53 == new_ptr_44_value ? ghv_83 : _GEN_7297; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7299 = 8'h54 == new_ptr_44_value ? ghv_84 : _GEN_7298; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7300 = 8'h55 == new_ptr_44_value ? ghv_85 : _GEN_7299; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7301 = 8'h56 == new_ptr_44_value ? ghv_86 : _GEN_7300; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7302 = 8'h57 == new_ptr_44_value ? ghv_87 : _GEN_7301; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7303 = 8'h58 == new_ptr_44_value ? ghv_88 : _GEN_7302; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7304 = 8'h59 == new_ptr_44_value ? ghv_89 : _GEN_7303; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7305 = 8'h5a == new_ptr_44_value ? ghv_90 : _GEN_7304; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7306 = 8'h5b == new_ptr_44_value ? ghv_91 : _GEN_7305; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7307 = 8'h5c == new_ptr_44_value ? ghv_92 : _GEN_7306; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7308 = 8'h5d == new_ptr_44_value ? ghv_93 : _GEN_7307; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7309 = 8'h5e == new_ptr_44_value ? ghv_94 : _GEN_7308; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7310 = 8'h5f == new_ptr_44_value ? ghv_95 : _GEN_7309; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7311 = 8'h60 == new_ptr_44_value ? ghv_96 : _GEN_7310; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7312 = 8'h61 == new_ptr_44_value ? ghv_97 : _GEN_7311; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7313 = 8'h62 == new_ptr_44_value ? ghv_98 : _GEN_7312; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7314 = 8'h63 == new_ptr_44_value ? ghv_99 : _GEN_7313; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7315 = 8'h64 == new_ptr_44_value ? ghv_100 : _GEN_7314; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7316 = 8'h65 == new_ptr_44_value ? ghv_101 : _GEN_7315; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7317 = 8'h66 == new_ptr_44_value ? ghv_102 : _GEN_7316; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7318 = 8'h67 == new_ptr_44_value ? ghv_103 : _GEN_7317; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7319 = 8'h68 == new_ptr_44_value ? ghv_104 : _GEN_7318; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7320 = 8'h69 == new_ptr_44_value ? ghv_105 : _GEN_7319; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7321 = 8'h6a == new_ptr_44_value ? ghv_106 : _GEN_7320; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7322 = 8'h6b == new_ptr_44_value ? ghv_107 : _GEN_7321; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7323 = 8'h6c == new_ptr_44_value ? ghv_108 : _GEN_7322; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7324 = 8'h6d == new_ptr_44_value ? ghv_109 : _GEN_7323; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7325 = 8'h6e == new_ptr_44_value ? ghv_110 : _GEN_7324; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7326 = 8'h6f == new_ptr_44_value ? ghv_111 : _GEN_7325; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7327 = 8'h70 == new_ptr_44_value ? ghv_112 : _GEN_7326; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7328 = 8'h71 == new_ptr_44_value ? ghv_113 : _GEN_7327; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7329 = 8'h72 == new_ptr_44_value ? ghv_114 : _GEN_7328; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7330 = 8'h73 == new_ptr_44_value ? ghv_115 : _GEN_7329; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7331 = 8'h74 == new_ptr_44_value ? ghv_116 : _GEN_7330; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7332 = 8'h75 == new_ptr_44_value ? ghv_117 : _GEN_7331; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7333 = 8'h76 == new_ptr_44_value ? ghv_118 : _GEN_7332; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7334 = 8'h77 == new_ptr_44_value ? ghv_119 : _GEN_7333; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7335 = 8'h78 == new_ptr_44_value ? ghv_120 : _GEN_7334; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7336 = 8'h79 == new_ptr_44_value ? ghv_121 : _GEN_7335; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7337 = 8'h7a == new_ptr_44_value ? ghv_122 : _GEN_7336; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7338 = 8'h7b == new_ptr_44_value ? ghv_123 : _GEN_7337; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7339 = 8'h7c == new_ptr_44_value ? ghv_124 : _GEN_7338; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7340 = 8'h7d == new_ptr_44_value ? ghv_125 : _GEN_7339; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7341 = 8'h7e == new_ptr_44_value ? ghv_126 : _GEN_7340; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7342 = 8'h7f == new_ptr_44_value ? ghv_127 : _GEN_7341; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7343 = 8'h80 == new_ptr_44_value ? ghv_128 : _GEN_7342; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7344 = 8'h81 == new_ptr_44_value ? ghv_129 : _GEN_7343; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7345 = 8'h82 == new_ptr_44_value ? ghv_130 : _GEN_7344; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7346 = 8'h83 == new_ptr_44_value ? ghv_131 : _GEN_7345; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7347 = 8'h84 == new_ptr_44_value ? ghv_132 : _GEN_7346; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7348 = 8'h85 == new_ptr_44_value ? ghv_133 : _GEN_7347; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7349 = 8'h86 == new_ptr_44_value ? ghv_134 : _GEN_7348; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7350 = 8'h87 == new_ptr_44_value ? ghv_135 : _GEN_7349; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7351 = 8'h88 == new_ptr_44_value ? ghv_136 : _GEN_7350; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7352 = 8'h89 == new_ptr_44_value ? ghv_137 : _GEN_7351; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7353 = 8'h8a == new_ptr_44_value ? ghv_138 : _GEN_7352; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7354 = 8'h8b == new_ptr_44_value ? ghv_139 : _GEN_7353; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7355 = 8'h8c == new_ptr_44_value ? ghv_140 : _GEN_7354; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7356 = 8'h8d == new_ptr_44_value ? ghv_141 : _GEN_7355; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7357 = 8'h8e == new_ptr_44_value ? ghv_142 : _GEN_7356; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_48_value = _new_ptr_value_T_97[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_7360 = 8'h1 == new_ptr_48_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7361 = 8'h2 == new_ptr_48_value ? ghv_2 : _GEN_7360; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7362 = 8'h3 == new_ptr_48_value ? ghv_3 : _GEN_7361; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7363 = 8'h4 == new_ptr_48_value ? ghv_4 : _GEN_7362; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7364 = 8'h5 == new_ptr_48_value ? ghv_5 : _GEN_7363; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7365 = 8'h6 == new_ptr_48_value ? ghv_6 : _GEN_7364; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7366 = 8'h7 == new_ptr_48_value ? ghv_7 : _GEN_7365; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7367 = 8'h8 == new_ptr_48_value ? ghv_8 : _GEN_7366; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7368 = 8'h9 == new_ptr_48_value ? ghv_9 : _GEN_7367; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7369 = 8'ha == new_ptr_48_value ? ghv_10 : _GEN_7368; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7370 = 8'hb == new_ptr_48_value ? ghv_11 : _GEN_7369; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7371 = 8'hc == new_ptr_48_value ? ghv_12 : _GEN_7370; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7372 = 8'hd == new_ptr_48_value ? ghv_13 : _GEN_7371; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7373 = 8'he == new_ptr_48_value ? ghv_14 : _GEN_7372; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7374 = 8'hf == new_ptr_48_value ? ghv_15 : _GEN_7373; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7375 = 8'h10 == new_ptr_48_value ? ghv_16 : _GEN_7374; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7376 = 8'h11 == new_ptr_48_value ? ghv_17 : _GEN_7375; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7377 = 8'h12 == new_ptr_48_value ? ghv_18 : _GEN_7376; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7378 = 8'h13 == new_ptr_48_value ? ghv_19 : _GEN_7377; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7379 = 8'h14 == new_ptr_48_value ? ghv_20 : _GEN_7378; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7380 = 8'h15 == new_ptr_48_value ? ghv_21 : _GEN_7379; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7381 = 8'h16 == new_ptr_48_value ? ghv_22 : _GEN_7380; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7382 = 8'h17 == new_ptr_48_value ? ghv_23 : _GEN_7381; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7383 = 8'h18 == new_ptr_48_value ? ghv_24 : _GEN_7382; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7384 = 8'h19 == new_ptr_48_value ? ghv_25 : _GEN_7383; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7385 = 8'h1a == new_ptr_48_value ? ghv_26 : _GEN_7384; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7386 = 8'h1b == new_ptr_48_value ? ghv_27 : _GEN_7385; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7387 = 8'h1c == new_ptr_48_value ? ghv_28 : _GEN_7386; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7388 = 8'h1d == new_ptr_48_value ? ghv_29 : _GEN_7387; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7389 = 8'h1e == new_ptr_48_value ? ghv_30 : _GEN_7388; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7390 = 8'h1f == new_ptr_48_value ? ghv_31 : _GEN_7389; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7391 = 8'h20 == new_ptr_48_value ? ghv_32 : _GEN_7390; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7392 = 8'h21 == new_ptr_48_value ? ghv_33 : _GEN_7391; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7393 = 8'h22 == new_ptr_48_value ? ghv_34 : _GEN_7392; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7394 = 8'h23 == new_ptr_48_value ? ghv_35 : _GEN_7393; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7395 = 8'h24 == new_ptr_48_value ? ghv_36 : _GEN_7394; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7396 = 8'h25 == new_ptr_48_value ? ghv_37 : _GEN_7395; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7397 = 8'h26 == new_ptr_48_value ? ghv_38 : _GEN_7396; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7398 = 8'h27 == new_ptr_48_value ? ghv_39 : _GEN_7397; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7399 = 8'h28 == new_ptr_48_value ? ghv_40 : _GEN_7398; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7400 = 8'h29 == new_ptr_48_value ? ghv_41 : _GEN_7399; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7401 = 8'h2a == new_ptr_48_value ? ghv_42 : _GEN_7400; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7402 = 8'h2b == new_ptr_48_value ? ghv_43 : _GEN_7401; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7403 = 8'h2c == new_ptr_48_value ? ghv_44 : _GEN_7402; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7404 = 8'h2d == new_ptr_48_value ? ghv_45 : _GEN_7403; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7405 = 8'h2e == new_ptr_48_value ? ghv_46 : _GEN_7404; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7406 = 8'h2f == new_ptr_48_value ? ghv_47 : _GEN_7405; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7407 = 8'h30 == new_ptr_48_value ? ghv_48 : _GEN_7406; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7408 = 8'h31 == new_ptr_48_value ? ghv_49 : _GEN_7407; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7409 = 8'h32 == new_ptr_48_value ? ghv_50 : _GEN_7408; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7410 = 8'h33 == new_ptr_48_value ? ghv_51 : _GEN_7409; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7411 = 8'h34 == new_ptr_48_value ? ghv_52 : _GEN_7410; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7412 = 8'h35 == new_ptr_48_value ? ghv_53 : _GEN_7411; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7413 = 8'h36 == new_ptr_48_value ? ghv_54 : _GEN_7412; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7414 = 8'h37 == new_ptr_48_value ? ghv_55 : _GEN_7413; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7415 = 8'h38 == new_ptr_48_value ? ghv_56 : _GEN_7414; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7416 = 8'h39 == new_ptr_48_value ? ghv_57 : _GEN_7415; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7417 = 8'h3a == new_ptr_48_value ? ghv_58 : _GEN_7416; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7418 = 8'h3b == new_ptr_48_value ? ghv_59 : _GEN_7417; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7419 = 8'h3c == new_ptr_48_value ? ghv_60 : _GEN_7418; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7420 = 8'h3d == new_ptr_48_value ? ghv_61 : _GEN_7419; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7421 = 8'h3e == new_ptr_48_value ? ghv_62 : _GEN_7420; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7422 = 8'h3f == new_ptr_48_value ? ghv_63 : _GEN_7421; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7423 = 8'h40 == new_ptr_48_value ? ghv_64 : _GEN_7422; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7424 = 8'h41 == new_ptr_48_value ? ghv_65 : _GEN_7423; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7425 = 8'h42 == new_ptr_48_value ? ghv_66 : _GEN_7424; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7426 = 8'h43 == new_ptr_48_value ? ghv_67 : _GEN_7425; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7427 = 8'h44 == new_ptr_48_value ? ghv_68 : _GEN_7426; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7428 = 8'h45 == new_ptr_48_value ? ghv_69 : _GEN_7427; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7429 = 8'h46 == new_ptr_48_value ? ghv_70 : _GEN_7428; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7430 = 8'h47 == new_ptr_48_value ? ghv_71 : _GEN_7429; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7431 = 8'h48 == new_ptr_48_value ? ghv_72 : _GEN_7430; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7432 = 8'h49 == new_ptr_48_value ? ghv_73 : _GEN_7431; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7433 = 8'h4a == new_ptr_48_value ? ghv_74 : _GEN_7432; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7434 = 8'h4b == new_ptr_48_value ? ghv_75 : _GEN_7433; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7435 = 8'h4c == new_ptr_48_value ? ghv_76 : _GEN_7434; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7436 = 8'h4d == new_ptr_48_value ? ghv_77 : _GEN_7435; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7437 = 8'h4e == new_ptr_48_value ? ghv_78 : _GEN_7436; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7438 = 8'h4f == new_ptr_48_value ? ghv_79 : _GEN_7437; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7439 = 8'h50 == new_ptr_48_value ? ghv_80 : _GEN_7438; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7440 = 8'h51 == new_ptr_48_value ? ghv_81 : _GEN_7439; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7441 = 8'h52 == new_ptr_48_value ? ghv_82 : _GEN_7440; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7442 = 8'h53 == new_ptr_48_value ? ghv_83 : _GEN_7441; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7443 = 8'h54 == new_ptr_48_value ? ghv_84 : _GEN_7442; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7444 = 8'h55 == new_ptr_48_value ? ghv_85 : _GEN_7443; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7445 = 8'h56 == new_ptr_48_value ? ghv_86 : _GEN_7444; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7446 = 8'h57 == new_ptr_48_value ? ghv_87 : _GEN_7445; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7447 = 8'h58 == new_ptr_48_value ? ghv_88 : _GEN_7446; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7448 = 8'h59 == new_ptr_48_value ? ghv_89 : _GEN_7447; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7449 = 8'h5a == new_ptr_48_value ? ghv_90 : _GEN_7448; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7450 = 8'h5b == new_ptr_48_value ? ghv_91 : _GEN_7449; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7451 = 8'h5c == new_ptr_48_value ? ghv_92 : _GEN_7450; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7452 = 8'h5d == new_ptr_48_value ? ghv_93 : _GEN_7451; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7453 = 8'h5e == new_ptr_48_value ? ghv_94 : _GEN_7452; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7454 = 8'h5f == new_ptr_48_value ? ghv_95 : _GEN_7453; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7455 = 8'h60 == new_ptr_48_value ? ghv_96 : _GEN_7454; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7456 = 8'h61 == new_ptr_48_value ? ghv_97 : _GEN_7455; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7457 = 8'h62 == new_ptr_48_value ? ghv_98 : _GEN_7456; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7458 = 8'h63 == new_ptr_48_value ? ghv_99 : _GEN_7457; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7459 = 8'h64 == new_ptr_48_value ? ghv_100 : _GEN_7458; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7460 = 8'h65 == new_ptr_48_value ? ghv_101 : _GEN_7459; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7461 = 8'h66 == new_ptr_48_value ? ghv_102 : _GEN_7460; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7462 = 8'h67 == new_ptr_48_value ? ghv_103 : _GEN_7461; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7463 = 8'h68 == new_ptr_48_value ? ghv_104 : _GEN_7462; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7464 = 8'h69 == new_ptr_48_value ? ghv_105 : _GEN_7463; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7465 = 8'h6a == new_ptr_48_value ? ghv_106 : _GEN_7464; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7466 = 8'h6b == new_ptr_48_value ? ghv_107 : _GEN_7465; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7467 = 8'h6c == new_ptr_48_value ? ghv_108 : _GEN_7466; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7468 = 8'h6d == new_ptr_48_value ? ghv_109 : _GEN_7467; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7469 = 8'h6e == new_ptr_48_value ? ghv_110 : _GEN_7468; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7470 = 8'h6f == new_ptr_48_value ? ghv_111 : _GEN_7469; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7471 = 8'h70 == new_ptr_48_value ? ghv_112 : _GEN_7470; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7472 = 8'h71 == new_ptr_48_value ? ghv_113 : _GEN_7471; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7473 = 8'h72 == new_ptr_48_value ? ghv_114 : _GEN_7472; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7474 = 8'h73 == new_ptr_48_value ? ghv_115 : _GEN_7473; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7475 = 8'h74 == new_ptr_48_value ? ghv_116 : _GEN_7474; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7476 = 8'h75 == new_ptr_48_value ? ghv_117 : _GEN_7475; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7477 = 8'h76 == new_ptr_48_value ? ghv_118 : _GEN_7476; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7478 = 8'h77 == new_ptr_48_value ? ghv_119 : _GEN_7477; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7479 = 8'h78 == new_ptr_48_value ? ghv_120 : _GEN_7478; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7480 = 8'h79 == new_ptr_48_value ? ghv_121 : _GEN_7479; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7481 = 8'h7a == new_ptr_48_value ? ghv_122 : _GEN_7480; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7482 = 8'h7b == new_ptr_48_value ? ghv_123 : _GEN_7481; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7483 = 8'h7c == new_ptr_48_value ? ghv_124 : _GEN_7482; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7484 = 8'h7d == new_ptr_48_value ? ghv_125 : _GEN_7483; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7485 = 8'h7e == new_ptr_48_value ? ghv_126 : _GEN_7484; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7486 = 8'h7f == new_ptr_48_value ? ghv_127 : _GEN_7485; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7487 = 8'h80 == new_ptr_48_value ? ghv_128 : _GEN_7486; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7488 = 8'h81 == new_ptr_48_value ? ghv_129 : _GEN_7487; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7489 = 8'h82 == new_ptr_48_value ? ghv_130 : _GEN_7488; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7490 = 8'h83 == new_ptr_48_value ? ghv_131 : _GEN_7489; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7491 = 8'h84 == new_ptr_48_value ? ghv_132 : _GEN_7490; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7492 = 8'h85 == new_ptr_48_value ? ghv_133 : _GEN_7491; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7493 = 8'h86 == new_ptr_48_value ? ghv_134 : _GEN_7492; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7494 = 8'h87 == new_ptr_48_value ? ghv_135 : _GEN_7493; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7495 = 8'h88 == new_ptr_48_value ? ghv_136 : _GEN_7494; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7496 = 8'h89 == new_ptr_48_value ? ghv_137 : _GEN_7495; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7497 = 8'h8a == new_ptr_48_value ? ghv_138 : _GEN_7496; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7498 = 8'h8b == new_ptr_48_value ? ghv_139 : _GEN_7497; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7499 = 8'h8c == new_ptr_48_value ? ghv_140 : _GEN_7498; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7500 = 8'h8d == new_ptr_48_value ? ghv_141 : _GEN_7499; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7501 = 8'h8e == new_ptr_48_value ? ghv_142 : _GEN_7500; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_59_value = _new_ptr_value_T_119[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_7504 = 8'h1 == new_ptr_59_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7505 = 8'h2 == new_ptr_59_value ? ghv_2 : _GEN_7504; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7506 = 8'h3 == new_ptr_59_value ? ghv_3 : _GEN_7505; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7507 = 8'h4 == new_ptr_59_value ? ghv_4 : _GEN_7506; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7508 = 8'h5 == new_ptr_59_value ? ghv_5 : _GEN_7507; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7509 = 8'h6 == new_ptr_59_value ? ghv_6 : _GEN_7508; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7510 = 8'h7 == new_ptr_59_value ? ghv_7 : _GEN_7509; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7511 = 8'h8 == new_ptr_59_value ? ghv_8 : _GEN_7510; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7512 = 8'h9 == new_ptr_59_value ? ghv_9 : _GEN_7511; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7513 = 8'ha == new_ptr_59_value ? ghv_10 : _GEN_7512; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7514 = 8'hb == new_ptr_59_value ? ghv_11 : _GEN_7513; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7515 = 8'hc == new_ptr_59_value ? ghv_12 : _GEN_7514; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7516 = 8'hd == new_ptr_59_value ? ghv_13 : _GEN_7515; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7517 = 8'he == new_ptr_59_value ? ghv_14 : _GEN_7516; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7518 = 8'hf == new_ptr_59_value ? ghv_15 : _GEN_7517; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7519 = 8'h10 == new_ptr_59_value ? ghv_16 : _GEN_7518; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7520 = 8'h11 == new_ptr_59_value ? ghv_17 : _GEN_7519; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7521 = 8'h12 == new_ptr_59_value ? ghv_18 : _GEN_7520; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7522 = 8'h13 == new_ptr_59_value ? ghv_19 : _GEN_7521; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7523 = 8'h14 == new_ptr_59_value ? ghv_20 : _GEN_7522; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7524 = 8'h15 == new_ptr_59_value ? ghv_21 : _GEN_7523; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7525 = 8'h16 == new_ptr_59_value ? ghv_22 : _GEN_7524; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7526 = 8'h17 == new_ptr_59_value ? ghv_23 : _GEN_7525; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7527 = 8'h18 == new_ptr_59_value ? ghv_24 : _GEN_7526; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7528 = 8'h19 == new_ptr_59_value ? ghv_25 : _GEN_7527; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7529 = 8'h1a == new_ptr_59_value ? ghv_26 : _GEN_7528; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7530 = 8'h1b == new_ptr_59_value ? ghv_27 : _GEN_7529; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7531 = 8'h1c == new_ptr_59_value ? ghv_28 : _GEN_7530; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7532 = 8'h1d == new_ptr_59_value ? ghv_29 : _GEN_7531; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7533 = 8'h1e == new_ptr_59_value ? ghv_30 : _GEN_7532; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7534 = 8'h1f == new_ptr_59_value ? ghv_31 : _GEN_7533; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7535 = 8'h20 == new_ptr_59_value ? ghv_32 : _GEN_7534; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7536 = 8'h21 == new_ptr_59_value ? ghv_33 : _GEN_7535; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7537 = 8'h22 == new_ptr_59_value ? ghv_34 : _GEN_7536; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7538 = 8'h23 == new_ptr_59_value ? ghv_35 : _GEN_7537; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7539 = 8'h24 == new_ptr_59_value ? ghv_36 : _GEN_7538; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7540 = 8'h25 == new_ptr_59_value ? ghv_37 : _GEN_7539; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7541 = 8'h26 == new_ptr_59_value ? ghv_38 : _GEN_7540; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7542 = 8'h27 == new_ptr_59_value ? ghv_39 : _GEN_7541; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7543 = 8'h28 == new_ptr_59_value ? ghv_40 : _GEN_7542; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7544 = 8'h29 == new_ptr_59_value ? ghv_41 : _GEN_7543; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7545 = 8'h2a == new_ptr_59_value ? ghv_42 : _GEN_7544; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7546 = 8'h2b == new_ptr_59_value ? ghv_43 : _GEN_7545; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7547 = 8'h2c == new_ptr_59_value ? ghv_44 : _GEN_7546; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7548 = 8'h2d == new_ptr_59_value ? ghv_45 : _GEN_7547; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7549 = 8'h2e == new_ptr_59_value ? ghv_46 : _GEN_7548; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7550 = 8'h2f == new_ptr_59_value ? ghv_47 : _GEN_7549; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7551 = 8'h30 == new_ptr_59_value ? ghv_48 : _GEN_7550; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7552 = 8'h31 == new_ptr_59_value ? ghv_49 : _GEN_7551; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7553 = 8'h32 == new_ptr_59_value ? ghv_50 : _GEN_7552; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7554 = 8'h33 == new_ptr_59_value ? ghv_51 : _GEN_7553; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7555 = 8'h34 == new_ptr_59_value ? ghv_52 : _GEN_7554; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7556 = 8'h35 == new_ptr_59_value ? ghv_53 : _GEN_7555; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7557 = 8'h36 == new_ptr_59_value ? ghv_54 : _GEN_7556; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7558 = 8'h37 == new_ptr_59_value ? ghv_55 : _GEN_7557; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7559 = 8'h38 == new_ptr_59_value ? ghv_56 : _GEN_7558; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7560 = 8'h39 == new_ptr_59_value ? ghv_57 : _GEN_7559; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7561 = 8'h3a == new_ptr_59_value ? ghv_58 : _GEN_7560; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7562 = 8'h3b == new_ptr_59_value ? ghv_59 : _GEN_7561; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7563 = 8'h3c == new_ptr_59_value ? ghv_60 : _GEN_7562; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7564 = 8'h3d == new_ptr_59_value ? ghv_61 : _GEN_7563; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7565 = 8'h3e == new_ptr_59_value ? ghv_62 : _GEN_7564; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7566 = 8'h3f == new_ptr_59_value ? ghv_63 : _GEN_7565; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7567 = 8'h40 == new_ptr_59_value ? ghv_64 : _GEN_7566; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7568 = 8'h41 == new_ptr_59_value ? ghv_65 : _GEN_7567; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7569 = 8'h42 == new_ptr_59_value ? ghv_66 : _GEN_7568; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7570 = 8'h43 == new_ptr_59_value ? ghv_67 : _GEN_7569; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7571 = 8'h44 == new_ptr_59_value ? ghv_68 : _GEN_7570; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7572 = 8'h45 == new_ptr_59_value ? ghv_69 : _GEN_7571; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7573 = 8'h46 == new_ptr_59_value ? ghv_70 : _GEN_7572; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7574 = 8'h47 == new_ptr_59_value ? ghv_71 : _GEN_7573; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7575 = 8'h48 == new_ptr_59_value ? ghv_72 : _GEN_7574; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7576 = 8'h49 == new_ptr_59_value ? ghv_73 : _GEN_7575; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7577 = 8'h4a == new_ptr_59_value ? ghv_74 : _GEN_7576; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7578 = 8'h4b == new_ptr_59_value ? ghv_75 : _GEN_7577; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7579 = 8'h4c == new_ptr_59_value ? ghv_76 : _GEN_7578; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7580 = 8'h4d == new_ptr_59_value ? ghv_77 : _GEN_7579; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7581 = 8'h4e == new_ptr_59_value ? ghv_78 : _GEN_7580; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7582 = 8'h4f == new_ptr_59_value ? ghv_79 : _GEN_7581; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7583 = 8'h50 == new_ptr_59_value ? ghv_80 : _GEN_7582; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7584 = 8'h51 == new_ptr_59_value ? ghv_81 : _GEN_7583; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7585 = 8'h52 == new_ptr_59_value ? ghv_82 : _GEN_7584; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7586 = 8'h53 == new_ptr_59_value ? ghv_83 : _GEN_7585; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7587 = 8'h54 == new_ptr_59_value ? ghv_84 : _GEN_7586; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7588 = 8'h55 == new_ptr_59_value ? ghv_85 : _GEN_7587; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7589 = 8'h56 == new_ptr_59_value ? ghv_86 : _GEN_7588; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7590 = 8'h57 == new_ptr_59_value ? ghv_87 : _GEN_7589; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7591 = 8'h58 == new_ptr_59_value ? ghv_88 : _GEN_7590; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7592 = 8'h59 == new_ptr_59_value ? ghv_89 : _GEN_7591; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7593 = 8'h5a == new_ptr_59_value ? ghv_90 : _GEN_7592; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7594 = 8'h5b == new_ptr_59_value ? ghv_91 : _GEN_7593; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7595 = 8'h5c == new_ptr_59_value ? ghv_92 : _GEN_7594; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7596 = 8'h5d == new_ptr_59_value ? ghv_93 : _GEN_7595; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7597 = 8'h5e == new_ptr_59_value ? ghv_94 : _GEN_7596; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7598 = 8'h5f == new_ptr_59_value ? ghv_95 : _GEN_7597; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7599 = 8'h60 == new_ptr_59_value ? ghv_96 : _GEN_7598; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7600 = 8'h61 == new_ptr_59_value ? ghv_97 : _GEN_7599; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7601 = 8'h62 == new_ptr_59_value ? ghv_98 : _GEN_7600; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7602 = 8'h63 == new_ptr_59_value ? ghv_99 : _GEN_7601; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7603 = 8'h64 == new_ptr_59_value ? ghv_100 : _GEN_7602; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7604 = 8'h65 == new_ptr_59_value ? ghv_101 : _GEN_7603; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7605 = 8'h66 == new_ptr_59_value ? ghv_102 : _GEN_7604; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7606 = 8'h67 == new_ptr_59_value ? ghv_103 : _GEN_7605; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7607 = 8'h68 == new_ptr_59_value ? ghv_104 : _GEN_7606; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7608 = 8'h69 == new_ptr_59_value ? ghv_105 : _GEN_7607; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7609 = 8'h6a == new_ptr_59_value ? ghv_106 : _GEN_7608; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7610 = 8'h6b == new_ptr_59_value ? ghv_107 : _GEN_7609; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7611 = 8'h6c == new_ptr_59_value ? ghv_108 : _GEN_7610; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7612 = 8'h6d == new_ptr_59_value ? ghv_109 : _GEN_7611; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7613 = 8'h6e == new_ptr_59_value ? ghv_110 : _GEN_7612; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7614 = 8'h6f == new_ptr_59_value ? ghv_111 : _GEN_7613; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7615 = 8'h70 == new_ptr_59_value ? ghv_112 : _GEN_7614; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7616 = 8'h71 == new_ptr_59_value ? ghv_113 : _GEN_7615; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7617 = 8'h72 == new_ptr_59_value ? ghv_114 : _GEN_7616; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7618 = 8'h73 == new_ptr_59_value ? ghv_115 : _GEN_7617; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7619 = 8'h74 == new_ptr_59_value ? ghv_116 : _GEN_7618; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7620 = 8'h75 == new_ptr_59_value ? ghv_117 : _GEN_7619; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7621 = 8'h76 == new_ptr_59_value ? ghv_118 : _GEN_7620; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7622 = 8'h77 == new_ptr_59_value ? ghv_119 : _GEN_7621; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7623 = 8'h78 == new_ptr_59_value ? ghv_120 : _GEN_7622; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7624 = 8'h79 == new_ptr_59_value ? ghv_121 : _GEN_7623; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7625 = 8'h7a == new_ptr_59_value ? ghv_122 : _GEN_7624; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7626 = 8'h7b == new_ptr_59_value ? ghv_123 : _GEN_7625; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7627 = 8'h7c == new_ptr_59_value ? ghv_124 : _GEN_7626; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7628 = 8'h7d == new_ptr_59_value ? ghv_125 : _GEN_7627; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7629 = 8'h7e == new_ptr_59_value ? ghv_126 : _GEN_7628; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7630 = 8'h7f == new_ptr_59_value ? ghv_127 : _GEN_7629; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7631 = 8'h80 == new_ptr_59_value ? ghv_128 : _GEN_7630; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7632 = 8'h81 == new_ptr_59_value ? ghv_129 : _GEN_7631; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7633 = 8'h82 == new_ptr_59_value ? ghv_130 : _GEN_7632; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7634 = 8'h83 == new_ptr_59_value ? ghv_131 : _GEN_7633; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7635 = 8'h84 == new_ptr_59_value ? ghv_132 : _GEN_7634; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7636 = 8'h85 == new_ptr_59_value ? ghv_133 : _GEN_7635; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7637 = 8'h86 == new_ptr_59_value ? ghv_134 : _GEN_7636; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7638 = 8'h87 == new_ptr_59_value ? ghv_135 : _GEN_7637; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7639 = 8'h88 == new_ptr_59_value ? ghv_136 : _GEN_7638; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7640 = 8'h89 == new_ptr_59_value ? ghv_137 : _GEN_7639; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7641 = 8'h8a == new_ptr_59_value ? ghv_138 : _GEN_7640; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7642 = 8'h8b == new_ptr_59_value ? ghv_139 : _GEN_7641; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7643 = 8'h8c == new_ptr_59_value ? ghv_140 : _GEN_7642; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7644 = 8'h8d == new_ptr_59_value ? ghv_141 : _GEN_7643; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7645 = 8'h8e == new_ptr_59_value ? ghv_142 : _GEN_7644; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_43_value = _new_ptr_value_T_87[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_7648 = 8'h1 == new_ptr_43_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7649 = 8'h2 == new_ptr_43_value ? ghv_2 : _GEN_7648; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7650 = 8'h3 == new_ptr_43_value ? ghv_3 : _GEN_7649; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7651 = 8'h4 == new_ptr_43_value ? ghv_4 : _GEN_7650; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7652 = 8'h5 == new_ptr_43_value ? ghv_5 : _GEN_7651; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7653 = 8'h6 == new_ptr_43_value ? ghv_6 : _GEN_7652; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7654 = 8'h7 == new_ptr_43_value ? ghv_7 : _GEN_7653; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7655 = 8'h8 == new_ptr_43_value ? ghv_8 : _GEN_7654; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7656 = 8'h9 == new_ptr_43_value ? ghv_9 : _GEN_7655; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7657 = 8'ha == new_ptr_43_value ? ghv_10 : _GEN_7656; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7658 = 8'hb == new_ptr_43_value ? ghv_11 : _GEN_7657; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7659 = 8'hc == new_ptr_43_value ? ghv_12 : _GEN_7658; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7660 = 8'hd == new_ptr_43_value ? ghv_13 : _GEN_7659; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7661 = 8'he == new_ptr_43_value ? ghv_14 : _GEN_7660; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7662 = 8'hf == new_ptr_43_value ? ghv_15 : _GEN_7661; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7663 = 8'h10 == new_ptr_43_value ? ghv_16 : _GEN_7662; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7664 = 8'h11 == new_ptr_43_value ? ghv_17 : _GEN_7663; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7665 = 8'h12 == new_ptr_43_value ? ghv_18 : _GEN_7664; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7666 = 8'h13 == new_ptr_43_value ? ghv_19 : _GEN_7665; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7667 = 8'h14 == new_ptr_43_value ? ghv_20 : _GEN_7666; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7668 = 8'h15 == new_ptr_43_value ? ghv_21 : _GEN_7667; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7669 = 8'h16 == new_ptr_43_value ? ghv_22 : _GEN_7668; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7670 = 8'h17 == new_ptr_43_value ? ghv_23 : _GEN_7669; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7671 = 8'h18 == new_ptr_43_value ? ghv_24 : _GEN_7670; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7672 = 8'h19 == new_ptr_43_value ? ghv_25 : _GEN_7671; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7673 = 8'h1a == new_ptr_43_value ? ghv_26 : _GEN_7672; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7674 = 8'h1b == new_ptr_43_value ? ghv_27 : _GEN_7673; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7675 = 8'h1c == new_ptr_43_value ? ghv_28 : _GEN_7674; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7676 = 8'h1d == new_ptr_43_value ? ghv_29 : _GEN_7675; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7677 = 8'h1e == new_ptr_43_value ? ghv_30 : _GEN_7676; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7678 = 8'h1f == new_ptr_43_value ? ghv_31 : _GEN_7677; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7679 = 8'h20 == new_ptr_43_value ? ghv_32 : _GEN_7678; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7680 = 8'h21 == new_ptr_43_value ? ghv_33 : _GEN_7679; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7681 = 8'h22 == new_ptr_43_value ? ghv_34 : _GEN_7680; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7682 = 8'h23 == new_ptr_43_value ? ghv_35 : _GEN_7681; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7683 = 8'h24 == new_ptr_43_value ? ghv_36 : _GEN_7682; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7684 = 8'h25 == new_ptr_43_value ? ghv_37 : _GEN_7683; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7685 = 8'h26 == new_ptr_43_value ? ghv_38 : _GEN_7684; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7686 = 8'h27 == new_ptr_43_value ? ghv_39 : _GEN_7685; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7687 = 8'h28 == new_ptr_43_value ? ghv_40 : _GEN_7686; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7688 = 8'h29 == new_ptr_43_value ? ghv_41 : _GEN_7687; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7689 = 8'h2a == new_ptr_43_value ? ghv_42 : _GEN_7688; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7690 = 8'h2b == new_ptr_43_value ? ghv_43 : _GEN_7689; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7691 = 8'h2c == new_ptr_43_value ? ghv_44 : _GEN_7690; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7692 = 8'h2d == new_ptr_43_value ? ghv_45 : _GEN_7691; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7693 = 8'h2e == new_ptr_43_value ? ghv_46 : _GEN_7692; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7694 = 8'h2f == new_ptr_43_value ? ghv_47 : _GEN_7693; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7695 = 8'h30 == new_ptr_43_value ? ghv_48 : _GEN_7694; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7696 = 8'h31 == new_ptr_43_value ? ghv_49 : _GEN_7695; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7697 = 8'h32 == new_ptr_43_value ? ghv_50 : _GEN_7696; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7698 = 8'h33 == new_ptr_43_value ? ghv_51 : _GEN_7697; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7699 = 8'h34 == new_ptr_43_value ? ghv_52 : _GEN_7698; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7700 = 8'h35 == new_ptr_43_value ? ghv_53 : _GEN_7699; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7701 = 8'h36 == new_ptr_43_value ? ghv_54 : _GEN_7700; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7702 = 8'h37 == new_ptr_43_value ? ghv_55 : _GEN_7701; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7703 = 8'h38 == new_ptr_43_value ? ghv_56 : _GEN_7702; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7704 = 8'h39 == new_ptr_43_value ? ghv_57 : _GEN_7703; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7705 = 8'h3a == new_ptr_43_value ? ghv_58 : _GEN_7704; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7706 = 8'h3b == new_ptr_43_value ? ghv_59 : _GEN_7705; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7707 = 8'h3c == new_ptr_43_value ? ghv_60 : _GEN_7706; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7708 = 8'h3d == new_ptr_43_value ? ghv_61 : _GEN_7707; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7709 = 8'h3e == new_ptr_43_value ? ghv_62 : _GEN_7708; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7710 = 8'h3f == new_ptr_43_value ? ghv_63 : _GEN_7709; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7711 = 8'h40 == new_ptr_43_value ? ghv_64 : _GEN_7710; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7712 = 8'h41 == new_ptr_43_value ? ghv_65 : _GEN_7711; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7713 = 8'h42 == new_ptr_43_value ? ghv_66 : _GEN_7712; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7714 = 8'h43 == new_ptr_43_value ? ghv_67 : _GEN_7713; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7715 = 8'h44 == new_ptr_43_value ? ghv_68 : _GEN_7714; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7716 = 8'h45 == new_ptr_43_value ? ghv_69 : _GEN_7715; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7717 = 8'h46 == new_ptr_43_value ? ghv_70 : _GEN_7716; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7718 = 8'h47 == new_ptr_43_value ? ghv_71 : _GEN_7717; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7719 = 8'h48 == new_ptr_43_value ? ghv_72 : _GEN_7718; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7720 = 8'h49 == new_ptr_43_value ? ghv_73 : _GEN_7719; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7721 = 8'h4a == new_ptr_43_value ? ghv_74 : _GEN_7720; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7722 = 8'h4b == new_ptr_43_value ? ghv_75 : _GEN_7721; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7723 = 8'h4c == new_ptr_43_value ? ghv_76 : _GEN_7722; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7724 = 8'h4d == new_ptr_43_value ? ghv_77 : _GEN_7723; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7725 = 8'h4e == new_ptr_43_value ? ghv_78 : _GEN_7724; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7726 = 8'h4f == new_ptr_43_value ? ghv_79 : _GEN_7725; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7727 = 8'h50 == new_ptr_43_value ? ghv_80 : _GEN_7726; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7728 = 8'h51 == new_ptr_43_value ? ghv_81 : _GEN_7727; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7729 = 8'h52 == new_ptr_43_value ? ghv_82 : _GEN_7728; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7730 = 8'h53 == new_ptr_43_value ? ghv_83 : _GEN_7729; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7731 = 8'h54 == new_ptr_43_value ? ghv_84 : _GEN_7730; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7732 = 8'h55 == new_ptr_43_value ? ghv_85 : _GEN_7731; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7733 = 8'h56 == new_ptr_43_value ? ghv_86 : _GEN_7732; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7734 = 8'h57 == new_ptr_43_value ? ghv_87 : _GEN_7733; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7735 = 8'h58 == new_ptr_43_value ? ghv_88 : _GEN_7734; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7736 = 8'h59 == new_ptr_43_value ? ghv_89 : _GEN_7735; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7737 = 8'h5a == new_ptr_43_value ? ghv_90 : _GEN_7736; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7738 = 8'h5b == new_ptr_43_value ? ghv_91 : _GEN_7737; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7739 = 8'h5c == new_ptr_43_value ? ghv_92 : _GEN_7738; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7740 = 8'h5d == new_ptr_43_value ? ghv_93 : _GEN_7739; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7741 = 8'h5e == new_ptr_43_value ? ghv_94 : _GEN_7740; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7742 = 8'h5f == new_ptr_43_value ? ghv_95 : _GEN_7741; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7743 = 8'h60 == new_ptr_43_value ? ghv_96 : _GEN_7742; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7744 = 8'h61 == new_ptr_43_value ? ghv_97 : _GEN_7743; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7745 = 8'h62 == new_ptr_43_value ? ghv_98 : _GEN_7744; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7746 = 8'h63 == new_ptr_43_value ? ghv_99 : _GEN_7745; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7747 = 8'h64 == new_ptr_43_value ? ghv_100 : _GEN_7746; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7748 = 8'h65 == new_ptr_43_value ? ghv_101 : _GEN_7747; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7749 = 8'h66 == new_ptr_43_value ? ghv_102 : _GEN_7748; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7750 = 8'h67 == new_ptr_43_value ? ghv_103 : _GEN_7749; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7751 = 8'h68 == new_ptr_43_value ? ghv_104 : _GEN_7750; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7752 = 8'h69 == new_ptr_43_value ? ghv_105 : _GEN_7751; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7753 = 8'h6a == new_ptr_43_value ? ghv_106 : _GEN_7752; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7754 = 8'h6b == new_ptr_43_value ? ghv_107 : _GEN_7753; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7755 = 8'h6c == new_ptr_43_value ? ghv_108 : _GEN_7754; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7756 = 8'h6d == new_ptr_43_value ? ghv_109 : _GEN_7755; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7757 = 8'h6e == new_ptr_43_value ? ghv_110 : _GEN_7756; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7758 = 8'h6f == new_ptr_43_value ? ghv_111 : _GEN_7757; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7759 = 8'h70 == new_ptr_43_value ? ghv_112 : _GEN_7758; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7760 = 8'h71 == new_ptr_43_value ? ghv_113 : _GEN_7759; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7761 = 8'h72 == new_ptr_43_value ? ghv_114 : _GEN_7760; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7762 = 8'h73 == new_ptr_43_value ? ghv_115 : _GEN_7761; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7763 = 8'h74 == new_ptr_43_value ? ghv_116 : _GEN_7762; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7764 = 8'h75 == new_ptr_43_value ? ghv_117 : _GEN_7763; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7765 = 8'h76 == new_ptr_43_value ? ghv_118 : _GEN_7764; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7766 = 8'h77 == new_ptr_43_value ? ghv_119 : _GEN_7765; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7767 = 8'h78 == new_ptr_43_value ? ghv_120 : _GEN_7766; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7768 = 8'h79 == new_ptr_43_value ? ghv_121 : _GEN_7767; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7769 = 8'h7a == new_ptr_43_value ? ghv_122 : _GEN_7768; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7770 = 8'h7b == new_ptr_43_value ? ghv_123 : _GEN_7769; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7771 = 8'h7c == new_ptr_43_value ? ghv_124 : _GEN_7770; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7772 = 8'h7d == new_ptr_43_value ? ghv_125 : _GEN_7771; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7773 = 8'h7e == new_ptr_43_value ? ghv_126 : _GEN_7772; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7774 = 8'h7f == new_ptr_43_value ? ghv_127 : _GEN_7773; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7775 = 8'h80 == new_ptr_43_value ? ghv_128 : _GEN_7774; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7776 = 8'h81 == new_ptr_43_value ? ghv_129 : _GEN_7775; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7777 = 8'h82 == new_ptr_43_value ? ghv_130 : _GEN_7776; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7778 = 8'h83 == new_ptr_43_value ? ghv_131 : _GEN_7777; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7779 = 8'h84 == new_ptr_43_value ? ghv_132 : _GEN_7778; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7780 = 8'h85 == new_ptr_43_value ? ghv_133 : _GEN_7779; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7781 = 8'h86 == new_ptr_43_value ? ghv_134 : _GEN_7780; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7782 = 8'h87 == new_ptr_43_value ? ghv_135 : _GEN_7781; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7783 = 8'h88 == new_ptr_43_value ? ghv_136 : _GEN_7782; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7784 = 8'h89 == new_ptr_43_value ? ghv_137 : _GEN_7783; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7785 = 8'h8a == new_ptr_43_value ? ghv_138 : _GEN_7784; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7786 = 8'h8b == new_ptr_43_value ? ghv_139 : _GEN_7785; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7787 = 8'h8c == new_ptr_43_value ? ghv_140 : _GEN_7786; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7788 = 8'h8d == new_ptr_43_value ? ghv_141 : _GEN_7787; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7789 = 8'h8e == new_ptr_43_value ? ghv_142 : _GEN_7788; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_50_value = _new_ptr_value_T_101[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_7792 = 8'h1 == new_ptr_50_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7793 = 8'h2 == new_ptr_50_value ? ghv_2 : _GEN_7792; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7794 = 8'h3 == new_ptr_50_value ? ghv_3 : _GEN_7793; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7795 = 8'h4 == new_ptr_50_value ? ghv_4 : _GEN_7794; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7796 = 8'h5 == new_ptr_50_value ? ghv_5 : _GEN_7795; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7797 = 8'h6 == new_ptr_50_value ? ghv_6 : _GEN_7796; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7798 = 8'h7 == new_ptr_50_value ? ghv_7 : _GEN_7797; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7799 = 8'h8 == new_ptr_50_value ? ghv_8 : _GEN_7798; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7800 = 8'h9 == new_ptr_50_value ? ghv_9 : _GEN_7799; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7801 = 8'ha == new_ptr_50_value ? ghv_10 : _GEN_7800; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7802 = 8'hb == new_ptr_50_value ? ghv_11 : _GEN_7801; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7803 = 8'hc == new_ptr_50_value ? ghv_12 : _GEN_7802; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7804 = 8'hd == new_ptr_50_value ? ghv_13 : _GEN_7803; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7805 = 8'he == new_ptr_50_value ? ghv_14 : _GEN_7804; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7806 = 8'hf == new_ptr_50_value ? ghv_15 : _GEN_7805; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7807 = 8'h10 == new_ptr_50_value ? ghv_16 : _GEN_7806; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7808 = 8'h11 == new_ptr_50_value ? ghv_17 : _GEN_7807; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7809 = 8'h12 == new_ptr_50_value ? ghv_18 : _GEN_7808; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7810 = 8'h13 == new_ptr_50_value ? ghv_19 : _GEN_7809; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7811 = 8'h14 == new_ptr_50_value ? ghv_20 : _GEN_7810; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7812 = 8'h15 == new_ptr_50_value ? ghv_21 : _GEN_7811; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7813 = 8'h16 == new_ptr_50_value ? ghv_22 : _GEN_7812; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7814 = 8'h17 == new_ptr_50_value ? ghv_23 : _GEN_7813; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7815 = 8'h18 == new_ptr_50_value ? ghv_24 : _GEN_7814; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7816 = 8'h19 == new_ptr_50_value ? ghv_25 : _GEN_7815; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7817 = 8'h1a == new_ptr_50_value ? ghv_26 : _GEN_7816; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7818 = 8'h1b == new_ptr_50_value ? ghv_27 : _GEN_7817; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7819 = 8'h1c == new_ptr_50_value ? ghv_28 : _GEN_7818; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7820 = 8'h1d == new_ptr_50_value ? ghv_29 : _GEN_7819; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7821 = 8'h1e == new_ptr_50_value ? ghv_30 : _GEN_7820; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7822 = 8'h1f == new_ptr_50_value ? ghv_31 : _GEN_7821; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7823 = 8'h20 == new_ptr_50_value ? ghv_32 : _GEN_7822; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7824 = 8'h21 == new_ptr_50_value ? ghv_33 : _GEN_7823; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7825 = 8'h22 == new_ptr_50_value ? ghv_34 : _GEN_7824; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7826 = 8'h23 == new_ptr_50_value ? ghv_35 : _GEN_7825; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7827 = 8'h24 == new_ptr_50_value ? ghv_36 : _GEN_7826; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7828 = 8'h25 == new_ptr_50_value ? ghv_37 : _GEN_7827; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7829 = 8'h26 == new_ptr_50_value ? ghv_38 : _GEN_7828; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7830 = 8'h27 == new_ptr_50_value ? ghv_39 : _GEN_7829; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7831 = 8'h28 == new_ptr_50_value ? ghv_40 : _GEN_7830; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7832 = 8'h29 == new_ptr_50_value ? ghv_41 : _GEN_7831; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7833 = 8'h2a == new_ptr_50_value ? ghv_42 : _GEN_7832; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7834 = 8'h2b == new_ptr_50_value ? ghv_43 : _GEN_7833; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7835 = 8'h2c == new_ptr_50_value ? ghv_44 : _GEN_7834; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7836 = 8'h2d == new_ptr_50_value ? ghv_45 : _GEN_7835; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7837 = 8'h2e == new_ptr_50_value ? ghv_46 : _GEN_7836; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7838 = 8'h2f == new_ptr_50_value ? ghv_47 : _GEN_7837; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7839 = 8'h30 == new_ptr_50_value ? ghv_48 : _GEN_7838; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7840 = 8'h31 == new_ptr_50_value ? ghv_49 : _GEN_7839; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7841 = 8'h32 == new_ptr_50_value ? ghv_50 : _GEN_7840; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7842 = 8'h33 == new_ptr_50_value ? ghv_51 : _GEN_7841; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7843 = 8'h34 == new_ptr_50_value ? ghv_52 : _GEN_7842; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7844 = 8'h35 == new_ptr_50_value ? ghv_53 : _GEN_7843; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7845 = 8'h36 == new_ptr_50_value ? ghv_54 : _GEN_7844; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7846 = 8'h37 == new_ptr_50_value ? ghv_55 : _GEN_7845; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7847 = 8'h38 == new_ptr_50_value ? ghv_56 : _GEN_7846; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7848 = 8'h39 == new_ptr_50_value ? ghv_57 : _GEN_7847; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7849 = 8'h3a == new_ptr_50_value ? ghv_58 : _GEN_7848; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7850 = 8'h3b == new_ptr_50_value ? ghv_59 : _GEN_7849; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7851 = 8'h3c == new_ptr_50_value ? ghv_60 : _GEN_7850; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7852 = 8'h3d == new_ptr_50_value ? ghv_61 : _GEN_7851; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7853 = 8'h3e == new_ptr_50_value ? ghv_62 : _GEN_7852; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7854 = 8'h3f == new_ptr_50_value ? ghv_63 : _GEN_7853; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7855 = 8'h40 == new_ptr_50_value ? ghv_64 : _GEN_7854; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7856 = 8'h41 == new_ptr_50_value ? ghv_65 : _GEN_7855; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7857 = 8'h42 == new_ptr_50_value ? ghv_66 : _GEN_7856; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7858 = 8'h43 == new_ptr_50_value ? ghv_67 : _GEN_7857; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7859 = 8'h44 == new_ptr_50_value ? ghv_68 : _GEN_7858; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7860 = 8'h45 == new_ptr_50_value ? ghv_69 : _GEN_7859; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7861 = 8'h46 == new_ptr_50_value ? ghv_70 : _GEN_7860; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7862 = 8'h47 == new_ptr_50_value ? ghv_71 : _GEN_7861; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7863 = 8'h48 == new_ptr_50_value ? ghv_72 : _GEN_7862; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7864 = 8'h49 == new_ptr_50_value ? ghv_73 : _GEN_7863; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7865 = 8'h4a == new_ptr_50_value ? ghv_74 : _GEN_7864; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7866 = 8'h4b == new_ptr_50_value ? ghv_75 : _GEN_7865; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7867 = 8'h4c == new_ptr_50_value ? ghv_76 : _GEN_7866; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7868 = 8'h4d == new_ptr_50_value ? ghv_77 : _GEN_7867; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7869 = 8'h4e == new_ptr_50_value ? ghv_78 : _GEN_7868; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7870 = 8'h4f == new_ptr_50_value ? ghv_79 : _GEN_7869; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7871 = 8'h50 == new_ptr_50_value ? ghv_80 : _GEN_7870; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7872 = 8'h51 == new_ptr_50_value ? ghv_81 : _GEN_7871; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7873 = 8'h52 == new_ptr_50_value ? ghv_82 : _GEN_7872; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7874 = 8'h53 == new_ptr_50_value ? ghv_83 : _GEN_7873; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7875 = 8'h54 == new_ptr_50_value ? ghv_84 : _GEN_7874; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7876 = 8'h55 == new_ptr_50_value ? ghv_85 : _GEN_7875; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7877 = 8'h56 == new_ptr_50_value ? ghv_86 : _GEN_7876; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7878 = 8'h57 == new_ptr_50_value ? ghv_87 : _GEN_7877; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7879 = 8'h58 == new_ptr_50_value ? ghv_88 : _GEN_7878; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7880 = 8'h59 == new_ptr_50_value ? ghv_89 : _GEN_7879; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7881 = 8'h5a == new_ptr_50_value ? ghv_90 : _GEN_7880; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7882 = 8'h5b == new_ptr_50_value ? ghv_91 : _GEN_7881; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7883 = 8'h5c == new_ptr_50_value ? ghv_92 : _GEN_7882; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7884 = 8'h5d == new_ptr_50_value ? ghv_93 : _GEN_7883; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7885 = 8'h5e == new_ptr_50_value ? ghv_94 : _GEN_7884; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7886 = 8'h5f == new_ptr_50_value ? ghv_95 : _GEN_7885; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7887 = 8'h60 == new_ptr_50_value ? ghv_96 : _GEN_7886; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7888 = 8'h61 == new_ptr_50_value ? ghv_97 : _GEN_7887; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7889 = 8'h62 == new_ptr_50_value ? ghv_98 : _GEN_7888; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7890 = 8'h63 == new_ptr_50_value ? ghv_99 : _GEN_7889; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7891 = 8'h64 == new_ptr_50_value ? ghv_100 : _GEN_7890; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7892 = 8'h65 == new_ptr_50_value ? ghv_101 : _GEN_7891; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7893 = 8'h66 == new_ptr_50_value ? ghv_102 : _GEN_7892; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7894 = 8'h67 == new_ptr_50_value ? ghv_103 : _GEN_7893; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7895 = 8'h68 == new_ptr_50_value ? ghv_104 : _GEN_7894; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7896 = 8'h69 == new_ptr_50_value ? ghv_105 : _GEN_7895; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7897 = 8'h6a == new_ptr_50_value ? ghv_106 : _GEN_7896; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7898 = 8'h6b == new_ptr_50_value ? ghv_107 : _GEN_7897; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7899 = 8'h6c == new_ptr_50_value ? ghv_108 : _GEN_7898; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7900 = 8'h6d == new_ptr_50_value ? ghv_109 : _GEN_7899; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7901 = 8'h6e == new_ptr_50_value ? ghv_110 : _GEN_7900; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7902 = 8'h6f == new_ptr_50_value ? ghv_111 : _GEN_7901; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7903 = 8'h70 == new_ptr_50_value ? ghv_112 : _GEN_7902; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7904 = 8'h71 == new_ptr_50_value ? ghv_113 : _GEN_7903; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7905 = 8'h72 == new_ptr_50_value ? ghv_114 : _GEN_7904; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7906 = 8'h73 == new_ptr_50_value ? ghv_115 : _GEN_7905; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7907 = 8'h74 == new_ptr_50_value ? ghv_116 : _GEN_7906; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7908 = 8'h75 == new_ptr_50_value ? ghv_117 : _GEN_7907; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7909 = 8'h76 == new_ptr_50_value ? ghv_118 : _GEN_7908; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7910 = 8'h77 == new_ptr_50_value ? ghv_119 : _GEN_7909; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7911 = 8'h78 == new_ptr_50_value ? ghv_120 : _GEN_7910; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7912 = 8'h79 == new_ptr_50_value ? ghv_121 : _GEN_7911; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7913 = 8'h7a == new_ptr_50_value ? ghv_122 : _GEN_7912; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7914 = 8'h7b == new_ptr_50_value ? ghv_123 : _GEN_7913; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7915 = 8'h7c == new_ptr_50_value ? ghv_124 : _GEN_7914; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7916 = 8'h7d == new_ptr_50_value ? ghv_125 : _GEN_7915; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7917 = 8'h7e == new_ptr_50_value ? ghv_126 : _GEN_7916; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7918 = 8'h7f == new_ptr_50_value ? ghv_127 : _GEN_7917; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7919 = 8'h80 == new_ptr_50_value ? ghv_128 : _GEN_7918; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7920 = 8'h81 == new_ptr_50_value ? ghv_129 : _GEN_7919; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7921 = 8'h82 == new_ptr_50_value ? ghv_130 : _GEN_7920; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7922 = 8'h83 == new_ptr_50_value ? ghv_131 : _GEN_7921; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7923 = 8'h84 == new_ptr_50_value ? ghv_132 : _GEN_7922; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7924 = 8'h85 == new_ptr_50_value ? ghv_133 : _GEN_7923; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7925 = 8'h86 == new_ptr_50_value ? ghv_134 : _GEN_7924; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7926 = 8'h87 == new_ptr_50_value ? ghv_135 : _GEN_7925; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7927 = 8'h88 == new_ptr_50_value ? ghv_136 : _GEN_7926; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7928 = 8'h89 == new_ptr_50_value ? ghv_137 : _GEN_7927; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7929 = 8'h8a == new_ptr_50_value ? ghv_138 : _GEN_7928; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7930 = 8'h8b == new_ptr_50_value ? ghv_139 : _GEN_7929; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7931 = 8'h8c == new_ptr_50_value ? ghv_140 : _GEN_7930; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7932 = 8'h8d == new_ptr_50_value ? ghv_141 : _GEN_7931; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7933 = 8'h8e == new_ptr_50_value ? ghv_142 : _GEN_7932; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_41_value = _new_ptr_value_T_83[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_7936 = 8'h1 == new_ptr_41_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7937 = 8'h2 == new_ptr_41_value ? ghv_2 : _GEN_7936; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7938 = 8'h3 == new_ptr_41_value ? ghv_3 : _GEN_7937; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7939 = 8'h4 == new_ptr_41_value ? ghv_4 : _GEN_7938; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7940 = 8'h5 == new_ptr_41_value ? ghv_5 : _GEN_7939; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7941 = 8'h6 == new_ptr_41_value ? ghv_6 : _GEN_7940; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7942 = 8'h7 == new_ptr_41_value ? ghv_7 : _GEN_7941; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7943 = 8'h8 == new_ptr_41_value ? ghv_8 : _GEN_7942; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7944 = 8'h9 == new_ptr_41_value ? ghv_9 : _GEN_7943; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7945 = 8'ha == new_ptr_41_value ? ghv_10 : _GEN_7944; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7946 = 8'hb == new_ptr_41_value ? ghv_11 : _GEN_7945; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7947 = 8'hc == new_ptr_41_value ? ghv_12 : _GEN_7946; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7948 = 8'hd == new_ptr_41_value ? ghv_13 : _GEN_7947; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7949 = 8'he == new_ptr_41_value ? ghv_14 : _GEN_7948; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7950 = 8'hf == new_ptr_41_value ? ghv_15 : _GEN_7949; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7951 = 8'h10 == new_ptr_41_value ? ghv_16 : _GEN_7950; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7952 = 8'h11 == new_ptr_41_value ? ghv_17 : _GEN_7951; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7953 = 8'h12 == new_ptr_41_value ? ghv_18 : _GEN_7952; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7954 = 8'h13 == new_ptr_41_value ? ghv_19 : _GEN_7953; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7955 = 8'h14 == new_ptr_41_value ? ghv_20 : _GEN_7954; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7956 = 8'h15 == new_ptr_41_value ? ghv_21 : _GEN_7955; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7957 = 8'h16 == new_ptr_41_value ? ghv_22 : _GEN_7956; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7958 = 8'h17 == new_ptr_41_value ? ghv_23 : _GEN_7957; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7959 = 8'h18 == new_ptr_41_value ? ghv_24 : _GEN_7958; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7960 = 8'h19 == new_ptr_41_value ? ghv_25 : _GEN_7959; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7961 = 8'h1a == new_ptr_41_value ? ghv_26 : _GEN_7960; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7962 = 8'h1b == new_ptr_41_value ? ghv_27 : _GEN_7961; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7963 = 8'h1c == new_ptr_41_value ? ghv_28 : _GEN_7962; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7964 = 8'h1d == new_ptr_41_value ? ghv_29 : _GEN_7963; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7965 = 8'h1e == new_ptr_41_value ? ghv_30 : _GEN_7964; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7966 = 8'h1f == new_ptr_41_value ? ghv_31 : _GEN_7965; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7967 = 8'h20 == new_ptr_41_value ? ghv_32 : _GEN_7966; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7968 = 8'h21 == new_ptr_41_value ? ghv_33 : _GEN_7967; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7969 = 8'h22 == new_ptr_41_value ? ghv_34 : _GEN_7968; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7970 = 8'h23 == new_ptr_41_value ? ghv_35 : _GEN_7969; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7971 = 8'h24 == new_ptr_41_value ? ghv_36 : _GEN_7970; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7972 = 8'h25 == new_ptr_41_value ? ghv_37 : _GEN_7971; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7973 = 8'h26 == new_ptr_41_value ? ghv_38 : _GEN_7972; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7974 = 8'h27 == new_ptr_41_value ? ghv_39 : _GEN_7973; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7975 = 8'h28 == new_ptr_41_value ? ghv_40 : _GEN_7974; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7976 = 8'h29 == new_ptr_41_value ? ghv_41 : _GEN_7975; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7977 = 8'h2a == new_ptr_41_value ? ghv_42 : _GEN_7976; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7978 = 8'h2b == new_ptr_41_value ? ghv_43 : _GEN_7977; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7979 = 8'h2c == new_ptr_41_value ? ghv_44 : _GEN_7978; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7980 = 8'h2d == new_ptr_41_value ? ghv_45 : _GEN_7979; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7981 = 8'h2e == new_ptr_41_value ? ghv_46 : _GEN_7980; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7982 = 8'h2f == new_ptr_41_value ? ghv_47 : _GEN_7981; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7983 = 8'h30 == new_ptr_41_value ? ghv_48 : _GEN_7982; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7984 = 8'h31 == new_ptr_41_value ? ghv_49 : _GEN_7983; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7985 = 8'h32 == new_ptr_41_value ? ghv_50 : _GEN_7984; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7986 = 8'h33 == new_ptr_41_value ? ghv_51 : _GEN_7985; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7987 = 8'h34 == new_ptr_41_value ? ghv_52 : _GEN_7986; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7988 = 8'h35 == new_ptr_41_value ? ghv_53 : _GEN_7987; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7989 = 8'h36 == new_ptr_41_value ? ghv_54 : _GEN_7988; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7990 = 8'h37 == new_ptr_41_value ? ghv_55 : _GEN_7989; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7991 = 8'h38 == new_ptr_41_value ? ghv_56 : _GEN_7990; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7992 = 8'h39 == new_ptr_41_value ? ghv_57 : _GEN_7991; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7993 = 8'h3a == new_ptr_41_value ? ghv_58 : _GEN_7992; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7994 = 8'h3b == new_ptr_41_value ? ghv_59 : _GEN_7993; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7995 = 8'h3c == new_ptr_41_value ? ghv_60 : _GEN_7994; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7996 = 8'h3d == new_ptr_41_value ? ghv_61 : _GEN_7995; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7997 = 8'h3e == new_ptr_41_value ? ghv_62 : _GEN_7996; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7998 = 8'h3f == new_ptr_41_value ? ghv_63 : _GEN_7997; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_7999 = 8'h40 == new_ptr_41_value ? ghv_64 : _GEN_7998; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8000 = 8'h41 == new_ptr_41_value ? ghv_65 : _GEN_7999; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8001 = 8'h42 == new_ptr_41_value ? ghv_66 : _GEN_8000; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8002 = 8'h43 == new_ptr_41_value ? ghv_67 : _GEN_8001; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8003 = 8'h44 == new_ptr_41_value ? ghv_68 : _GEN_8002; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8004 = 8'h45 == new_ptr_41_value ? ghv_69 : _GEN_8003; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8005 = 8'h46 == new_ptr_41_value ? ghv_70 : _GEN_8004; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8006 = 8'h47 == new_ptr_41_value ? ghv_71 : _GEN_8005; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8007 = 8'h48 == new_ptr_41_value ? ghv_72 : _GEN_8006; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8008 = 8'h49 == new_ptr_41_value ? ghv_73 : _GEN_8007; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8009 = 8'h4a == new_ptr_41_value ? ghv_74 : _GEN_8008; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8010 = 8'h4b == new_ptr_41_value ? ghv_75 : _GEN_8009; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8011 = 8'h4c == new_ptr_41_value ? ghv_76 : _GEN_8010; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8012 = 8'h4d == new_ptr_41_value ? ghv_77 : _GEN_8011; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8013 = 8'h4e == new_ptr_41_value ? ghv_78 : _GEN_8012; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8014 = 8'h4f == new_ptr_41_value ? ghv_79 : _GEN_8013; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8015 = 8'h50 == new_ptr_41_value ? ghv_80 : _GEN_8014; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8016 = 8'h51 == new_ptr_41_value ? ghv_81 : _GEN_8015; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8017 = 8'h52 == new_ptr_41_value ? ghv_82 : _GEN_8016; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8018 = 8'h53 == new_ptr_41_value ? ghv_83 : _GEN_8017; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8019 = 8'h54 == new_ptr_41_value ? ghv_84 : _GEN_8018; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8020 = 8'h55 == new_ptr_41_value ? ghv_85 : _GEN_8019; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8021 = 8'h56 == new_ptr_41_value ? ghv_86 : _GEN_8020; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8022 = 8'h57 == new_ptr_41_value ? ghv_87 : _GEN_8021; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8023 = 8'h58 == new_ptr_41_value ? ghv_88 : _GEN_8022; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8024 = 8'h59 == new_ptr_41_value ? ghv_89 : _GEN_8023; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8025 = 8'h5a == new_ptr_41_value ? ghv_90 : _GEN_8024; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8026 = 8'h5b == new_ptr_41_value ? ghv_91 : _GEN_8025; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8027 = 8'h5c == new_ptr_41_value ? ghv_92 : _GEN_8026; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8028 = 8'h5d == new_ptr_41_value ? ghv_93 : _GEN_8027; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8029 = 8'h5e == new_ptr_41_value ? ghv_94 : _GEN_8028; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8030 = 8'h5f == new_ptr_41_value ? ghv_95 : _GEN_8029; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8031 = 8'h60 == new_ptr_41_value ? ghv_96 : _GEN_8030; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8032 = 8'h61 == new_ptr_41_value ? ghv_97 : _GEN_8031; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8033 = 8'h62 == new_ptr_41_value ? ghv_98 : _GEN_8032; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8034 = 8'h63 == new_ptr_41_value ? ghv_99 : _GEN_8033; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8035 = 8'h64 == new_ptr_41_value ? ghv_100 : _GEN_8034; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8036 = 8'h65 == new_ptr_41_value ? ghv_101 : _GEN_8035; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8037 = 8'h66 == new_ptr_41_value ? ghv_102 : _GEN_8036; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8038 = 8'h67 == new_ptr_41_value ? ghv_103 : _GEN_8037; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8039 = 8'h68 == new_ptr_41_value ? ghv_104 : _GEN_8038; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8040 = 8'h69 == new_ptr_41_value ? ghv_105 : _GEN_8039; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8041 = 8'h6a == new_ptr_41_value ? ghv_106 : _GEN_8040; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8042 = 8'h6b == new_ptr_41_value ? ghv_107 : _GEN_8041; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8043 = 8'h6c == new_ptr_41_value ? ghv_108 : _GEN_8042; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8044 = 8'h6d == new_ptr_41_value ? ghv_109 : _GEN_8043; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8045 = 8'h6e == new_ptr_41_value ? ghv_110 : _GEN_8044; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8046 = 8'h6f == new_ptr_41_value ? ghv_111 : _GEN_8045; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8047 = 8'h70 == new_ptr_41_value ? ghv_112 : _GEN_8046; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8048 = 8'h71 == new_ptr_41_value ? ghv_113 : _GEN_8047; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8049 = 8'h72 == new_ptr_41_value ? ghv_114 : _GEN_8048; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8050 = 8'h73 == new_ptr_41_value ? ghv_115 : _GEN_8049; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8051 = 8'h74 == new_ptr_41_value ? ghv_116 : _GEN_8050; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8052 = 8'h75 == new_ptr_41_value ? ghv_117 : _GEN_8051; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8053 = 8'h76 == new_ptr_41_value ? ghv_118 : _GEN_8052; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8054 = 8'h77 == new_ptr_41_value ? ghv_119 : _GEN_8053; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8055 = 8'h78 == new_ptr_41_value ? ghv_120 : _GEN_8054; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8056 = 8'h79 == new_ptr_41_value ? ghv_121 : _GEN_8055; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8057 = 8'h7a == new_ptr_41_value ? ghv_122 : _GEN_8056; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8058 = 8'h7b == new_ptr_41_value ? ghv_123 : _GEN_8057; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8059 = 8'h7c == new_ptr_41_value ? ghv_124 : _GEN_8058; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8060 = 8'h7d == new_ptr_41_value ? ghv_125 : _GEN_8059; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8061 = 8'h7e == new_ptr_41_value ? ghv_126 : _GEN_8060; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8062 = 8'h7f == new_ptr_41_value ? ghv_127 : _GEN_8061; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8063 = 8'h80 == new_ptr_41_value ? ghv_128 : _GEN_8062; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8064 = 8'h81 == new_ptr_41_value ? ghv_129 : _GEN_8063; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8065 = 8'h82 == new_ptr_41_value ? ghv_130 : _GEN_8064; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8066 = 8'h83 == new_ptr_41_value ? ghv_131 : _GEN_8065; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8067 = 8'h84 == new_ptr_41_value ? ghv_132 : _GEN_8066; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8068 = 8'h85 == new_ptr_41_value ? ghv_133 : _GEN_8067; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8069 = 8'h86 == new_ptr_41_value ? ghv_134 : _GEN_8068; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8070 = 8'h87 == new_ptr_41_value ? ghv_135 : _GEN_8069; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8071 = 8'h88 == new_ptr_41_value ? ghv_136 : _GEN_8070; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8072 = 8'h89 == new_ptr_41_value ? ghv_137 : _GEN_8071; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8073 = 8'h8a == new_ptr_41_value ? ghv_138 : _GEN_8072; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8074 = 8'h8b == new_ptr_41_value ? ghv_139 : _GEN_8073; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8075 = 8'h8c == new_ptr_41_value ? ghv_140 : _GEN_8074; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8076 = 8'h8d == new_ptr_41_value ? ghv_141 : _GEN_8075; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8077 = 8'h8e == new_ptr_41_value ? ghv_142 : _GEN_8076; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_58_value = _new_ptr_value_T_117[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_8080 = 8'h1 == new_ptr_58_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8081 = 8'h2 == new_ptr_58_value ? ghv_2 : _GEN_8080; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8082 = 8'h3 == new_ptr_58_value ? ghv_3 : _GEN_8081; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8083 = 8'h4 == new_ptr_58_value ? ghv_4 : _GEN_8082; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8084 = 8'h5 == new_ptr_58_value ? ghv_5 : _GEN_8083; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8085 = 8'h6 == new_ptr_58_value ? ghv_6 : _GEN_8084; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8086 = 8'h7 == new_ptr_58_value ? ghv_7 : _GEN_8085; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8087 = 8'h8 == new_ptr_58_value ? ghv_8 : _GEN_8086; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8088 = 8'h9 == new_ptr_58_value ? ghv_9 : _GEN_8087; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8089 = 8'ha == new_ptr_58_value ? ghv_10 : _GEN_8088; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8090 = 8'hb == new_ptr_58_value ? ghv_11 : _GEN_8089; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8091 = 8'hc == new_ptr_58_value ? ghv_12 : _GEN_8090; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8092 = 8'hd == new_ptr_58_value ? ghv_13 : _GEN_8091; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8093 = 8'he == new_ptr_58_value ? ghv_14 : _GEN_8092; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8094 = 8'hf == new_ptr_58_value ? ghv_15 : _GEN_8093; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8095 = 8'h10 == new_ptr_58_value ? ghv_16 : _GEN_8094; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8096 = 8'h11 == new_ptr_58_value ? ghv_17 : _GEN_8095; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8097 = 8'h12 == new_ptr_58_value ? ghv_18 : _GEN_8096; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8098 = 8'h13 == new_ptr_58_value ? ghv_19 : _GEN_8097; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8099 = 8'h14 == new_ptr_58_value ? ghv_20 : _GEN_8098; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8100 = 8'h15 == new_ptr_58_value ? ghv_21 : _GEN_8099; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8101 = 8'h16 == new_ptr_58_value ? ghv_22 : _GEN_8100; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8102 = 8'h17 == new_ptr_58_value ? ghv_23 : _GEN_8101; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8103 = 8'h18 == new_ptr_58_value ? ghv_24 : _GEN_8102; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8104 = 8'h19 == new_ptr_58_value ? ghv_25 : _GEN_8103; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8105 = 8'h1a == new_ptr_58_value ? ghv_26 : _GEN_8104; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8106 = 8'h1b == new_ptr_58_value ? ghv_27 : _GEN_8105; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8107 = 8'h1c == new_ptr_58_value ? ghv_28 : _GEN_8106; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8108 = 8'h1d == new_ptr_58_value ? ghv_29 : _GEN_8107; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8109 = 8'h1e == new_ptr_58_value ? ghv_30 : _GEN_8108; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8110 = 8'h1f == new_ptr_58_value ? ghv_31 : _GEN_8109; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8111 = 8'h20 == new_ptr_58_value ? ghv_32 : _GEN_8110; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8112 = 8'h21 == new_ptr_58_value ? ghv_33 : _GEN_8111; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8113 = 8'h22 == new_ptr_58_value ? ghv_34 : _GEN_8112; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8114 = 8'h23 == new_ptr_58_value ? ghv_35 : _GEN_8113; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8115 = 8'h24 == new_ptr_58_value ? ghv_36 : _GEN_8114; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8116 = 8'h25 == new_ptr_58_value ? ghv_37 : _GEN_8115; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8117 = 8'h26 == new_ptr_58_value ? ghv_38 : _GEN_8116; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8118 = 8'h27 == new_ptr_58_value ? ghv_39 : _GEN_8117; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8119 = 8'h28 == new_ptr_58_value ? ghv_40 : _GEN_8118; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8120 = 8'h29 == new_ptr_58_value ? ghv_41 : _GEN_8119; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8121 = 8'h2a == new_ptr_58_value ? ghv_42 : _GEN_8120; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8122 = 8'h2b == new_ptr_58_value ? ghv_43 : _GEN_8121; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8123 = 8'h2c == new_ptr_58_value ? ghv_44 : _GEN_8122; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8124 = 8'h2d == new_ptr_58_value ? ghv_45 : _GEN_8123; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8125 = 8'h2e == new_ptr_58_value ? ghv_46 : _GEN_8124; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8126 = 8'h2f == new_ptr_58_value ? ghv_47 : _GEN_8125; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8127 = 8'h30 == new_ptr_58_value ? ghv_48 : _GEN_8126; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8128 = 8'h31 == new_ptr_58_value ? ghv_49 : _GEN_8127; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8129 = 8'h32 == new_ptr_58_value ? ghv_50 : _GEN_8128; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8130 = 8'h33 == new_ptr_58_value ? ghv_51 : _GEN_8129; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8131 = 8'h34 == new_ptr_58_value ? ghv_52 : _GEN_8130; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8132 = 8'h35 == new_ptr_58_value ? ghv_53 : _GEN_8131; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8133 = 8'h36 == new_ptr_58_value ? ghv_54 : _GEN_8132; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8134 = 8'h37 == new_ptr_58_value ? ghv_55 : _GEN_8133; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8135 = 8'h38 == new_ptr_58_value ? ghv_56 : _GEN_8134; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8136 = 8'h39 == new_ptr_58_value ? ghv_57 : _GEN_8135; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8137 = 8'h3a == new_ptr_58_value ? ghv_58 : _GEN_8136; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8138 = 8'h3b == new_ptr_58_value ? ghv_59 : _GEN_8137; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8139 = 8'h3c == new_ptr_58_value ? ghv_60 : _GEN_8138; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8140 = 8'h3d == new_ptr_58_value ? ghv_61 : _GEN_8139; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8141 = 8'h3e == new_ptr_58_value ? ghv_62 : _GEN_8140; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8142 = 8'h3f == new_ptr_58_value ? ghv_63 : _GEN_8141; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8143 = 8'h40 == new_ptr_58_value ? ghv_64 : _GEN_8142; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8144 = 8'h41 == new_ptr_58_value ? ghv_65 : _GEN_8143; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8145 = 8'h42 == new_ptr_58_value ? ghv_66 : _GEN_8144; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8146 = 8'h43 == new_ptr_58_value ? ghv_67 : _GEN_8145; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8147 = 8'h44 == new_ptr_58_value ? ghv_68 : _GEN_8146; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8148 = 8'h45 == new_ptr_58_value ? ghv_69 : _GEN_8147; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8149 = 8'h46 == new_ptr_58_value ? ghv_70 : _GEN_8148; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8150 = 8'h47 == new_ptr_58_value ? ghv_71 : _GEN_8149; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8151 = 8'h48 == new_ptr_58_value ? ghv_72 : _GEN_8150; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8152 = 8'h49 == new_ptr_58_value ? ghv_73 : _GEN_8151; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8153 = 8'h4a == new_ptr_58_value ? ghv_74 : _GEN_8152; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8154 = 8'h4b == new_ptr_58_value ? ghv_75 : _GEN_8153; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8155 = 8'h4c == new_ptr_58_value ? ghv_76 : _GEN_8154; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8156 = 8'h4d == new_ptr_58_value ? ghv_77 : _GEN_8155; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8157 = 8'h4e == new_ptr_58_value ? ghv_78 : _GEN_8156; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8158 = 8'h4f == new_ptr_58_value ? ghv_79 : _GEN_8157; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8159 = 8'h50 == new_ptr_58_value ? ghv_80 : _GEN_8158; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8160 = 8'h51 == new_ptr_58_value ? ghv_81 : _GEN_8159; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8161 = 8'h52 == new_ptr_58_value ? ghv_82 : _GEN_8160; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8162 = 8'h53 == new_ptr_58_value ? ghv_83 : _GEN_8161; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8163 = 8'h54 == new_ptr_58_value ? ghv_84 : _GEN_8162; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8164 = 8'h55 == new_ptr_58_value ? ghv_85 : _GEN_8163; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8165 = 8'h56 == new_ptr_58_value ? ghv_86 : _GEN_8164; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8166 = 8'h57 == new_ptr_58_value ? ghv_87 : _GEN_8165; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8167 = 8'h58 == new_ptr_58_value ? ghv_88 : _GEN_8166; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8168 = 8'h59 == new_ptr_58_value ? ghv_89 : _GEN_8167; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8169 = 8'h5a == new_ptr_58_value ? ghv_90 : _GEN_8168; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8170 = 8'h5b == new_ptr_58_value ? ghv_91 : _GEN_8169; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8171 = 8'h5c == new_ptr_58_value ? ghv_92 : _GEN_8170; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8172 = 8'h5d == new_ptr_58_value ? ghv_93 : _GEN_8171; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8173 = 8'h5e == new_ptr_58_value ? ghv_94 : _GEN_8172; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8174 = 8'h5f == new_ptr_58_value ? ghv_95 : _GEN_8173; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8175 = 8'h60 == new_ptr_58_value ? ghv_96 : _GEN_8174; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8176 = 8'h61 == new_ptr_58_value ? ghv_97 : _GEN_8175; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8177 = 8'h62 == new_ptr_58_value ? ghv_98 : _GEN_8176; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8178 = 8'h63 == new_ptr_58_value ? ghv_99 : _GEN_8177; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8179 = 8'h64 == new_ptr_58_value ? ghv_100 : _GEN_8178; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8180 = 8'h65 == new_ptr_58_value ? ghv_101 : _GEN_8179; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8181 = 8'h66 == new_ptr_58_value ? ghv_102 : _GEN_8180; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8182 = 8'h67 == new_ptr_58_value ? ghv_103 : _GEN_8181; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8183 = 8'h68 == new_ptr_58_value ? ghv_104 : _GEN_8182; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8184 = 8'h69 == new_ptr_58_value ? ghv_105 : _GEN_8183; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8185 = 8'h6a == new_ptr_58_value ? ghv_106 : _GEN_8184; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8186 = 8'h6b == new_ptr_58_value ? ghv_107 : _GEN_8185; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8187 = 8'h6c == new_ptr_58_value ? ghv_108 : _GEN_8186; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8188 = 8'h6d == new_ptr_58_value ? ghv_109 : _GEN_8187; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8189 = 8'h6e == new_ptr_58_value ? ghv_110 : _GEN_8188; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8190 = 8'h6f == new_ptr_58_value ? ghv_111 : _GEN_8189; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8191 = 8'h70 == new_ptr_58_value ? ghv_112 : _GEN_8190; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8192 = 8'h71 == new_ptr_58_value ? ghv_113 : _GEN_8191; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8193 = 8'h72 == new_ptr_58_value ? ghv_114 : _GEN_8192; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8194 = 8'h73 == new_ptr_58_value ? ghv_115 : _GEN_8193; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8195 = 8'h74 == new_ptr_58_value ? ghv_116 : _GEN_8194; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8196 = 8'h75 == new_ptr_58_value ? ghv_117 : _GEN_8195; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8197 = 8'h76 == new_ptr_58_value ? ghv_118 : _GEN_8196; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8198 = 8'h77 == new_ptr_58_value ? ghv_119 : _GEN_8197; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8199 = 8'h78 == new_ptr_58_value ? ghv_120 : _GEN_8198; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8200 = 8'h79 == new_ptr_58_value ? ghv_121 : _GEN_8199; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8201 = 8'h7a == new_ptr_58_value ? ghv_122 : _GEN_8200; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8202 = 8'h7b == new_ptr_58_value ? ghv_123 : _GEN_8201; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8203 = 8'h7c == new_ptr_58_value ? ghv_124 : _GEN_8202; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8204 = 8'h7d == new_ptr_58_value ? ghv_125 : _GEN_8203; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8205 = 8'h7e == new_ptr_58_value ? ghv_126 : _GEN_8204; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8206 = 8'h7f == new_ptr_58_value ? ghv_127 : _GEN_8205; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8207 = 8'h80 == new_ptr_58_value ? ghv_128 : _GEN_8206; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8208 = 8'h81 == new_ptr_58_value ? ghv_129 : _GEN_8207; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8209 = 8'h82 == new_ptr_58_value ? ghv_130 : _GEN_8208; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8210 = 8'h83 == new_ptr_58_value ? ghv_131 : _GEN_8209; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8211 = 8'h84 == new_ptr_58_value ? ghv_132 : _GEN_8210; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8212 = 8'h85 == new_ptr_58_value ? ghv_133 : _GEN_8211; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8213 = 8'h86 == new_ptr_58_value ? ghv_134 : _GEN_8212; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8214 = 8'h87 == new_ptr_58_value ? ghv_135 : _GEN_8213; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8215 = 8'h88 == new_ptr_58_value ? ghv_136 : _GEN_8214; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8216 = 8'h89 == new_ptr_58_value ? ghv_137 : _GEN_8215; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8217 = 8'h8a == new_ptr_58_value ? ghv_138 : _GEN_8216; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8218 = 8'h8b == new_ptr_58_value ? ghv_139 : _GEN_8217; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8219 = 8'h8c == new_ptr_58_value ? ghv_140 : _GEN_8218; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8220 = 8'h8d == new_ptr_58_value ? ghv_141 : _GEN_8219; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8221 = 8'h8e == new_ptr_58_value ? ghv_142 : _GEN_8220; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_51_value = _new_ptr_value_T_103[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_8224 = 8'h1 == new_ptr_51_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8225 = 8'h2 == new_ptr_51_value ? ghv_2 : _GEN_8224; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8226 = 8'h3 == new_ptr_51_value ? ghv_3 : _GEN_8225; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8227 = 8'h4 == new_ptr_51_value ? ghv_4 : _GEN_8226; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8228 = 8'h5 == new_ptr_51_value ? ghv_5 : _GEN_8227; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8229 = 8'h6 == new_ptr_51_value ? ghv_6 : _GEN_8228; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8230 = 8'h7 == new_ptr_51_value ? ghv_7 : _GEN_8229; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8231 = 8'h8 == new_ptr_51_value ? ghv_8 : _GEN_8230; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8232 = 8'h9 == new_ptr_51_value ? ghv_9 : _GEN_8231; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8233 = 8'ha == new_ptr_51_value ? ghv_10 : _GEN_8232; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8234 = 8'hb == new_ptr_51_value ? ghv_11 : _GEN_8233; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8235 = 8'hc == new_ptr_51_value ? ghv_12 : _GEN_8234; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8236 = 8'hd == new_ptr_51_value ? ghv_13 : _GEN_8235; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8237 = 8'he == new_ptr_51_value ? ghv_14 : _GEN_8236; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8238 = 8'hf == new_ptr_51_value ? ghv_15 : _GEN_8237; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8239 = 8'h10 == new_ptr_51_value ? ghv_16 : _GEN_8238; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8240 = 8'h11 == new_ptr_51_value ? ghv_17 : _GEN_8239; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8241 = 8'h12 == new_ptr_51_value ? ghv_18 : _GEN_8240; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8242 = 8'h13 == new_ptr_51_value ? ghv_19 : _GEN_8241; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8243 = 8'h14 == new_ptr_51_value ? ghv_20 : _GEN_8242; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8244 = 8'h15 == new_ptr_51_value ? ghv_21 : _GEN_8243; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8245 = 8'h16 == new_ptr_51_value ? ghv_22 : _GEN_8244; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8246 = 8'h17 == new_ptr_51_value ? ghv_23 : _GEN_8245; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8247 = 8'h18 == new_ptr_51_value ? ghv_24 : _GEN_8246; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8248 = 8'h19 == new_ptr_51_value ? ghv_25 : _GEN_8247; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8249 = 8'h1a == new_ptr_51_value ? ghv_26 : _GEN_8248; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8250 = 8'h1b == new_ptr_51_value ? ghv_27 : _GEN_8249; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8251 = 8'h1c == new_ptr_51_value ? ghv_28 : _GEN_8250; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8252 = 8'h1d == new_ptr_51_value ? ghv_29 : _GEN_8251; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8253 = 8'h1e == new_ptr_51_value ? ghv_30 : _GEN_8252; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8254 = 8'h1f == new_ptr_51_value ? ghv_31 : _GEN_8253; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8255 = 8'h20 == new_ptr_51_value ? ghv_32 : _GEN_8254; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8256 = 8'h21 == new_ptr_51_value ? ghv_33 : _GEN_8255; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8257 = 8'h22 == new_ptr_51_value ? ghv_34 : _GEN_8256; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8258 = 8'h23 == new_ptr_51_value ? ghv_35 : _GEN_8257; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8259 = 8'h24 == new_ptr_51_value ? ghv_36 : _GEN_8258; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8260 = 8'h25 == new_ptr_51_value ? ghv_37 : _GEN_8259; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8261 = 8'h26 == new_ptr_51_value ? ghv_38 : _GEN_8260; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8262 = 8'h27 == new_ptr_51_value ? ghv_39 : _GEN_8261; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8263 = 8'h28 == new_ptr_51_value ? ghv_40 : _GEN_8262; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8264 = 8'h29 == new_ptr_51_value ? ghv_41 : _GEN_8263; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8265 = 8'h2a == new_ptr_51_value ? ghv_42 : _GEN_8264; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8266 = 8'h2b == new_ptr_51_value ? ghv_43 : _GEN_8265; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8267 = 8'h2c == new_ptr_51_value ? ghv_44 : _GEN_8266; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8268 = 8'h2d == new_ptr_51_value ? ghv_45 : _GEN_8267; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8269 = 8'h2e == new_ptr_51_value ? ghv_46 : _GEN_8268; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8270 = 8'h2f == new_ptr_51_value ? ghv_47 : _GEN_8269; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8271 = 8'h30 == new_ptr_51_value ? ghv_48 : _GEN_8270; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8272 = 8'h31 == new_ptr_51_value ? ghv_49 : _GEN_8271; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8273 = 8'h32 == new_ptr_51_value ? ghv_50 : _GEN_8272; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8274 = 8'h33 == new_ptr_51_value ? ghv_51 : _GEN_8273; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8275 = 8'h34 == new_ptr_51_value ? ghv_52 : _GEN_8274; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8276 = 8'h35 == new_ptr_51_value ? ghv_53 : _GEN_8275; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8277 = 8'h36 == new_ptr_51_value ? ghv_54 : _GEN_8276; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8278 = 8'h37 == new_ptr_51_value ? ghv_55 : _GEN_8277; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8279 = 8'h38 == new_ptr_51_value ? ghv_56 : _GEN_8278; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8280 = 8'h39 == new_ptr_51_value ? ghv_57 : _GEN_8279; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8281 = 8'h3a == new_ptr_51_value ? ghv_58 : _GEN_8280; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8282 = 8'h3b == new_ptr_51_value ? ghv_59 : _GEN_8281; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8283 = 8'h3c == new_ptr_51_value ? ghv_60 : _GEN_8282; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8284 = 8'h3d == new_ptr_51_value ? ghv_61 : _GEN_8283; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8285 = 8'h3e == new_ptr_51_value ? ghv_62 : _GEN_8284; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8286 = 8'h3f == new_ptr_51_value ? ghv_63 : _GEN_8285; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8287 = 8'h40 == new_ptr_51_value ? ghv_64 : _GEN_8286; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8288 = 8'h41 == new_ptr_51_value ? ghv_65 : _GEN_8287; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8289 = 8'h42 == new_ptr_51_value ? ghv_66 : _GEN_8288; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8290 = 8'h43 == new_ptr_51_value ? ghv_67 : _GEN_8289; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8291 = 8'h44 == new_ptr_51_value ? ghv_68 : _GEN_8290; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8292 = 8'h45 == new_ptr_51_value ? ghv_69 : _GEN_8291; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8293 = 8'h46 == new_ptr_51_value ? ghv_70 : _GEN_8292; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8294 = 8'h47 == new_ptr_51_value ? ghv_71 : _GEN_8293; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8295 = 8'h48 == new_ptr_51_value ? ghv_72 : _GEN_8294; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8296 = 8'h49 == new_ptr_51_value ? ghv_73 : _GEN_8295; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8297 = 8'h4a == new_ptr_51_value ? ghv_74 : _GEN_8296; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8298 = 8'h4b == new_ptr_51_value ? ghv_75 : _GEN_8297; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8299 = 8'h4c == new_ptr_51_value ? ghv_76 : _GEN_8298; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8300 = 8'h4d == new_ptr_51_value ? ghv_77 : _GEN_8299; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8301 = 8'h4e == new_ptr_51_value ? ghv_78 : _GEN_8300; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8302 = 8'h4f == new_ptr_51_value ? ghv_79 : _GEN_8301; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8303 = 8'h50 == new_ptr_51_value ? ghv_80 : _GEN_8302; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8304 = 8'h51 == new_ptr_51_value ? ghv_81 : _GEN_8303; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8305 = 8'h52 == new_ptr_51_value ? ghv_82 : _GEN_8304; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8306 = 8'h53 == new_ptr_51_value ? ghv_83 : _GEN_8305; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8307 = 8'h54 == new_ptr_51_value ? ghv_84 : _GEN_8306; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8308 = 8'h55 == new_ptr_51_value ? ghv_85 : _GEN_8307; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8309 = 8'h56 == new_ptr_51_value ? ghv_86 : _GEN_8308; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8310 = 8'h57 == new_ptr_51_value ? ghv_87 : _GEN_8309; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8311 = 8'h58 == new_ptr_51_value ? ghv_88 : _GEN_8310; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8312 = 8'h59 == new_ptr_51_value ? ghv_89 : _GEN_8311; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8313 = 8'h5a == new_ptr_51_value ? ghv_90 : _GEN_8312; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8314 = 8'h5b == new_ptr_51_value ? ghv_91 : _GEN_8313; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8315 = 8'h5c == new_ptr_51_value ? ghv_92 : _GEN_8314; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8316 = 8'h5d == new_ptr_51_value ? ghv_93 : _GEN_8315; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8317 = 8'h5e == new_ptr_51_value ? ghv_94 : _GEN_8316; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8318 = 8'h5f == new_ptr_51_value ? ghv_95 : _GEN_8317; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8319 = 8'h60 == new_ptr_51_value ? ghv_96 : _GEN_8318; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8320 = 8'h61 == new_ptr_51_value ? ghv_97 : _GEN_8319; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8321 = 8'h62 == new_ptr_51_value ? ghv_98 : _GEN_8320; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8322 = 8'h63 == new_ptr_51_value ? ghv_99 : _GEN_8321; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8323 = 8'h64 == new_ptr_51_value ? ghv_100 : _GEN_8322; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8324 = 8'h65 == new_ptr_51_value ? ghv_101 : _GEN_8323; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8325 = 8'h66 == new_ptr_51_value ? ghv_102 : _GEN_8324; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8326 = 8'h67 == new_ptr_51_value ? ghv_103 : _GEN_8325; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8327 = 8'h68 == new_ptr_51_value ? ghv_104 : _GEN_8326; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8328 = 8'h69 == new_ptr_51_value ? ghv_105 : _GEN_8327; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8329 = 8'h6a == new_ptr_51_value ? ghv_106 : _GEN_8328; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8330 = 8'h6b == new_ptr_51_value ? ghv_107 : _GEN_8329; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8331 = 8'h6c == new_ptr_51_value ? ghv_108 : _GEN_8330; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8332 = 8'h6d == new_ptr_51_value ? ghv_109 : _GEN_8331; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8333 = 8'h6e == new_ptr_51_value ? ghv_110 : _GEN_8332; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8334 = 8'h6f == new_ptr_51_value ? ghv_111 : _GEN_8333; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8335 = 8'h70 == new_ptr_51_value ? ghv_112 : _GEN_8334; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8336 = 8'h71 == new_ptr_51_value ? ghv_113 : _GEN_8335; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8337 = 8'h72 == new_ptr_51_value ? ghv_114 : _GEN_8336; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8338 = 8'h73 == new_ptr_51_value ? ghv_115 : _GEN_8337; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8339 = 8'h74 == new_ptr_51_value ? ghv_116 : _GEN_8338; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8340 = 8'h75 == new_ptr_51_value ? ghv_117 : _GEN_8339; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8341 = 8'h76 == new_ptr_51_value ? ghv_118 : _GEN_8340; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8342 = 8'h77 == new_ptr_51_value ? ghv_119 : _GEN_8341; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8343 = 8'h78 == new_ptr_51_value ? ghv_120 : _GEN_8342; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8344 = 8'h79 == new_ptr_51_value ? ghv_121 : _GEN_8343; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8345 = 8'h7a == new_ptr_51_value ? ghv_122 : _GEN_8344; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8346 = 8'h7b == new_ptr_51_value ? ghv_123 : _GEN_8345; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8347 = 8'h7c == new_ptr_51_value ? ghv_124 : _GEN_8346; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8348 = 8'h7d == new_ptr_51_value ? ghv_125 : _GEN_8347; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8349 = 8'h7e == new_ptr_51_value ? ghv_126 : _GEN_8348; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8350 = 8'h7f == new_ptr_51_value ? ghv_127 : _GEN_8349; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8351 = 8'h80 == new_ptr_51_value ? ghv_128 : _GEN_8350; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8352 = 8'h81 == new_ptr_51_value ? ghv_129 : _GEN_8351; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8353 = 8'h82 == new_ptr_51_value ? ghv_130 : _GEN_8352; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8354 = 8'h83 == new_ptr_51_value ? ghv_131 : _GEN_8353; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8355 = 8'h84 == new_ptr_51_value ? ghv_132 : _GEN_8354; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8356 = 8'h85 == new_ptr_51_value ? ghv_133 : _GEN_8355; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8357 = 8'h86 == new_ptr_51_value ? ghv_134 : _GEN_8356; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8358 = 8'h87 == new_ptr_51_value ? ghv_135 : _GEN_8357; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8359 = 8'h88 == new_ptr_51_value ? ghv_136 : _GEN_8358; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8360 = 8'h89 == new_ptr_51_value ? ghv_137 : _GEN_8359; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8361 = 8'h8a == new_ptr_51_value ? ghv_138 : _GEN_8360; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8362 = 8'h8b == new_ptr_51_value ? ghv_139 : _GEN_8361; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8363 = 8'h8c == new_ptr_51_value ? ghv_140 : _GEN_8362; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8364 = 8'h8d == new_ptr_51_value ? ghv_141 : _GEN_8363; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8365 = 8'h8e == new_ptr_51_value ? ghv_142 : _GEN_8364; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_47_value = _new_ptr_value_T_95[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_8368 = 8'h1 == new_ptr_47_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8369 = 8'h2 == new_ptr_47_value ? ghv_2 : _GEN_8368; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8370 = 8'h3 == new_ptr_47_value ? ghv_3 : _GEN_8369; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8371 = 8'h4 == new_ptr_47_value ? ghv_4 : _GEN_8370; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8372 = 8'h5 == new_ptr_47_value ? ghv_5 : _GEN_8371; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8373 = 8'h6 == new_ptr_47_value ? ghv_6 : _GEN_8372; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8374 = 8'h7 == new_ptr_47_value ? ghv_7 : _GEN_8373; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8375 = 8'h8 == new_ptr_47_value ? ghv_8 : _GEN_8374; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8376 = 8'h9 == new_ptr_47_value ? ghv_9 : _GEN_8375; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8377 = 8'ha == new_ptr_47_value ? ghv_10 : _GEN_8376; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8378 = 8'hb == new_ptr_47_value ? ghv_11 : _GEN_8377; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8379 = 8'hc == new_ptr_47_value ? ghv_12 : _GEN_8378; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8380 = 8'hd == new_ptr_47_value ? ghv_13 : _GEN_8379; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8381 = 8'he == new_ptr_47_value ? ghv_14 : _GEN_8380; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8382 = 8'hf == new_ptr_47_value ? ghv_15 : _GEN_8381; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8383 = 8'h10 == new_ptr_47_value ? ghv_16 : _GEN_8382; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8384 = 8'h11 == new_ptr_47_value ? ghv_17 : _GEN_8383; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8385 = 8'h12 == new_ptr_47_value ? ghv_18 : _GEN_8384; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8386 = 8'h13 == new_ptr_47_value ? ghv_19 : _GEN_8385; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8387 = 8'h14 == new_ptr_47_value ? ghv_20 : _GEN_8386; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8388 = 8'h15 == new_ptr_47_value ? ghv_21 : _GEN_8387; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8389 = 8'h16 == new_ptr_47_value ? ghv_22 : _GEN_8388; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8390 = 8'h17 == new_ptr_47_value ? ghv_23 : _GEN_8389; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8391 = 8'h18 == new_ptr_47_value ? ghv_24 : _GEN_8390; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8392 = 8'h19 == new_ptr_47_value ? ghv_25 : _GEN_8391; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8393 = 8'h1a == new_ptr_47_value ? ghv_26 : _GEN_8392; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8394 = 8'h1b == new_ptr_47_value ? ghv_27 : _GEN_8393; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8395 = 8'h1c == new_ptr_47_value ? ghv_28 : _GEN_8394; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8396 = 8'h1d == new_ptr_47_value ? ghv_29 : _GEN_8395; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8397 = 8'h1e == new_ptr_47_value ? ghv_30 : _GEN_8396; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8398 = 8'h1f == new_ptr_47_value ? ghv_31 : _GEN_8397; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8399 = 8'h20 == new_ptr_47_value ? ghv_32 : _GEN_8398; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8400 = 8'h21 == new_ptr_47_value ? ghv_33 : _GEN_8399; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8401 = 8'h22 == new_ptr_47_value ? ghv_34 : _GEN_8400; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8402 = 8'h23 == new_ptr_47_value ? ghv_35 : _GEN_8401; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8403 = 8'h24 == new_ptr_47_value ? ghv_36 : _GEN_8402; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8404 = 8'h25 == new_ptr_47_value ? ghv_37 : _GEN_8403; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8405 = 8'h26 == new_ptr_47_value ? ghv_38 : _GEN_8404; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8406 = 8'h27 == new_ptr_47_value ? ghv_39 : _GEN_8405; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8407 = 8'h28 == new_ptr_47_value ? ghv_40 : _GEN_8406; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8408 = 8'h29 == new_ptr_47_value ? ghv_41 : _GEN_8407; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8409 = 8'h2a == new_ptr_47_value ? ghv_42 : _GEN_8408; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8410 = 8'h2b == new_ptr_47_value ? ghv_43 : _GEN_8409; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8411 = 8'h2c == new_ptr_47_value ? ghv_44 : _GEN_8410; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8412 = 8'h2d == new_ptr_47_value ? ghv_45 : _GEN_8411; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8413 = 8'h2e == new_ptr_47_value ? ghv_46 : _GEN_8412; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8414 = 8'h2f == new_ptr_47_value ? ghv_47 : _GEN_8413; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8415 = 8'h30 == new_ptr_47_value ? ghv_48 : _GEN_8414; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8416 = 8'h31 == new_ptr_47_value ? ghv_49 : _GEN_8415; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8417 = 8'h32 == new_ptr_47_value ? ghv_50 : _GEN_8416; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8418 = 8'h33 == new_ptr_47_value ? ghv_51 : _GEN_8417; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8419 = 8'h34 == new_ptr_47_value ? ghv_52 : _GEN_8418; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8420 = 8'h35 == new_ptr_47_value ? ghv_53 : _GEN_8419; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8421 = 8'h36 == new_ptr_47_value ? ghv_54 : _GEN_8420; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8422 = 8'h37 == new_ptr_47_value ? ghv_55 : _GEN_8421; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8423 = 8'h38 == new_ptr_47_value ? ghv_56 : _GEN_8422; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8424 = 8'h39 == new_ptr_47_value ? ghv_57 : _GEN_8423; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8425 = 8'h3a == new_ptr_47_value ? ghv_58 : _GEN_8424; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8426 = 8'h3b == new_ptr_47_value ? ghv_59 : _GEN_8425; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8427 = 8'h3c == new_ptr_47_value ? ghv_60 : _GEN_8426; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8428 = 8'h3d == new_ptr_47_value ? ghv_61 : _GEN_8427; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8429 = 8'h3e == new_ptr_47_value ? ghv_62 : _GEN_8428; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8430 = 8'h3f == new_ptr_47_value ? ghv_63 : _GEN_8429; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8431 = 8'h40 == new_ptr_47_value ? ghv_64 : _GEN_8430; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8432 = 8'h41 == new_ptr_47_value ? ghv_65 : _GEN_8431; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8433 = 8'h42 == new_ptr_47_value ? ghv_66 : _GEN_8432; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8434 = 8'h43 == new_ptr_47_value ? ghv_67 : _GEN_8433; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8435 = 8'h44 == new_ptr_47_value ? ghv_68 : _GEN_8434; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8436 = 8'h45 == new_ptr_47_value ? ghv_69 : _GEN_8435; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8437 = 8'h46 == new_ptr_47_value ? ghv_70 : _GEN_8436; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8438 = 8'h47 == new_ptr_47_value ? ghv_71 : _GEN_8437; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8439 = 8'h48 == new_ptr_47_value ? ghv_72 : _GEN_8438; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8440 = 8'h49 == new_ptr_47_value ? ghv_73 : _GEN_8439; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8441 = 8'h4a == new_ptr_47_value ? ghv_74 : _GEN_8440; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8442 = 8'h4b == new_ptr_47_value ? ghv_75 : _GEN_8441; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8443 = 8'h4c == new_ptr_47_value ? ghv_76 : _GEN_8442; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8444 = 8'h4d == new_ptr_47_value ? ghv_77 : _GEN_8443; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8445 = 8'h4e == new_ptr_47_value ? ghv_78 : _GEN_8444; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8446 = 8'h4f == new_ptr_47_value ? ghv_79 : _GEN_8445; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8447 = 8'h50 == new_ptr_47_value ? ghv_80 : _GEN_8446; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8448 = 8'h51 == new_ptr_47_value ? ghv_81 : _GEN_8447; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8449 = 8'h52 == new_ptr_47_value ? ghv_82 : _GEN_8448; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8450 = 8'h53 == new_ptr_47_value ? ghv_83 : _GEN_8449; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8451 = 8'h54 == new_ptr_47_value ? ghv_84 : _GEN_8450; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8452 = 8'h55 == new_ptr_47_value ? ghv_85 : _GEN_8451; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8453 = 8'h56 == new_ptr_47_value ? ghv_86 : _GEN_8452; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8454 = 8'h57 == new_ptr_47_value ? ghv_87 : _GEN_8453; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8455 = 8'h58 == new_ptr_47_value ? ghv_88 : _GEN_8454; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8456 = 8'h59 == new_ptr_47_value ? ghv_89 : _GEN_8455; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8457 = 8'h5a == new_ptr_47_value ? ghv_90 : _GEN_8456; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8458 = 8'h5b == new_ptr_47_value ? ghv_91 : _GEN_8457; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8459 = 8'h5c == new_ptr_47_value ? ghv_92 : _GEN_8458; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8460 = 8'h5d == new_ptr_47_value ? ghv_93 : _GEN_8459; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8461 = 8'h5e == new_ptr_47_value ? ghv_94 : _GEN_8460; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8462 = 8'h5f == new_ptr_47_value ? ghv_95 : _GEN_8461; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8463 = 8'h60 == new_ptr_47_value ? ghv_96 : _GEN_8462; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8464 = 8'h61 == new_ptr_47_value ? ghv_97 : _GEN_8463; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8465 = 8'h62 == new_ptr_47_value ? ghv_98 : _GEN_8464; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8466 = 8'h63 == new_ptr_47_value ? ghv_99 : _GEN_8465; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8467 = 8'h64 == new_ptr_47_value ? ghv_100 : _GEN_8466; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8468 = 8'h65 == new_ptr_47_value ? ghv_101 : _GEN_8467; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8469 = 8'h66 == new_ptr_47_value ? ghv_102 : _GEN_8468; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8470 = 8'h67 == new_ptr_47_value ? ghv_103 : _GEN_8469; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8471 = 8'h68 == new_ptr_47_value ? ghv_104 : _GEN_8470; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8472 = 8'h69 == new_ptr_47_value ? ghv_105 : _GEN_8471; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8473 = 8'h6a == new_ptr_47_value ? ghv_106 : _GEN_8472; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8474 = 8'h6b == new_ptr_47_value ? ghv_107 : _GEN_8473; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8475 = 8'h6c == new_ptr_47_value ? ghv_108 : _GEN_8474; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8476 = 8'h6d == new_ptr_47_value ? ghv_109 : _GEN_8475; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8477 = 8'h6e == new_ptr_47_value ? ghv_110 : _GEN_8476; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8478 = 8'h6f == new_ptr_47_value ? ghv_111 : _GEN_8477; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8479 = 8'h70 == new_ptr_47_value ? ghv_112 : _GEN_8478; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8480 = 8'h71 == new_ptr_47_value ? ghv_113 : _GEN_8479; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8481 = 8'h72 == new_ptr_47_value ? ghv_114 : _GEN_8480; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8482 = 8'h73 == new_ptr_47_value ? ghv_115 : _GEN_8481; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8483 = 8'h74 == new_ptr_47_value ? ghv_116 : _GEN_8482; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8484 = 8'h75 == new_ptr_47_value ? ghv_117 : _GEN_8483; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8485 = 8'h76 == new_ptr_47_value ? ghv_118 : _GEN_8484; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8486 = 8'h77 == new_ptr_47_value ? ghv_119 : _GEN_8485; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8487 = 8'h78 == new_ptr_47_value ? ghv_120 : _GEN_8486; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8488 = 8'h79 == new_ptr_47_value ? ghv_121 : _GEN_8487; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8489 = 8'h7a == new_ptr_47_value ? ghv_122 : _GEN_8488; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8490 = 8'h7b == new_ptr_47_value ? ghv_123 : _GEN_8489; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8491 = 8'h7c == new_ptr_47_value ? ghv_124 : _GEN_8490; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8492 = 8'h7d == new_ptr_47_value ? ghv_125 : _GEN_8491; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8493 = 8'h7e == new_ptr_47_value ? ghv_126 : _GEN_8492; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8494 = 8'h7f == new_ptr_47_value ? ghv_127 : _GEN_8493; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8495 = 8'h80 == new_ptr_47_value ? ghv_128 : _GEN_8494; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8496 = 8'h81 == new_ptr_47_value ? ghv_129 : _GEN_8495; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8497 = 8'h82 == new_ptr_47_value ? ghv_130 : _GEN_8496; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8498 = 8'h83 == new_ptr_47_value ? ghv_131 : _GEN_8497; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8499 = 8'h84 == new_ptr_47_value ? ghv_132 : _GEN_8498; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8500 = 8'h85 == new_ptr_47_value ? ghv_133 : _GEN_8499; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8501 = 8'h86 == new_ptr_47_value ? ghv_134 : _GEN_8500; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8502 = 8'h87 == new_ptr_47_value ? ghv_135 : _GEN_8501; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8503 = 8'h88 == new_ptr_47_value ? ghv_136 : _GEN_8502; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8504 = 8'h89 == new_ptr_47_value ? ghv_137 : _GEN_8503; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8505 = 8'h8a == new_ptr_47_value ? ghv_138 : _GEN_8504; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8506 = 8'h8b == new_ptr_47_value ? ghv_139 : _GEN_8505; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8507 = 8'h8c == new_ptr_47_value ? ghv_140 : _GEN_8506; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8508 = 8'h8d == new_ptr_47_value ? ghv_141 : _GEN_8507; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8509 = 8'h8e == new_ptr_47_value ? ghv_142 : _GEN_8508; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_45_value = _new_ptr_value_T_91[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_8512 = 8'h1 == new_ptr_45_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8513 = 8'h2 == new_ptr_45_value ? ghv_2 : _GEN_8512; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8514 = 8'h3 == new_ptr_45_value ? ghv_3 : _GEN_8513; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8515 = 8'h4 == new_ptr_45_value ? ghv_4 : _GEN_8514; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8516 = 8'h5 == new_ptr_45_value ? ghv_5 : _GEN_8515; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8517 = 8'h6 == new_ptr_45_value ? ghv_6 : _GEN_8516; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8518 = 8'h7 == new_ptr_45_value ? ghv_7 : _GEN_8517; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8519 = 8'h8 == new_ptr_45_value ? ghv_8 : _GEN_8518; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8520 = 8'h9 == new_ptr_45_value ? ghv_9 : _GEN_8519; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8521 = 8'ha == new_ptr_45_value ? ghv_10 : _GEN_8520; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8522 = 8'hb == new_ptr_45_value ? ghv_11 : _GEN_8521; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8523 = 8'hc == new_ptr_45_value ? ghv_12 : _GEN_8522; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8524 = 8'hd == new_ptr_45_value ? ghv_13 : _GEN_8523; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8525 = 8'he == new_ptr_45_value ? ghv_14 : _GEN_8524; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8526 = 8'hf == new_ptr_45_value ? ghv_15 : _GEN_8525; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8527 = 8'h10 == new_ptr_45_value ? ghv_16 : _GEN_8526; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8528 = 8'h11 == new_ptr_45_value ? ghv_17 : _GEN_8527; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8529 = 8'h12 == new_ptr_45_value ? ghv_18 : _GEN_8528; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8530 = 8'h13 == new_ptr_45_value ? ghv_19 : _GEN_8529; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8531 = 8'h14 == new_ptr_45_value ? ghv_20 : _GEN_8530; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8532 = 8'h15 == new_ptr_45_value ? ghv_21 : _GEN_8531; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8533 = 8'h16 == new_ptr_45_value ? ghv_22 : _GEN_8532; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8534 = 8'h17 == new_ptr_45_value ? ghv_23 : _GEN_8533; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8535 = 8'h18 == new_ptr_45_value ? ghv_24 : _GEN_8534; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8536 = 8'h19 == new_ptr_45_value ? ghv_25 : _GEN_8535; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8537 = 8'h1a == new_ptr_45_value ? ghv_26 : _GEN_8536; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8538 = 8'h1b == new_ptr_45_value ? ghv_27 : _GEN_8537; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8539 = 8'h1c == new_ptr_45_value ? ghv_28 : _GEN_8538; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8540 = 8'h1d == new_ptr_45_value ? ghv_29 : _GEN_8539; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8541 = 8'h1e == new_ptr_45_value ? ghv_30 : _GEN_8540; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8542 = 8'h1f == new_ptr_45_value ? ghv_31 : _GEN_8541; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8543 = 8'h20 == new_ptr_45_value ? ghv_32 : _GEN_8542; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8544 = 8'h21 == new_ptr_45_value ? ghv_33 : _GEN_8543; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8545 = 8'h22 == new_ptr_45_value ? ghv_34 : _GEN_8544; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8546 = 8'h23 == new_ptr_45_value ? ghv_35 : _GEN_8545; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8547 = 8'h24 == new_ptr_45_value ? ghv_36 : _GEN_8546; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8548 = 8'h25 == new_ptr_45_value ? ghv_37 : _GEN_8547; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8549 = 8'h26 == new_ptr_45_value ? ghv_38 : _GEN_8548; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8550 = 8'h27 == new_ptr_45_value ? ghv_39 : _GEN_8549; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8551 = 8'h28 == new_ptr_45_value ? ghv_40 : _GEN_8550; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8552 = 8'h29 == new_ptr_45_value ? ghv_41 : _GEN_8551; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8553 = 8'h2a == new_ptr_45_value ? ghv_42 : _GEN_8552; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8554 = 8'h2b == new_ptr_45_value ? ghv_43 : _GEN_8553; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8555 = 8'h2c == new_ptr_45_value ? ghv_44 : _GEN_8554; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8556 = 8'h2d == new_ptr_45_value ? ghv_45 : _GEN_8555; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8557 = 8'h2e == new_ptr_45_value ? ghv_46 : _GEN_8556; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8558 = 8'h2f == new_ptr_45_value ? ghv_47 : _GEN_8557; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8559 = 8'h30 == new_ptr_45_value ? ghv_48 : _GEN_8558; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8560 = 8'h31 == new_ptr_45_value ? ghv_49 : _GEN_8559; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8561 = 8'h32 == new_ptr_45_value ? ghv_50 : _GEN_8560; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8562 = 8'h33 == new_ptr_45_value ? ghv_51 : _GEN_8561; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8563 = 8'h34 == new_ptr_45_value ? ghv_52 : _GEN_8562; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8564 = 8'h35 == new_ptr_45_value ? ghv_53 : _GEN_8563; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8565 = 8'h36 == new_ptr_45_value ? ghv_54 : _GEN_8564; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8566 = 8'h37 == new_ptr_45_value ? ghv_55 : _GEN_8565; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8567 = 8'h38 == new_ptr_45_value ? ghv_56 : _GEN_8566; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8568 = 8'h39 == new_ptr_45_value ? ghv_57 : _GEN_8567; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8569 = 8'h3a == new_ptr_45_value ? ghv_58 : _GEN_8568; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8570 = 8'h3b == new_ptr_45_value ? ghv_59 : _GEN_8569; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8571 = 8'h3c == new_ptr_45_value ? ghv_60 : _GEN_8570; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8572 = 8'h3d == new_ptr_45_value ? ghv_61 : _GEN_8571; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8573 = 8'h3e == new_ptr_45_value ? ghv_62 : _GEN_8572; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8574 = 8'h3f == new_ptr_45_value ? ghv_63 : _GEN_8573; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8575 = 8'h40 == new_ptr_45_value ? ghv_64 : _GEN_8574; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8576 = 8'h41 == new_ptr_45_value ? ghv_65 : _GEN_8575; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8577 = 8'h42 == new_ptr_45_value ? ghv_66 : _GEN_8576; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8578 = 8'h43 == new_ptr_45_value ? ghv_67 : _GEN_8577; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8579 = 8'h44 == new_ptr_45_value ? ghv_68 : _GEN_8578; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8580 = 8'h45 == new_ptr_45_value ? ghv_69 : _GEN_8579; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8581 = 8'h46 == new_ptr_45_value ? ghv_70 : _GEN_8580; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8582 = 8'h47 == new_ptr_45_value ? ghv_71 : _GEN_8581; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8583 = 8'h48 == new_ptr_45_value ? ghv_72 : _GEN_8582; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8584 = 8'h49 == new_ptr_45_value ? ghv_73 : _GEN_8583; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8585 = 8'h4a == new_ptr_45_value ? ghv_74 : _GEN_8584; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8586 = 8'h4b == new_ptr_45_value ? ghv_75 : _GEN_8585; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8587 = 8'h4c == new_ptr_45_value ? ghv_76 : _GEN_8586; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8588 = 8'h4d == new_ptr_45_value ? ghv_77 : _GEN_8587; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8589 = 8'h4e == new_ptr_45_value ? ghv_78 : _GEN_8588; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8590 = 8'h4f == new_ptr_45_value ? ghv_79 : _GEN_8589; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8591 = 8'h50 == new_ptr_45_value ? ghv_80 : _GEN_8590; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8592 = 8'h51 == new_ptr_45_value ? ghv_81 : _GEN_8591; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8593 = 8'h52 == new_ptr_45_value ? ghv_82 : _GEN_8592; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8594 = 8'h53 == new_ptr_45_value ? ghv_83 : _GEN_8593; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8595 = 8'h54 == new_ptr_45_value ? ghv_84 : _GEN_8594; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8596 = 8'h55 == new_ptr_45_value ? ghv_85 : _GEN_8595; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8597 = 8'h56 == new_ptr_45_value ? ghv_86 : _GEN_8596; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8598 = 8'h57 == new_ptr_45_value ? ghv_87 : _GEN_8597; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8599 = 8'h58 == new_ptr_45_value ? ghv_88 : _GEN_8598; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8600 = 8'h59 == new_ptr_45_value ? ghv_89 : _GEN_8599; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8601 = 8'h5a == new_ptr_45_value ? ghv_90 : _GEN_8600; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8602 = 8'h5b == new_ptr_45_value ? ghv_91 : _GEN_8601; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8603 = 8'h5c == new_ptr_45_value ? ghv_92 : _GEN_8602; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8604 = 8'h5d == new_ptr_45_value ? ghv_93 : _GEN_8603; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8605 = 8'h5e == new_ptr_45_value ? ghv_94 : _GEN_8604; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8606 = 8'h5f == new_ptr_45_value ? ghv_95 : _GEN_8605; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8607 = 8'h60 == new_ptr_45_value ? ghv_96 : _GEN_8606; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8608 = 8'h61 == new_ptr_45_value ? ghv_97 : _GEN_8607; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8609 = 8'h62 == new_ptr_45_value ? ghv_98 : _GEN_8608; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8610 = 8'h63 == new_ptr_45_value ? ghv_99 : _GEN_8609; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8611 = 8'h64 == new_ptr_45_value ? ghv_100 : _GEN_8610; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8612 = 8'h65 == new_ptr_45_value ? ghv_101 : _GEN_8611; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8613 = 8'h66 == new_ptr_45_value ? ghv_102 : _GEN_8612; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8614 = 8'h67 == new_ptr_45_value ? ghv_103 : _GEN_8613; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8615 = 8'h68 == new_ptr_45_value ? ghv_104 : _GEN_8614; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8616 = 8'h69 == new_ptr_45_value ? ghv_105 : _GEN_8615; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8617 = 8'h6a == new_ptr_45_value ? ghv_106 : _GEN_8616; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8618 = 8'h6b == new_ptr_45_value ? ghv_107 : _GEN_8617; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8619 = 8'h6c == new_ptr_45_value ? ghv_108 : _GEN_8618; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8620 = 8'h6d == new_ptr_45_value ? ghv_109 : _GEN_8619; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8621 = 8'h6e == new_ptr_45_value ? ghv_110 : _GEN_8620; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8622 = 8'h6f == new_ptr_45_value ? ghv_111 : _GEN_8621; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8623 = 8'h70 == new_ptr_45_value ? ghv_112 : _GEN_8622; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8624 = 8'h71 == new_ptr_45_value ? ghv_113 : _GEN_8623; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8625 = 8'h72 == new_ptr_45_value ? ghv_114 : _GEN_8624; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8626 = 8'h73 == new_ptr_45_value ? ghv_115 : _GEN_8625; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8627 = 8'h74 == new_ptr_45_value ? ghv_116 : _GEN_8626; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8628 = 8'h75 == new_ptr_45_value ? ghv_117 : _GEN_8627; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8629 = 8'h76 == new_ptr_45_value ? ghv_118 : _GEN_8628; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8630 = 8'h77 == new_ptr_45_value ? ghv_119 : _GEN_8629; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8631 = 8'h78 == new_ptr_45_value ? ghv_120 : _GEN_8630; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8632 = 8'h79 == new_ptr_45_value ? ghv_121 : _GEN_8631; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8633 = 8'h7a == new_ptr_45_value ? ghv_122 : _GEN_8632; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8634 = 8'h7b == new_ptr_45_value ? ghv_123 : _GEN_8633; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8635 = 8'h7c == new_ptr_45_value ? ghv_124 : _GEN_8634; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8636 = 8'h7d == new_ptr_45_value ? ghv_125 : _GEN_8635; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8637 = 8'h7e == new_ptr_45_value ? ghv_126 : _GEN_8636; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8638 = 8'h7f == new_ptr_45_value ? ghv_127 : _GEN_8637; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8639 = 8'h80 == new_ptr_45_value ? ghv_128 : _GEN_8638; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8640 = 8'h81 == new_ptr_45_value ? ghv_129 : _GEN_8639; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8641 = 8'h82 == new_ptr_45_value ? ghv_130 : _GEN_8640; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8642 = 8'h83 == new_ptr_45_value ? ghv_131 : _GEN_8641; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8643 = 8'h84 == new_ptr_45_value ? ghv_132 : _GEN_8642; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8644 = 8'h85 == new_ptr_45_value ? ghv_133 : _GEN_8643; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8645 = 8'h86 == new_ptr_45_value ? ghv_134 : _GEN_8644; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8646 = 8'h87 == new_ptr_45_value ? ghv_135 : _GEN_8645; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8647 = 8'h88 == new_ptr_45_value ? ghv_136 : _GEN_8646; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8648 = 8'h89 == new_ptr_45_value ? ghv_137 : _GEN_8647; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8649 = 8'h8a == new_ptr_45_value ? ghv_138 : _GEN_8648; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8650 = 8'h8b == new_ptr_45_value ? ghv_139 : _GEN_8649; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8651 = 8'h8c == new_ptr_45_value ? ghv_140 : _GEN_8650; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8652 = 8'h8d == new_ptr_45_value ? ghv_141 : _GEN_8651; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8653 = 8'h8e == new_ptr_45_value ? ghv_142 : _GEN_8652; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_40_value = _new_ptr_value_T_81[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_8656 = 8'h1 == new_ptr_40_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8657 = 8'h2 == new_ptr_40_value ? ghv_2 : _GEN_8656; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8658 = 8'h3 == new_ptr_40_value ? ghv_3 : _GEN_8657; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8659 = 8'h4 == new_ptr_40_value ? ghv_4 : _GEN_8658; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8660 = 8'h5 == new_ptr_40_value ? ghv_5 : _GEN_8659; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8661 = 8'h6 == new_ptr_40_value ? ghv_6 : _GEN_8660; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8662 = 8'h7 == new_ptr_40_value ? ghv_7 : _GEN_8661; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8663 = 8'h8 == new_ptr_40_value ? ghv_8 : _GEN_8662; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8664 = 8'h9 == new_ptr_40_value ? ghv_9 : _GEN_8663; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8665 = 8'ha == new_ptr_40_value ? ghv_10 : _GEN_8664; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8666 = 8'hb == new_ptr_40_value ? ghv_11 : _GEN_8665; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8667 = 8'hc == new_ptr_40_value ? ghv_12 : _GEN_8666; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8668 = 8'hd == new_ptr_40_value ? ghv_13 : _GEN_8667; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8669 = 8'he == new_ptr_40_value ? ghv_14 : _GEN_8668; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8670 = 8'hf == new_ptr_40_value ? ghv_15 : _GEN_8669; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8671 = 8'h10 == new_ptr_40_value ? ghv_16 : _GEN_8670; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8672 = 8'h11 == new_ptr_40_value ? ghv_17 : _GEN_8671; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8673 = 8'h12 == new_ptr_40_value ? ghv_18 : _GEN_8672; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8674 = 8'h13 == new_ptr_40_value ? ghv_19 : _GEN_8673; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8675 = 8'h14 == new_ptr_40_value ? ghv_20 : _GEN_8674; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8676 = 8'h15 == new_ptr_40_value ? ghv_21 : _GEN_8675; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8677 = 8'h16 == new_ptr_40_value ? ghv_22 : _GEN_8676; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8678 = 8'h17 == new_ptr_40_value ? ghv_23 : _GEN_8677; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8679 = 8'h18 == new_ptr_40_value ? ghv_24 : _GEN_8678; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8680 = 8'h19 == new_ptr_40_value ? ghv_25 : _GEN_8679; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8681 = 8'h1a == new_ptr_40_value ? ghv_26 : _GEN_8680; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8682 = 8'h1b == new_ptr_40_value ? ghv_27 : _GEN_8681; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8683 = 8'h1c == new_ptr_40_value ? ghv_28 : _GEN_8682; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8684 = 8'h1d == new_ptr_40_value ? ghv_29 : _GEN_8683; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8685 = 8'h1e == new_ptr_40_value ? ghv_30 : _GEN_8684; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8686 = 8'h1f == new_ptr_40_value ? ghv_31 : _GEN_8685; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8687 = 8'h20 == new_ptr_40_value ? ghv_32 : _GEN_8686; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8688 = 8'h21 == new_ptr_40_value ? ghv_33 : _GEN_8687; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8689 = 8'h22 == new_ptr_40_value ? ghv_34 : _GEN_8688; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8690 = 8'h23 == new_ptr_40_value ? ghv_35 : _GEN_8689; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8691 = 8'h24 == new_ptr_40_value ? ghv_36 : _GEN_8690; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8692 = 8'h25 == new_ptr_40_value ? ghv_37 : _GEN_8691; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8693 = 8'h26 == new_ptr_40_value ? ghv_38 : _GEN_8692; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8694 = 8'h27 == new_ptr_40_value ? ghv_39 : _GEN_8693; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8695 = 8'h28 == new_ptr_40_value ? ghv_40 : _GEN_8694; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8696 = 8'h29 == new_ptr_40_value ? ghv_41 : _GEN_8695; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8697 = 8'h2a == new_ptr_40_value ? ghv_42 : _GEN_8696; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8698 = 8'h2b == new_ptr_40_value ? ghv_43 : _GEN_8697; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8699 = 8'h2c == new_ptr_40_value ? ghv_44 : _GEN_8698; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8700 = 8'h2d == new_ptr_40_value ? ghv_45 : _GEN_8699; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8701 = 8'h2e == new_ptr_40_value ? ghv_46 : _GEN_8700; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8702 = 8'h2f == new_ptr_40_value ? ghv_47 : _GEN_8701; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8703 = 8'h30 == new_ptr_40_value ? ghv_48 : _GEN_8702; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8704 = 8'h31 == new_ptr_40_value ? ghv_49 : _GEN_8703; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8705 = 8'h32 == new_ptr_40_value ? ghv_50 : _GEN_8704; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8706 = 8'h33 == new_ptr_40_value ? ghv_51 : _GEN_8705; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8707 = 8'h34 == new_ptr_40_value ? ghv_52 : _GEN_8706; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8708 = 8'h35 == new_ptr_40_value ? ghv_53 : _GEN_8707; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8709 = 8'h36 == new_ptr_40_value ? ghv_54 : _GEN_8708; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8710 = 8'h37 == new_ptr_40_value ? ghv_55 : _GEN_8709; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8711 = 8'h38 == new_ptr_40_value ? ghv_56 : _GEN_8710; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8712 = 8'h39 == new_ptr_40_value ? ghv_57 : _GEN_8711; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8713 = 8'h3a == new_ptr_40_value ? ghv_58 : _GEN_8712; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8714 = 8'h3b == new_ptr_40_value ? ghv_59 : _GEN_8713; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8715 = 8'h3c == new_ptr_40_value ? ghv_60 : _GEN_8714; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8716 = 8'h3d == new_ptr_40_value ? ghv_61 : _GEN_8715; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8717 = 8'h3e == new_ptr_40_value ? ghv_62 : _GEN_8716; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8718 = 8'h3f == new_ptr_40_value ? ghv_63 : _GEN_8717; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8719 = 8'h40 == new_ptr_40_value ? ghv_64 : _GEN_8718; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8720 = 8'h41 == new_ptr_40_value ? ghv_65 : _GEN_8719; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8721 = 8'h42 == new_ptr_40_value ? ghv_66 : _GEN_8720; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8722 = 8'h43 == new_ptr_40_value ? ghv_67 : _GEN_8721; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8723 = 8'h44 == new_ptr_40_value ? ghv_68 : _GEN_8722; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8724 = 8'h45 == new_ptr_40_value ? ghv_69 : _GEN_8723; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8725 = 8'h46 == new_ptr_40_value ? ghv_70 : _GEN_8724; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8726 = 8'h47 == new_ptr_40_value ? ghv_71 : _GEN_8725; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8727 = 8'h48 == new_ptr_40_value ? ghv_72 : _GEN_8726; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8728 = 8'h49 == new_ptr_40_value ? ghv_73 : _GEN_8727; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8729 = 8'h4a == new_ptr_40_value ? ghv_74 : _GEN_8728; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8730 = 8'h4b == new_ptr_40_value ? ghv_75 : _GEN_8729; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8731 = 8'h4c == new_ptr_40_value ? ghv_76 : _GEN_8730; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8732 = 8'h4d == new_ptr_40_value ? ghv_77 : _GEN_8731; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8733 = 8'h4e == new_ptr_40_value ? ghv_78 : _GEN_8732; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8734 = 8'h4f == new_ptr_40_value ? ghv_79 : _GEN_8733; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8735 = 8'h50 == new_ptr_40_value ? ghv_80 : _GEN_8734; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8736 = 8'h51 == new_ptr_40_value ? ghv_81 : _GEN_8735; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8737 = 8'h52 == new_ptr_40_value ? ghv_82 : _GEN_8736; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8738 = 8'h53 == new_ptr_40_value ? ghv_83 : _GEN_8737; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8739 = 8'h54 == new_ptr_40_value ? ghv_84 : _GEN_8738; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8740 = 8'h55 == new_ptr_40_value ? ghv_85 : _GEN_8739; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8741 = 8'h56 == new_ptr_40_value ? ghv_86 : _GEN_8740; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8742 = 8'h57 == new_ptr_40_value ? ghv_87 : _GEN_8741; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8743 = 8'h58 == new_ptr_40_value ? ghv_88 : _GEN_8742; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8744 = 8'h59 == new_ptr_40_value ? ghv_89 : _GEN_8743; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8745 = 8'h5a == new_ptr_40_value ? ghv_90 : _GEN_8744; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8746 = 8'h5b == new_ptr_40_value ? ghv_91 : _GEN_8745; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8747 = 8'h5c == new_ptr_40_value ? ghv_92 : _GEN_8746; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8748 = 8'h5d == new_ptr_40_value ? ghv_93 : _GEN_8747; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8749 = 8'h5e == new_ptr_40_value ? ghv_94 : _GEN_8748; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8750 = 8'h5f == new_ptr_40_value ? ghv_95 : _GEN_8749; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8751 = 8'h60 == new_ptr_40_value ? ghv_96 : _GEN_8750; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8752 = 8'h61 == new_ptr_40_value ? ghv_97 : _GEN_8751; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8753 = 8'h62 == new_ptr_40_value ? ghv_98 : _GEN_8752; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8754 = 8'h63 == new_ptr_40_value ? ghv_99 : _GEN_8753; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8755 = 8'h64 == new_ptr_40_value ? ghv_100 : _GEN_8754; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8756 = 8'h65 == new_ptr_40_value ? ghv_101 : _GEN_8755; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8757 = 8'h66 == new_ptr_40_value ? ghv_102 : _GEN_8756; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8758 = 8'h67 == new_ptr_40_value ? ghv_103 : _GEN_8757; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8759 = 8'h68 == new_ptr_40_value ? ghv_104 : _GEN_8758; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8760 = 8'h69 == new_ptr_40_value ? ghv_105 : _GEN_8759; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8761 = 8'h6a == new_ptr_40_value ? ghv_106 : _GEN_8760; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8762 = 8'h6b == new_ptr_40_value ? ghv_107 : _GEN_8761; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8763 = 8'h6c == new_ptr_40_value ? ghv_108 : _GEN_8762; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8764 = 8'h6d == new_ptr_40_value ? ghv_109 : _GEN_8763; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8765 = 8'h6e == new_ptr_40_value ? ghv_110 : _GEN_8764; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8766 = 8'h6f == new_ptr_40_value ? ghv_111 : _GEN_8765; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8767 = 8'h70 == new_ptr_40_value ? ghv_112 : _GEN_8766; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8768 = 8'h71 == new_ptr_40_value ? ghv_113 : _GEN_8767; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8769 = 8'h72 == new_ptr_40_value ? ghv_114 : _GEN_8768; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8770 = 8'h73 == new_ptr_40_value ? ghv_115 : _GEN_8769; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8771 = 8'h74 == new_ptr_40_value ? ghv_116 : _GEN_8770; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8772 = 8'h75 == new_ptr_40_value ? ghv_117 : _GEN_8771; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8773 = 8'h76 == new_ptr_40_value ? ghv_118 : _GEN_8772; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8774 = 8'h77 == new_ptr_40_value ? ghv_119 : _GEN_8773; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8775 = 8'h78 == new_ptr_40_value ? ghv_120 : _GEN_8774; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8776 = 8'h79 == new_ptr_40_value ? ghv_121 : _GEN_8775; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8777 = 8'h7a == new_ptr_40_value ? ghv_122 : _GEN_8776; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8778 = 8'h7b == new_ptr_40_value ? ghv_123 : _GEN_8777; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8779 = 8'h7c == new_ptr_40_value ? ghv_124 : _GEN_8778; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8780 = 8'h7d == new_ptr_40_value ? ghv_125 : _GEN_8779; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8781 = 8'h7e == new_ptr_40_value ? ghv_126 : _GEN_8780; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8782 = 8'h7f == new_ptr_40_value ? ghv_127 : _GEN_8781; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8783 = 8'h80 == new_ptr_40_value ? ghv_128 : _GEN_8782; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8784 = 8'h81 == new_ptr_40_value ? ghv_129 : _GEN_8783; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8785 = 8'h82 == new_ptr_40_value ? ghv_130 : _GEN_8784; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8786 = 8'h83 == new_ptr_40_value ? ghv_131 : _GEN_8785; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8787 = 8'h84 == new_ptr_40_value ? ghv_132 : _GEN_8786; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8788 = 8'h85 == new_ptr_40_value ? ghv_133 : _GEN_8787; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8789 = 8'h86 == new_ptr_40_value ? ghv_134 : _GEN_8788; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8790 = 8'h87 == new_ptr_40_value ? ghv_135 : _GEN_8789; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8791 = 8'h88 == new_ptr_40_value ? ghv_136 : _GEN_8790; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8792 = 8'h89 == new_ptr_40_value ? ghv_137 : _GEN_8791; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8793 = 8'h8a == new_ptr_40_value ? ghv_138 : _GEN_8792; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8794 = 8'h8b == new_ptr_40_value ? ghv_139 : _GEN_8793; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8795 = 8'h8c == new_ptr_40_value ? ghv_140 : _GEN_8794; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8796 = 8'h8d == new_ptr_40_value ? ghv_141 : _GEN_8795; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8797 = 8'h8e == new_ptr_40_value ? ghv_142 : _GEN_8796; // @[FrontendBundle.scala 329:{20,20}]
  wire  _s3_ghv_wens_T_26 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_0_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_53 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_1_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_0_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_1_value & _s3_predicted_ghist_ptr_T_45 & s3_redirect
    ; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_80 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_1_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_1_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_1_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_107 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_3_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_1_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_3_value & _s3_predicted_ghist_ptr_T_45 & s3_redirect
    ; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_134 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_3_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_2_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_3_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_161 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_5_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_2_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_5_value & _s3_predicted_ghist_ptr_T_45 & s3_redirect
    ; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_188 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_5_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_3_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_5_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_215 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_7_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_3_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_7_value & _s3_predicted_ghist_ptr_T_45 & s3_redirect
    ; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_242 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_7_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_4_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_7_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_269 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_9_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_4_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_9_value & _s3_predicted_ghist_ptr_T_45 & s3_redirect
    ; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_296 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_9_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_5_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_9_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_323 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_11_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_5_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_11_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_350 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_11_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_6_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_11_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_377 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_13_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_6_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_13_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_404 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_13_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_7_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_13_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_431 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_15_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_7_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_15_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_458 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_15_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_8_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_15_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_485 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_17_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_8_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_17_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_512 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_17_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_9_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_17_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_539 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_19_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_9_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_19_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_566 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_19_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_10_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_19_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_593 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_21_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_10_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_21_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_620 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_21_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_11_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_21_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_647 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_23_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_11_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_23_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_674 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_23_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_12_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_23_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_701 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_25_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_12_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_25_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_728 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_25_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_13_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_25_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_755 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_27_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_13_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_27_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_782 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_27_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_14_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_27_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_809 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_29_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_14_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_29_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_836 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_29_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_15_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_29_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_863 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_31_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_15_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_31_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_890 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_31_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_16_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_31_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_917 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_33_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_16_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_33_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_944 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_33_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_17_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_33_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_971 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_35_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_17_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_35_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_998 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_35_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_18_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_35_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_1025 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_37_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_18_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_37_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_1052 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_37_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_19_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_37_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_1079 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_39_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_19_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_39_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_1106 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_39_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_20_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_39_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_1133 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_41_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_20_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_41_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_1160 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_41_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_21_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_41_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_1187 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_43_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_21_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_43_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_1214 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_43_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_22_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_43_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_1241 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_45_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_22_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_45_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_1268 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_45_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_23_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_45_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_1295 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_47_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_23_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_47_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_1322 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_47_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_24_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_47_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_1349 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_49_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_24_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_49_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_1376 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_49_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_25_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_49_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_1403 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_51_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_25_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_51_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_1430 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_51_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_26_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_51_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_1457 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_53_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_26_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_53_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_1484 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_53_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_27_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_53_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_1511 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_55_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_27_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_55_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_1538 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_55_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_28_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_55_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_1565 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_57_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_28_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_57_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_1592 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_57_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_29_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_57_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_1619 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_59_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_29_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_59_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_1646 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_59_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_30_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_59_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_1673 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_61_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_30_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_61_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_1700 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_61_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_31_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_61_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_1727 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_63_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_31_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_63_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_1754 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_63_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_32_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_63_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_1781 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_65_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_32_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_65_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_1808 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_65_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_33_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_65_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_1835 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_67_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_33_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_67_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_1862 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_67_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_34_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_67_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_1889 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_69_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_34_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_69_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_1916 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_69_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_35_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_69_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_1943 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_71_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_35_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_71_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_1970 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_71_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_36_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_71_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_1997 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_73_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_36_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_73_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_2024 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_73_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_37_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_73_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_2051 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_75_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_37_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_75_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_2078 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_75_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_38_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_75_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_2105 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_77_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_38_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_77_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_2132 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_77_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_39_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_77_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_2159 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_79_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_39_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_79_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_2186 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_79_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_40_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_79_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_2213 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_81_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_40_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_81_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_2240 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_81_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_41_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_81_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_2267 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_83_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_41_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_83_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_2294 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_83_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_42_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_83_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_2321 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_85_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_42_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_85_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_2348 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_85_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_43_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_85_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_2375 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_87_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_43_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_87_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_2402 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_87_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_44_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_87_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_2429 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_89_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_44_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_89_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_2456 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_89_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_45_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_89_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_2483 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_91_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_45_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_91_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_2510 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_91_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_46_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_91_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_2537 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_93_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_46_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_93_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_2564 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_93_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_47_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_93_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_2591 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_95_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_47_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_95_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_2618 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_95_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_48_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_95_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_2645 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_97_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_48_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_97_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_2672 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_97_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_49_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_97_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_2699 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_99_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_49_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_99_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_2726 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_99_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_50_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_99_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_2753 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_101_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_50_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_101_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_2780 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_101_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_51_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_101_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_2807 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_103_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_51_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_103_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_2834 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_103_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_52_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_103_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_2861 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_105_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_52_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_105_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_2888 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_105_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_53_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_105_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_2915 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_107_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_53_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_107_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_2942 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_107_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_54_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_107_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_2969 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_109_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_54_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_109_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_2996 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_109_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_55_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_109_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_3023 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_111_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_55_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_111_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_3050 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_111_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_56_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_111_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_3077 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_113_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_56_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_113_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_3104 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_113_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_57_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_113_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_3131 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_115_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_57_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_115_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_3158 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_115_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_58_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_115_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_3185 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_117_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_58_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_117_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_3212 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_117_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_59_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_117_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_3239 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_119_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_59_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_119_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_3266 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_119_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_60_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_119_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_3293 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_121_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_60_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_121_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_3320 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_121_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_61_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_121_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_3347 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_123_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_61_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_123_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_3374 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_123_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_62_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_123_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_3401 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_125_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_62_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_125_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_3428 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_125_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_63_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_125_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_3455 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_127_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_63_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_127_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_3482 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_127_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_64_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_127_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_3509 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_129_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_64_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_129_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_3536 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_129_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_65_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_129_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_3563 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_131_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_65_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_131_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_3590 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_131_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_66_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_131_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_3617 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_133_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_66_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_133_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_3644 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_133_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_67_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_133_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_3671 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_135_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_67_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_135_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_3698 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_135_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_68_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_135_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_3725 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_137_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_68_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_137_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_3752 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_137_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_69_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_137_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_3779 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_139_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_69_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_139_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_3806 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_139_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_70_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_139_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_3833 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_141_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_70_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_141_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_3860 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_141_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_71_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_141_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_3887 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_143_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_71_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_143_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_3914 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_143_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_72_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_143_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_3941 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_145_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_72_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_145_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_3968 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_145_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_73_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_145_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_3995 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_147_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_73_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_147_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_4022 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_147_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_74_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_147_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_4049 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_149_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_74_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_149_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_4076 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_149_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_75_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_149_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_4103 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_151_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_75_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_151_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_4130 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_151_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_76_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_151_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_4157 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_153_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_76_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_153_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_4184 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_153_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_77_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_153_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_4211 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_155_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_77_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_155_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_4238 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_155_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_78_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_155_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_4265 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_157_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_78_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_157_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_4292 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_157_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_79_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_157_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_4319 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_159_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_79_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_159_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_4346 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_159_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_80_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_159_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_4373 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_161_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_80_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_161_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_4400 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_161_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_81_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_161_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_4427 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_163_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_81_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_163_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_4454 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_163_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_82_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_163_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_4481 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_165_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_82_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_165_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_4508 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_165_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_83_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_165_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_4535 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_167_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_83_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_167_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_4562 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_167_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_84_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_167_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_4589 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_169_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_84_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_169_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_4616 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_169_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_85_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_169_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_4643 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_171_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_85_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_171_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_4670 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_171_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_86_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_171_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_4697 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_173_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_86_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_173_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_4724 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_173_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_87_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_173_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_4751 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_175_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_87_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_175_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_4778 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_175_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_88_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_175_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_4805 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_177_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_88_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_177_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_4832 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_177_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_89_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_177_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_4859 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_179_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_89_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_179_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_4886 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_179_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_90_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_179_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_4913 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_181_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_90_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_181_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_4940 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_181_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_91_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_181_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_4967 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_183_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_91_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_183_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_4994 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_183_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_92_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_183_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_5021 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_185_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_92_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_185_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_5048 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_185_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_93_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_185_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_5075 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_187_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_93_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_187_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_5102 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_187_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_94_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_187_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_5129 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_189_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_94_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_189_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_5156 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_189_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_95_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_189_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_5183 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_191_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_95_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_191_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_5210 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_191_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_96_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_191_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_5237 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_193_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_96_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_193_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_5264 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_193_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_97_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_193_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_5291 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_195_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_97_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_195_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_5318 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_195_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_98_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_195_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_5345 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_197_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_98_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_197_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_5372 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_197_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_99_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_197_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_5399 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_199_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_99_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_199_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_5426 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_199_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_100_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_199_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_5453 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_201_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_100_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_201_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_5480 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_201_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_101_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_201_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_5507 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_203_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_101_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_203_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_5534 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_203_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_102_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_203_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_5561 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_205_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_102_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_205_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_5588 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_205_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_103_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_205_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_5615 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_207_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_103_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_207_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_5642 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_207_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_104_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_207_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_5669 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_209_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_104_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_209_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_5696 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_209_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_105_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_209_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_5723 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_211_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_105_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_211_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_5750 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_211_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_106_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_211_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_5777 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_213_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_106_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_213_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_5804 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_213_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_107_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_213_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_5831 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_215_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_107_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_215_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_5858 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_215_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_108_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_215_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_5885 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_217_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_108_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_217_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_5912 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_217_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_109_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_217_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_5939 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_219_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_109_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_219_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_5966 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_219_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_110_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_219_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_5993 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_221_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_110_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_221_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_6020 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_221_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_111_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_221_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_6047 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_223_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_111_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_223_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_6074 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_223_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_112_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_223_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_6101 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_225_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_112_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_225_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_6128 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_225_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_113_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_225_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_6155 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_227_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_113_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_227_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_6182 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_227_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_114_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_227_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_6209 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_229_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_114_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_229_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_6236 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_229_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_115_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_229_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_6263 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_231_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_115_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_231_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_6290 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_231_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_116_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_231_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_6317 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_233_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_116_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_233_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_6344 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_233_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_117_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_233_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_6371 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_235_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_117_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_235_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_6398 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_235_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_118_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_235_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_6425 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_237_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_118_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_237_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_6452 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_237_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_119_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_237_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_6479 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_239_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_119_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_239_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_6506 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_239_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_120_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_239_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_6533 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_241_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_120_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_241_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_6560 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_241_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_121_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_241_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_6587 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_243_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_121_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_243_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_6614 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_243_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_122_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_243_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_6641 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_245_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_122_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_245_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_6668 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_245_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_123_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_245_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_6695 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_247_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_123_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_247_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_6722 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_247_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_124_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_247_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_6749 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_249_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_124_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_249_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_6776 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_249_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_125_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_249_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_6803 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_251_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_125_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_251_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_6830 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_251_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_126_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_251_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_6857 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_253_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_126_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_253_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_6884 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_253_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_127_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_253_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_6911 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_255_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_127_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_255_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_6938 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_255_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_128_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_255_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_6965 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_257_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_128_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_257_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_6992 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_257_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_129_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_257_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_7019 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_259_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_129_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_259_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_7046 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_259_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_130_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_259_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_7073 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_261_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_130_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_261_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_7100 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_261_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_131_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_261_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_7127 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_263_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_131_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_263_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_7154 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_263_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_132_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_263_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_7181 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_265_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_132_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_265_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_7208 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_265_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_133_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_265_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_7235 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_267_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_133_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_267_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_7262 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_267_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_134_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_267_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_7289 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_269_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_134_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_269_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_7316 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_269_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_135_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_269_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_7343 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_271_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_135_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_271_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_7370 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_271_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_136_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_271_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_7397 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_273_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_136_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_273_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_7424 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_273_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_137_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_273_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_7451 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_275_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_137_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_275_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_7478 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_275_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_138_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_275_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_7505 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_277_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_138_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_277_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_7532 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_277_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_139_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_277_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_7559 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_279_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_139_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_279_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_7586 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_279_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_140_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_279_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_7613 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_281_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_140_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_281_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_7640 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_281_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_141_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_281_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_7667 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_283_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_141_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_283_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_7694 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_283_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_142_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_283_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_7721 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_285_value & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_142_1 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_285_value & _s3_predicted_ghist_ptr_T_45 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_7748 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_285_value & _s3_predicted_ghist_ptr_WIRE__0; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_143_0 = s3_ghist_ptr_value == s1_ghv_wens_new_ptr_285_value & _s3_predicted_ghist_ptr_WIRE__0 &
    s3_redirect; // @[BPU.scala 551:119]
  wire  _s3_ghv_wens_T_7775 = s3_ghist_ptr_value == 8'h0 & _s3_predicted_ghist_ptr_T_45; // @[BPU.scala 551:90]
  wire  s3_ghv_wens_143_1 = s3_ghist_ptr_value == 8'h0 & _s3_predicted_ghist_ptr_T_45 & s3_redirect; // @[BPU.scala 551:119]
  wire [1:0] hi_2 = {_s3_predicted_ghist_ptr_T_60,_s3_predicted_ghist_ptr_T_32}; // @[BPU.scala 579:60]
  wire  _T_666 = s3_ghv_wens_0_0 | s3_ghv_wens_0_1; // @[BPU.scala 582:26]
  wire  _T_667 = s3_ghv_wens_1_0 | s3_ghv_wens_1_1; // @[BPU.scala 582:26]
  wire  _T_668 = s3_ghv_wens_2_0 | s3_ghv_wens_2_1; // @[BPU.scala 582:26]
  wire  _T_669 = s3_ghv_wens_3_0 | s3_ghv_wens_3_1; // @[BPU.scala 582:26]
  wire  _T_670 = s3_ghv_wens_4_0 | s3_ghv_wens_4_1; // @[BPU.scala 582:26]
  wire  _T_671 = s3_ghv_wens_5_0 | s3_ghv_wens_5_1; // @[BPU.scala 582:26]
  wire  _T_672 = s3_ghv_wens_6_0 | s3_ghv_wens_6_1; // @[BPU.scala 582:26]
  wire  _T_673 = s3_ghv_wens_7_0 | s3_ghv_wens_7_1; // @[BPU.scala 582:26]
  wire  _T_674 = s3_ghv_wens_8_0 | s3_ghv_wens_8_1; // @[BPU.scala 582:26]
  wire  _T_675 = s3_ghv_wens_9_0 | s3_ghv_wens_9_1; // @[BPU.scala 582:26]
  wire  _T_676 = s3_ghv_wens_10_0 | s3_ghv_wens_10_1; // @[BPU.scala 582:26]
  wire  _T_677 = s3_ghv_wens_11_0 | s3_ghv_wens_11_1; // @[BPU.scala 582:26]
  wire  _T_678 = s3_ghv_wens_12_0 | s3_ghv_wens_12_1; // @[BPU.scala 582:26]
  wire  _T_679 = s3_ghv_wens_13_0 | s3_ghv_wens_13_1; // @[BPU.scala 582:26]
  wire  _T_680 = s3_ghv_wens_14_0 | s3_ghv_wens_14_1; // @[BPU.scala 582:26]
  wire  _T_681 = s3_ghv_wens_15_0 | s3_ghv_wens_15_1; // @[BPU.scala 582:26]
  wire  _T_682 = s3_ghv_wens_16_0 | s3_ghv_wens_16_1; // @[BPU.scala 582:26]
  wire  _T_683 = s3_ghv_wens_17_0 | s3_ghv_wens_17_1; // @[BPU.scala 582:26]
  wire  _T_684 = s3_ghv_wens_18_0 | s3_ghv_wens_18_1; // @[BPU.scala 582:26]
  wire  _T_685 = s3_ghv_wens_19_0 | s3_ghv_wens_19_1; // @[BPU.scala 582:26]
  wire  _T_686 = s3_ghv_wens_20_0 | s3_ghv_wens_20_1; // @[BPU.scala 582:26]
  wire  _T_687 = s3_ghv_wens_21_0 | s3_ghv_wens_21_1; // @[BPU.scala 582:26]
  wire  _T_688 = s3_ghv_wens_22_0 | s3_ghv_wens_22_1; // @[BPU.scala 582:26]
  wire  _T_689 = s3_ghv_wens_23_0 | s3_ghv_wens_23_1; // @[BPU.scala 582:26]
  wire  _T_690 = s3_ghv_wens_24_0 | s3_ghv_wens_24_1; // @[BPU.scala 582:26]
  wire  _T_691 = s3_ghv_wens_25_0 | s3_ghv_wens_25_1; // @[BPU.scala 582:26]
  wire  _T_692 = s3_ghv_wens_26_0 | s3_ghv_wens_26_1; // @[BPU.scala 582:26]
  wire  _T_693 = s3_ghv_wens_27_0 | s3_ghv_wens_27_1; // @[BPU.scala 582:26]
  wire  _T_694 = s3_ghv_wens_28_0 | s3_ghv_wens_28_1; // @[BPU.scala 582:26]
  wire  _T_695 = s3_ghv_wens_29_0 | s3_ghv_wens_29_1; // @[BPU.scala 582:26]
  wire  _T_696 = s3_ghv_wens_30_0 | s3_ghv_wens_30_1; // @[BPU.scala 582:26]
  wire  _T_697 = s3_ghv_wens_31_0 | s3_ghv_wens_31_1; // @[BPU.scala 582:26]
  wire  _T_698 = s3_ghv_wens_32_0 | s3_ghv_wens_32_1; // @[BPU.scala 582:26]
  wire  _T_699 = s3_ghv_wens_33_0 | s3_ghv_wens_33_1; // @[BPU.scala 582:26]
  wire  _T_700 = s3_ghv_wens_34_0 | s3_ghv_wens_34_1; // @[BPU.scala 582:26]
  wire  _T_701 = s3_ghv_wens_35_0 | s3_ghv_wens_35_1; // @[BPU.scala 582:26]
  wire  _T_702 = s3_ghv_wens_36_0 | s3_ghv_wens_36_1; // @[BPU.scala 582:26]
  wire  _T_703 = s3_ghv_wens_37_0 | s3_ghv_wens_37_1; // @[BPU.scala 582:26]
  wire  _T_704 = s3_ghv_wens_38_0 | s3_ghv_wens_38_1; // @[BPU.scala 582:26]
  wire  _T_705 = s3_ghv_wens_39_0 | s3_ghv_wens_39_1; // @[BPU.scala 582:26]
  wire  _T_706 = s3_ghv_wens_40_0 | s3_ghv_wens_40_1; // @[BPU.scala 582:26]
  wire  _T_707 = s3_ghv_wens_41_0 | s3_ghv_wens_41_1; // @[BPU.scala 582:26]
  wire  _T_708 = s3_ghv_wens_42_0 | s3_ghv_wens_42_1; // @[BPU.scala 582:26]
  wire  _T_709 = s3_ghv_wens_43_0 | s3_ghv_wens_43_1; // @[BPU.scala 582:26]
  wire  _T_710 = s3_ghv_wens_44_0 | s3_ghv_wens_44_1; // @[BPU.scala 582:26]
  wire  _T_711 = s3_ghv_wens_45_0 | s3_ghv_wens_45_1; // @[BPU.scala 582:26]
  wire  _T_712 = s3_ghv_wens_46_0 | s3_ghv_wens_46_1; // @[BPU.scala 582:26]
  wire  _T_713 = s3_ghv_wens_47_0 | s3_ghv_wens_47_1; // @[BPU.scala 582:26]
  wire  _T_714 = s3_ghv_wens_48_0 | s3_ghv_wens_48_1; // @[BPU.scala 582:26]
  wire  _T_715 = s3_ghv_wens_49_0 | s3_ghv_wens_49_1; // @[BPU.scala 582:26]
  wire  _T_716 = s3_ghv_wens_50_0 | s3_ghv_wens_50_1; // @[BPU.scala 582:26]
  wire  _T_717 = s3_ghv_wens_51_0 | s3_ghv_wens_51_1; // @[BPU.scala 582:26]
  wire  _T_718 = s3_ghv_wens_52_0 | s3_ghv_wens_52_1; // @[BPU.scala 582:26]
  wire  _T_719 = s3_ghv_wens_53_0 | s3_ghv_wens_53_1; // @[BPU.scala 582:26]
  wire  _T_720 = s3_ghv_wens_54_0 | s3_ghv_wens_54_1; // @[BPU.scala 582:26]
  wire  _T_721 = s3_ghv_wens_55_0 | s3_ghv_wens_55_1; // @[BPU.scala 582:26]
  wire  _T_722 = s3_ghv_wens_56_0 | s3_ghv_wens_56_1; // @[BPU.scala 582:26]
  wire  _T_723 = s3_ghv_wens_57_0 | s3_ghv_wens_57_1; // @[BPU.scala 582:26]
  wire  _T_724 = s3_ghv_wens_58_0 | s3_ghv_wens_58_1; // @[BPU.scala 582:26]
  wire  _T_725 = s3_ghv_wens_59_0 | s3_ghv_wens_59_1; // @[BPU.scala 582:26]
  wire  _T_726 = s3_ghv_wens_60_0 | s3_ghv_wens_60_1; // @[BPU.scala 582:26]
  wire  _T_727 = s3_ghv_wens_61_0 | s3_ghv_wens_61_1; // @[BPU.scala 582:26]
  wire  _T_728 = s3_ghv_wens_62_0 | s3_ghv_wens_62_1; // @[BPU.scala 582:26]
  wire  _T_729 = s3_ghv_wens_63_0 | s3_ghv_wens_63_1; // @[BPU.scala 582:26]
  wire  _T_730 = s3_ghv_wens_64_0 | s3_ghv_wens_64_1; // @[BPU.scala 582:26]
  wire  _T_731 = s3_ghv_wens_65_0 | s3_ghv_wens_65_1; // @[BPU.scala 582:26]
  wire  _T_732 = s3_ghv_wens_66_0 | s3_ghv_wens_66_1; // @[BPU.scala 582:26]
  wire  _T_733 = s3_ghv_wens_67_0 | s3_ghv_wens_67_1; // @[BPU.scala 582:26]
  wire  _T_734 = s3_ghv_wens_68_0 | s3_ghv_wens_68_1; // @[BPU.scala 582:26]
  wire  _T_735 = s3_ghv_wens_69_0 | s3_ghv_wens_69_1; // @[BPU.scala 582:26]
  wire  _T_736 = s3_ghv_wens_70_0 | s3_ghv_wens_70_1; // @[BPU.scala 582:26]
  wire  _T_737 = s3_ghv_wens_71_0 | s3_ghv_wens_71_1; // @[BPU.scala 582:26]
  wire  _T_738 = s3_ghv_wens_72_0 | s3_ghv_wens_72_1; // @[BPU.scala 582:26]
  wire  _T_739 = s3_ghv_wens_73_0 | s3_ghv_wens_73_1; // @[BPU.scala 582:26]
  wire  _T_740 = s3_ghv_wens_74_0 | s3_ghv_wens_74_1; // @[BPU.scala 582:26]
  wire  _T_741 = s3_ghv_wens_75_0 | s3_ghv_wens_75_1; // @[BPU.scala 582:26]
  wire  _T_742 = s3_ghv_wens_76_0 | s3_ghv_wens_76_1; // @[BPU.scala 582:26]
  wire  _T_743 = s3_ghv_wens_77_0 | s3_ghv_wens_77_1; // @[BPU.scala 582:26]
  wire  _T_744 = s3_ghv_wens_78_0 | s3_ghv_wens_78_1; // @[BPU.scala 582:26]
  wire  _T_745 = s3_ghv_wens_79_0 | s3_ghv_wens_79_1; // @[BPU.scala 582:26]
  wire  _T_746 = s3_ghv_wens_80_0 | s3_ghv_wens_80_1; // @[BPU.scala 582:26]
  wire  _T_747 = s3_ghv_wens_81_0 | s3_ghv_wens_81_1; // @[BPU.scala 582:26]
  wire  _T_748 = s3_ghv_wens_82_0 | s3_ghv_wens_82_1; // @[BPU.scala 582:26]
  wire  _T_749 = s3_ghv_wens_83_0 | s3_ghv_wens_83_1; // @[BPU.scala 582:26]
  wire  _T_750 = s3_ghv_wens_84_0 | s3_ghv_wens_84_1; // @[BPU.scala 582:26]
  wire  _T_751 = s3_ghv_wens_85_0 | s3_ghv_wens_85_1; // @[BPU.scala 582:26]
  wire  _T_752 = s3_ghv_wens_86_0 | s3_ghv_wens_86_1; // @[BPU.scala 582:26]
  wire  _T_753 = s3_ghv_wens_87_0 | s3_ghv_wens_87_1; // @[BPU.scala 582:26]
  wire  _T_754 = s3_ghv_wens_88_0 | s3_ghv_wens_88_1; // @[BPU.scala 582:26]
  wire  _T_755 = s3_ghv_wens_89_0 | s3_ghv_wens_89_1; // @[BPU.scala 582:26]
  wire  _T_756 = s3_ghv_wens_90_0 | s3_ghv_wens_90_1; // @[BPU.scala 582:26]
  wire  _T_757 = s3_ghv_wens_91_0 | s3_ghv_wens_91_1; // @[BPU.scala 582:26]
  wire  _T_758 = s3_ghv_wens_92_0 | s3_ghv_wens_92_1; // @[BPU.scala 582:26]
  wire  _T_759 = s3_ghv_wens_93_0 | s3_ghv_wens_93_1; // @[BPU.scala 582:26]
  wire  _T_760 = s3_ghv_wens_94_0 | s3_ghv_wens_94_1; // @[BPU.scala 582:26]
  wire  _T_761 = s3_ghv_wens_95_0 | s3_ghv_wens_95_1; // @[BPU.scala 582:26]
  wire  _T_762 = s3_ghv_wens_96_0 | s3_ghv_wens_96_1; // @[BPU.scala 582:26]
  wire  _T_763 = s3_ghv_wens_97_0 | s3_ghv_wens_97_1; // @[BPU.scala 582:26]
  wire  _T_764 = s3_ghv_wens_98_0 | s3_ghv_wens_98_1; // @[BPU.scala 582:26]
  wire  _T_765 = s3_ghv_wens_99_0 | s3_ghv_wens_99_1; // @[BPU.scala 582:26]
  wire  _T_766 = s3_ghv_wens_100_0 | s3_ghv_wens_100_1; // @[BPU.scala 582:26]
  wire  _T_767 = s3_ghv_wens_101_0 | s3_ghv_wens_101_1; // @[BPU.scala 582:26]
  wire  _T_768 = s3_ghv_wens_102_0 | s3_ghv_wens_102_1; // @[BPU.scala 582:26]
  wire  _T_769 = s3_ghv_wens_103_0 | s3_ghv_wens_103_1; // @[BPU.scala 582:26]
  wire  _T_770 = s3_ghv_wens_104_0 | s3_ghv_wens_104_1; // @[BPU.scala 582:26]
  wire  _T_771 = s3_ghv_wens_105_0 | s3_ghv_wens_105_1; // @[BPU.scala 582:26]
  wire  _T_772 = s3_ghv_wens_106_0 | s3_ghv_wens_106_1; // @[BPU.scala 582:26]
  wire  _T_773 = s3_ghv_wens_107_0 | s3_ghv_wens_107_1; // @[BPU.scala 582:26]
  wire  _T_774 = s3_ghv_wens_108_0 | s3_ghv_wens_108_1; // @[BPU.scala 582:26]
  wire  _T_775 = s3_ghv_wens_109_0 | s3_ghv_wens_109_1; // @[BPU.scala 582:26]
  wire  _T_776 = s3_ghv_wens_110_0 | s3_ghv_wens_110_1; // @[BPU.scala 582:26]
  wire  _T_777 = s3_ghv_wens_111_0 | s3_ghv_wens_111_1; // @[BPU.scala 582:26]
  wire  _T_778 = s3_ghv_wens_112_0 | s3_ghv_wens_112_1; // @[BPU.scala 582:26]
  wire  _T_779 = s3_ghv_wens_113_0 | s3_ghv_wens_113_1; // @[BPU.scala 582:26]
  wire  _T_780 = s3_ghv_wens_114_0 | s3_ghv_wens_114_1; // @[BPU.scala 582:26]
  wire  _T_781 = s3_ghv_wens_115_0 | s3_ghv_wens_115_1; // @[BPU.scala 582:26]
  wire  _T_782 = s3_ghv_wens_116_0 | s3_ghv_wens_116_1; // @[BPU.scala 582:26]
  wire  _T_783 = s3_ghv_wens_117_0 | s3_ghv_wens_117_1; // @[BPU.scala 582:26]
  wire  _T_784 = s3_ghv_wens_118_0 | s3_ghv_wens_118_1; // @[BPU.scala 582:26]
  wire  _T_785 = s3_ghv_wens_119_0 | s3_ghv_wens_119_1; // @[BPU.scala 582:26]
  wire  _T_786 = s3_ghv_wens_120_0 | s3_ghv_wens_120_1; // @[BPU.scala 582:26]
  wire  _T_787 = s3_ghv_wens_121_0 | s3_ghv_wens_121_1; // @[BPU.scala 582:26]
  wire  _T_788 = s3_ghv_wens_122_0 | s3_ghv_wens_122_1; // @[BPU.scala 582:26]
  wire  _T_789 = s3_ghv_wens_123_0 | s3_ghv_wens_123_1; // @[BPU.scala 582:26]
  wire  _T_790 = s3_ghv_wens_124_0 | s3_ghv_wens_124_1; // @[BPU.scala 582:26]
  wire  _T_791 = s3_ghv_wens_125_0 | s3_ghv_wens_125_1; // @[BPU.scala 582:26]
  wire  _T_792 = s3_ghv_wens_126_0 | s3_ghv_wens_126_1; // @[BPU.scala 582:26]
  wire  _T_793 = s3_ghv_wens_127_0 | s3_ghv_wens_127_1; // @[BPU.scala 582:26]
  wire  _T_794 = s3_ghv_wens_128_0 | s3_ghv_wens_128_1; // @[BPU.scala 582:26]
  wire  _T_795 = s3_ghv_wens_129_0 | s3_ghv_wens_129_1; // @[BPU.scala 582:26]
  wire  _T_796 = s3_ghv_wens_130_0 | s3_ghv_wens_130_1; // @[BPU.scala 582:26]
  wire  _T_797 = s3_ghv_wens_131_0 | s3_ghv_wens_131_1; // @[BPU.scala 582:26]
  wire  _T_798 = s3_ghv_wens_132_0 | s3_ghv_wens_132_1; // @[BPU.scala 582:26]
  wire  _T_799 = s3_ghv_wens_133_0 | s3_ghv_wens_133_1; // @[BPU.scala 582:26]
  wire  _T_800 = s3_ghv_wens_134_0 | s3_ghv_wens_134_1; // @[BPU.scala 582:26]
  wire  _T_801 = s3_ghv_wens_135_0 | s3_ghv_wens_135_1; // @[BPU.scala 582:26]
  wire  _T_802 = s3_ghv_wens_136_0 | s3_ghv_wens_136_1; // @[BPU.scala 582:26]
  wire  _T_803 = s3_ghv_wens_137_0 | s3_ghv_wens_137_1; // @[BPU.scala 582:26]
  wire  _T_804 = s3_ghv_wens_138_0 | s3_ghv_wens_138_1; // @[BPU.scala 582:26]
  wire  _T_805 = s3_ghv_wens_139_0 | s3_ghv_wens_139_1; // @[BPU.scala 582:26]
  wire  _T_806 = s3_ghv_wens_140_0 | s3_ghv_wens_140_1; // @[BPU.scala 582:26]
  wire  _T_807 = s3_ghv_wens_141_0 | s3_ghv_wens_141_1; // @[BPU.scala 582:26]
  wire  _T_808 = s3_ghv_wens_142_0 | s3_ghv_wens_142_1; // @[BPU.scala 582:26]
  wire  _T_809 = s3_ghv_wens_143_0 | s3_ghv_wens_143_1; // @[BPU.scala 582:26]
  reg  s2_ftq_idx_flag; // @[Reg.scala 16:16]
  reg [2:0] s2_ftq_idx_value; // @[Reg.scala 16:16]
  reg  s3_ftq_idx_flag; // @[Reg.scala 16:16]
  reg [2:0] s3_ftq_idx_value; // @[Reg.scala 16:16]
  reg  predictors_io_update_REG_valid; // @[BPU.scala 601:34]
  reg [38:0] predictors_io_update_REG_bits_pc; // @[BPU.scala 601:34]
  reg [7:0] predictors_io_update_REG_bits_spec_info_folded_hist_hist_17_folded_hist; // @[BPU.scala 601:34]
  reg [7:0] predictors_io_update_REG_bits_spec_info_folded_hist_hist_16_folded_hist; // @[BPU.scala 601:34]
  reg [10:0] predictors_io_update_REG_bits_spec_info_folded_hist_hist_15_folded_hist; // @[BPU.scala 601:34]
  reg [6:0] predictors_io_update_REG_bits_spec_info_folded_hist_hist_14_folded_hist; // @[BPU.scala 601:34]
  reg [6:0] predictors_io_update_REG_bits_spec_info_folded_hist_hist_13_folded_hist; // @[BPU.scala 601:34]
  reg [6:0] predictors_io_update_REG_bits_spec_info_folded_hist_hist_12_folded_hist; // @[BPU.scala 601:34]
  reg [8:0] predictors_io_update_REG_bits_spec_info_folded_hist_hist_10_folded_hist; // @[BPU.scala 601:34]
  reg [6:0] predictors_io_update_REG_bits_spec_info_folded_hist_hist_9_folded_hist; // @[BPU.scala 601:34]
  reg [7:0] predictors_io_update_REG_bits_spec_info_folded_hist_hist_8_folded_hist; // @[BPU.scala 601:34]
  reg [8:0] predictors_io_update_REG_bits_spec_info_folded_hist_hist_7_folded_hist; // @[BPU.scala 601:34]
  reg [8:0] predictors_io_update_REG_bits_spec_info_folded_hist_hist_6_folded_hist; // @[BPU.scala 601:34]
  reg [10:0] predictors_io_update_REG_bits_spec_info_folded_hist_hist_5_folded_hist; // @[BPU.scala 601:34]
  reg [3:0] predictors_io_update_REG_bits_spec_info_folded_hist_hist_4_folded_hist; // @[BPU.scala 601:34]
  reg [10:0] predictors_io_update_REG_bits_spec_info_folded_hist_hist_3_folded_hist; // @[BPU.scala 601:34]
  reg [7:0] predictors_io_update_REG_bits_spec_info_folded_hist_hist_2_folded_hist; // @[BPU.scala 601:34]
  reg [7:0] predictors_io_update_REG_bits_spec_info_folded_hist_hist_1_folded_hist; // @[BPU.scala 601:34]
  reg [7:0] predictors_io_update_REG_bits_spec_info_folded_hist_hist_0_folded_hist; // @[BPU.scala 601:34]
  reg  predictors_io_update_REG_bits_ftb_entry_valid; // @[BPU.scala 601:34]
  reg [2:0] predictors_io_update_REG_bits_ftb_entry_brSlots_0_offset; // @[BPU.scala 601:34]
  reg [11:0] predictors_io_update_REG_bits_ftb_entry_brSlots_0_lower; // @[BPU.scala 601:34]
  reg [1:0] predictors_io_update_REG_bits_ftb_entry_brSlots_0_tarStat; // @[BPU.scala 601:34]
  reg  predictors_io_update_REG_bits_ftb_entry_brSlots_0_sharing; // @[BPU.scala 601:34]
  reg  predictors_io_update_REG_bits_ftb_entry_brSlots_0_valid; // @[BPU.scala 601:34]
  reg [2:0] predictors_io_update_REG_bits_ftb_entry_tailSlot_offset; // @[BPU.scala 601:34]
  reg [19:0] predictors_io_update_REG_bits_ftb_entry_tailSlot_lower; // @[BPU.scala 601:34]
  reg [1:0] predictors_io_update_REG_bits_ftb_entry_tailSlot_tarStat; // @[BPU.scala 601:34]
  reg  predictors_io_update_REG_bits_ftb_entry_tailSlot_sharing; // @[BPU.scala 601:34]
  reg  predictors_io_update_REG_bits_ftb_entry_tailSlot_valid; // @[BPU.scala 601:34]
  reg [2:0] predictors_io_update_REG_bits_ftb_entry_pftAddr; // @[BPU.scala 601:34]
  reg  predictors_io_update_REG_bits_ftb_entry_carry; // @[BPU.scala 601:34]
  reg  predictors_io_update_REG_bits_ftb_entry_isCall; // @[BPU.scala 601:34]
  reg  predictors_io_update_REG_bits_ftb_entry_isRet; // @[BPU.scala 601:34]
  reg  predictors_io_update_REG_bits_ftb_entry_isJalr; // @[BPU.scala 601:34]
  reg  predictors_io_update_REG_bits_ftb_entry_last_may_be_rvi_call; // @[BPU.scala 601:34]
  reg  predictors_io_update_REG_bits_ftb_entry_always_taken_0; // @[BPU.scala 601:34]
  reg  predictors_io_update_REG_bits_ftb_entry_always_taken_1; // @[BPU.scala 601:34]
  reg  predictors_io_update_REG_bits_br_taken_mask_0; // @[BPU.scala 601:34]
  reg  predictors_io_update_REG_bits_br_taken_mask_1; // @[BPU.scala 601:34]
  reg  predictors_io_update_REG_bits_jmp_taken; // @[BPU.scala 601:34]
  reg  predictors_io_update_REG_bits_mispred_mask_0; // @[BPU.scala 601:34]
  reg  predictors_io_update_REG_bits_mispred_mask_1; // @[BPU.scala 601:34]
  reg  predictors_io_update_REG_bits_mispred_mask_2; // @[BPU.scala 601:34]
  reg  predictors_io_update_REG_bits_old_entry; // @[BPU.scala 601:34]
  reg [255:0] predictors_io_update_REG_bits_meta; // @[BPU.scala 601:34]
  reg [38:0] predictors_io_update_REG_bits_full_target; // @[BPU.scala 601:34]
  wire [1:0] _shouldShiftVec_T_2 = do_redirect_bits_cfiUpdate_shift - 2'h1; // @[BPU.scala 609:129]
  wire [3:0] _shouldShiftVec_T_3 = 4'h1 << _shouldShiftVec_T_2; // @[BPU.scala 609:120]
  wire [3:0] _GEN_11931 = {{1'd0}, _shouldShiftVec_T_3[3:1]}; // @[ParallelMux.scala 36:53]
  wire [3:0] _shouldShiftVec_T_8 = _shouldShiftVec_T_3 | _GEN_11931; // @[ParallelMux.scala 36:53]
  wire [1:0] _GEN_11932 = {{1'd0}, _shouldShiftVec_T_3[3]}; // @[ParallelMux.scala 36:53]
  wire [1:0] _shouldShiftVec_T_9 = _shouldShiftVec_T_3[3:2] | _GEN_11932; // @[ParallelMux.scala 36:53]
  wire [3:0] _shouldShiftVec_WIRE_2 = {{2'd0}, _shouldShiftVec_T_9}; // @[ParallelMux.scala 36:{73,73}]
  wire [3:0] _shouldShiftVec_T_10 = _shouldShiftVec_T_8 | _shouldShiftVec_WIRE_2; // @[ParallelMux.scala 36:53]
  wire  shouldShiftVec_0 = do_redirect_bits_cfiUpdate_shift == 2'h0 ? 1'h0 : _shouldShiftVec_T_10[0]; // @[BPU.scala 609:27]
  wire  shouldShiftVec_1 = do_redirect_bits_cfiUpdate_shift == 2'h0 ? 1'h0 : _shouldShiftVec_T_10[1]; // @[BPU.scala 609:27]
  wire  real_br_taken_mask_0 = do_redirect_bits_cfiUpdate_shift == 2'h1 & do_redirect_bits_cfiUpdate_taken &
    do_redirect_bits_cfiUpdate_addIntoHist; // @[BPU.scala 617:80]
  wire  real_br_taken_mask_1 = do_redirect_bits_cfiUpdate_shift == 2'h2 & do_redirect_bits_cfiUpdate_taken &
    do_redirect_bits_cfiUpdate_addIntoHist; // @[BPU.scala 617:80]
  wire [7:0] _GEN_11933 = {{6'd0}, do_redirect_bits_cfiUpdate_shift}; // @[CircularQueuePtr.scala 54:50]
  wire [7:0] _updated_ptr_flipped_new_ptr_T_1 = 8'h90 - _GEN_11933; // @[CircularQueuePtr.scala 54:50]
  wire [8:0] updated_ptr_flipped_new_ptr_new_value = do_redirect_bits_cfiUpdate_histPtr_value +
    _updated_ptr_flipped_new_ptr_T_1; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _updated_ptr_flipped_new_ptr_diff_T_1 = {1'h0,updated_ptr_flipped_new_ptr_new_value}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] updated_ptr_flipped_new_ptr_diff = $signed(_updated_ptr_flipped_new_ptr_diff_T_1) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  updated_ptr_flipped_new_ptr_reverse_flag = $signed(updated_ptr_flipped_new_ptr_diff) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire  updated_ptr_flipped_new_ptr_flag = updated_ptr_flipped_new_ptr_reverse_flag ? ~
    do_redirect_bits_cfiUpdate_histPtr_flag : do_redirect_bits_cfiUpdate_histPtr_flag; // @[CircularQueuePtr.scala 44:26]
  wire [9:0] _updated_ptr_flipped_new_ptr_new_ptr_value_T = $signed(_updated_ptr_flipped_new_ptr_diff_T_1) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _updated_ptr_flipped_new_ptr_new_ptr_value_T_1 = updated_ptr_flipped_new_ptr_reverse_flag ?
    _updated_ptr_flipped_new_ptr_new_ptr_value_T : {{1'd0}, updated_ptr_flipped_new_ptr_new_value}; // @[CircularQueuePtr.scala 45:27]
  wire  _updated_fh_T = do_redirect_bits_cfiUpdate_taken & do_redirect_bits_cfiUpdate_addIntoHist; // @[BPU.scala 622:92]
  wire  updated_fh_ob__0 = do_redirect_bits_cfiUpdate_lastBrNumOH[0] & do_redirect_bits_cfiUpdate_afhob_afhob_3_bits_0
     | do_redirect_bits_cfiUpdate_lastBrNumOH[1] & do_redirect_bits_cfiUpdate_afhob_afhob_3_bits_1 |
    do_redirect_bits_cfiUpdate_lastBrNumOH[2] & do_redirect_bits_cfiUpdate_afhob_afhob_3_bits_2; // @[Mux.scala 27:73]
  wire  updated_fh_ob__1 = do_redirect_bits_cfiUpdate_lastBrNumOH[0] & do_redirect_bits_cfiUpdate_afhob_afhob_3_bits_1
     | do_redirect_bits_cfiUpdate_lastBrNumOH[1] & do_redirect_bits_cfiUpdate_afhob_afhob_3_bits_2 |
    do_redirect_bits_cfiUpdate_lastBrNumOH[2] & do_redirect_bits_cfiUpdate_afhob_afhob_3_bits_3; // @[Mux.scala 27:73]
  wire  updated_fh_res_hist_0_new_folded_hist_original_bits_masked__0 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_0_folded_hist[0]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_0_new_folded_hist_original_bits_masked__1 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_0_folded_hist[1]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_0_new_folded_hist_original_bits_masked__2 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_0_folded_hist[2]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_0_new_folded_hist_original_bits_masked__3 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_0_folded_hist[3]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_0_new_folded_hist_original_bits_masked__4 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_0_folded_hist[4]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_0_new_folded_hist_original_bits_masked__5 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_0_folded_hist[5]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_0_new_folded_hist_original_bits_masked__6 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_0_folded_hist[6]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_0_new_folded_hist_original_bits_masked__7 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_0_folded_hist[7]; // @[FrontendBundle.scala 280:54]
  wire [7:0] updated_fh_res_hist_0_new_folded_hist_xored = {
    updated_fh_res_hist_0_new_folded_hist_original_bits_masked__7,
    updated_fh_res_hist_0_new_folded_hist_original_bits_masked__6,
    updated_fh_res_hist_0_new_folded_hist_original_bits_masked__5,
    updated_fh_res_hist_0_new_folded_hist_original_bits_masked__4,
    updated_fh_res_hist_0_new_folded_hist_original_bits_masked__3,
    updated_fh_res_hist_0_new_folded_hist_original_bits_masked__2,
    updated_fh_res_hist_0_new_folded_hist_original_bits_masked__1,
    updated_fh_res_hist_0_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [15:0] updated_fh_res_hist_0_new_folded_hist_src_doubled = {
    updated_fh_res_hist_0_new_folded_hist_original_bits_masked__7,
    updated_fh_res_hist_0_new_folded_hist_original_bits_masked__6,
    updated_fh_res_hist_0_new_folded_hist_original_bits_masked__5,
    updated_fh_res_hist_0_new_folded_hist_original_bits_masked__4,
    updated_fh_res_hist_0_new_folded_hist_original_bits_masked__3,
    updated_fh_res_hist_0_new_folded_hist_original_bits_masked__2,
    updated_fh_res_hist_0_new_folded_hist_original_bits_masked__1,
    updated_fh_res_hist_0_new_folded_hist_original_bits_masked__0,updated_fh_res_hist_0_new_folded_hist_xored}; // @[Cat.scala 31:58]
  wire [7:0] updated_fh_res_hist_0_new_folded_hist = updated_fh_res_hist_0_new_folded_hist_src_doubled[15:8]; // @[FrontendBundle.scala 221:30]
  wire  updated_fh_ob_1_0 = do_redirect_bits_cfiUpdate_lastBrNumOH[0] & do_redirect_bits_cfiUpdate_afhob_afhob_2_bits_0
     | do_redirect_bits_cfiUpdate_lastBrNumOH[1] & do_redirect_bits_cfiUpdate_afhob_afhob_2_bits_1 |
    do_redirect_bits_cfiUpdate_lastBrNumOH[2] & do_redirect_bits_cfiUpdate_afhob_afhob_2_bits_2; // @[Mux.scala 27:73]
  wire  updated_fh_ob_1_1 = do_redirect_bits_cfiUpdate_lastBrNumOH[0] & do_redirect_bits_cfiUpdate_afhob_afhob_2_bits_1
     | do_redirect_bits_cfiUpdate_lastBrNumOH[1] & do_redirect_bits_cfiUpdate_afhob_afhob_2_bits_2 |
    do_redirect_bits_cfiUpdate_lastBrNumOH[2] & do_redirect_bits_cfiUpdate_afhob_afhob_2_bits_3; // @[Mux.scala 27:73]
  wire  updated_fh_res_hist_1_new_folded_hist_original_bits_masked__0 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_1_folded_hist[0]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_1_new_folded_hist_original_bits_masked__1 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_1_folded_hist[1]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_1_new_folded_hist_original_bits_masked__2 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_1_folded_hist[2]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_1_new_folded_hist_original_bits_masked__3 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_1_folded_hist[3]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_1_new_folded_hist_original_bits_masked__4 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_1_folded_hist[4]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_1_new_folded_hist_original_bits_masked__5 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_1_folded_hist[5]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_1_new_folded_hist_original_bits_masked__6 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_1_folded_hist[6]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_1_new_folded_hist_original_bits_masked__7 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_1_folded_hist[7]; // @[FrontendBundle.scala 280:54]
  wire [7:0] updated_fh_res_hist_1_new_folded_hist_xored = {
    updated_fh_res_hist_1_new_folded_hist_original_bits_masked__7,
    updated_fh_res_hist_1_new_folded_hist_original_bits_masked__6,
    updated_fh_res_hist_1_new_folded_hist_original_bits_masked__5,
    updated_fh_res_hist_1_new_folded_hist_original_bits_masked__4,
    updated_fh_res_hist_1_new_folded_hist_original_bits_masked__3,
    updated_fh_res_hist_1_new_folded_hist_original_bits_masked__2,
    updated_fh_res_hist_1_new_folded_hist_original_bits_masked__1,
    updated_fh_res_hist_1_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [15:0] updated_fh_res_hist_1_new_folded_hist_src_doubled = {
    updated_fh_res_hist_1_new_folded_hist_original_bits_masked__7,
    updated_fh_res_hist_1_new_folded_hist_original_bits_masked__6,
    updated_fh_res_hist_1_new_folded_hist_original_bits_masked__5,
    updated_fh_res_hist_1_new_folded_hist_original_bits_masked__4,
    updated_fh_res_hist_1_new_folded_hist_original_bits_masked__3,
    updated_fh_res_hist_1_new_folded_hist_original_bits_masked__2,
    updated_fh_res_hist_1_new_folded_hist_original_bits_masked__1,
    updated_fh_res_hist_1_new_folded_hist_original_bits_masked__0,updated_fh_res_hist_1_new_folded_hist_xored}; // @[Cat.scala 31:58]
  wire [7:0] updated_fh_res_hist_1_new_folded_hist = updated_fh_res_hist_1_new_folded_hist_src_doubled[15:8]; // @[FrontendBundle.scala 221:30]
  wire  updated_fh_ob_2_0 = do_redirect_bits_cfiUpdate_lastBrNumOH[0] & do_redirect_bits_cfiUpdate_afhob_afhob_5_bits_0
     | do_redirect_bits_cfiUpdate_lastBrNumOH[1] & do_redirect_bits_cfiUpdate_afhob_afhob_5_bits_1 |
    do_redirect_bits_cfiUpdate_lastBrNumOH[2] & do_redirect_bits_cfiUpdate_afhob_afhob_5_bits_2; // @[Mux.scala 27:73]
  wire  updated_fh_ob_2_1 = do_redirect_bits_cfiUpdate_lastBrNumOH[0] & do_redirect_bits_cfiUpdate_afhob_afhob_5_bits_1
     | do_redirect_bits_cfiUpdate_lastBrNumOH[1] & do_redirect_bits_cfiUpdate_afhob_afhob_5_bits_2 |
    do_redirect_bits_cfiUpdate_lastBrNumOH[2] & do_redirect_bits_cfiUpdate_afhob_afhob_5_bits_3; // @[Mux.scala 27:73]
  wire  updated_fh_res_hist_2_new_folded_hist_original_bits_masked__0 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_2_folded_hist[0]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_2_new_folded_hist_original_bits_masked__1 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_2_folded_hist[1]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_2_new_folded_hist_original_bits_masked__2 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_2_folded_hist[2]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_2_new_folded_hist_original_bits_masked__3 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_2_folded_hist[3]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_2_new_folded_hist_original_bits_masked__4 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_2_folded_hist[4]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_2_new_folded_hist_original_bits_masked__5 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_2_folded_hist[5]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_2_new_folded_hist_original_bits_masked__6 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_2_folded_hist[6]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_2_new_folded_hist_original_bits_masked__7 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_2_folded_hist[7]; // @[FrontendBundle.scala 280:54]
  wire [7:0] updated_fh_res_hist_2_new_folded_hist_xored = {
    updated_fh_res_hist_2_new_folded_hist_original_bits_masked__7,
    updated_fh_res_hist_2_new_folded_hist_original_bits_masked__6,
    updated_fh_res_hist_2_new_folded_hist_original_bits_masked__5,
    updated_fh_res_hist_2_new_folded_hist_original_bits_masked__4,
    updated_fh_res_hist_2_new_folded_hist_original_bits_masked__3,
    updated_fh_res_hist_2_new_folded_hist_original_bits_masked__2,
    updated_fh_res_hist_2_new_folded_hist_original_bits_masked__1,
    updated_fh_res_hist_2_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [15:0] updated_fh_res_hist_2_new_folded_hist_src_doubled = {
    updated_fh_res_hist_2_new_folded_hist_original_bits_masked__7,
    updated_fh_res_hist_2_new_folded_hist_original_bits_masked__6,
    updated_fh_res_hist_2_new_folded_hist_original_bits_masked__5,
    updated_fh_res_hist_2_new_folded_hist_original_bits_masked__4,
    updated_fh_res_hist_2_new_folded_hist_original_bits_masked__3,
    updated_fh_res_hist_2_new_folded_hist_original_bits_masked__2,
    updated_fh_res_hist_2_new_folded_hist_original_bits_masked__1,
    updated_fh_res_hist_2_new_folded_hist_original_bits_masked__0,updated_fh_res_hist_2_new_folded_hist_xored}; // @[Cat.scala 31:58]
  wire [7:0] updated_fh_res_hist_2_new_folded_hist = updated_fh_res_hist_2_new_folded_hist_src_doubled[15:8]; // @[FrontendBundle.scala 221:30]
  wire  updated_fh_res_hist_3_new_folded_hist_original_bits_masked__0 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_3_folded_hist[0]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_3_new_folded_hist_original_bits_masked__1 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_3_folded_hist[1]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_3_new_folded_hist_original_bits_masked__2 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_3_folded_hist[2]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_3_new_folded_hist_original_bits_masked__3 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_3_folded_hist[3]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_3_new_folded_hist_original_bits_masked__4 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_3_folded_hist[4]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_3_new_folded_hist_original_bits_masked__5 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_3_folded_hist[5]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_3_new_folded_hist_original_bits_masked__6 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_3_folded_hist[6]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_3_new_folded_hist_original_bits_masked__7 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_3_folded_hist[7]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_3_new_folded_hist_original_bits_masked__8 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_3_folded_hist[8]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_3_new_folded_hist_original_bits_masked__9 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_3_folded_hist[9]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_3_new_folded_hist_original_bits_masked__10 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_3_folded_hist[10]; // @[FrontendBundle.scala 280:54]
  wire [4:0] updated_fh_res_hist_3_new_folded_hist_xored_lo = {
    updated_fh_res_hist_3_new_folded_hist_original_bits_masked__4,
    updated_fh_res_hist_3_new_folded_hist_original_bits_masked__3,
    updated_fh_res_hist_3_new_folded_hist_original_bits_masked__2,
    updated_fh_res_hist_3_new_folded_hist_original_bits_masked__1,
    updated_fh_res_hist_3_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [10:0] updated_fh_res_hist_3_new_folded_hist_xored = {
    updated_fh_res_hist_3_new_folded_hist_original_bits_masked__10,
    updated_fh_res_hist_3_new_folded_hist_original_bits_masked__9,
    updated_fh_res_hist_3_new_folded_hist_original_bits_masked__8,
    updated_fh_res_hist_3_new_folded_hist_original_bits_masked__7,
    updated_fh_res_hist_3_new_folded_hist_original_bits_masked__6,
    updated_fh_res_hist_3_new_folded_hist_original_bits_masked__5,updated_fh_res_hist_3_new_folded_hist_xored_lo}; // @[FrontendBundle.scala 258:11]
  wire [21:0] updated_fh_res_hist_3_new_folded_hist_src_doubled = {
    updated_fh_res_hist_3_new_folded_hist_original_bits_masked__10,
    updated_fh_res_hist_3_new_folded_hist_original_bits_masked__9,
    updated_fh_res_hist_3_new_folded_hist_original_bits_masked__8,
    updated_fh_res_hist_3_new_folded_hist_original_bits_masked__7,
    updated_fh_res_hist_3_new_folded_hist_original_bits_masked__6,
    updated_fh_res_hist_3_new_folded_hist_original_bits_masked__5,updated_fh_res_hist_3_new_folded_hist_xored_lo,
    updated_fh_res_hist_3_new_folded_hist_xored}; // @[Cat.scala 31:58]
  wire [10:0] updated_fh_res_hist_3_new_folded_hist = updated_fh_res_hist_3_new_folded_hist_src_doubled[21:11]; // @[FrontendBundle.scala 221:30]
  wire [3:0] _GEN_11934 = {{3'd0}, _updated_fh_T}; // @[FrontendBundle.scala 290:29]
  wire [3:0] updated_fh_res_hist_4_new_folded_hist = do_redirect_bits_cfiUpdate_folded_hist_hist_4_folded_hist |
    _GEN_11934; // @[FrontendBundle.scala 290:29]
  wire  updated_fh_ob_4_0 = do_redirect_bits_cfiUpdate_lastBrNumOH[0] & do_redirect_bits_cfiUpdate_afhob_afhob_1_bits_0
     | do_redirect_bits_cfiUpdate_lastBrNumOH[1] & do_redirect_bits_cfiUpdate_afhob_afhob_1_bits_1 |
    do_redirect_bits_cfiUpdate_lastBrNumOH[2] & do_redirect_bits_cfiUpdate_afhob_afhob_1_bits_2; // @[Mux.scala 27:73]
  wire  updated_fh_ob_4_1 = do_redirect_bits_cfiUpdate_lastBrNumOH[0] & do_redirect_bits_cfiUpdate_afhob_afhob_1_bits_1
     | do_redirect_bits_cfiUpdate_lastBrNumOH[1] & do_redirect_bits_cfiUpdate_afhob_afhob_1_bits_2 |
    do_redirect_bits_cfiUpdate_lastBrNumOH[2] & do_redirect_bits_cfiUpdate_afhob_afhob_1_bits_3; // @[Mux.scala 27:73]
  wire  updated_fh_res_hist_5_new_folded_hist_original_bits_masked__0 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_5_folded_hist[0]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_5_new_folded_hist_original_bits_masked__1 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_5_folded_hist[1]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_5_new_folded_hist_original_bits_masked__2 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_5_folded_hist[2]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_5_new_folded_hist_original_bits_masked__3 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_5_folded_hist[3]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_5_new_folded_hist_original_bits_masked__4 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_5_folded_hist[4]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_5_new_folded_hist_original_bits_masked__5 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_5_folded_hist[5]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_5_new_folded_hist_original_bits_masked__6 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_5_folded_hist[6]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_5_new_folded_hist_original_bits_masked__7 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_5_folded_hist[7]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_5_new_folded_hist_original_bits_masked__8 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_5_folded_hist[8]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_5_new_folded_hist_original_bits_masked__9 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_5_folded_hist[9]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_5_new_folded_hist_original_bits_masked__10 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_5_folded_hist[10]; // @[FrontendBundle.scala 280:54]
  wire [4:0] updated_fh_res_hist_5_new_folded_hist_xored_lo = {
    updated_fh_res_hist_5_new_folded_hist_original_bits_masked__4,
    updated_fh_res_hist_5_new_folded_hist_original_bits_masked__3,
    updated_fh_res_hist_5_new_folded_hist_original_bits_masked__2,
    updated_fh_res_hist_5_new_folded_hist_original_bits_masked__1,
    updated_fh_res_hist_5_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [10:0] updated_fh_res_hist_5_new_folded_hist_xored = {
    updated_fh_res_hist_5_new_folded_hist_original_bits_masked__10,
    updated_fh_res_hist_5_new_folded_hist_original_bits_masked__9,
    updated_fh_res_hist_5_new_folded_hist_original_bits_masked__8,
    updated_fh_res_hist_5_new_folded_hist_original_bits_masked__7,
    updated_fh_res_hist_5_new_folded_hist_original_bits_masked__6,
    updated_fh_res_hist_5_new_folded_hist_original_bits_masked__5,updated_fh_res_hist_5_new_folded_hist_xored_lo}; // @[FrontendBundle.scala 258:11]
  wire [21:0] updated_fh_res_hist_5_new_folded_hist_src_doubled = {
    updated_fh_res_hist_5_new_folded_hist_original_bits_masked__10,
    updated_fh_res_hist_5_new_folded_hist_original_bits_masked__9,
    updated_fh_res_hist_5_new_folded_hist_original_bits_masked__8,
    updated_fh_res_hist_5_new_folded_hist_original_bits_masked__7,
    updated_fh_res_hist_5_new_folded_hist_original_bits_masked__6,
    updated_fh_res_hist_5_new_folded_hist_original_bits_masked__5,updated_fh_res_hist_5_new_folded_hist_xored_lo,
    updated_fh_res_hist_5_new_folded_hist_xored}; // @[Cat.scala 31:58]
  wire [10:0] updated_fh_res_hist_5_new_folded_hist = updated_fh_res_hist_5_new_folded_hist_src_doubled[21:11]; // @[FrontendBundle.scala 221:30]
  wire  updated_fh_res_hist_6_new_folded_hist_original_bits_masked__0 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_6_folded_hist[0]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_6_new_folded_hist_original_bits_masked__1 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_6_folded_hist[1]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_6_new_folded_hist_original_bits_masked__2 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_6_folded_hist[2]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_6_new_folded_hist_original_bits_masked__3 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_6_folded_hist[3]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_6_new_folded_hist_original_bits_masked__4 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_6_folded_hist[4]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_6_new_folded_hist_original_bits_masked__5 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_6_folded_hist[5]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_6_new_folded_hist_original_bits_masked__6 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_6_folded_hist[6]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_6_new_folded_hist_original_bits_masked__7 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_6_folded_hist[7]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_6_new_folded_hist_original_bits_masked__8 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_6_folded_hist[8]; // @[FrontendBundle.scala 280:54]
  wire [8:0] updated_fh_res_hist_6_new_folded_hist_xored = {
    updated_fh_res_hist_6_new_folded_hist_original_bits_masked__8,
    updated_fh_res_hist_6_new_folded_hist_original_bits_masked__7,
    updated_fh_res_hist_6_new_folded_hist_original_bits_masked__6,
    updated_fh_res_hist_6_new_folded_hist_original_bits_masked__5,
    updated_fh_res_hist_6_new_folded_hist_original_bits_masked__4,
    updated_fh_res_hist_6_new_folded_hist_original_bits_masked__3,
    updated_fh_res_hist_6_new_folded_hist_original_bits_masked__2,
    updated_fh_res_hist_6_new_folded_hist_original_bits_masked__1,
    updated_fh_res_hist_6_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [17:0] updated_fh_res_hist_6_new_folded_hist_src_doubled = {
    updated_fh_res_hist_6_new_folded_hist_original_bits_masked__8,
    updated_fh_res_hist_6_new_folded_hist_original_bits_masked__7,
    updated_fh_res_hist_6_new_folded_hist_original_bits_masked__6,
    updated_fh_res_hist_6_new_folded_hist_original_bits_masked__5,
    updated_fh_res_hist_6_new_folded_hist_original_bits_masked__4,
    updated_fh_res_hist_6_new_folded_hist_original_bits_masked__3,
    updated_fh_res_hist_6_new_folded_hist_original_bits_masked__2,
    updated_fh_res_hist_6_new_folded_hist_original_bits_masked__1,
    updated_fh_res_hist_6_new_folded_hist_original_bits_masked__0,updated_fh_res_hist_6_new_folded_hist_xored}; // @[Cat.scala 31:58]
  wire [8:0] updated_fh_res_hist_6_new_folded_hist = updated_fh_res_hist_6_new_folded_hist_src_doubled[17:9]; // @[FrontendBundle.scala 221:30]
  wire  updated_fh_res_hist_7_new_folded_hist_original_bits_masked__0 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_7_folded_hist[0]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_7_new_folded_hist_original_bits_masked__1 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_7_folded_hist[1]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_7_new_folded_hist_original_bits_masked__2 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_7_folded_hist[2]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_7_new_folded_hist_original_bits_masked__3 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_7_folded_hist[3]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_7_new_folded_hist_original_bits_masked__4 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_7_folded_hist[4]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_7_new_folded_hist_original_bits_masked__5 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_7_folded_hist[5]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_7_new_folded_hist_original_bits_masked__6 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_7_folded_hist[6]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_7_new_folded_hist_original_bits_masked__7 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_7_folded_hist[7]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_7_new_folded_hist_original_bits_masked__8 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_7_folded_hist[8]; // @[FrontendBundle.scala 280:54]
  wire [8:0] updated_fh_res_hist_7_new_folded_hist_xored = {
    updated_fh_res_hist_7_new_folded_hist_original_bits_masked__8,
    updated_fh_res_hist_7_new_folded_hist_original_bits_masked__7,
    updated_fh_res_hist_7_new_folded_hist_original_bits_masked__6,
    updated_fh_res_hist_7_new_folded_hist_original_bits_masked__5,
    updated_fh_res_hist_7_new_folded_hist_original_bits_masked__4,
    updated_fh_res_hist_7_new_folded_hist_original_bits_masked__3,
    updated_fh_res_hist_7_new_folded_hist_original_bits_masked__2,
    updated_fh_res_hist_7_new_folded_hist_original_bits_masked__1,
    updated_fh_res_hist_7_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [17:0] updated_fh_res_hist_7_new_folded_hist_src_doubled = {
    updated_fh_res_hist_7_new_folded_hist_original_bits_masked__8,
    updated_fh_res_hist_7_new_folded_hist_original_bits_masked__7,
    updated_fh_res_hist_7_new_folded_hist_original_bits_masked__6,
    updated_fh_res_hist_7_new_folded_hist_original_bits_masked__5,
    updated_fh_res_hist_7_new_folded_hist_original_bits_masked__4,
    updated_fh_res_hist_7_new_folded_hist_original_bits_masked__3,
    updated_fh_res_hist_7_new_folded_hist_original_bits_masked__2,
    updated_fh_res_hist_7_new_folded_hist_original_bits_masked__1,
    updated_fh_res_hist_7_new_folded_hist_original_bits_masked__0,updated_fh_res_hist_7_new_folded_hist_xored}; // @[Cat.scala 31:58]
  wire [8:0] updated_fh_res_hist_7_new_folded_hist = updated_fh_res_hist_7_new_folded_hist_src_doubled[17:9]; // @[FrontendBundle.scala 221:30]
  wire [7:0] _GEN_11935 = {{7'd0}, _updated_fh_T}; // @[FrontendBundle.scala 290:29]
  wire [7:0] updated_fh_res_hist_8_new_folded_hist = do_redirect_bits_cfiUpdate_folded_hist_hist_8_folded_hist |
    _GEN_11935; // @[FrontendBundle.scala 290:29]
  wire  updated_fh_res_hist_9_new_folded_hist_original_bits_masked__0 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_9_folded_hist[0]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_9_new_folded_hist_original_bits_masked__1 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_9_folded_hist[1]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_9_new_folded_hist_original_bits_masked__2 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_9_folded_hist[2]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_9_new_folded_hist_original_bits_masked__3 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_9_folded_hist[3]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_9_new_folded_hist_original_bits_masked__4 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_9_folded_hist[4]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_9_new_folded_hist_original_bits_masked__5 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_9_folded_hist[5]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_9_new_folded_hist_original_bits_masked__6 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_9_folded_hist[6]; // @[FrontendBundle.scala 280:54]
  wire [6:0] updated_fh_res_hist_9_new_folded_hist_xored = {
    updated_fh_res_hist_9_new_folded_hist_original_bits_masked__6,
    updated_fh_res_hist_9_new_folded_hist_original_bits_masked__5,
    updated_fh_res_hist_9_new_folded_hist_original_bits_masked__4,
    updated_fh_res_hist_9_new_folded_hist_original_bits_masked__3,
    updated_fh_res_hist_9_new_folded_hist_original_bits_masked__2,
    updated_fh_res_hist_9_new_folded_hist_original_bits_masked__1,
    updated_fh_res_hist_9_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [13:0] updated_fh_res_hist_9_new_folded_hist_src_doubled = {
    updated_fh_res_hist_9_new_folded_hist_original_bits_masked__6,
    updated_fh_res_hist_9_new_folded_hist_original_bits_masked__5,
    updated_fh_res_hist_9_new_folded_hist_original_bits_masked__4,
    updated_fh_res_hist_9_new_folded_hist_original_bits_masked__3,
    updated_fh_res_hist_9_new_folded_hist_original_bits_masked__2,
    updated_fh_res_hist_9_new_folded_hist_original_bits_masked__1,
    updated_fh_res_hist_9_new_folded_hist_original_bits_masked__0,updated_fh_res_hist_9_new_folded_hist_xored}; // @[Cat.scala 31:58]
  wire [6:0] updated_fh_res_hist_9_new_folded_hist = updated_fh_res_hist_9_new_folded_hist_src_doubled[13:7]; // @[FrontendBundle.scala 221:30]
  wire  updated_fh_res_hist_10_new_folded_hist_original_bits_masked__0 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_10_folded_hist[0]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_10_new_folded_hist_original_bits_masked__1 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_10_folded_hist[1]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_10_new_folded_hist_original_bits_masked__2 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_10_folded_hist[2]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_10_new_folded_hist_original_bits_masked__3 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_10_folded_hist[3]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_10_new_folded_hist_original_bits_masked__4 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_10_folded_hist[4]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_10_new_folded_hist_original_bits_masked__5 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_10_folded_hist[5]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_10_new_folded_hist_original_bits_masked__6 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_10_folded_hist[6]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_10_new_folded_hist_original_bits_masked__7 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_10_folded_hist[7]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_10_new_folded_hist_original_bits_masked__8 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_10_folded_hist[8]; // @[FrontendBundle.scala 280:54]
  wire [8:0] updated_fh_res_hist_10_new_folded_hist_xored = {
    updated_fh_res_hist_10_new_folded_hist_original_bits_masked__8,
    updated_fh_res_hist_10_new_folded_hist_original_bits_masked__7,
    updated_fh_res_hist_10_new_folded_hist_original_bits_masked__6,
    updated_fh_res_hist_10_new_folded_hist_original_bits_masked__5,
    updated_fh_res_hist_10_new_folded_hist_original_bits_masked__4,
    updated_fh_res_hist_10_new_folded_hist_original_bits_masked__3,
    updated_fh_res_hist_10_new_folded_hist_original_bits_masked__2,
    updated_fh_res_hist_10_new_folded_hist_original_bits_masked__1,
    updated_fh_res_hist_10_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [17:0] updated_fh_res_hist_10_new_folded_hist_src_doubled = {
    updated_fh_res_hist_10_new_folded_hist_original_bits_masked__8,
    updated_fh_res_hist_10_new_folded_hist_original_bits_masked__7,
    updated_fh_res_hist_10_new_folded_hist_original_bits_masked__6,
    updated_fh_res_hist_10_new_folded_hist_original_bits_masked__5,
    updated_fh_res_hist_10_new_folded_hist_original_bits_masked__4,
    updated_fh_res_hist_10_new_folded_hist_original_bits_masked__3,
    updated_fh_res_hist_10_new_folded_hist_original_bits_masked__2,
    updated_fh_res_hist_10_new_folded_hist_original_bits_masked__1,
    updated_fh_res_hist_10_new_folded_hist_original_bits_masked__0,updated_fh_res_hist_10_new_folded_hist_xored}; // @[Cat.scala 31:58]
  wire [8:0] updated_fh_res_hist_10_new_folded_hist = updated_fh_res_hist_10_new_folded_hist_src_doubled[17:9]; // @[FrontendBundle.scala 221:30]
  wire [7:0] updated_fh_res_hist_11_new_folded_hist = do_redirect_bits_cfiUpdate_folded_hist_hist_11_folded_hist |
    _GEN_11935; // @[FrontendBundle.scala 290:29]
  wire  updated_fh_res_hist_12_new_folded_hist_original_bits_masked__0 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_12_folded_hist[0]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_12_new_folded_hist_original_bits_masked__1 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_12_folded_hist[1]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_12_new_folded_hist_original_bits_masked__2 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_12_folded_hist[2]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_12_new_folded_hist_original_bits_masked__3 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_12_folded_hist[3]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_12_new_folded_hist_original_bits_masked__4 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_12_folded_hist[4]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_12_new_folded_hist_original_bits_masked__5 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_12_folded_hist[5]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_12_new_folded_hist_original_bits_masked__6 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_12_folded_hist[6]; // @[FrontendBundle.scala 280:54]
  wire [6:0] updated_fh_res_hist_12_new_folded_hist_xored = {
    updated_fh_res_hist_12_new_folded_hist_original_bits_masked__6,
    updated_fh_res_hist_12_new_folded_hist_original_bits_masked__5,
    updated_fh_res_hist_12_new_folded_hist_original_bits_masked__4,
    updated_fh_res_hist_12_new_folded_hist_original_bits_masked__3,
    updated_fh_res_hist_12_new_folded_hist_original_bits_masked__2,
    updated_fh_res_hist_12_new_folded_hist_original_bits_masked__1,
    updated_fh_res_hist_12_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [13:0] updated_fh_res_hist_12_new_folded_hist_src_doubled = {
    updated_fh_res_hist_12_new_folded_hist_original_bits_masked__6,
    updated_fh_res_hist_12_new_folded_hist_original_bits_masked__5,
    updated_fh_res_hist_12_new_folded_hist_original_bits_masked__4,
    updated_fh_res_hist_12_new_folded_hist_original_bits_masked__3,
    updated_fh_res_hist_12_new_folded_hist_original_bits_masked__2,
    updated_fh_res_hist_12_new_folded_hist_original_bits_masked__1,
    updated_fh_res_hist_12_new_folded_hist_original_bits_masked__0,updated_fh_res_hist_12_new_folded_hist_xored}; // @[Cat.scala 31:58]
  wire [6:0] updated_fh_res_hist_12_new_folded_hist = updated_fh_res_hist_12_new_folded_hist_src_doubled[13:7]; // @[FrontendBundle.scala 221:30]
  wire  updated_fh_ob_10_0 = do_redirect_bits_cfiUpdate_lastBrNumOH[0] & do_redirect_bits_cfiUpdate_afhob_afhob_4_bits_0
     | do_redirect_bits_cfiUpdate_lastBrNumOH[1] & do_redirect_bits_cfiUpdate_afhob_afhob_4_bits_1 |
    do_redirect_bits_cfiUpdate_lastBrNumOH[2] & do_redirect_bits_cfiUpdate_afhob_afhob_4_bits_2; // @[Mux.scala 27:73]
  wire  updated_fh_res_hist_13_new_folded_hist_original_bits_masked__0 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_13_folded_hist[0]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_13_new_folded_hist_original_bits_masked__1 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_13_folded_hist[1]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_13_new_folded_hist_original_bits_masked__2 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_13_folded_hist[2]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_13_new_folded_hist_original_bits_masked__3 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_13_folded_hist[3]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_13_new_folded_hist_original_bits_masked__4 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_13_folded_hist[4]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_13_new_folded_hist_original_bits_masked__5 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_13_folded_hist[5]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_13_new_folded_hist_original_bits_masked__6 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_13_folded_hist[6]; // @[FrontendBundle.scala 280:54]
  wire [6:0] updated_fh_res_hist_13_new_folded_hist_xored = {
    updated_fh_res_hist_13_new_folded_hist_original_bits_masked__6,
    updated_fh_res_hist_13_new_folded_hist_original_bits_masked__5,
    updated_fh_res_hist_13_new_folded_hist_original_bits_masked__4,
    updated_fh_res_hist_13_new_folded_hist_original_bits_masked__3,
    updated_fh_res_hist_13_new_folded_hist_original_bits_masked__2,
    updated_fh_res_hist_13_new_folded_hist_original_bits_masked__1,
    updated_fh_res_hist_13_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [13:0] updated_fh_res_hist_13_new_folded_hist_src_doubled = {
    updated_fh_res_hist_13_new_folded_hist_original_bits_masked__6,
    updated_fh_res_hist_13_new_folded_hist_original_bits_masked__5,
    updated_fh_res_hist_13_new_folded_hist_original_bits_masked__4,
    updated_fh_res_hist_13_new_folded_hist_original_bits_masked__3,
    updated_fh_res_hist_13_new_folded_hist_original_bits_masked__2,
    updated_fh_res_hist_13_new_folded_hist_original_bits_masked__1,
    updated_fh_res_hist_13_new_folded_hist_original_bits_masked__0,updated_fh_res_hist_13_new_folded_hist_xored}; // @[Cat.scala 31:58]
  wire [6:0] updated_fh_res_hist_13_new_folded_hist = updated_fh_res_hist_13_new_folded_hist_src_doubled[13:7]; // @[FrontendBundle.scala 221:30]
  wire  updated_fh_res_hist_14_new_folded_hist_original_bits_masked__0 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_14_folded_hist[0]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_14_new_folded_hist_original_bits_masked__1 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_14_folded_hist[1]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_14_new_folded_hist_original_bits_masked__2 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_14_folded_hist[2]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_14_new_folded_hist_original_bits_masked__3 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_14_folded_hist[3]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_14_new_folded_hist_original_bits_masked__4 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_14_folded_hist[4]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_14_new_folded_hist_original_bits_masked__5 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_14_folded_hist[5]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_14_new_folded_hist_original_bits_masked__6 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_14_folded_hist[6]; // @[FrontendBundle.scala 280:54]
  wire [6:0] updated_fh_res_hist_14_new_folded_hist_xored = {
    updated_fh_res_hist_14_new_folded_hist_original_bits_masked__6,
    updated_fh_res_hist_14_new_folded_hist_original_bits_masked__5,
    updated_fh_res_hist_14_new_folded_hist_original_bits_masked__4,
    updated_fh_res_hist_14_new_folded_hist_original_bits_masked__3,
    updated_fh_res_hist_14_new_folded_hist_original_bits_masked__2,
    updated_fh_res_hist_14_new_folded_hist_original_bits_masked__1,
    updated_fh_res_hist_14_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [13:0] updated_fh_res_hist_14_new_folded_hist_src_doubled = {
    updated_fh_res_hist_14_new_folded_hist_original_bits_masked__6,
    updated_fh_res_hist_14_new_folded_hist_original_bits_masked__5,
    updated_fh_res_hist_14_new_folded_hist_original_bits_masked__4,
    updated_fh_res_hist_14_new_folded_hist_original_bits_masked__3,
    updated_fh_res_hist_14_new_folded_hist_original_bits_masked__2,
    updated_fh_res_hist_14_new_folded_hist_original_bits_masked__1,
    updated_fh_res_hist_14_new_folded_hist_original_bits_masked__0,updated_fh_res_hist_14_new_folded_hist_xored}; // @[Cat.scala 31:58]
  wire [6:0] updated_fh_res_hist_14_new_folded_hist = updated_fh_res_hist_14_new_folded_hist_src_doubled[13:7]; // @[FrontendBundle.scala 221:30]
  wire  updated_fh_res_hist_15_new_folded_hist_original_bits_masked__0 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_15_folded_hist[0]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_15_new_folded_hist_original_bits_masked__1 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_15_folded_hist[1]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_15_new_folded_hist_original_bits_masked__2 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_15_folded_hist[2]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_15_new_folded_hist_original_bits_masked__3 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_15_folded_hist[3]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_15_new_folded_hist_original_bits_masked__4 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_15_folded_hist[4]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_15_new_folded_hist_original_bits_masked__5 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_15_folded_hist[5]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_15_new_folded_hist_original_bits_masked__6 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_15_folded_hist[6]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_15_new_folded_hist_original_bits_masked__7 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_15_folded_hist[7]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_15_new_folded_hist_original_bits_masked__8 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_15_folded_hist[8]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_15_new_folded_hist_original_bits_masked__9 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_15_folded_hist[9]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_15_new_folded_hist_original_bits_masked__10 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_15_folded_hist[10]; // @[FrontendBundle.scala 280:54]
  wire [4:0] updated_fh_res_hist_15_new_folded_hist_xored_lo = {
    updated_fh_res_hist_15_new_folded_hist_original_bits_masked__4,
    updated_fh_res_hist_15_new_folded_hist_original_bits_masked__3,
    updated_fh_res_hist_15_new_folded_hist_original_bits_masked__2,
    updated_fh_res_hist_15_new_folded_hist_original_bits_masked__1,
    updated_fh_res_hist_15_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [10:0] updated_fh_res_hist_15_new_folded_hist_xored = {
    updated_fh_res_hist_15_new_folded_hist_original_bits_masked__10,
    updated_fh_res_hist_15_new_folded_hist_original_bits_masked__9,
    updated_fh_res_hist_15_new_folded_hist_original_bits_masked__8,
    updated_fh_res_hist_15_new_folded_hist_original_bits_masked__7,
    updated_fh_res_hist_15_new_folded_hist_original_bits_masked__6,
    updated_fh_res_hist_15_new_folded_hist_original_bits_masked__5,updated_fh_res_hist_15_new_folded_hist_xored_lo}; // @[FrontendBundle.scala 258:11]
  wire [21:0] updated_fh_res_hist_15_new_folded_hist_src_doubled = {
    updated_fh_res_hist_15_new_folded_hist_original_bits_masked__10,
    updated_fh_res_hist_15_new_folded_hist_original_bits_masked__9,
    updated_fh_res_hist_15_new_folded_hist_original_bits_masked__8,
    updated_fh_res_hist_15_new_folded_hist_original_bits_masked__7,
    updated_fh_res_hist_15_new_folded_hist_original_bits_masked__6,
    updated_fh_res_hist_15_new_folded_hist_original_bits_masked__5,updated_fh_res_hist_15_new_folded_hist_xored_lo,
    updated_fh_res_hist_15_new_folded_hist_xored}; // @[Cat.scala 31:58]
  wire [10:0] updated_fh_res_hist_15_new_folded_hist = updated_fh_res_hist_15_new_folded_hist_src_doubled[21:11]; // @[FrontendBundle.scala 221:30]
  wire  updated_fh_ob_13_0 = do_redirect_bits_cfiUpdate_lastBrNumOH[0] & do_redirect_bits_cfiUpdate_afhob_afhob_0_bits_0
     | do_redirect_bits_cfiUpdate_lastBrNumOH[1] & do_redirect_bits_cfiUpdate_afhob_afhob_0_bits_1 |
    do_redirect_bits_cfiUpdate_lastBrNumOH[2] & do_redirect_bits_cfiUpdate_afhob_afhob_0_bits_2; // @[Mux.scala 27:73]
  wire  updated_fh_ob_13_1 = do_redirect_bits_cfiUpdate_lastBrNumOH[0] & do_redirect_bits_cfiUpdate_afhob_afhob_0_bits_1
     | do_redirect_bits_cfiUpdate_lastBrNumOH[1] & do_redirect_bits_cfiUpdate_afhob_afhob_0_bits_2 |
    do_redirect_bits_cfiUpdate_lastBrNumOH[2] & do_redirect_bits_cfiUpdate_afhob_afhob_0_bits_3; // @[Mux.scala 27:73]
  wire  updated_fh_res_hist_16_new_folded_hist_original_bits_masked__0 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_16_folded_hist[0]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_16_new_folded_hist_original_bits_masked__1 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_16_folded_hist[1]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_16_new_folded_hist_original_bits_masked__2 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_16_folded_hist[2]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_16_new_folded_hist_original_bits_masked__3 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_16_folded_hist[3]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_16_new_folded_hist_original_bits_masked__4 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_16_folded_hist[4]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_16_new_folded_hist_original_bits_masked__5 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_16_folded_hist[5]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_16_new_folded_hist_original_bits_masked__6 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_16_folded_hist[6]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_16_new_folded_hist_original_bits_masked__7 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_16_folded_hist[7]; // @[FrontendBundle.scala 280:54]
  wire [7:0] updated_fh_res_hist_16_new_folded_hist_xored = {
    updated_fh_res_hist_16_new_folded_hist_original_bits_masked__7,
    updated_fh_res_hist_16_new_folded_hist_original_bits_masked__6,
    updated_fh_res_hist_16_new_folded_hist_original_bits_masked__5,
    updated_fh_res_hist_16_new_folded_hist_original_bits_masked__4,
    updated_fh_res_hist_16_new_folded_hist_original_bits_masked__3,
    updated_fh_res_hist_16_new_folded_hist_original_bits_masked__2,
    updated_fh_res_hist_16_new_folded_hist_original_bits_masked__1,
    updated_fh_res_hist_16_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [15:0] updated_fh_res_hist_16_new_folded_hist_src_doubled = {
    updated_fh_res_hist_16_new_folded_hist_original_bits_masked__7,
    updated_fh_res_hist_16_new_folded_hist_original_bits_masked__6,
    updated_fh_res_hist_16_new_folded_hist_original_bits_masked__5,
    updated_fh_res_hist_16_new_folded_hist_original_bits_masked__4,
    updated_fh_res_hist_16_new_folded_hist_original_bits_masked__3,
    updated_fh_res_hist_16_new_folded_hist_original_bits_masked__2,
    updated_fh_res_hist_16_new_folded_hist_original_bits_masked__1,
    updated_fh_res_hist_16_new_folded_hist_original_bits_masked__0,updated_fh_res_hist_16_new_folded_hist_xored}; // @[Cat.scala 31:58]
  wire [7:0] updated_fh_res_hist_16_new_folded_hist = updated_fh_res_hist_16_new_folded_hist_src_doubled[15:8]; // @[FrontendBundle.scala 221:30]
  wire  updated_fh_res_hist_17_new_folded_hist_original_bits_masked__0 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_17_folded_hist[0]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_17_new_folded_hist_original_bits_masked__1 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_17_folded_hist[1]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_17_new_folded_hist_original_bits_masked__2 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_17_folded_hist[2]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_17_new_folded_hist_original_bits_masked__3 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_17_folded_hist[3]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_17_new_folded_hist_original_bits_masked__4 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_17_folded_hist[4]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_17_new_folded_hist_original_bits_masked__5 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_17_folded_hist[5]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_17_new_folded_hist_original_bits_masked__6 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_17_folded_hist[6]; // @[FrontendBundle.scala 280:54]
  wire  updated_fh_res_hist_17_new_folded_hist_original_bits_masked__7 =
    do_redirect_bits_cfiUpdate_folded_hist_hist_17_folded_hist[7]; // @[FrontendBundle.scala 280:54]
  wire [7:0] updated_fh_res_hist_17_new_folded_hist_xored = {
    updated_fh_res_hist_17_new_folded_hist_original_bits_masked__7,
    updated_fh_res_hist_17_new_folded_hist_original_bits_masked__6,
    updated_fh_res_hist_17_new_folded_hist_original_bits_masked__5,
    updated_fh_res_hist_17_new_folded_hist_original_bits_masked__4,
    updated_fh_res_hist_17_new_folded_hist_original_bits_masked__3,
    updated_fh_res_hist_17_new_folded_hist_original_bits_masked__2,
    updated_fh_res_hist_17_new_folded_hist_original_bits_masked__1,
    updated_fh_res_hist_17_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [15:0] updated_fh_res_hist_17_new_folded_hist_src_doubled = {
    updated_fh_res_hist_17_new_folded_hist_original_bits_masked__7,
    updated_fh_res_hist_17_new_folded_hist_original_bits_masked__6,
    updated_fh_res_hist_17_new_folded_hist_original_bits_masked__5,
    updated_fh_res_hist_17_new_folded_hist_original_bits_masked__4,
    updated_fh_res_hist_17_new_folded_hist_original_bits_masked__3,
    updated_fh_res_hist_17_new_folded_hist_original_bits_masked__2,
    updated_fh_res_hist_17_new_folded_hist_original_bits_masked__1,
    updated_fh_res_hist_17_new_folded_hist_original_bits_masked__0,updated_fh_res_hist_17_new_folded_hist_xored}; // @[Cat.scala 31:58]
  wire [7:0] updated_fh_res_hist_17_new_folded_hist = updated_fh_res_hist_17_new_folded_hist_src_doubled[15:8]; // @[FrontendBundle.scala 221:30]
  wire [1:0] updated_fh_res_hist_0_new_folded_hist_newest_bits_masked_1 = {1'h0,_updated_fh_T}; // @[FrontendBundle.scala 274:102]
  wire  updated_fh_res_hist_0_new_folded_hist_xored_res_1_6 = updated_fh_res_hist_0_new_folded_hist_newest_bits_masked_1
    [1] ^ updated_fh_res_hist_0_new_folded_hist_original_bits_masked__6; // @[FrontendBundle.scala 256:48]
  wire  updated_fh_res_hist_0_new_folded_hist_xored_res_1_7 = updated_fh_res_hist_0_new_folded_hist_newest_bits_masked_1
    [0] ^ updated_fh_ob__0 ^ updated_fh_res_hist_0_new_folded_hist_original_bits_masked__7; // @[FrontendBundle.scala 256:48]
  wire [7:0] updated_fh_res_hist_0_new_folded_hist_xored_1 = {updated_fh_res_hist_0_new_folded_hist_xored_res_1_7,
    updated_fh_res_hist_0_new_folded_hist_xored_res_1_6,updated_fh_res_hist_0_new_folded_hist_original_bits_masked__5,
    updated_fh_res_hist_0_new_folded_hist_original_bits_masked__4,
    updated_fh_res_hist_0_new_folded_hist_original_bits_masked__3,
    updated_fh_res_hist_0_new_folded_hist_original_bits_masked__2,
    updated_fh_res_hist_0_new_folded_hist_original_bits_masked__1,
    updated_fh_res_hist_0_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [15:0] updated_fh_res_hist_0_new_folded_hist_src_doubled_1 = {updated_fh_res_hist_0_new_folded_hist_xored_res_1_7
    ,updated_fh_res_hist_0_new_folded_hist_xored_res_1_6,updated_fh_res_hist_0_new_folded_hist_original_bits_masked__5,
    updated_fh_res_hist_0_new_folded_hist_original_bits_masked__4,
    updated_fh_res_hist_0_new_folded_hist_original_bits_masked__3,
    updated_fh_res_hist_0_new_folded_hist_original_bits_masked__2,
    updated_fh_res_hist_0_new_folded_hist_original_bits_masked__1,
    updated_fh_res_hist_0_new_folded_hist_original_bits_masked__0,updated_fh_res_hist_0_new_folded_hist_xored_1}; // @[Cat.scala 31:58]
  wire [7:0] updated_fh_res_hist_0_new_folded_hist_1 = updated_fh_res_hist_0_new_folded_hist_src_doubled_1[14:7]; // @[FrontendBundle.scala 221:30]
  wire  updated_fh_res_hist_1_new_folded_hist_xored_res_1_6 = updated_fh_res_hist_0_new_folded_hist_newest_bits_masked_1
    [1] ^ updated_fh_res_hist_1_new_folded_hist_original_bits_masked__6; // @[FrontendBundle.scala 256:48]
  wire  updated_fh_res_hist_1_new_folded_hist_xored_res_1_7 = updated_fh_res_hist_0_new_folded_hist_newest_bits_masked_1
    [0] ^ updated_fh_ob_1_0 ^ updated_fh_res_hist_1_new_folded_hist_original_bits_masked__7; // @[FrontendBundle.scala 256:48]
  wire [7:0] updated_fh_res_hist_1_new_folded_hist_xored_1 = {updated_fh_res_hist_1_new_folded_hist_xored_res_1_7,
    updated_fh_res_hist_1_new_folded_hist_xored_res_1_6,updated_fh_res_hist_1_new_folded_hist_original_bits_masked__5,
    updated_fh_res_hist_1_new_folded_hist_original_bits_masked__4,
    updated_fh_res_hist_1_new_folded_hist_original_bits_masked__3,
    updated_fh_res_hist_1_new_folded_hist_original_bits_masked__2,
    updated_fh_res_hist_1_new_folded_hist_original_bits_masked__1,
    updated_fh_res_hist_1_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [15:0] updated_fh_res_hist_1_new_folded_hist_src_doubled_1 = {updated_fh_res_hist_1_new_folded_hist_xored_res_1_7
    ,updated_fh_res_hist_1_new_folded_hist_xored_res_1_6,updated_fh_res_hist_1_new_folded_hist_original_bits_masked__5,
    updated_fh_res_hist_1_new_folded_hist_original_bits_masked__4,
    updated_fh_res_hist_1_new_folded_hist_original_bits_masked__3,
    updated_fh_res_hist_1_new_folded_hist_original_bits_masked__2,
    updated_fh_res_hist_1_new_folded_hist_original_bits_masked__1,
    updated_fh_res_hist_1_new_folded_hist_original_bits_masked__0,updated_fh_res_hist_1_new_folded_hist_xored_1}; // @[Cat.scala 31:58]
  wire [7:0] updated_fh_res_hist_1_new_folded_hist_1 = updated_fh_res_hist_1_new_folded_hist_src_doubled_1[14:7]; // @[FrontendBundle.scala 221:30]
  wire  updated_fh_res_hist_2_new_folded_hist_xored_res_1_6 = updated_fh_res_hist_0_new_folded_hist_newest_bits_masked_1
    [1] ^ updated_fh_ob_2_0 ^ updated_fh_res_hist_2_new_folded_hist_original_bits_masked__6; // @[FrontendBundle.scala 256:48]
  wire  updated_fh_res_hist_2_new_folded_hist_xored_res_1_7 = updated_fh_res_hist_0_new_folded_hist_newest_bits_masked_1
    [0] ^ updated_fh_res_hist_2_new_folded_hist_original_bits_masked__7; // @[FrontendBundle.scala 256:48]
  wire [7:0] updated_fh_res_hist_2_new_folded_hist_xored_1 = {updated_fh_res_hist_2_new_folded_hist_xored_res_1_7,
    updated_fh_res_hist_2_new_folded_hist_xored_res_1_6,updated_fh_res_hist_2_new_folded_hist_original_bits_masked__5,
    updated_fh_res_hist_2_new_folded_hist_original_bits_masked__4,
    updated_fh_res_hist_2_new_folded_hist_original_bits_masked__3,
    updated_fh_res_hist_2_new_folded_hist_original_bits_masked__2,
    updated_fh_res_hist_2_new_folded_hist_original_bits_masked__1,
    updated_fh_res_hist_2_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [15:0] updated_fh_res_hist_2_new_folded_hist_src_doubled_1 = {updated_fh_res_hist_2_new_folded_hist_xored_res_1_7
    ,updated_fh_res_hist_2_new_folded_hist_xored_res_1_6,updated_fh_res_hist_2_new_folded_hist_original_bits_masked__5,
    updated_fh_res_hist_2_new_folded_hist_original_bits_masked__4,
    updated_fh_res_hist_2_new_folded_hist_original_bits_masked__3,
    updated_fh_res_hist_2_new_folded_hist_original_bits_masked__2,
    updated_fh_res_hist_2_new_folded_hist_original_bits_masked__1,
    updated_fh_res_hist_2_new_folded_hist_original_bits_masked__0,updated_fh_res_hist_2_new_folded_hist_xored_1}; // @[Cat.scala 31:58]
  wire [7:0] updated_fh_res_hist_2_new_folded_hist_1 = updated_fh_res_hist_2_new_folded_hist_src_doubled_1[14:7]; // @[FrontendBundle.scala 221:30]
  wire  updated_fh_res_hist_3_new_folded_hist_xored_res_1_9 = updated_fh_res_hist_0_new_folded_hist_newest_bits_masked_1
    [1] ^ updated_fh_ob_1_0 ^ updated_fh_res_hist_3_new_folded_hist_original_bits_masked__9; // @[FrontendBundle.scala 256:48]
  wire  updated_fh_res_hist_3_new_folded_hist_xored_res_1_10 =
    updated_fh_res_hist_0_new_folded_hist_newest_bits_masked_1[0] ^
    updated_fh_res_hist_3_new_folded_hist_original_bits_masked__10; // @[FrontendBundle.scala 256:48]
  wire [10:0] updated_fh_res_hist_3_new_folded_hist_xored_1 = {updated_fh_res_hist_3_new_folded_hist_xored_res_1_10,
    updated_fh_res_hist_3_new_folded_hist_xored_res_1_9,updated_fh_res_hist_3_new_folded_hist_original_bits_masked__8,
    updated_fh_res_hist_3_new_folded_hist_original_bits_masked__7,
    updated_fh_res_hist_3_new_folded_hist_original_bits_masked__6,
    updated_fh_res_hist_3_new_folded_hist_original_bits_masked__5,updated_fh_res_hist_3_new_folded_hist_xored_lo}; // @[FrontendBundle.scala 258:11]
  wire [21:0] updated_fh_res_hist_3_new_folded_hist_src_doubled_1 = {
    updated_fh_res_hist_3_new_folded_hist_xored_res_1_10,updated_fh_res_hist_3_new_folded_hist_xored_res_1_9,
    updated_fh_res_hist_3_new_folded_hist_original_bits_masked__8,
    updated_fh_res_hist_3_new_folded_hist_original_bits_masked__7,
    updated_fh_res_hist_3_new_folded_hist_original_bits_masked__6,
    updated_fh_res_hist_3_new_folded_hist_original_bits_masked__5,updated_fh_res_hist_3_new_folded_hist_xored_lo,
    updated_fh_res_hist_3_new_folded_hist_xored_1}; // @[Cat.scala 31:58]
  wire [10:0] updated_fh_res_hist_3_new_folded_hist_1 = updated_fh_res_hist_3_new_folded_hist_src_doubled_1[20:10]; // @[FrontendBundle.scala 221:30]
  wire [4:0] _updated_fh_res_hist_4_new_folded_hist_T_2 = {do_redirect_bits_cfiUpdate_folded_hist_hist_4_folded_hist
    , 1'h0}; // @[FrontendBundle.scala 290:21]
  wire [4:0] _GEN_11937 = {{4'd0}, _updated_fh_T}; // @[FrontendBundle.scala 290:29]
  wire [4:0] _updated_fh_res_hist_4_new_folded_hist_T_3 = _updated_fh_res_hist_4_new_folded_hist_T_2 | _GEN_11937; // @[FrontendBundle.scala 290:29]
  wire [3:0] updated_fh_res_hist_4_new_folded_hist_1 = _updated_fh_res_hist_4_new_folded_hist_T_3[3:0]; // @[FrontendBundle.scala 290:37]
  wire  updated_fh_res_hist_5_new_folded_hist_xored_res_1_1 = updated_fh_ob_4_0 ^
    updated_fh_res_hist_5_new_folded_hist_original_bits_masked__1; // @[FrontendBundle.scala 256:48]
  wire  updated_fh_res_hist_5_new_folded_hist_xored_res_1_9 = updated_fh_res_hist_0_new_folded_hist_newest_bits_masked_1
    [1] ^ updated_fh_res_hist_5_new_folded_hist_original_bits_masked__9; // @[FrontendBundle.scala 256:48]
  wire  updated_fh_res_hist_5_new_folded_hist_xored_res_1_10 =
    updated_fh_res_hist_0_new_folded_hist_newest_bits_masked_1[0] ^
    updated_fh_res_hist_5_new_folded_hist_original_bits_masked__10; // @[FrontendBundle.scala 256:48]
  wire [4:0] updated_fh_res_hist_5_new_folded_hist_xored_lo_1 = {
    updated_fh_res_hist_5_new_folded_hist_original_bits_masked__4,
    updated_fh_res_hist_5_new_folded_hist_original_bits_masked__3,
    updated_fh_res_hist_5_new_folded_hist_original_bits_masked__2,updated_fh_res_hist_5_new_folded_hist_xored_res_1_1,
    updated_fh_res_hist_5_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [10:0] updated_fh_res_hist_5_new_folded_hist_xored_1 = {updated_fh_res_hist_5_new_folded_hist_xored_res_1_10,
    updated_fh_res_hist_5_new_folded_hist_xored_res_1_9,updated_fh_res_hist_5_new_folded_hist_original_bits_masked__8,
    updated_fh_res_hist_5_new_folded_hist_original_bits_masked__7,
    updated_fh_res_hist_5_new_folded_hist_original_bits_masked__6,
    updated_fh_res_hist_5_new_folded_hist_original_bits_masked__5,updated_fh_res_hist_5_new_folded_hist_xored_lo_1}; // @[FrontendBundle.scala 258:11]
  wire [21:0] updated_fh_res_hist_5_new_folded_hist_src_doubled_1 = {
    updated_fh_res_hist_5_new_folded_hist_xored_res_1_10,updated_fh_res_hist_5_new_folded_hist_xored_res_1_9,
    updated_fh_res_hist_5_new_folded_hist_original_bits_masked__8,
    updated_fh_res_hist_5_new_folded_hist_original_bits_masked__7,
    updated_fh_res_hist_5_new_folded_hist_original_bits_masked__6,
    updated_fh_res_hist_5_new_folded_hist_original_bits_masked__5,updated_fh_res_hist_5_new_folded_hist_xored_lo_1,
    updated_fh_res_hist_5_new_folded_hist_xored_1}; // @[Cat.scala 31:58]
  wire [10:0] updated_fh_res_hist_5_new_folded_hist_1 = updated_fh_res_hist_5_new_folded_hist_src_doubled_1[20:10]; // @[FrontendBundle.scala 221:30]
  wire  updated_fh_res_hist_6_new_folded_hist_xored_res_1_3 = updated_fh_ob_4_0 ^
    updated_fh_res_hist_6_new_folded_hist_original_bits_masked__3; // @[FrontendBundle.scala 256:48]
  wire  updated_fh_res_hist_6_new_folded_hist_xored_res_1_7 = updated_fh_res_hist_0_new_folded_hist_newest_bits_masked_1
    [1] ^ updated_fh_res_hist_6_new_folded_hist_original_bits_masked__7; // @[FrontendBundle.scala 256:48]
  wire  updated_fh_res_hist_6_new_folded_hist_xored_res_1_8 = updated_fh_res_hist_0_new_folded_hist_newest_bits_masked_1
    [0] ^ updated_fh_res_hist_6_new_folded_hist_original_bits_masked__8; // @[FrontendBundle.scala 256:48]
  wire [8:0] updated_fh_res_hist_6_new_folded_hist_xored_1 = {updated_fh_res_hist_6_new_folded_hist_xored_res_1_8,
    updated_fh_res_hist_6_new_folded_hist_xored_res_1_7,updated_fh_res_hist_6_new_folded_hist_original_bits_masked__6,
    updated_fh_res_hist_6_new_folded_hist_original_bits_masked__5,
    updated_fh_res_hist_6_new_folded_hist_original_bits_masked__4,updated_fh_res_hist_6_new_folded_hist_xored_res_1_3,
    updated_fh_res_hist_6_new_folded_hist_original_bits_masked__2,
    updated_fh_res_hist_6_new_folded_hist_original_bits_masked__1,
    updated_fh_res_hist_6_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [17:0] updated_fh_res_hist_6_new_folded_hist_src_doubled_1 = {updated_fh_res_hist_6_new_folded_hist_xored_res_1_8
    ,updated_fh_res_hist_6_new_folded_hist_xored_res_1_7,updated_fh_res_hist_6_new_folded_hist_original_bits_masked__6,
    updated_fh_res_hist_6_new_folded_hist_original_bits_masked__5,
    updated_fh_res_hist_6_new_folded_hist_original_bits_masked__4,updated_fh_res_hist_6_new_folded_hist_xored_res_1_3,
    updated_fh_res_hist_6_new_folded_hist_original_bits_masked__2,
    updated_fh_res_hist_6_new_folded_hist_original_bits_masked__1,
    updated_fh_res_hist_6_new_folded_hist_original_bits_masked__0,updated_fh_res_hist_6_new_folded_hist_xored_1}; // @[Cat.scala 31:58]
  wire [8:0] updated_fh_res_hist_6_new_folded_hist_1 = updated_fh_res_hist_6_new_folded_hist_src_doubled_1[16:8]; // @[FrontendBundle.scala 221:30]
  wire  updated_fh_res_hist_7_new_folded_hist_xored_res_1_6 = updated_fh_ob__0 ^
    updated_fh_res_hist_7_new_folded_hist_original_bits_masked__6; // @[FrontendBundle.scala 256:48]
  wire  updated_fh_res_hist_7_new_folded_hist_xored_res_1_7 = updated_fh_res_hist_0_new_folded_hist_newest_bits_masked_1
    [1] ^ updated_fh_res_hist_7_new_folded_hist_original_bits_masked__7; // @[FrontendBundle.scala 256:48]
  wire  updated_fh_res_hist_7_new_folded_hist_xored_res_1_8 = updated_fh_res_hist_0_new_folded_hist_newest_bits_masked_1
    [0] ^ updated_fh_res_hist_7_new_folded_hist_original_bits_masked__8; // @[FrontendBundle.scala 256:48]
  wire [8:0] updated_fh_res_hist_7_new_folded_hist_xored_1 = {updated_fh_res_hist_7_new_folded_hist_xored_res_1_8,
    updated_fh_res_hist_7_new_folded_hist_xored_res_1_7,updated_fh_res_hist_7_new_folded_hist_xored_res_1_6,
    updated_fh_res_hist_7_new_folded_hist_original_bits_masked__5,
    updated_fh_res_hist_7_new_folded_hist_original_bits_masked__4,
    updated_fh_res_hist_7_new_folded_hist_original_bits_masked__3,
    updated_fh_res_hist_7_new_folded_hist_original_bits_masked__2,
    updated_fh_res_hist_7_new_folded_hist_original_bits_masked__1,
    updated_fh_res_hist_7_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [17:0] updated_fh_res_hist_7_new_folded_hist_src_doubled_1 = {updated_fh_res_hist_7_new_folded_hist_xored_res_1_8
    ,updated_fh_res_hist_7_new_folded_hist_xored_res_1_7,updated_fh_res_hist_7_new_folded_hist_xored_res_1_6,
    updated_fh_res_hist_7_new_folded_hist_original_bits_masked__5,
    updated_fh_res_hist_7_new_folded_hist_original_bits_masked__4,
    updated_fh_res_hist_7_new_folded_hist_original_bits_masked__3,
    updated_fh_res_hist_7_new_folded_hist_original_bits_masked__2,
    updated_fh_res_hist_7_new_folded_hist_original_bits_masked__1,
    updated_fh_res_hist_7_new_folded_hist_original_bits_masked__0,updated_fh_res_hist_7_new_folded_hist_xored_1}; // @[Cat.scala 31:58]
  wire [8:0] updated_fh_res_hist_7_new_folded_hist_1 = updated_fh_res_hist_7_new_folded_hist_src_doubled_1[16:8]; // @[FrontendBundle.scala 221:30]
  wire [8:0] _updated_fh_res_hist_8_new_folded_hist_T_2 = {do_redirect_bits_cfiUpdate_folded_hist_hist_8_folded_hist
    , 1'h0}; // @[FrontendBundle.scala 290:21]
  wire [8:0] _GEN_11938 = {{8'd0}, _updated_fh_T}; // @[FrontendBundle.scala 290:29]
  wire [8:0] _updated_fh_res_hist_8_new_folded_hist_T_3 = _updated_fh_res_hist_8_new_folded_hist_T_2 | _GEN_11938; // @[FrontendBundle.scala 290:29]
  wire [7:0] updated_fh_res_hist_8_new_folded_hist_1 = _updated_fh_res_hist_8_new_folded_hist_T_3[7:0]; // @[FrontendBundle.scala 290:37]
  wire  updated_fh_res_hist_9_new_folded_hist_xored_res_1_3 = updated_fh_ob_1_0 ^
    updated_fh_res_hist_9_new_folded_hist_original_bits_masked__3; // @[FrontendBundle.scala 256:48]
  wire  updated_fh_res_hist_9_new_folded_hist_xored_res_1_5 = updated_fh_res_hist_0_new_folded_hist_newest_bits_masked_1
    [1] ^ updated_fh_res_hist_9_new_folded_hist_original_bits_masked__5; // @[FrontendBundle.scala 256:48]
  wire  updated_fh_res_hist_9_new_folded_hist_xored_res_1_6 = updated_fh_res_hist_0_new_folded_hist_newest_bits_masked_1
    [0] ^ updated_fh_res_hist_9_new_folded_hist_original_bits_masked__6; // @[FrontendBundle.scala 256:48]
  wire [6:0] updated_fh_res_hist_9_new_folded_hist_xored_1 = {updated_fh_res_hist_9_new_folded_hist_xored_res_1_6,
    updated_fh_res_hist_9_new_folded_hist_xored_res_1_5,updated_fh_res_hist_9_new_folded_hist_original_bits_masked__4,
    updated_fh_res_hist_9_new_folded_hist_xored_res_1_3,updated_fh_res_hist_9_new_folded_hist_original_bits_masked__2,
    updated_fh_res_hist_9_new_folded_hist_original_bits_masked__1,
    updated_fh_res_hist_9_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [13:0] updated_fh_res_hist_9_new_folded_hist_src_doubled_1 = {updated_fh_res_hist_9_new_folded_hist_xored_res_1_6
    ,updated_fh_res_hist_9_new_folded_hist_xored_res_1_5,updated_fh_res_hist_9_new_folded_hist_original_bits_masked__4,
    updated_fh_res_hist_9_new_folded_hist_xored_res_1_3,updated_fh_res_hist_9_new_folded_hist_original_bits_masked__2,
    updated_fh_res_hist_9_new_folded_hist_original_bits_masked__1,
    updated_fh_res_hist_9_new_folded_hist_original_bits_masked__0,updated_fh_res_hist_9_new_folded_hist_xored_1}; // @[Cat.scala 31:58]
  wire [6:0] updated_fh_res_hist_9_new_folded_hist_1 = updated_fh_res_hist_9_new_folded_hist_src_doubled_1[12:6]; // @[FrontendBundle.scala 221:30]
  wire  updated_fh_res_hist_10_new_folded_hist_xored_res_1_4 = updated_fh_ob_1_0 ^
    updated_fh_res_hist_10_new_folded_hist_original_bits_masked__4; // @[FrontendBundle.scala 256:48]
  wire  updated_fh_res_hist_10_new_folded_hist_xored_res_1_7 =
    updated_fh_res_hist_0_new_folded_hist_newest_bits_masked_1[1] ^
    updated_fh_res_hist_10_new_folded_hist_original_bits_masked__7; // @[FrontendBundle.scala 256:48]
  wire  updated_fh_res_hist_10_new_folded_hist_xored_res_1_8 =
    updated_fh_res_hist_0_new_folded_hist_newest_bits_masked_1[0] ^
    updated_fh_res_hist_10_new_folded_hist_original_bits_masked__8; // @[FrontendBundle.scala 256:48]
  wire [8:0] updated_fh_res_hist_10_new_folded_hist_xored_1 = {updated_fh_res_hist_10_new_folded_hist_xored_res_1_8,
    updated_fh_res_hist_10_new_folded_hist_xored_res_1_7,updated_fh_res_hist_10_new_folded_hist_original_bits_masked__6,
    updated_fh_res_hist_10_new_folded_hist_original_bits_masked__5,updated_fh_res_hist_10_new_folded_hist_xored_res_1_4,
    updated_fh_res_hist_10_new_folded_hist_original_bits_masked__3,
    updated_fh_res_hist_10_new_folded_hist_original_bits_masked__2,
    updated_fh_res_hist_10_new_folded_hist_original_bits_masked__1,
    updated_fh_res_hist_10_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [17:0] updated_fh_res_hist_10_new_folded_hist_src_doubled_1 = {
    updated_fh_res_hist_10_new_folded_hist_xored_res_1_8,updated_fh_res_hist_10_new_folded_hist_xored_res_1_7,
    updated_fh_res_hist_10_new_folded_hist_original_bits_masked__6,
    updated_fh_res_hist_10_new_folded_hist_original_bits_masked__5,updated_fh_res_hist_10_new_folded_hist_xored_res_1_4,
    updated_fh_res_hist_10_new_folded_hist_original_bits_masked__3,
    updated_fh_res_hist_10_new_folded_hist_original_bits_masked__2,
    updated_fh_res_hist_10_new_folded_hist_original_bits_masked__1,
    updated_fh_res_hist_10_new_folded_hist_original_bits_masked__0,updated_fh_res_hist_10_new_folded_hist_xored_1}; // @[Cat.scala 31:58]
  wire [8:0] updated_fh_res_hist_10_new_folded_hist_1 = updated_fh_res_hist_10_new_folded_hist_src_doubled_1[16:8]; // @[FrontendBundle.scala 221:30]
  wire [8:0] _updated_fh_res_hist_11_new_folded_hist_T_2 = {do_redirect_bits_cfiUpdate_folded_hist_hist_11_folded_hist
    , 1'h0}; // @[FrontendBundle.scala 290:21]
  wire [8:0] _updated_fh_res_hist_11_new_folded_hist_T_3 = _updated_fh_res_hist_11_new_folded_hist_T_2 | _GEN_11938; // @[FrontendBundle.scala 290:29]
  wire [7:0] updated_fh_res_hist_11_new_folded_hist_1 = _updated_fh_res_hist_11_new_folded_hist_T_3[7:0]; // @[FrontendBundle.scala 290:37]
  wire  updated_fh_res_hist_12_new_folded_hist_xored_res_1_5 =
    updated_fh_res_hist_0_new_folded_hist_newest_bits_masked_1[1] ^ updated_fh_ob_4_0 ^
    updated_fh_res_hist_12_new_folded_hist_original_bits_masked__5; // @[FrontendBundle.scala 256:48]
  wire  updated_fh_res_hist_12_new_folded_hist_xored_res_1_6 =
    updated_fh_res_hist_0_new_folded_hist_newest_bits_masked_1[0] ^
    updated_fh_res_hist_12_new_folded_hist_original_bits_masked__6; // @[FrontendBundle.scala 256:48]
  wire [6:0] updated_fh_res_hist_12_new_folded_hist_xored_1 = {updated_fh_res_hist_12_new_folded_hist_xored_res_1_6,
    updated_fh_res_hist_12_new_folded_hist_xored_res_1_5,updated_fh_res_hist_12_new_folded_hist_original_bits_masked__4,
    updated_fh_res_hist_12_new_folded_hist_original_bits_masked__3,
    updated_fh_res_hist_12_new_folded_hist_original_bits_masked__2,
    updated_fh_res_hist_12_new_folded_hist_original_bits_masked__1,
    updated_fh_res_hist_12_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [13:0] updated_fh_res_hist_12_new_folded_hist_src_doubled_1 = {
    updated_fh_res_hist_12_new_folded_hist_xored_res_1_6,updated_fh_res_hist_12_new_folded_hist_xored_res_1_5,
    updated_fh_res_hist_12_new_folded_hist_original_bits_masked__4,
    updated_fh_res_hist_12_new_folded_hist_original_bits_masked__3,
    updated_fh_res_hist_12_new_folded_hist_original_bits_masked__2,
    updated_fh_res_hist_12_new_folded_hist_original_bits_masked__1,
    updated_fh_res_hist_12_new_folded_hist_original_bits_masked__0,updated_fh_res_hist_12_new_folded_hist_xored_1}; // @[Cat.scala 31:58]
  wire [6:0] updated_fh_res_hist_12_new_folded_hist_1 = updated_fh_res_hist_12_new_folded_hist_src_doubled_1[12:6]; // @[FrontendBundle.scala 221:30]
  wire  updated_fh_res_hist_13_new_folded_hist_xored_res_1_0 = updated_fh_ob_10_0 ^
    updated_fh_res_hist_13_new_folded_hist_original_bits_masked__0; // @[FrontendBundle.scala 256:48]
  wire  updated_fh_res_hist_13_new_folded_hist_xored_res_1_5 =
    updated_fh_res_hist_0_new_folded_hist_newest_bits_masked_1[1] ^
    updated_fh_res_hist_13_new_folded_hist_original_bits_masked__5; // @[FrontendBundle.scala 256:48]
  wire  updated_fh_res_hist_13_new_folded_hist_xored_res_1_6 =
    updated_fh_res_hist_0_new_folded_hist_newest_bits_masked_1[0] ^
    updated_fh_res_hist_13_new_folded_hist_original_bits_masked__6; // @[FrontendBundle.scala 256:48]
  wire [6:0] updated_fh_res_hist_13_new_folded_hist_xored_1 = {updated_fh_res_hist_13_new_folded_hist_xored_res_1_6,
    updated_fh_res_hist_13_new_folded_hist_xored_res_1_5,updated_fh_res_hist_13_new_folded_hist_original_bits_masked__4,
    updated_fh_res_hist_13_new_folded_hist_original_bits_masked__3,
    updated_fh_res_hist_13_new_folded_hist_original_bits_masked__2,
    updated_fh_res_hist_13_new_folded_hist_original_bits_masked__1,updated_fh_res_hist_13_new_folded_hist_xored_res_1_0}
    ; // @[FrontendBundle.scala 258:11]
  wire [13:0] updated_fh_res_hist_13_new_folded_hist_src_doubled_1 = {
    updated_fh_res_hist_13_new_folded_hist_xored_res_1_6,updated_fh_res_hist_13_new_folded_hist_xored_res_1_5,
    updated_fh_res_hist_13_new_folded_hist_original_bits_masked__4,
    updated_fh_res_hist_13_new_folded_hist_original_bits_masked__3,
    updated_fh_res_hist_13_new_folded_hist_original_bits_masked__2,
    updated_fh_res_hist_13_new_folded_hist_original_bits_masked__1,updated_fh_res_hist_13_new_folded_hist_xored_res_1_0,
    updated_fh_res_hist_13_new_folded_hist_xored_1}; // @[Cat.scala 31:58]
  wire [6:0] updated_fh_res_hist_13_new_folded_hist_1 = updated_fh_res_hist_13_new_folded_hist_src_doubled_1[12:6]; // @[FrontendBundle.scala 221:30]
  wire  updated_fh_res_hist_14_new_folded_hist_xored_res_1_5 =
    updated_fh_res_hist_0_new_folded_hist_newest_bits_masked_1[1] ^
    updated_fh_res_hist_14_new_folded_hist_original_bits_masked__5; // @[FrontendBundle.scala 256:48]
  wire  updated_fh_res_hist_14_new_folded_hist_xored_res_1_6 =
    updated_fh_res_hist_0_new_folded_hist_newest_bits_masked_1[0] ^ updated_fh_ob_2_0 ^
    updated_fh_res_hist_14_new_folded_hist_original_bits_masked__6; // @[FrontendBundle.scala 256:48]
  wire [6:0] updated_fh_res_hist_14_new_folded_hist_xored_1 = {updated_fh_res_hist_14_new_folded_hist_xored_res_1_6,
    updated_fh_res_hist_14_new_folded_hist_xored_res_1_5,updated_fh_res_hist_14_new_folded_hist_original_bits_masked__4,
    updated_fh_res_hist_14_new_folded_hist_original_bits_masked__3,
    updated_fh_res_hist_14_new_folded_hist_original_bits_masked__2,
    updated_fh_res_hist_14_new_folded_hist_original_bits_masked__1,
    updated_fh_res_hist_14_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [13:0] updated_fh_res_hist_14_new_folded_hist_src_doubled_1 = {
    updated_fh_res_hist_14_new_folded_hist_xored_res_1_6,updated_fh_res_hist_14_new_folded_hist_xored_res_1_5,
    updated_fh_res_hist_14_new_folded_hist_original_bits_masked__4,
    updated_fh_res_hist_14_new_folded_hist_original_bits_masked__3,
    updated_fh_res_hist_14_new_folded_hist_original_bits_masked__2,
    updated_fh_res_hist_14_new_folded_hist_original_bits_masked__1,
    updated_fh_res_hist_14_new_folded_hist_original_bits_masked__0,updated_fh_res_hist_14_new_folded_hist_xored_1}; // @[Cat.scala 31:58]
  wire [6:0] updated_fh_res_hist_14_new_folded_hist_1 = updated_fh_res_hist_14_new_folded_hist_src_doubled_1[12:6]; // @[FrontendBundle.scala 221:30]
  wire  updated_fh_res_hist_15_new_folded_hist_xored_res_1_8 = updated_fh_ob_2_0 ^
    updated_fh_res_hist_15_new_folded_hist_original_bits_masked__8; // @[FrontendBundle.scala 256:48]
  wire  updated_fh_res_hist_15_new_folded_hist_xored_res_1_9 =
    updated_fh_res_hist_0_new_folded_hist_newest_bits_masked_1[1] ^
    updated_fh_res_hist_15_new_folded_hist_original_bits_masked__9; // @[FrontendBundle.scala 256:48]
  wire  updated_fh_res_hist_15_new_folded_hist_xored_res_1_10 =
    updated_fh_res_hist_0_new_folded_hist_newest_bits_masked_1[0] ^
    updated_fh_res_hist_15_new_folded_hist_original_bits_masked__10; // @[FrontendBundle.scala 256:48]
  wire [10:0] updated_fh_res_hist_15_new_folded_hist_xored_1 = {updated_fh_res_hist_15_new_folded_hist_xored_res_1_10,
    updated_fh_res_hist_15_new_folded_hist_xored_res_1_9,updated_fh_res_hist_15_new_folded_hist_xored_res_1_8,
    updated_fh_res_hist_15_new_folded_hist_original_bits_masked__7,
    updated_fh_res_hist_15_new_folded_hist_original_bits_masked__6,
    updated_fh_res_hist_15_new_folded_hist_original_bits_masked__5,updated_fh_res_hist_15_new_folded_hist_xored_lo}; // @[FrontendBundle.scala 258:11]
  wire [21:0] updated_fh_res_hist_15_new_folded_hist_src_doubled_1 = {
    updated_fh_res_hist_15_new_folded_hist_xored_res_1_10,updated_fh_res_hist_15_new_folded_hist_xored_res_1_9,
    updated_fh_res_hist_15_new_folded_hist_xored_res_1_8,updated_fh_res_hist_15_new_folded_hist_original_bits_masked__7,
    updated_fh_res_hist_15_new_folded_hist_original_bits_masked__6,
    updated_fh_res_hist_15_new_folded_hist_original_bits_masked__5,updated_fh_res_hist_15_new_folded_hist_xored_lo,
    updated_fh_res_hist_15_new_folded_hist_xored_1}; // @[Cat.scala 31:58]
  wire [10:0] updated_fh_res_hist_15_new_folded_hist_1 = updated_fh_res_hist_15_new_folded_hist_src_doubled_1[20:10]; // @[FrontendBundle.scala 221:30]
  wire  updated_fh_res_hist_16_new_folded_hist_xored_res_1_1 = updated_fh_ob_13_0 ^
    updated_fh_res_hist_16_new_folded_hist_original_bits_masked__1; // @[FrontendBundle.scala 256:48]
  wire  updated_fh_res_hist_16_new_folded_hist_xored_res_1_6 =
    updated_fh_res_hist_0_new_folded_hist_newest_bits_masked_1[1] ^
    updated_fh_res_hist_16_new_folded_hist_original_bits_masked__6; // @[FrontendBundle.scala 256:48]
  wire  updated_fh_res_hist_16_new_folded_hist_xored_res_1_7 =
    updated_fh_res_hist_0_new_folded_hist_newest_bits_masked_1[0] ^
    updated_fh_res_hist_16_new_folded_hist_original_bits_masked__7; // @[FrontendBundle.scala 256:48]
  wire [7:0] updated_fh_res_hist_16_new_folded_hist_xored_1 = {updated_fh_res_hist_16_new_folded_hist_xored_res_1_7,
    updated_fh_res_hist_16_new_folded_hist_xored_res_1_6,updated_fh_res_hist_16_new_folded_hist_original_bits_masked__5,
    updated_fh_res_hist_16_new_folded_hist_original_bits_masked__4,
    updated_fh_res_hist_16_new_folded_hist_original_bits_masked__3,
    updated_fh_res_hist_16_new_folded_hist_original_bits_masked__2,updated_fh_res_hist_16_new_folded_hist_xored_res_1_1,
    updated_fh_res_hist_16_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [15:0] updated_fh_res_hist_16_new_folded_hist_src_doubled_1 = {
    updated_fh_res_hist_16_new_folded_hist_xored_res_1_7,updated_fh_res_hist_16_new_folded_hist_xored_res_1_6,
    updated_fh_res_hist_16_new_folded_hist_original_bits_masked__5,
    updated_fh_res_hist_16_new_folded_hist_original_bits_masked__4,
    updated_fh_res_hist_16_new_folded_hist_original_bits_masked__3,
    updated_fh_res_hist_16_new_folded_hist_original_bits_masked__2,updated_fh_res_hist_16_new_folded_hist_xored_res_1_1,
    updated_fh_res_hist_16_new_folded_hist_original_bits_masked__0,updated_fh_res_hist_16_new_folded_hist_xored_1}; // @[Cat.scala 31:58]
  wire [7:0] updated_fh_res_hist_16_new_folded_hist_1 = updated_fh_res_hist_16_new_folded_hist_src_doubled_1[14:7]; // @[FrontendBundle.scala 221:30]
  wire  updated_fh_res_hist_17_new_folded_hist_xored_res_1_4 = updated_fh_ob_4_0 ^
    updated_fh_res_hist_17_new_folded_hist_original_bits_masked__4; // @[FrontendBundle.scala 256:48]
  wire  updated_fh_res_hist_17_new_folded_hist_xored_res_1_6 =
    updated_fh_res_hist_0_new_folded_hist_newest_bits_masked_1[1] ^
    updated_fh_res_hist_17_new_folded_hist_original_bits_masked__6; // @[FrontendBundle.scala 256:48]
  wire  updated_fh_res_hist_17_new_folded_hist_xored_res_1_7 =
    updated_fh_res_hist_0_new_folded_hist_newest_bits_masked_1[0] ^
    updated_fh_res_hist_17_new_folded_hist_original_bits_masked__7; // @[FrontendBundle.scala 256:48]
  wire [7:0] updated_fh_res_hist_17_new_folded_hist_xored_1 = {updated_fh_res_hist_17_new_folded_hist_xored_res_1_7,
    updated_fh_res_hist_17_new_folded_hist_xored_res_1_6,updated_fh_res_hist_17_new_folded_hist_original_bits_masked__5,
    updated_fh_res_hist_17_new_folded_hist_xored_res_1_4,updated_fh_res_hist_17_new_folded_hist_original_bits_masked__3,
    updated_fh_res_hist_17_new_folded_hist_original_bits_masked__2,
    updated_fh_res_hist_17_new_folded_hist_original_bits_masked__1,
    updated_fh_res_hist_17_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [15:0] updated_fh_res_hist_17_new_folded_hist_src_doubled_1 = {
    updated_fh_res_hist_17_new_folded_hist_xored_res_1_7,updated_fh_res_hist_17_new_folded_hist_xored_res_1_6,
    updated_fh_res_hist_17_new_folded_hist_original_bits_masked__5,updated_fh_res_hist_17_new_folded_hist_xored_res_1_4,
    updated_fh_res_hist_17_new_folded_hist_original_bits_masked__3,
    updated_fh_res_hist_17_new_folded_hist_original_bits_masked__2,
    updated_fh_res_hist_17_new_folded_hist_original_bits_masked__1,
    updated_fh_res_hist_17_new_folded_hist_original_bits_masked__0,updated_fh_res_hist_17_new_folded_hist_xored_1}; // @[Cat.scala 31:58]
  wire [7:0] updated_fh_res_hist_17_new_folded_hist_1 = updated_fh_res_hist_17_new_folded_hist_src_doubled_1[14:7]; // @[FrontendBundle.scala 221:30]
  wire [1:0] updated_fh_res_hist_0_new_folded_hist_newest_bits_masked_2 = {_updated_fh_T,1'h0}; // @[FrontendBundle.scala 274:102]
  wire  updated_fh_res_hist_0_new_folded_hist_xored_res_2_6 = updated_fh_res_hist_0_new_folded_hist_newest_bits_masked_2
    [1] ^ updated_fh_ob__1 ^ updated_fh_res_hist_0_new_folded_hist_original_bits_masked__6; // @[FrontendBundle.scala 256:48]
  wire  updated_fh_res_hist_0_new_folded_hist_xored_res_2_7 = updated_fh_res_hist_0_new_folded_hist_newest_bits_masked_2
    [0] ^ updated_fh_ob__0 ^ updated_fh_res_hist_0_new_folded_hist_original_bits_masked__7; // @[FrontendBundle.scala 256:48]
  wire [7:0] updated_fh_res_hist_0_new_folded_hist_xored_2 = {updated_fh_res_hist_0_new_folded_hist_xored_res_2_7,
    updated_fh_res_hist_0_new_folded_hist_xored_res_2_6,updated_fh_res_hist_0_new_folded_hist_original_bits_masked__5,
    updated_fh_res_hist_0_new_folded_hist_original_bits_masked__4,
    updated_fh_res_hist_0_new_folded_hist_original_bits_masked__3,
    updated_fh_res_hist_0_new_folded_hist_original_bits_masked__2,
    updated_fh_res_hist_0_new_folded_hist_original_bits_masked__1,
    updated_fh_res_hist_0_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [15:0] updated_fh_res_hist_0_new_folded_hist_src_doubled_2 = {updated_fh_res_hist_0_new_folded_hist_xored_res_2_7
    ,updated_fh_res_hist_0_new_folded_hist_xored_res_2_6,updated_fh_res_hist_0_new_folded_hist_original_bits_masked__5,
    updated_fh_res_hist_0_new_folded_hist_original_bits_masked__4,
    updated_fh_res_hist_0_new_folded_hist_original_bits_masked__3,
    updated_fh_res_hist_0_new_folded_hist_original_bits_masked__2,
    updated_fh_res_hist_0_new_folded_hist_original_bits_masked__1,
    updated_fh_res_hist_0_new_folded_hist_original_bits_masked__0,updated_fh_res_hist_0_new_folded_hist_xored_2}; // @[Cat.scala 31:58]
  wire [7:0] updated_fh_res_hist_0_new_folded_hist_2 = updated_fh_res_hist_0_new_folded_hist_src_doubled_2[13:6]; // @[FrontendBundle.scala 221:30]
  wire  updated_fh_res_hist_1_new_folded_hist_xored_res_2_6 = updated_fh_res_hist_0_new_folded_hist_newest_bits_masked_2
    [1] ^ updated_fh_ob_1_1 ^ updated_fh_res_hist_1_new_folded_hist_original_bits_masked__6; // @[FrontendBundle.scala 256:48]
  wire  updated_fh_res_hist_1_new_folded_hist_xored_res_2_7 = updated_fh_res_hist_0_new_folded_hist_newest_bits_masked_2
    [0] ^ updated_fh_ob_1_0 ^ updated_fh_res_hist_1_new_folded_hist_original_bits_masked__7; // @[FrontendBundle.scala 256:48]
  wire [7:0] updated_fh_res_hist_1_new_folded_hist_xored_2 = {updated_fh_res_hist_1_new_folded_hist_xored_res_2_7,
    updated_fh_res_hist_1_new_folded_hist_xored_res_2_6,updated_fh_res_hist_1_new_folded_hist_original_bits_masked__5,
    updated_fh_res_hist_1_new_folded_hist_original_bits_masked__4,
    updated_fh_res_hist_1_new_folded_hist_original_bits_masked__3,
    updated_fh_res_hist_1_new_folded_hist_original_bits_masked__2,
    updated_fh_res_hist_1_new_folded_hist_original_bits_masked__1,
    updated_fh_res_hist_1_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [15:0] updated_fh_res_hist_1_new_folded_hist_src_doubled_2 = {updated_fh_res_hist_1_new_folded_hist_xored_res_2_7
    ,updated_fh_res_hist_1_new_folded_hist_xored_res_2_6,updated_fh_res_hist_1_new_folded_hist_original_bits_masked__5,
    updated_fh_res_hist_1_new_folded_hist_original_bits_masked__4,
    updated_fh_res_hist_1_new_folded_hist_original_bits_masked__3,
    updated_fh_res_hist_1_new_folded_hist_original_bits_masked__2,
    updated_fh_res_hist_1_new_folded_hist_original_bits_masked__1,
    updated_fh_res_hist_1_new_folded_hist_original_bits_masked__0,updated_fh_res_hist_1_new_folded_hist_xored_2}; // @[Cat.scala 31:58]
  wire [7:0] updated_fh_res_hist_1_new_folded_hist_2 = updated_fh_res_hist_1_new_folded_hist_src_doubled_2[13:6]; // @[FrontendBundle.scala 221:30]
  wire  updated_fh_res_hist_2_new_folded_hist_xored_res_2_5 = updated_fh_ob_2_1 ^
    updated_fh_res_hist_2_new_folded_hist_original_bits_masked__5; // @[FrontendBundle.scala 256:48]
  wire  updated_fh_res_hist_2_new_folded_hist_xored_res_2_6 = updated_fh_res_hist_0_new_folded_hist_newest_bits_masked_2
    [1] ^ updated_fh_ob_2_0 ^ updated_fh_res_hist_2_new_folded_hist_original_bits_masked__6; // @[FrontendBundle.scala 256:48]
  wire  updated_fh_res_hist_2_new_folded_hist_xored_res_2_7 = updated_fh_res_hist_0_new_folded_hist_newest_bits_masked_2
    [0] ^ updated_fh_res_hist_2_new_folded_hist_original_bits_masked__7; // @[FrontendBundle.scala 256:48]
  wire [7:0] updated_fh_res_hist_2_new_folded_hist_xored_2 = {updated_fh_res_hist_2_new_folded_hist_xored_res_2_7,
    updated_fh_res_hist_2_new_folded_hist_xored_res_2_6,updated_fh_res_hist_2_new_folded_hist_xored_res_2_5,
    updated_fh_res_hist_2_new_folded_hist_original_bits_masked__4,
    updated_fh_res_hist_2_new_folded_hist_original_bits_masked__3,
    updated_fh_res_hist_2_new_folded_hist_original_bits_masked__2,
    updated_fh_res_hist_2_new_folded_hist_original_bits_masked__1,
    updated_fh_res_hist_2_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [15:0] updated_fh_res_hist_2_new_folded_hist_src_doubled_2 = {updated_fh_res_hist_2_new_folded_hist_xored_res_2_7
    ,updated_fh_res_hist_2_new_folded_hist_xored_res_2_6,updated_fh_res_hist_2_new_folded_hist_xored_res_2_5,
    updated_fh_res_hist_2_new_folded_hist_original_bits_masked__4,
    updated_fh_res_hist_2_new_folded_hist_original_bits_masked__3,
    updated_fh_res_hist_2_new_folded_hist_original_bits_masked__2,
    updated_fh_res_hist_2_new_folded_hist_original_bits_masked__1,
    updated_fh_res_hist_2_new_folded_hist_original_bits_masked__0,updated_fh_res_hist_2_new_folded_hist_xored_2}; // @[Cat.scala 31:58]
  wire [7:0] updated_fh_res_hist_2_new_folded_hist_2 = updated_fh_res_hist_2_new_folded_hist_src_doubled_2[13:6]; // @[FrontendBundle.scala 221:30]
  wire  updated_fh_res_hist_3_new_folded_hist_xored_res_2_8 = updated_fh_ob_1_1 ^
    updated_fh_res_hist_3_new_folded_hist_original_bits_masked__8; // @[FrontendBundle.scala 256:48]
  wire  updated_fh_res_hist_3_new_folded_hist_xored_res_2_9 = updated_fh_res_hist_0_new_folded_hist_newest_bits_masked_2
    [1] ^ updated_fh_ob_1_0 ^ updated_fh_res_hist_3_new_folded_hist_original_bits_masked__9; // @[FrontendBundle.scala 256:48]
  wire  updated_fh_res_hist_3_new_folded_hist_xored_res_2_10 =
    updated_fh_res_hist_0_new_folded_hist_newest_bits_masked_2[0] ^
    updated_fh_res_hist_3_new_folded_hist_original_bits_masked__10; // @[FrontendBundle.scala 256:48]
  wire [10:0] updated_fh_res_hist_3_new_folded_hist_xored_2 = {updated_fh_res_hist_3_new_folded_hist_xored_res_2_10,
    updated_fh_res_hist_3_new_folded_hist_xored_res_2_9,updated_fh_res_hist_3_new_folded_hist_xored_res_2_8,
    updated_fh_res_hist_3_new_folded_hist_original_bits_masked__7,
    updated_fh_res_hist_3_new_folded_hist_original_bits_masked__6,
    updated_fh_res_hist_3_new_folded_hist_original_bits_masked__5,updated_fh_res_hist_3_new_folded_hist_xored_lo}; // @[FrontendBundle.scala 258:11]
  wire [21:0] updated_fh_res_hist_3_new_folded_hist_src_doubled_2 = {
    updated_fh_res_hist_3_new_folded_hist_xored_res_2_10,updated_fh_res_hist_3_new_folded_hist_xored_res_2_9,
    updated_fh_res_hist_3_new_folded_hist_xored_res_2_8,updated_fh_res_hist_3_new_folded_hist_original_bits_masked__7,
    updated_fh_res_hist_3_new_folded_hist_original_bits_masked__6,
    updated_fh_res_hist_3_new_folded_hist_original_bits_masked__5,updated_fh_res_hist_3_new_folded_hist_xored_lo,
    updated_fh_res_hist_3_new_folded_hist_xored_2}; // @[Cat.scala 31:58]
  wire [10:0] updated_fh_res_hist_3_new_folded_hist_2 = updated_fh_res_hist_3_new_folded_hist_src_doubled_2[19:9]; // @[FrontendBundle.scala 221:30]
  wire [5:0] _updated_fh_res_hist_4_new_folded_hist_T_4 = {do_redirect_bits_cfiUpdate_folded_hist_hist_4_folded_hist
    , 2'h0}; // @[FrontendBundle.scala 290:21]
  wire [5:0] _GEN_11940 = {{5'd0}, _updated_fh_T}; // @[FrontendBundle.scala 290:29]
  wire [5:0] _updated_fh_res_hist_4_new_folded_hist_T_5 = _updated_fh_res_hist_4_new_folded_hist_T_4 | _GEN_11940; // @[FrontendBundle.scala 290:29]
  wire [3:0] updated_fh_res_hist_4_new_folded_hist_2 = _updated_fh_res_hist_4_new_folded_hist_T_5[3:0]; // @[FrontendBundle.scala 290:37]
  wire  updated_fh_res_hist_5_new_folded_hist_xored_res_2_0 = updated_fh_ob_4_1 ^
    updated_fh_res_hist_5_new_folded_hist_original_bits_masked__0; // @[FrontendBundle.scala 256:48]
  wire  updated_fh_res_hist_5_new_folded_hist_xored_res_2_9 = updated_fh_res_hist_0_new_folded_hist_newest_bits_masked_2
    [1] ^ updated_fh_res_hist_5_new_folded_hist_original_bits_masked__9; // @[FrontendBundle.scala 256:48]
  wire  updated_fh_res_hist_5_new_folded_hist_xored_res_2_10 =
    updated_fh_res_hist_0_new_folded_hist_newest_bits_masked_2[0] ^
    updated_fh_res_hist_5_new_folded_hist_original_bits_masked__10; // @[FrontendBundle.scala 256:48]
  wire [4:0] updated_fh_res_hist_5_new_folded_hist_xored_lo_2 = {
    updated_fh_res_hist_5_new_folded_hist_original_bits_masked__4,
    updated_fh_res_hist_5_new_folded_hist_original_bits_masked__3,
    updated_fh_res_hist_5_new_folded_hist_original_bits_masked__2,updated_fh_res_hist_5_new_folded_hist_xored_res_1_1,
    updated_fh_res_hist_5_new_folded_hist_xored_res_2_0}; // @[FrontendBundle.scala 258:11]
  wire [10:0] updated_fh_res_hist_5_new_folded_hist_xored_2 = {updated_fh_res_hist_5_new_folded_hist_xored_res_2_10,
    updated_fh_res_hist_5_new_folded_hist_xored_res_2_9,updated_fh_res_hist_5_new_folded_hist_original_bits_masked__8,
    updated_fh_res_hist_5_new_folded_hist_original_bits_masked__7,
    updated_fh_res_hist_5_new_folded_hist_original_bits_masked__6,
    updated_fh_res_hist_5_new_folded_hist_original_bits_masked__5,updated_fh_res_hist_5_new_folded_hist_xored_lo_2}; // @[FrontendBundle.scala 258:11]
  wire [21:0] updated_fh_res_hist_5_new_folded_hist_src_doubled_2 = {
    updated_fh_res_hist_5_new_folded_hist_xored_res_2_10,updated_fh_res_hist_5_new_folded_hist_xored_res_2_9,
    updated_fh_res_hist_5_new_folded_hist_original_bits_masked__8,
    updated_fh_res_hist_5_new_folded_hist_original_bits_masked__7,
    updated_fh_res_hist_5_new_folded_hist_original_bits_masked__6,
    updated_fh_res_hist_5_new_folded_hist_original_bits_masked__5,updated_fh_res_hist_5_new_folded_hist_xored_lo_2,
    updated_fh_res_hist_5_new_folded_hist_xored_2}; // @[Cat.scala 31:58]
  wire [10:0] updated_fh_res_hist_5_new_folded_hist_2 = updated_fh_res_hist_5_new_folded_hist_src_doubled_2[19:9]; // @[FrontendBundle.scala 221:30]
  wire  updated_fh_res_hist_6_new_folded_hist_xored_res_2_2 = updated_fh_ob_4_1 ^
    updated_fh_res_hist_6_new_folded_hist_original_bits_masked__2; // @[FrontendBundle.scala 256:48]
  wire  updated_fh_res_hist_6_new_folded_hist_xored_res_2_7 = updated_fh_res_hist_0_new_folded_hist_newest_bits_masked_2
    [1] ^ updated_fh_res_hist_6_new_folded_hist_original_bits_masked__7; // @[FrontendBundle.scala 256:48]
  wire  updated_fh_res_hist_6_new_folded_hist_xored_res_2_8 = updated_fh_res_hist_0_new_folded_hist_newest_bits_masked_2
    [0] ^ updated_fh_res_hist_6_new_folded_hist_original_bits_masked__8; // @[FrontendBundle.scala 256:48]
  wire [8:0] updated_fh_res_hist_6_new_folded_hist_xored_2 = {updated_fh_res_hist_6_new_folded_hist_xored_res_2_8,
    updated_fh_res_hist_6_new_folded_hist_xored_res_2_7,updated_fh_res_hist_6_new_folded_hist_original_bits_masked__6,
    updated_fh_res_hist_6_new_folded_hist_original_bits_masked__5,
    updated_fh_res_hist_6_new_folded_hist_original_bits_masked__4,updated_fh_res_hist_6_new_folded_hist_xored_res_1_3,
    updated_fh_res_hist_6_new_folded_hist_xored_res_2_2,updated_fh_res_hist_6_new_folded_hist_original_bits_masked__1,
    updated_fh_res_hist_6_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [17:0] updated_fh_res_hist_6_new_folded_hist_src_doubled_2 = {updated_fh_res_hist_6_new_folded_hist_xored_res_2_8
    ,updated_fh_res_hist_6_new_folded_hist_xored_res_2_7,updated_fh_res_hist_6_new_folded_hist_original_bits_masked__6,
    updated_fh_res_hist_6_new_folded_hist_original_bits_masked__5,
    updated_fh_res_hist_6_new_folded_hist_original_bits_masked__4,updated_fh_res_hist_6_new_folded_hist_xored_res_1_3,
    updated_fh_res_hist_6_new_folded_hist_xored_res_2_2,updated_fh_res_hist_6_new_folded_hist_original_bits_masked__1,
    updated_fh_res_hist_6_new_folded_hist_original_bits_masked__0,updated_fh_res_hist_6_new_folded_hist_xored_2}; // @[Cat.scala 31:58]
  wire [8:0] updated_fh_res_hist_6_new_folded_hist_2 = updated_fh_res_hist_6_new_folded_hist_src_doubled_2[15:7]; // @[FrontendBundle.scala 221:30]
  wire  updated_fh_res_hist_7_new_folded_hist_xored_res_2_5 = updated_fh_ob__1 ^
    updated_fh_res_hist_7_new_folded_hist_original_bits_masked__5; // @[FrontendBundle.scala 256:48]
  wire  updated_fh_res_hist_7_new_folded_hist_xored_res_2_7 = updated_fh_res_hist_0_new_folded_hist_newest_bits_masked_2
    [1] ^ updated_fh_res_hist_7_new_folded_hist_original_bits_masked__7; // @[FrontendBundle.scala 256:48]
  wire  updated_fh_res_hist_7_new_folded_hist_xored_res_2_8 = updated_fh_res_hist_0_new_folded_hist_newest_bits_masked_2
    [0] ^ updated_fh_res_hist_7_new_folded_hist_original_bits_masked__8; // @[FrontendBundle.scala 256:48]
  wire [8:0] updated_fh_res_hist_7_new_folded_hist_xored_2 = {updated_fh_res_hist_7_new_folded_hist_xored_res_2_8,
    updated_fh_res_hist_7_new_folded_hist_xored_res_2_7,updated_fh_res_hist_7_new_folded_hist_xored_res_1_6,
    updated_fh_res_hist_7_new_folded_hist_xored_res_2_5,updated_fh_res_hist_7_new_folded_hist_original_bits_masked__4,
    updated_fh_res_hist_7_new_folded_hist_original_bits_masked__3,
    updated_fh_res_hist_7_new_folded_hist_original_bits_masked__2,
    updated_fh_res_hist_7_new_folded_hist_original_bits_masked__1,
    updated_fh_res_hist_7_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [17:0] updated_fh_res_hist_7_new_folded_hist_src_doubled_2 = {updated_fh_res_hist_7_new_folded_hist_xored_res_2_8
    ,updated_fh_res_hist_7_new_folded_hist_xored_res_2_7,updated_fh_res_hist_7_new_folded_hist_xored_res_1_6,
    updated_fh_res_hist_7_new_folded_hist_xored_res_2_5,updated_fh_res_hist_7_new_folded_hist_original_bits_masked__4,
    updated_fh_res_hist_7_new_folded_hist_original_bits_masked__3,
    updated_fh_res_hist_7_new_folded_hist_original_bits_masked__2,
    updated_fh_res_hist_7_new_folded_hist_original_bits_masked__1,
    updated_fh_res_hist_7_new_folded_hist_original_bits_masked__0,updated_fh_res_hist_7_new_folded_hist_xored_2}; // @[Cat.scala 31:58]
  wire [8:0] updated_fh_res_hist_7_new_folded_hist_2 = updated_fh_res_hist_7_new_folded_hist_src_doubled_2[15:7]; // @[FrontendBundle.scala 221:30]
  wire [9:0] _updated_fh_res_hist_8_new_folded_hist_T_4 = {do_redirect_bits_cfiUpdate_folded_hist_hist_8_folded_hist
    , 2'h0}; // @[FrontendBundle.scala 290:21]
  wire [9:0] _GEN_11941 = {{9'd0}, _updated_fh_T}; // @[FrontendBundle.scala 290:29]
  wire [9:0] _updated_fh_res_hist_8_new_folded_hist_T_5 = _updated_fh_res_hist_8_new_folded_hist_T_4 | _GEN_11941; // @[FrontendBundle.scala 290:29]
  wire [7:0] updated_fh_res_hist_8_new_folded_hist_2 = _updated_fh_res_hist_8_new_folded_hist_T_5[7:0]; // @[FrontendBundle.scala 290:37]
  wire  updated_fh_res_hist_9_new_folded_hist_xored_res_2_2 = updated_fh_ob_1_1 ^
    updated_fh_res_hist_9_new_folded_hist_original_bits_masked__2; // @[FrontendBundle.scala 256:48]
  wire  updated_fh_res_hist_9_new_folded_hist_xored_res_2_5 = updated_fh_res_hist_0_new_folded_hist_newest_bits_masked_2
    [1] ^ updated_fh_res_hist_9_new_folded_hist_original_bits_masked__5; // @[FrontendBundle.scala 256:48]
  wire  updated_fh_res_hist_9_new_folded_hist_xored_res_2_6 = updated_fh_res_hist_0_new_folded_hist_newest_bits_masked_2
    [0] ^ updated_fh_res_hist_9_new_folded_hist_original_bits_masked__6; // @[FrontendBundle.scala 256:48]
  wire [6:0] updated_fh_res_hist_9_new_folded_hist_xored_2 = {updated_fh_res_hist_9_new_folded_hist_xored_res_2_6,
    updated_fh_res_hist_9_new_folded_hist_xored_res_2_5,updated_fh_res_hist_9_new_folded_hist_original_bits_masked__4,
    updated_fh_res_hist_9_new_folded_hist_xored_res_1_3,updated_fh_res_hist_9_new_folded_hist_xored_res_2_2,
    updated_fh_res_hist_9_new_folded_hist_original_bits_masked__1,
    updated_fh_res_hist_9_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [13:0] updated_fh_res_hist_9_new_folded_hist_src_doubled_2 = {updated_fh_res_hist_9_new_folded_hist_xored_res_2_6
    ,updated_fh_res_hist_9_new_folded_hist_xored_res_2_5,updated_fh_res_hist_9_new_folded_hist_original_bits_masked__4,
    updated_fh_res_hist_9_new_folded_hist_xored_res_1_3,updated_fh_res_hist_9_new_folded_hist_xored_res_2_2,
    updated_fh_res_hist_9_new_folded_hist_original_bits_masked__1,
    updated_fh_res_hist_9_new_folded_hist_original_bits_masked__0,updated_fh_res_hist_9_new_folded_hist_xored_2}; // @[Cat.scala 31:58]
  wire [6:0] updated_fh_res_hist_9_new_folded_hist_2 = updated_fh_res_hist_9_new_folded_hist_src_doubled_2[11:5]; // @[FrontendBundle.scala 221:30]
  wire  updated_fh_res_hist_10_new_folded_hist_xored_res_2_3 = updated_fh_ob_1_1 ^
    updated_fh_res_hist_10_new_folded_hist_original_bits_masked__3; // @[FrontendBundle.scala 256:48]
  wire  updated_fh_res_hist_10_new_folded_hist_xored_res_2_7 =
    updated_fh_res_hist_0_new_folded_hist_newest_bits_masked_2[1] ^
    updated_fh_res_hist_10_new_folded_hist_original_bits_masked__7; // @[FrontendBundle.scala 256:48]
  wire  updated_fh_res_hist_10_new_folded_hist_xored_res_2_8 =
    updated_fh_res_hist_0_new_folded_hist_newest_bits_masked_2[0] ^
    updated_fh_res_hist_10_new_folded_hist_original_bits_masked__8; // @[FrontendBundle.scala 256:48]
  wire [8:0] updated_fh_res_hist_10_new_folded_hist_xored_2 = {updated_fh_res_hist_10_new_folded_hist_xored_res_2_8,
    updated_fh_res_hist_10_new_folded_hist_xored_res_2_7,updated_fh_res_hist_10_new_folded_hist_original_bits_masked__6,
    updated_fh_res_hist_10_new_folded_hist_original_bits_masked__5,updated_fh_res_hist_10_new_folded_hist_xored_res_1_4,
    updated_fh_res_hist_10_new_folded_hist_xored_res_2_3,updated_fh_res_hist_10_new_folded_hist_original_bits_masked__2,
    updated_fh_res_hist_10_new_folded_hist_original_bits_masked__1,
    updated_fh_res_hist_10_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [17:0] updated_fh_res_hist_10_new_folded_hist_src_doubled_2 = {
    updated_fh_res_hist_10_new_folded_hist_xored_res_2_8,updated_fh_res_hist_10_new_folded_hist_xored_res_2_7,
    updated_fh_res_hist_10_new_folded_hist_original_bits_masked__6,
    updated_fh_res_hist_10_new_folded_hist_original_bits_masked__5,updated_fh_res_hist_10_new_folded_hist_xored_res_1_4,
    updated_fh_res_hist_10_new_folded_hist_xored_res_2_3,updated_fh_res_hist_10_new_folded_hist_original_bits_masked__2,
    updated_fh_res_hist_10_new_folded_hist_original_bits_masked__1,
    updated_fh_res_hist_10_new_folded_hist_original_bits_masked__0,updated_fh_res_hist_10_new_folded_hist_xored_2}; // @[Cat.scala 31:58]
  wire [8:0] updated_fh_res_hist_10_new_folded_hist_2 = updated_fh_res_hist_10_new_folded_hist_src_doubled_2[15:7]; // @[FrontendBundle.scala 221:30]
  wire [9:0] _updated_fh_res_hist_11_new_folded_hist_T_4 = {do_redirect_bits_cfiUpdate_folded_hist_hist_11_folded_hist
    , 2'h0}; // @[FrontendBundle.scala 290:21]
  wire [9:0] _updated_fh_res_hist_11_new_folded_hist_T_5 = _updated_fh_res_hist_11_new_folded_hist_T_4 | _GEN_11941; // @[FrontendBundle.scala 290:29]
  wire [7:0] updated_fh_res_hist_11_new_folded_hist_2 = _updated_fh_res_hist_11_new_folded_hist_T_5[7:0]; // @[FrontendBundle.scala 290:37]
  wire  updated_fh_res_hist_12_new_folded_hist_xored_res_2_4 = updated_fh_ob_4_1 ^
    updated_fh_res_hist_12_new_folded_hist_original_bits_masked__4; // @[FrontendBundle.scala 256:48]
  wire  updated_fh_res_hist_12_new_folded_hist_xored_res_2_5 =
    updated_fh_res_hist_0_new_folded_hist_newest_bits_masked_2[1] ^ updated_fh_ob_4_0 ^
    updated_fh_res_hist_12_new_folded_hist_original_bits_masked__5; // @[FrontendBundle.scala 256:48]
  wire  updated_fh_res_hist_12_new_folded_hist_xored_res_2_6 =
    updated_fh_res_hist_0_new_folded_hist_newest_bits_masked_2[0] ^
    updated_fh_res_hist_12_new_folded_hist_original_bits_masked__6; // @[FrontendBundle.scala 256:48]
  wire [6:0] updated_fh_res_hist_12_new_folded_hist_xored_2 = {updated_fh_res_hist_12_new_folded_hist_xored_res_2_6,
    updated_fh_res_hist_12_new_folded_hist_xored_res_2_5,updated_fh_res_hist_12_new_folded_hist_xored_res_2_4,
    updated_fh_res_hist_12_new_folded_hist_original_bits_masked__3,
    updated_fh_res_hist_12_new_folded_hist_original_bits_masked__2,
    updated_fh_res_hist_12_new_folded_hist_original_bits_masked__1,
    updated_fh_res_hist_12_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [13:0] updated_fh_res_hist_12_new_folded_hist_src_doubled_2 = {
    updated_fh_res_hist_12_new_folded_hist_xored_res_2_6,updated_fh_res_hist_12_new_folded_hist_xored_res_2_5,
    updated_fh_res_hist_12_new_folded_hist_xored_res_2_4,updated_fh_res_hist_12_new_folded_hist_original_bits_masked__3,
    updated_fh_res_hist_12_new_folded_hist_original_bits_masked__2,
    updated_fh_res_hist_12_new_folded_hist_original_bits_masked__1,
    updated_fh_res_hist_12_new_folded_hist_original_bits_masked__0,updated_fh_res_hist_12_new_folded_hist_xored_2}; // @[Cat.scala 31:58]
  wire [6:0] updated_fh_res_hist_12_new_folded_hist_2 = updated_fh_res_hist_12_new_folded_hist_src_doubled_2[11:5]; // @[FrontendBundle.scala 221:30]
  wire  updated_fh_res_hist_13_new_folded_hist_xored_res_2_5 =
    updated_fh_res_hist_0_new_folded_hist_newest_bits_masked_2[1] ^
    updated_fh_res_hist_13_new_folded_hist_original_bits_masked__5; // @[FrontendBundle.scala 256:48]
  wire [6:0] updated_fh_res_hist_13_new_folded_hist_xored_2 = {
    updated_fh_res_hist_0_new_folded_hist_newest_bits_masked_2[0],updated_fh_res_hist_13_new_folded_hist_xored_res_2_5,
    updated_fh_res_hist_13_new_folded_hist_original_bits_masked__4,
    updated_fh_res_hist_13_new_folded_hist_original_bits_masked__3,
    updated_fh_res_hist_13_new_folded_hist_original_bits_masked__2,
    updated_fh_res_hist_13_new_folded_hist_original_bits_masked__1,updated_fh_res_hist_13_new_folded_hist_xored_res_1_0}
    ; // @[FrontendBundle.scala 258:11]
  wire [13:0] updated_fh_res_hist_13_new_folded_hist_src_doubled_2 = {
    updated_fh_res_hist_0_new_folded_hist_newest_bits_masked_2[0],updated_fh_res_hist_13_new_folded_hist_xored_res_2_5,
    updated_fh_res_hist_13_new_folded_hist_original_bits_masked__4,
    updated_fh_res_hist_13_new_folded_hist_original_bits_masked__3,
    updated_fh_res_hist_13_new_folded_hist_original_bits_masked__2,
    updated_fh_res_hist_13_new_folded_hist_original_bits_masked__1,updated_fh_res_hist_13_new_folded_hist_xored_res_1_0,
    updated_fh_res_hist_13_new_folded_hist_xored_2}; // @[Cat.scala 31:58]
  wire [6:0] updated_fh_res_hist_13_new_folded_hist_2 = updated_fh_res_hist_13_new_folded_hist_src_doubled_2[11:5]; // @[FrontendBundle.scala 221:30]
  wire  updated_fh_res_hist_14_new_folded_hist_xored_res_2_5 =
    updated_fh_res_hist_0_new_folded_hist_newest_bits_masked_2[1] ^ updated_fh_ob_2_1 ^
    updated_fh_res_hist_14_new_folded_hist_original_bits_masked__5; // @[FrontendBundle.scala 256:48]
  wire  updated_fh_res_hist_14_new_folded_hist_xored_res_2_6 =
    updated_fh_res_hist_0_new_folded_hist_newest_bits_masked_2[0] ^ updated_fh_ob_2_0 ^
    updated_fh_res_hist_14_new_folded_hist_original_bits_masked__6; // @[FrontendBundle.scala 256:48]
  wire [6:0] updated_fh_res_hist_14_new_folded_hist_xored_2 = {updated_fh_res_hist_14_new_folded_hist_xored_res_2_6,
    updated_fh_res_hist_14_new_folded_hist_xored_res_2_5,updated_fh_res_hist_14_new_folded_hist_original_bits_masked__4,
    updated_fh_res_hist_14_new_folded_hist_original_bits_masked__3,
    updated_fh_res_hist_14_new_folded_hist_original_bits_masked__2,
    updated_fh_res_hist_14_new_folded_hist_original_bits_masked__1,
    updated_fh_res_hist_14_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [13:0] updated_fh_res_hist_14_new_folded_hist_src_doubled_2 = {
    updated_fh_res_hist_14_new_folded_hist_xored_res_2_6,updated_fh_res_hist_14_new_folded_hist_xored_res_2_5,
    updated_fh_res_hist_14_new_folded_hist_original_bits_masked__4,
    updated_fh_res_hist_14_new_folded_hist_original_bits_masked__3,
    updated_fh_res_hist_14_new_folded_hist_original_bits_masked__2,
    updated_fh_res_hist_14_new_folded_hist_original_bits_masked__1,
    updated_fh_res_hist_14_new_folded_hist_original_bits_masked__0,updated_fh_res_hist_14_new_folded_hist_xored_2}; // @[Cat.scala 31:58]
  wire [6:0] updated_fh_res_hist_14_new_folded_hist_2 = updated_fh_res_hist_14_new_folded_hist_src_doubled_2[11:5]; // @[FrontendBundle.scala 221:30]
  wire  updated_fh_res_hist_15_new_folded_hist_xored_res_2_7 = updated_fh_ob_2_1 ^
    updated_fh_res_hist_15_new_folded_hist_original_bits_masked__7; // @[FrontendBundle.scala 256:48]
  wire  updated_fh_res_hist_15_new_folded_hist_xored_res_2_9 =
    updated_fh_res_hist_0_new_folded_hist_newest_bits_masked_2[1] ^
    updated_fh_res_hist_15_new_folded_hist_original_bits_masked__9; // @[FrontendBundle.scala 256:48]
  wire  updated_fh_res_hist_15_new_folded_hist_xored_res_2_10 =
    updated_fh_res_hist_0_new_folded_hist_newest_bits_masked_2[0] ^
    updated_fh_res_hist_15_new_folded_hist_original_bits_masked__10; // @[FrontendBundle.scala 256:48]
  wire [10:0] updated_fh_res_hist_15_new_folded_hist_xored_2 = {updated_fh_res_hist_15_new_folded_hist_xored_res_2_10,
    updated_fh_res_hist_15_new_folded_hist_xored_res_2_9,updated_fh_res_hist_15_new_folded_hist_xored_res_1_8,
    updated_fh_res_hist_15_new_folded_hist_xored_res_2_7,updated_fh_res_hist_15_new_folded_hist_original_bits_masked__6,
    updated_fh_res_hist_15_new_folded_hist_original_bits_masked__5,updated_fh_res_hist_15_new_folded_hist_xored_lo}; // @[FrontendBundle.scala 258:11]
  wire [21:0] updated_fh_res_hist_15_new_folded_hist_src_doubled_2 = {
    updated_fh_res_hist_15_new_folded_hist_xored_res_2_10,updated_fh_res_hist_15_new_folded_hist_xored_res_2_9,
    updated_fh_res_hist_15_new_folded_hist_xored_res_1_8,updated_fh_res_hist_15_new_folded_hist_xored_res_2_7,
    updated_fh_res_hist_15_new_folded_hist_original_bits_masked__6,
    updated_fh_res_hist_15_new_folded_hist_original_bits_masked__5,updated_fh_res_hist_15_new_folded_hist_xored_lo,
    updated_fh_res_hist_15_new_folded_hist_xored_2}; // @[Cat.scala 31:58]
  wire [10:0] updated_fh_res_hist_15_new_folded_hist_2 = updated_fh_res_hist_15_new_folded_hist_src_doubled_2[19:9]; // @[FrontendBundle.scala 221:30]
  wire  updated_fh_res_hist_16_new_folded_hist_xored_res_2_0 = updated_fh_ob_13_1 ^
    updated_fh_res_hist_16_new_folded_hist_original_bits_masked__0; // @[FrontendBundle.scala 256:48]
  wire  updated_fh_res_hist_16_new_folded_hist_xored_res_2_6 =
    updated_fh_res_hist_0_new_folded_hist_newest_bits_masked_2[1] ^
    updated_fh_res_hist_16_new_folded_hist_original_bits_masked__6; // @[FrontendBundle.scala 256:48]
  wire  updated_fh_res_hist_16_new_folded_hist_xored_res_2_7 =
    updated_fh_res_hist_0_new_folded_hist_newest_bits_masked_2[0] ^
    updated_fh_res_hist_16_new_folded_hist_original_bits_masked__7; // @[FrontendBundle.scala 256:48]
  wire [7:0] updated_fh_res_hist_16_new_folded_hist_xored_2 = {updated_fh_res_hist_16_new_folded_hist_xored_res_2_7,
    updated_fh_res_hist_16_new_folded_hist_xored_res_2_6,updated_fh_res_hist_16_new_folded_hist_original_bits_masked__5,
    updated_fh_res_hist_16_new_folded_hist_original_bits_masked__4,
    updated_fh_res_hist_16_new_folded_hist_original_bits_masked__3,
    updated_fh_res_hist_16_new_folded_hist_original_bits_masked__2,updated_fh_res_hist_16_new_folded_hist_xored_res_1_1,
    updated_fh_res_hist_16_new_folded_hist_xored_res_2_0}; // @[FrontendBundle.scala 258:11]
  wire [15:0] updated_fh_res_hist_16_new_folded_hist_src_doubled_2 = {
    updated_fh_res_hist_16_new_folded_hist_xored_res_2_7,updated_fh_res_hist_16_new_folded_hist_xored_res_2_6,
    updated_fh_res_hist_16_new_folded_hist_original_bits_masked__5,
    updated_fh_res_hist_16_new_folded_hist_original_bits_masked__4,
    updated_fh_res_hist_16_new_folded_hist_original_bits_masked__3,
    updated_fh_res_hist_16_new_folded_hist_original_bits_masked__2,updated_fh_res_hist_16_new_folded_hist_xored_res_1_1,
    updated_fh_res_hist_16_new_folded_hist_xored_res_2_0,updated_fh_res_hist_16_new_folded_hist_xored_2}; // @[Cat.scala 31:58]
  wire [7:0] updated_fh_res_hist_16_new_folded_hist_2 = updated_fh_res_hist_16_new_folded_hist_src_doubled_2[13:6]; // @[FrontendBundle.scala 221:30]
  wire  updated_fh_res_hist_17_new_folded_hist_xored_res_2_3 = updated_fh_ob_4_1 ^
    updated_fh_res_hist_17_new_folded_hist_original_bits_masked__3; // @[FrontendBundle.scala 256:48]
  wire  updated_fh_res_hist_17_new_folded_hist_xored_res_2_6 =
    updated_fh_res_hist_0_new_folded_hist_newest_bits_masked_2[1] ^
    updated_fh_res_hist_17_new_folded_hist_original_bits_masked__6; // @[FrontendBundle.scala 256:48]
  wire  updated_fh_res_hist_17_new_folded_hist_xored_res_2_7 =
    updated_fh_res_hist_0_new_folded_hist_newest_bits_masked_2[0] ^
    updated_fh_res_hist_17_new_folded_hist_original_bits_masked__7; // @[FrontendBundle.scala 256:48]
  wire [7:0] updated_fh_res_hist_17_new_folded_hist_xored_2 = {updated_fh_res_hist_17_new_folded_hist_xored_res_2_7,
    updated_fh_res_hist_17_new_folded_hist_xored_res_2_6,updated_fh_res_hist_17_new_folded_hist_original_bits_masked__5,
    updated_fh_res_hist_17_new_folded_hist_xored_res_1_4,updated_fh_res_hist_17_new_folded_hist_xored_res_2_3,
    updated_fh_res_hist_17_new_folded_hist_original_bits_masked__2,
    updated_fh_res_hist_17_new_folded_hist_original_bits_masked__1,
    updated_fh_res_hist_17_new_folded_hist_original_bits_masked__0}; // @[FrontendBundle.scala 258:11]
  wire [15:0] updated_fh_res_hist_17_new_folded_hist_src_doubled_2 = {
    updated_fh_res_hist_17_new_folded_hist_xored_res_2_7,updated_fh_res_hist_17_new_folded_hist_xored_res_2_6,
    updated_fh_res_hist_17_new_folded_hist_original_bits_masked__5,updated_fh_res_hist_17_new_folded_hist_xored_res_1_4,
    updated_fh_res_hist_17_new_folded_hist_xored_res_2_3,updated_fh_res_hist_17_new_folded_hist_original_bits_masked__2,
    updated_fh_res_hist_17_new_folded_hist_original_bits_masked__1,
    updated_fh_res_hist_17_new_folded_hist_original_bits_masked__0,updated_fh_res_hist_17_new_folded_hist_xored_2}; // @[Cat.scala 31:58]
  wire [7:0] updated_fh_res_hist_17_new_folded_hist_2 = updated_fh_res_hist_17_new_folded_hist_src_doubled_2[13:6]; // @[FrontendBundle.scala 221:30]
  wire [3:0] _thisBrNumOH_T = 4'h1 << do_redirect_bits_cfiUpdate_shift; // @[OneHot.scala 64:12]
  wire [8:0] new_value_60 = do_redirect_bits_cfiUpdate_histPtr_value + 8'h74; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_361 = {1'h0,new_value_60}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_60 = $signed(_diff_T_361) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_60 = $signed(diff_60) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_120 = $signed(_diff_T_361) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_121 = reverse_flag_60 ? _new_ptr_value_T_120 : {{1'd0}, new_value_60}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_61 = do_redirect_bits_cfiUpdate_histPtr_value + 8'h6; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_367 = {1'h0,new_value_61}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_61 = $signed(_diff_T_367) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_61 = $signed(diff_61) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_122 = $signed(_diff_T_367) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_123 = reverse_flag_61 ? _new_ptr_value_T_122 : {{1'd0}, new_value_61}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_62 = do_redirect_bits_cfiUpdate_histPtr_value + 8'hb; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_373 = {1'h0,new_value_62}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_62 = $signed(_diff_T_373) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_62 = $signed(diff_62) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_124 = $signed(_diff_T_373) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_125 = reverse_flag_62 ? _new_ptr_value_T_124 : {{1'd0}, new_value_62}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_63 = do_redirect_bits_cfiUpdate_histPtr_value + 8'hf; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_379 = {1'h0,new_value_63}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_63 = $signed(_diff_T_379) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_63 = $signed(diff_63) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_126 = $signed(_diff_T_379) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_127 = reverse_flag_63 ? _new_ptr_value_T_126 : {{1'd0}, new_value_63}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_64 = do_redirect_bits_cfiUpdate_histPtr_value + 8'h1e; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_385 = {1'h0,new_value_64}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_64 = $signed(_diff_T_385) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_64 = $signed(diff_64) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_128 = $signed(_diff_T_385) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_129 = reverse_flag_64 ? _new_ptr_value_T_128 : {{1'd0}, new_value_64}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_65 = do_redirect_bits_cfiUpdate_histPtr_value + 8'h75; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_391 = {1'h0,new_value_65}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_65 = $signed(_diff_T_391) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_65 = $signed(diff_65) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_130 = $signed(_diff_T_391) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_131 = reverse_flag_65 ? _new_ptr_value_T_130 : {{1'd0}, new_value_65}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_66 = do_redirect_bits_cfiUpdate_histPtr_value + 8'h7; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_397 = {1'h0,new_value_66}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_66 = $signed(_diff_T_397) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_66 = $signed(diff_66) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_132 = $signed(_diff_T_397) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_133 = reverse_flag_66 ? _new_ptr_value_T_132 : {{1'd0}, new_value_66}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_67 = do_redirect_bits_cfiUpdate_histPtr_value + 8'h76; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_403 = {1'h0,new_value_67}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_67 = $signed(_diff_T_403) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_67 = $signed(diff_67) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_134 = $signed(_diff_T_403) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_135 = reverse_flag_67 ? _new_ptr_value_T_134 : {{1'd0}, new_value_67}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_68 = do_redirect_bits_cfiUpdate_histPtr_value + 8'h1d; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_409 = {1'h0,new_value_68}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_68 = $signed(_diff_T_409) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_68 = $signed(diff_68) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_136 = $signed(_diff_T_409) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_137 = reverse_flag_68 ? _new_ptr_value_T_136 : {{1'd0}, new_value_68}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_69 = do_redirect_bits_cfiUpdate_histPtr_value + 8'ha; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_415 = {1'h0,new_value_69}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_69 = $signed(_diff_T_415) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_69 = $signed(diff_69) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_138 = $signed(_diff_T_415) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_139 = reverse_flag_69 ? _new_ptr_value_T_138 : {{1'd0}, new_value_69}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_70 = do_redirect_bits_cfiUpdate_histPtr_value + 8'he; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_421 = {1'h0,new_value_70}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_70 = $signed(_diff_T_421) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_70 = $signed(diff_70) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_140 = $signed(_diff_T_421) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_141 = reverse_flag_70 ? _new_ptr_value_T_140 : {{1'd0}, new_value_70}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_71 = do_redirect_bits_cfiUpdate_histPtr_value + 8'h77; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_427 = {1'h0,new_value_71}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_71 = $signed(_diff_T_427) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_71 = $signed(diff_71) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_142 = $signed(_diff_T_427) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_143 = reverse_flag_71 ? _new_ptr_value_T_142 : {{1'd0}, new_value_71}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_72 = do_redirect_bits_cfiUpdate_histPtr_value + 8'hd; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_433 = {1'h0,new_value_72}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_72 = $signed(_diff_T_433) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_72 = $signed(diff_72) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_144 = $signed(_diff_T_433) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_145 = reverse_flag_72 ? _new_ptr_value_T_144 : {{1'd0}, new_value_72}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_73 = do_redirect_bits_cfiUpdate_histPtr_value + 8'h8; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_439 = {1'h0,new_value_73}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_73 = $signed(_diff_T_439) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_73 = $signed(diff_73) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_146 = $signed(_diff_T_439) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_147 = reverse_flag_73 ? _new_ptr_value_T_146 : {{1'd0}, new_value_73}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_74 = do_redirect_bits_cfiUpdate_histPtr_value + 8'h20; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_445 = {1'h0,new_value_74}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_74 = $signed(_diff_T_445) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_74 = $signed(diff_74) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_148 = $signed(_diff_T_445) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_149 = reverse_flag_74 ? _new_ptr_value_T_148 : {{1'd0}, new_value_74}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_75 = do_redirect_bits_cfiUpdate_histPtr_value + 8'hc; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_451 = {1'h0,new_value_75}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_75 = $signed(_diff_T_451) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_75 = $signed(diff_75) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_150 = $signed(_diff_T_451) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_151 = reverse_flag_75 ? _new_ptr_value_T_150 : {{1'd0}, new_value_75}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_76 = do_redirect_bits_cfiUpdate_histPtr_value + 8'h9; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_457 = {1'h0,new_value_76}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_76 = $signed(_diff_T_457) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_76 = $signed(diff_76) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_152 = $signed(_diff_T_457) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_153 = reverse_flag_76 ? _new_ptr_value_T_152 : {{1'd0}, new_value_76}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_77 = do_redirect_bits_cfiUpdate_histPtr_value + 8'h1f; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_463 = {1'h0,new_value_77}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_77 = $signed(_diff_T_463) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_77 = $signed(diff_77) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_154 = $signed(_diff_T_463) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_155 = reverse_flag_77 ? _new_ptr_value_T_154 : {{1'd0}, new_value_77}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_78 = do_redirect_bits_cfiUpdate_histPtr_value + 8'h5; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_469 = {1'h0,new_value_78}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_78 = $signed(_diff_T_469) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_78 = $signed(diff_78) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_156 = $signed(_diff_T_469) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_157 = reverse_flag_78 ? _new_ptr_value_T_156 : {{1'd0}, new_value_78}; // @[CircularQueuePtr.scala 45:27]
  wire [8:0] new_value_79 = do_redirect_bits_cfiUpdate_histPtr_value + 8'h10; // @[CircularQueuePtr.scala 41:34]
  wire [9:0] _diff_T_475 = {1'h0,new_value_79}; // @[CircularQueuePtr.scala 42:49]
  wire [9:0] diff_79 = $signed(_diff_T_475) - 10'sh90; // @[CircularQueuePtr.scala 42:52]
  wire  reverse_flag_79 = $signed(diff_79) >= 10'sh0; // @[CircularQueuePtr.scala 43:31]
  wire [9:0] _new_ptr_value_T_158 = $signed(_diff_T_475) - 10'sh90; // @[CircularQueuePtr.scala 46:20]
  wire [9:0] _new_ptr_value_T_159 = reverse_flag_79 ? _new_ptr_value_T_158 : {{1'd0}, new_value_79}; // @[CircularQueuePtr.scala 45:27]
  wire [7:0] new_ptr_69_value = _new_ptr_value_T_139[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_8830 = 8'h1 == new_ptr_69_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8831 = 8'h2 == new_ptr_69_value ? ghv_2 : _GEN_8830; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8832 = 8'h3 == new_ptr_69_value ? ghv_3 : _GEN_8831; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8833 = 8'h4 == new_ptr_69_value ? ghv_4 : _GEN_8832; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8834 = 8'h5 == new_ptr_69_value ? ghv_5 : _GEN_8833; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8835 = 8'h6 == new_ptr_69_value ? ghv_6 : _GEN_8834; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8836 = 8'h7 == new_ptr_69_value ? ghv_7 : _GEN_8835; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8837 = 8'h8 == new_ptr_69_value ? ghv_8 : _GEN_8836; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8838 = 8'h9 == new_ptr_69_value ? ghv_9 : _GEN_8837; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8839 = 8'ha == new_ptr_69_value ? ghv_10 : _GEN_8838; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8840 = 8'hb == new_ptr_69_value ? ghv_11 : _GEN_8839; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8841 = 8'hc == new_ptr_69_value ? ghv_12 : _GEN_8840; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8842 = 8'hd == new_ptr_69_value ? ghv_13 : _GEN_8841; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8843 = 8'he == new_ptr_69_value ? ghv_14 : _GEN_8842; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8844 = 8'hf == new_ptr_69_value ? ghv_15 : _GEN_8843; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8845 = 8'h10 == new_ptr_69_value ? ghv_16 : _GEN_8844; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8846 = 8'h11 == new_ptr_69_value ? ghv_17 : _GEN_8845; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8847 = 8'h12 == new_ptr_69_value ? ghv_18 : _GEN_8846; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8848 = 8'h13 == new_ptr_69_value ? ghv_19 : _GEN_8847; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8849 = 8'h14 == new_ptr_69_value ? ghv_20 : _GEN_8848; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8850 = 8'h15 == new_ptr_69_value ? ghv_21 : _GEN_8849; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8851 = 8'h16 == new_ptr_69_value ? ghv_22 : _GEN_8850; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8852 = 8'h17 == new_ptr_69_value ? ghv_23 : _GEN_8851; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8853 = 8'h18 == new_ptr_69_value ? ghv_24 : _GEN_8852; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8854 = 8'h19 == new_ptr_69_value ? ghv_25 : _GEN_8853; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8855 = 8'h1a == new_ptr_69_value ? ghv_26 : _GEN_8854; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8856 = 8'h1b == new_ptr_69_value ? ghv_27 : _GEN_8855; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8857 = 8'h1c == new_ptr_69_value ? ghv_28 : _GEN_8856; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8858 = 8'h1d == new_ptr_69_value ? ghv_29 : _GEN_8857; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8859 = 8'h1e == new_ptr_69_value ? ghv_30 : _GEN_8858; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8860 = 8'h1f == new_ptr_69_value ? ghv_31 : _GEN_8859; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8861 = 8'h20 == new_ptr_69_value ? ghv_32 : _GEN_8860; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8862 = 8'h21 == new_ptr_69_value ? ghv_33 : _GEN_8861; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8863 = 8'h22 == new_ptr_69_value ? ghv_34 : _GEN_8862; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8864 = 8'h23 == new_ptr_69_value ? ghv_35 : _GEN_8863; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8865 = 8'h24 == new_ptr_69_value ? ghv_36 : _GEN_8864; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8866 = 8'h25 == new_ptr_69_value ? ghv_37 : _GEN_8865; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8867 = 8'h26 == new_ptr_69_value ? ghv_38 : _GEN_8866; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8868 = 8'h27 == new_ptr_69_value ? ghv_39 : _GEN_8867; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8869 = 8'h28 == new_ptr_69_value ? ghv_40 : _GEN_8868; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8870 = 8'h29 == new_ptr_69_value ? ghv_41 : _GEN_8869; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8871 = 8'h2a == new_ptr_69_value ? ghv_42 : _GEN_8870; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8872 = 8'h2b == new_ptr_69_value ? ghv_43 : _GEN_8871; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8873 = 8'h2c == new_ptr_69_value ? ghv_44 : _GEN_8872; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8874 = 8'h2d == new_ptr_69_value ? ghv_45 : _GEN_8873; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8875 = 8'h2e == new_ptr_69_value ? ghv_46 : _GEN_8874; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8876 = 8'h2f == new_ptr_69_value ? ghv_47 : _GEN_8875; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8877 = 8'h30 == new_ptr_69_value ? ghv_48 : _GEN_8876; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8878 = 8'h31 == new_ptr_69_value ? ghv_49 : _GEN_8877; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8879 = 8'h32 == new_ptr_69_value ? ghv_50 : _GEN_8878; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8880 = 8'h33 == new_ptr_69_value ? ghv_51 : _GEN_8879; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8881 = 8'h34 == new_ptr_69_value ? ghv_52 : _GEN_8880; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8882 = 8'h35 == new_ptr_69_value ? ghv_53 : _GEN_8881; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8883 = 8'h36 == new_ptr_69_value ? ghv_54 : _GEN_8882; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8884 = 8'h37 == new_ptr_69_value ? ghv_55 : _GEN_8883; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8885 = 8'h38 == new_ptr_69_value ? ghv_56 : _GEN_8884; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8886 = 8'h39 == new_ptr_69_value ? ghv_57 : _GEN_8885; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8887 = 8'h3a == new_ptr_69_value ? ghv_58 : _GEN_8886; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8888 = 8'h3b == new_ptr_69_value ? ghv_59 : _GEN_8887; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8889 = 8'h3c == new_ptr_69_value ? ghv_60 : _GEN_8888; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8890 = 8'h3d == new_ptr_69_value ? ghv_61 : _GEN_8889; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8891 = 8'h3e == new_ptr_69_value ? ghv_62 : _GEN_8890; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8892 = 8'h3f == new_ptr_69_value ? ghv_63 : _GEN_8891; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8893 = 8'h40 == new_ptr_69_value ? ghv_64 : _GEN_8892; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8894 = 8'h41 == new_ptr_69_value ? ghv_65 : _GEN_8893; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8895 = 8'h42 == new_ptr_69_value ? ghv_66 : _GEN_8894; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8896 = 8'h43 == new_ptr_69_value ? ghv_67 : _GEN_8895; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8897 = 8'h44 == new_ptr_69_value ? ghv_68 : _GEN_8896; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8898 = 8'h45 == new_ptr_69_value ? ghv_69 : _GEN_8897; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8899 = 8'h46 == new_ptr_69_value ? ghv_70 : _GEN_8898; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8900 = 8'h47 == new_ptr_69_value ? ghv_71 : _GEN_8899; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8901 = 8'h48 == new_ptr_69_value ? ghv_72 : _GEN_8900; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8902 = 8'h49 == new_ptr_69_value ? ghv_73 : _GEN_8901; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8903 = 8'h4a == new_ptr_69_value ? ghv_74 : _GEN_8902; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8904 = 8'h4b == new_ptr_69_value ? ghv_75 : _GEN_8903; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8905 = 8'h4c == new_ptr_69_value ? ghv_76 : _GEN_8904; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8906 = 8'h4d == new_ptr_69_value ? ghv_77 : _GEN_8905; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8907 = 8'h4e == new_ptr_69_value ? ghv_78 : _GEN_8906; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8908 = 8'h4f == new_ptr_69_value ? ghv_79 : _GEN_8907; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8909 = 8'h50 == new_ptr_69_value ? ghv_80 : _GEN_8908; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8910 = 8'h51 == new_ptr_69_value ? ghv_81 : _GEN_8909; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8911 = 8'h52 == new_ptr_69_value ? ghv_82 : _GEN_8910; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8912 = 8'h53 == new_ptr_69_value ? ghv_83 : _GEN_8911; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8913 = 8'h54 == new_ptr_69_value ? ghv_84 : _GEN_8912; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8914 = 8'h55 == new_ptr_69_value ? ghv_85 : _GEN_8913; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8915 = 8'h56 == new_ptr_69_value ? ghv_86 : _GEN_8914; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8916 = 8'h57 == new_ptr_69_value ? ghv_87 : _GEN_8915; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8917 = 8'h58 == new_ptr_69_value ? ghv_88 : _GEN_8916; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8918 = 8'h59 == new_ptr_69_value ? ghv_89 : _GEN_8917; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8919 = 8'h5a == new_ptr_69_value ? ghv_90 : _GEN_8918; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8920 = 8'h5b == new_ptr_69_value ? ghv_91 : _GEN_8919; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8921 = 8'h5c == new_ptr_69_value ? ghv_92 : _GEN_8920; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8922 = 8'h5d == new_ptr_69_value ? ghv_93 : _GEN_8921; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8923 = 8'h5e == new_ptr_69_value ? ghv_94 : _GEN_8922; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8924 = 8'h5f == new_ptr_69_value ? ghv_95 : _GEN_8923; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8925 = 8'h60 == new_ptr_69_value ? ghv_96 : _GEN_8924; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8926 = 8'h61 == new_ptr_69_value ? ghv_97 : _GEN_8925; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8927 = 8'h62 == new_ptr_69_value ? ghv_98 : _GEN_8926; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8928 = 8'h63 == new_ptr_69_value ? ghv_99 : _GEN_8927; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8929 = 8'h64 == new_ptr_69_value ? ghv_100 : _GEN_8928; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8930 = 8'h65 == new_ptr_69_value ? ghv_101 : _GEN_8929; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8931 = 8'h66 == new_ptr_69_value ? ghv_102 : _GEN_8930; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8932 = 8'h67 == new_ptr_69_value ? ghv_103 : _GEN_8931; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8933 = 8'h68 == new_ptr_69_value ? ghv_104 : _GEN_8932; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8934 = 8'h69 == new_ptr_69_value ? ghv_105 : _GEN_8933; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8935 = 8'h6a == new_ptr_69_value ? ghv_106 : _GEN_8934; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8936 = 8'h6b == new_ptr_69_value ? ghv_107 : _GEN_8935; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8937 = 8'h6c == new_ptr_69_value ? ghv_108 : _GEN_8936; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8938 = 8'h6d == new_ptr_69_value ? ghv_109 : _GEN_8937; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8939 = 8'h6e == new_ptr_69_value ? ghv_110 : _GEN_8938; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8940 = 8'h6f == new_ptr_69_value ? ghv_111 : _GEN_8939; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8941 = 8'h70 == new_ptr_69_value ? ghv_112 : _GEN_8940; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8942 = 8'h71 == new_ptr_69_value ? ghv_113 : _GEN_8941; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8943 = 8'h72 == new_ptr_69_value ? ghv_114 : _GEN_8942; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8944 = 8'h73 == new_ptr_69_value ? ghv_115 : _GEN_8943; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8945 = 8'h74 == new_ptr_69_value ? ghv_116 : _GEN_8944; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8946 = 8'h75 == new_ptr_69_value ? ghv_117 : _GEN_8945; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8947 = 8'h76 == new_ptr_69_value ? ghv_118 : _GEN_8946; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8948 = 8'h77 == new_ptr_69_value ? ghv_119 : _GEN_8947; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8949 = 8'h78 == new_ptr_69_value ? ghv_120 : _GEN_8948; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8950 = 8'h79 == new_ptr_69_value ? ghv_121 : _GEN_8949; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8951 = 8'h7a == new_ptr_69_value ? ghv_122 : _GEN_8950; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8952 = 8'h7b == new_ptr_69_value ? ghv_123 : _GEN_8951; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8953 = 8'h7c == new_ptr_69_value ? ghv_124 : _GEN_8952; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8954 = 8'h7d == new_ptr_69_value ? ghv_125 : _GEN_8953; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8955 = 8'h7e == new_ptr_69_value ? ghv_126 : _GEN_8954; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8956 = 8'h7f == new_ptr_69_value ? ghv_127 : _GEN_8955; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8957 = 8'h80 == new_ptr_69_value ? ghv_128 : _GEN_8956; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8958 = 8'h81 == new_ptr_69_value ? ghv_129 : _GEN_8957; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8959 = 8'h82 == new_ptr_69_value ? ghv_130 : _GEN_8958; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8960 = 8'h83 == new_ptr_69_value ? ghv_131 : _GEN_8959; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8961 = 8'h84 == new_ptr_69_value ? ghv_132 : _GEN_8960; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8962 = 8'h85 == new_ptr_69_value ? ghv_133 : _GEN_8961; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8963 = 8'h86 == new_ptr_69_value ? ghv_134 : _GEN_8962; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8964 = 8'h87 == new_ptr_69_value ? ghv_135 : _GEN_8963; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8965 = 8'h88 == new_ptr_69_value ? ghv_136 : _GEN_8964; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8966 = 8'h89 == new_ptr_69_value ? ghv_137 : _GEN_8965; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8967 = 8'h8a == new_ptr_69_value ? ghv_138 : _GEN_8966; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8968 = 8'h8b == new_ptr_69_value ? ghv_139 : _GEN_8967; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8969 = 8'h8c == new_ptr_69_value ? ghv_140 : _GEN_8968; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8970 = 8'h8d == new_ptr_69_value ? ghv_141 : _GEN_8969; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8971 = 8'h8e == new_ptr_69_value ? ghv_142 : _GEN_8970; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_76_value = _new_ptr_value_T_153[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_8974 = 8'h1 == new_ptr_76_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8975 = 8'h2 == new_ptr_76_value ? ghv_2 : _GEN_8974; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8976 = 8'h3 == new_ptr_76_value ? ghv_3 : _GEN_8975; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8977 = 8'h4 == new_ptr_76_value ? ghv_4 : _GEN_8976; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8978 = 8'h5 == new_ptr_76_value ? ghv_5 : _GEN_8977; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8979 = 8'h6 == new_ptr_76_value ? ghv_6 : _GEN_8978; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8980 = 8'h7 == new_ptr_76_value ? ghv_7 : _GEN_8979; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8981 = 8'h8 == new_ptr_76_value ? ghv_8 : _GEN_8980; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8982 = 8'h9 == new_ptr_76_value ? ghv_9 : _GEN_8981; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8983 = 8'ha == new_ptr_76_value ? ghv_10 : _GEN_8982; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8984 = 8'hb == new_ptr_76_value ? ghv_11 : _GEN_8983; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8985 = 8'hc == new_ptr_76_value ? ghv_12 : _GEN_8984; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8986 = 8'hd == new_ptr_76_value ? ghv_13 : _GEN_8985; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8987 = 8'he == new_ptr_76_value ? ghv_14 : _GEN_8986; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8988 = 8'hf == new_ptr_76_value ? ghv_15 : _GEN_8987; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8989 = 8'h10 == new_ptr_76_value ? ghv_16 : _GEN_8988; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8990 = 8'h11 == new_ptr_76_value ? ghv_17 : _GEN_8989; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8991 = 8'h12 == new_ptr_76_value ? ghv_18 : _GEN_8990; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8992 = 8'h13 == new_ptr_76_value ? ghv_19 : _GEN_8991; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8993 = 8'h14 == new_ptr_76_value ? ghv_20 : _GEN_8992; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8994 = 8'h15 == new_ptr_76_value ? ghv_21 : _GEN_8993; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8995 = 8'h16 == new_ptr_76_value ? ghv_22 : _GEN_8994; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8996 = 8'h17 == new_ptr_76_value ? ghv_23 : _GEN_8995; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8997 = 8'h18 == new_ptr_76_value ? ghv_24 : _GEN_8996; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8998 = 8'h19 == new_ptr_76_value ? ghv_25 : _GEN_8997; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_8999 = 8'h1a == new_ptr_76_value ? ghv_26 : _GEN_8998; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9000 = 8'h1b == new_ptr_76_value ? ghv_27 : _GEN_8999; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9001 = 8'h1c == new_ptr_76_value ? ghv_28 : _GEN_9000; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9002 = 8'h1d == new_ptr_76_value ? ghv_29 : _GEN_9001; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9003 = 8'h1e == new_ptr_76_value ? ghv_30 : _GEN_9002; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9004 = 8'h1f == new_ptr_76_value ? ghv_31 : _GEN_9003; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9005 = 8'h20 == new_ptr_76_value ? ghv_32 : _GEN_9004; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9006 = 8'h21 == new_ptr_76_value ? ghv_33 : _GEN_9005; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9007 = 8'h22 == new_ptr_76_value ? ghv_34 : _GEN_9006; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9008 = 8'h23 == new_ptr_76_value ? ghv_35 : _GEN_9007; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9009 = 8'h24 == new_ptr_76_value ? ghv_36 : _GEN_9008; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9010 = 8'h25 == new_ptr_76_value ? ghv_37 : _GEN_9009; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9011 = 8'h26 == new_ptr_76_value ? ghv_38 : _GEN_9010; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9012 = 8'h27 == new_ptr_76_value ? ghv_39 : _GEN_9011; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9013 = 8'h28 == new_ptr_76_value ? ghv_40 : _GEN_9012; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9014 = 8'h29 == new_ptr_76_value ? ghv_41 : _GEN_9013; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9015 = 8'h2a == new_ptr_76_value ? ghv_42 : _GEN_9014; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9016 = 8'h2b == new_ptr_76_value ? ghv_43 : _GEN_9015; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9017 = 8'h2c == new_ptr_76_value ? ghv_44 : _GEN_9016; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9018 = 8'h2d == new_ptr_76_value ? ghv_45 : _GEN_9017; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9019 = 8'h2e == new_ptr_76_value ? ghv_46 : _GEN_9018; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9020 = 8'h2f == new_ptr_76_value ? ghv_47 : _GEN_9019; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9021 = 8'h30 == new_ptr_76_value ? ghv_48 : _GEN_9020; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9022 = 8'h31 == new_ptr_76_value ? ghv_49 : _GEN_9021; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9023 = 8'h32 == new_ptr_76_value ? ghv_50 : _GEN_9022; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9024 = 8'h33 == new_ptr_76_value ? ghv_51 : _GEN_9023; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9025 = 8'h34 == new_ptr_76_value ? ghv_52 : _GEN_9024; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9026 = 8'h35 == new_ptr_76_value ? ghv_53 : _GEN_9025; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9027 = 8'h36 == new_ptr_76_value ? ghv_54 : _GEN_9026; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9028 = 8'h37 == new_ptr_76_value ? ghv_55 : _GEN_9027; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9029 = 8'h38 == new_ptr_76_value ? ghv_56 : _GEN_9028; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9030 = 8'h39 == new_ptr_76_value ? ghv_57 : _GEN_9029; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9031 = 8'h3a == new_ptr_76_value ? ghv_58 : _GEN_9030; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9032 = 8'h3b == new_ptr_76_value ? ghv_59 : _GEN_9031; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9033 = 8'h3c == new_ptr_76_value ? ghv_60 : _GEN_9032; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9034 = 8'h3d == new_ptr_76_value ? ghv_61 : _GEN_9033; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9035 = 8'h3e == new_ptr_76_value ? ghv_62 : _GEN_9034; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9036 = 8'h3f == new_ptr_76_value ? ghv_63 : _GEN_9035; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9037 = 8'h40 == new_ptr_76_value ? ghv_64 : _GEN_9036; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9038 = 8'h41 == new_ptr_76_value ? ghv_65 : _GEN_9037; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9039 = 8'h42 == new_ptr_76_value ? ghv_66 : _GEN_9038; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9040 = 8'h43 == new_ptr_76_value ? ghv_67 : _GEN_9039; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9041 = 8'h44 == new_ptr_76_value ? ghv_68 : _GEN_9040; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9042 = 8'h45 == new_ptr_76_value ? ghv_69 : _GEN_9041; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9043 = 8'h46 == new_ptr_76_value ? ghv_70 : _GEN_9042; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9044 = 8'h47 == new_ptr_76_value ? ghv_71 : _GEN_9043; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9045 = 8'h48 == new_ptr_76_value ? ghv_72 : _GEN_9044; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9046 = 8'h49 == new_ptr_76_value ? ghv_73 : _GEN_9045; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9047 = 8'h4a == new_ptr_76_value ? ghv_74 : _GEN_9046; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9048 = 8'h4b == new_ptr_76_value ? ghv_75 : _GEN_9047; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9049 = 8'h4c == new_ptr_76_value ? ghv_76 : _GEN_9048; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9050 = 8'h4d == new_ptr_76_value ? ghv_77 : _GEN_9049; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9051 = 8'h4e == new_ptr_76_value ? ghv_78 : _GEN_9050; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9052 = 8'h4f == new_ptr_76_value ? ghv_79 : _GEN_9051; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9053 = 8'h50 == new_ptr_76_value ? ghv_80 : _GEN_9052; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9054 = 8'h51 == new_ptr_76_value ? ghv_81 : _GEN_9053; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9055 = 8'h52 == new_ptr_76_value ? ghv_82 : _GEN_9054; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9056 = 8'h53 == new_ptr_76_value ? ghv_83 : _GEN_9055; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9057 = 8'h54 == new_ptr_76_value ? ghv_84 : _GEN_9056; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9058 = 8'h55 == new_ptr_76_value ? ghv_85 : _GEN_9057; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9059 = 8'h56 == new_ptr_76_value ? ghv_86 : _GEN_9058; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9060 = 8'h57 == new_ptr_76_value ? ghv_87 : _GEN_9059; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9061 = 8'h58 == new_ptr_76_value ? ghv_88 : _GEN_9060; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9062 = 8'h59 == new_ptr_76_value ? ghv_89 : _GEN_9061; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9063 = 8'h5a == new_ptr_76_value ? ghv_90 : _GEN_9062; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9064 = 8'h5b == new_ptr_76_value ? ghv_91 : _GEN_9063; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9065 = 8'h5c == new_ptr_76_value ? ghv_92 : _GEN_9064; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9066 = 8'h5d == new_ptr_76_value ? ghv_93 : _GEN_9065; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9067 = 8'h5e == new_ptr_76_value ? ghv_94 : _GEN_9066; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9068 = 8'h5f == new_ptr_76_value ? ghv_95 : _GEN_9067; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9069 = 8'h60 == new_ptr_76_value ? ghv_96 : _GEN_9068; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9070 = 8'h61 == new_ptr_76_value ? ghv_97 : _GEN_9069; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9071 = 8'h62 == new_ptr_76_value ? ghv_98 : _GEN_9070; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9072 = 8'h63 == new_ptr_76_value ? ghv_99 : _GEN_9071; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9073 = 8'h64 == new_ptr_76_value ? ghv_100 : _GEN_9072; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9074 = 8'h65 == new_ptr_76_value ? ghv_101 : _GEN_9073; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9075 = 8'h66 == new_ptr_76_value ? ghv_102 : _GEN_9074; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9076 = 8'h67 == new_ptr_76_value ? ghv_103 : _GEN_9075; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9077 = 8'h68 == new_ptr_76_value ? ghv_104 : _GEN_9076; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9078 = 8'h69 == new_ptr_76_value ? ghv_105 : _GEN_9077; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9079 = 8'h6a == new_ptr_76_value ? ghv_106 : _GEN_9078; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9080 = 8'h6b == new_ptr_76_value ? ghv_107 : _GEN_9079; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9081 = 8'h6c == new_ptr_76_value ? ghv_108 : _GEN_9080; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9082 = 8'h6d == new_ptr_76_value ? ghv_109 : _GEN_9081; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9083 = 8'h6e == new_ptr_76_value ? ghv_110 : _GEN_9082; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9084 = 8'h6f == new_ptr_76_value ? ghv_111 : _GEN_9083; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9085 = 8'h70 == new_ptr_76_value ? ghv_112 : _GEN_9084; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9086 = 8'h71 == new_ptr_76_value ? ghv_113 : _GEN_9085; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9087 = 8'h72 == new_ptr_76_value ? ghv_114 : _GEN_9086; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9088 = 8'h73 == new_ptr_76_value ? ghv_115 : _GEN_9087; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9089 = 8'h74 == new_ptr_76_value ? ghv_116 : _GEN_9088; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9090 = 8'h75 == new_ptr_76_value ? ghv_117 : _GEN_9089; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9091 = 8'h76 == new_ptr_76_value ? ghv_118 : _GEN_9090; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9092 = 8'h77 == new_ptr_76_value ? ghv_119 : _GEN_9091; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9093 = 8'h78 == new_ptr_76_value ? ghv_120 : _GEN_9092; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9094 = 8'h79 == new_ptr_76_value ? ghv_121 : _GEN_9093; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9095 = 8'h7a == new_ptr_76_value ? ghv_122 : _GEN_9094; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9096 = 8'h7b == new_ptr_76_value ? ghv_123 : _GEN_9095; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9097 = 8'h7c == new_ptr_76_value ? ghv_124 : _GEN_9096; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9098 = 8'h7d == new_ptr_76_value ? ghv_125 : _GEN_9097; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9099 = 8'h7e == new_ptr_76_value ? ghv_126 : _GEN_9098; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9100 = 8'h7f == new_ptr_76_value ? ghv_127 : _GEN_9099; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9101 = 8'h80 == new_ptr_76_value ? ghv_128 : _GEN_9100; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9102 = 8'h81 == new_ptr_76_value ? ghv_129 : _GEN_9101; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9103 = 8'h82 == new_ptr_76_value ? ghv_130 : _GEN_9102; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9104 = 8'h83 == new_ptr_76_value ? ghv_131 : _GEN_9103; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9105 = 8'h84 == new_ptr_76_value ? ghv_132 : _GEN_9104; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9106 = 8'h85 == new_ptr_76_value ? ghv_133 : _GEN_9105; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9107 = 8'h86 == new_ptr_76_value ? ghv_134 : _GEN_9106; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9108 = 8'h87 == new_ptr_76_value ? ghv_135 : _GEN_9107; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9109 = 8'h88 == new_ptr_76_value ? ghv_136 : _GEN_9108; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9110 = 8'h89 == new_ptr_76_value ? ghv_137 : _GEN_9109; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9111 = 8'h8a == new_ptr_76_value ? ghv_138 : _GEN_9110; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9112 = 8'h8b == new_ptr_76_value ? ghv_139 : _GEN_9111; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9113 = 8'h8c == new_ptr_76_value ? ghv_140 : _GEN_9112; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9114 = 8'h8d == new_ptr_76_value ? ghv_141 : _GEN_9113; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9115 = 8'h8e == new_ptr_76_value ? ghv_142 : _GEN_9114; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_73_value = _new_ptr_value_T_147[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_9118 = 8'h1 == new_ptr_73_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9119 = 8'h2 == new_ptr_73_value ? ghv_2 : _GEN_9118; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9120 = 8'h3 == new_ptr_73_value ? ghv_3 : _GEN_9119; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9121 = 8'h4 == new_ptr_73_value ? ghv_4 : _GEN_9120; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9122 = 8'h5 == new_ptr_73_value ? ghv_5 : _GEN_9121; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9123 = 8'h6 == new_ptr_73_value ? ghv_6 : _GEN_9122; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9124 = 8'h7 == new_ptr_73_value ? ghv_7 : _GEN_9123; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9125 = 8'h8 == new_ptr_73_value ? ghv_8 : _GEN_9124; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9126 = 8'h9 == new_ptr_73_value ? ghv_9 : _GEN_9125; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9127 = 8'ha == new_ptr_73_value ? ghv_10 : _GEN_9126; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9128 = 8'hb == new_ptr_73_value ? ghv_11 : _GEN_9127; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9129 = 8'hc == new_ptr_73_value ? ghv_12 : _GEN_9128; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9130 = 8'hd == new_ptr_73_value ? ghv_13 : _GEN_9129; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9131 = 8'he == new_ptr_73_value ? ghv_14 : _GEN_9130; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9132 = 8'hf == new_ptr_73_value ? ghv_15 : _GEN_9131; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9133 = 8'h10 == new_ptr_73_value ? ghv_16 : _GEN_9132; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9134 = 8'h11 == new_ptr_73_value ? ghv_17 : _GEN_9133; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9135 = 8'h12 == new_ptr_73_value ? ghv_18 : _GEN_9134; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9136 = 8'h13 == new_ptr_73_value ? ghv_19 : _GEN_9135; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9137 = 8'h14 == new_ptr_73_value ? ghv_20 : _GEN_9136; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9138 = 8'h15 == new_ptr_73_value ? ghv_21 : _GEN_9137; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9139 = 8'h16 == new_ptr_73_value ? ghv_22 : _GEN_9138; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9140 = 8'h17 == new_ptr_73_value ? ghv_23 : _GEN_9139; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9141 = 8'h18 == new_ptr_73_value ? ghv_24 : _GEN_9140; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9142 = 8'h19 == new_ptr_73_value ? ghv_25 : _GEN_9141; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9143 = 8'h1a == new_ptr_73_value ? ghv_26 : _GEN_9142; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9144 = 8'h1b == new_ptr_73_value ? ghv_27 : _GEN_9143; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9145 = 8'h1c == new_ptr_73_value ? ghv_28 : _GEN_9144; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9146 = 8'h1d == new_ptr_73_value ? ghv_29 : _GEN_9145; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9147 = 8'h1e == new_ptr_73_value ? ghv_30 : _GEN_9146; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9148 = 8'h1f == new_ptr_73_value ? ghv_31 : _GEN_9147; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9149 = 8'h20 == new_ptr_73_value ? ghv_32 : _GEN_9148; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9150 = 8'h21 == new_ptr_73_value ? ghv_33 : _GEN_9149; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9151 = 8'h22 == new_ptr_73_value ? ghv_34 : _GEN_9150; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9152 = 8'h23 == new_ptr_73_value ? ghv_35 : _GEN_9151; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9153 = 8'h24 == new_ptr_73_value ? ghv_36 : _GEN_9152; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9154 = 8'h25 == new_ptr_73_value ? ghv_37 : _GEN_9153; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9155 = 8'h26 == new_ptr_73_value ? ghv_38 : _GEN_9154; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9156 = 8'h27 == new_ptr_73_value ? ghv_39 : _GEN_9155; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9157 = 8'h28 == new_ptr_73_value ? ghv_40 : _GEN_9156; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9158 = 8'h29 == new_ptr_73_value ? ghv_41 : _GEN_9157; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9159 = 8'h2a == new_ptr_73_value ? ghv_42 : _GEN_9158; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9160 = 8'h2b == new_ptr_73_value ? ghv_43 : _GEN_9159; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9161 = 8'h2c == new_ptr_73_value ? ghv_44 : _GEN_9160; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9162 = 8'h2d == new_ptr_73_value ? ghv_45 : _GEN_9161; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9163 = 8'h2e == new_ptr_73_value ? ghv_46 : _GEN_9162; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9164 = 8'h2f == new_ptr_73_value ? ghv_47 : _GEN_9163; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9165 = 8'h30 == new_ptr_73_value ? ghv_48 : _GEN_9164; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9166 = 8'h31 == new_ptr_73_value ? ghv_49 : _GEN_9165; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9167 = 8'h32 == new_ptr_73_value ? ghv_50 : _GEN_9166; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9168 = 8'h33 == new_ptr_73_value ? ghv_51 : _GEN_9167; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9169 = 8'h34 == new_ptr_73_value ? ghv_52 : _GEN_9168; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9170 = 8'h35 == new_ptr_73_value ? ghv_53 : _GEN_9169; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9171 = 8'h36 == new_ptr_73_value ? ghv_54 : _GEN_9170; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9172 = 8'h37 == new_ptr_73_value ? ghv_55 : _GEN_9171; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9173 = 8'h38 == new_ptr_73_value ? ghv_56 : _GEN_9172; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9174 = 8'h39 == new_ptr_73_value ? ghv_57 : _GEN_9173; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9175 = 8'h3a == new_ptr_73_value ? ghv_58 : _GEN_9174; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9176 = 8'h3b == new_ptr_73_value ? ghv_59 : _GEN_9175; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9177 = 8'h3c == new_ptr_73_value ? ghv_60 : _GEN_9176; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9178 = 8'h3d == new_ptr_73_value ? ghv_61 : _GEN_9177; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9179 = 8'h3e == new_ptr_73_value ? ghv_62 : _GEN_9178; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9180 = 8'h3f == new_ptr_73_value ? ghv_63 : _GEN_9179; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9181 = 8'h40 == new_ptr_73_value ? ghv_64 : _GEN_9180; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9182 = 8'h41 == new_ptr_73_value ? ghv_65 : _GEN_9181; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9183 = 8'h42 == new_ptr_73_value ? ghv_66 : _GEN_9182; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9184 = 8'h43 == new_ptr_73_value ? ghv_67 : _GEN_9183; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9185 = 8'h44 == new_ptr_73_value ? ghv_68 : _GEN_9184; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9186 = 8'h45 == new_ptr_73_value ? ghv_69 : _GEN_9185; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9187 = 8'h46 == new_ptr_73_value ? ghv_70 : _GEN_9186; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9188 = 8'h47 == new_ptr_73_value ? ghv_71 : _GEN_9187; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9189 = 8'h48 == new_ptr_73_value ? ghv_72 : _GEN_9188; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9190 = 8'h49 == new_ptr_73_value ? ghv_73 : _GEN_9189; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9191 = 8'h4a == new_ptr_73_value ? ghv_74 : _GEN_9190; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9192 = 8'h4b == new_ptr_73_value ? ghv_75 : _GEN_9191; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9193 = 8'h4c == new_ptr_73_value ? ghv_76 : _GEN_9192; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9194 = 8'h4d == new_ptr_73_value ? ghv_77 : _GEN_9193; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9195 = 8'h4e == new_ptr_73_value ? ghv_78 : _GEN_9194; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9196 = 8'h4f == new_ptr_73_value ? ghv_79 : _GEN_9195; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9197 = 8'h50 == new_ptr_73_value ? ghv_80 : _GEN_9196; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9198 = 8'h51 == new_ptr_73_value ? ghv_81 : _GEN_9197; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9199 = 8'h52 == new_ptr_73_value ? ghv_82 : _GEN_9198; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9200 = 8'h53 == new_ptr_73_value ? ghv_83 : _GEN_9199; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9201 = 8'h54 == new_ptr_73_value ? ghv_84 : _GEN_9200; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9202 = 8'h55 == new_ptr_73_value ? ghv_85 : _GEN_9201; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9203 = 8'h56 == new_ptr_73_value ? ghv_86 : _GEN_9202; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9204 = 8'h57 == new_ptr_73_value ? ghv_87 : _GEN_9203; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9205 = 8'h58 == new_ptr_73_value ? ghv_88 : _GEN_9204; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9206 = 8'h59 == new_ptr_73_value ? ghv_89 : _GEN_9205; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9207 = 8'h5a == new_ptr_73_value ? ghv_90 : _GEN_9206; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9208 = 8'h5b == new_ptr_73_value ? ghv_91 : _GEN_9207; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9209 = 8'h5c == new_ptr_73_value ? ghv_92 : _GEN_9208; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9210 = 8'h5d == new_ptr_73_value ? ghv_93 : _GEN_9209; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9211 = 8'h5e == new_ptr_73_value ? ghv_94 : _GEN_9210; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9212 = 8'h5f == new_ptr_73_value ? ghv_95 : _GEN_9211; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9213 = 8'h60 == new_ptr_73_value ? ghv_96 : _GEN_9212; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9214 = 8'h61 == new_ptr_73_value ? ghv_97 : _GEN_9213; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9215 = 8'h62 == new_ptr_73_value ? ghv_98 : _GEN_9214; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9216 = 8'h63 == new_ptr_73_value ? ghv_99 : _GEN_9215; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9217 = 8'h64 == new_ptr_73_value ? ghv_100 : _GEN_9216; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9218 = 8'h65 == new_ptr_73_value ? ghv_101 : _GEN_9217; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9219 = 8'h66 == new_ptr_73_value ? ghv_102 : _GEN_9218; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9220 = 8'h67 == new_ptr_73_value ? ghv_103 : _GEN_9219; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9221 = 8'h68 == new_ptr_73_value ? ghv_104 : _GEN_9220; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9222 = 8'h69 == new_ptr_73_value ? ghv_105 : _GEN_9221; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9223 = 8'h6a == new_ptr_73_value ? ghv_106 : _GEN_9222; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9224 = 8'h6b == new_ptr_73_value ? ghv_107 : _GEN_9223; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9225 = 8'h6c == new_ptr_73_value ? ghv_108 : _GEN_9224; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9226 = 8'h6d == new_ptr_73_value ? ghv_109 : _GEN_9225; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9227 = 8'h6e == new_ptr_73_value ? ghv_110 : _GEN_9226; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9228 = 8'h6f == new_ptr_73_value ? ghv_111 : _GEN_9227; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9229 = 8'h70 == new_ptr_73_value ? ghv_112 : _GEN_9228; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9230 = 8'h71 == new_ptr_73_value ? ghv_113 : _GEN_9229; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9231 = 8'h72 == new_ptr_73_value ? ghv_114 : _GEN_9230; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9232 = 8'h73 == new_ptr_73_value ? ghv_115 : _GEN_9231; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9233 = 8'h74 == new_ptr_73_value ? ghv_116 : _GEN_9232; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9234 = 8'h75 == new_ptr_73_value ? ghv_117 : _GEN_9233; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9235 = 8'h76 == new_ptr_73_value ? ghv_118 : _GEN_9234; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9236 = 8'h77 == new_ptr_73_value ? ghv_119 : _GEN_9235; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9237 = 8'h78 == new_ptr_73_value ? ghv_120 : _GEN_9236; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9238 = 8'h79 == new_ptr_73_value ? ghv_121 : _GEN_9237; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9239 = 8'h7a == new_ptr_73_value ? ghv_122 : _GEN_9238; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9240 = 8'h7b == new_ptr_73_value ? ghv_123 : _GEN_9239; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9241 = 8'h7c == new_ptr_73_value ? ghv_124 : _GEN_9240; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9242 = 8'h7d == new_ptr_73_value ? ghv_125 : _GEN_9241; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9243 = 8'h7e == new_ptr_73_value ? ghv_126 : _GEN_9242; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9244 = 8'h7f == new_ptr_73_value ? ghv_127 : _GEN_9243; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9245 = 8'h80 == new_ptr_73_value ? ghv_128 : _GEN_9244; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9246 = 8'h81 == new_ptr_73_value ? ghv_129 : _GEN_9245; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9247 = 8'h82 == new_ptr_73_value ? ghv_130 : _GEN_9246; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9248 = 8'h83 == new_ptr_73_value ? ghv_131 : _GEN_9247; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9249 = 8'h84 == new_ptr_73_value ? ghv_132 : _GEN_9248; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9250 = 8'h85 == new_ptr_73_value ? ghv_133 : _GEN_9249; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9251 = 8'h86 == new_ptr_73_value ? ghv_134 : _GEN_9250; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9252 = 8'h87 == new_ptr_73_value ? ghv_135 : _GEN_9251; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9253 = 8'h88 == new_ptr_73_value ? ghv_136 : _GEN_9252; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9254 = 8'h89 == new_ptr_73_value ? ghv_137 : _GEN_9253; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9255 = 8'h8a == new_ptr_73_value ? ghv_138 : _GEN_9254; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9256 = 8'h8b == new_ptr_73_value ? ghv_139 : _GEN_9255; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9257 = 8'h8c == new_ptr_73_value ? ghv_140 : _GEN_9256; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9258 = 8'h8d == new_ptr_73_value ? ghv_141 : _GEN_9257; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9259 = 8'h8e == new_ptr_73_value ? ghv_142 : _GEN_9258; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_66_value = _new_ptr_value_T_133[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_9262 = 8'h1 == new_ptr_66_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9263 = 8'h2 == new_ptr_66_value ? ghv_2 : _GEN_9262; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9264 = 8'h3 == new_ptr_66_value ? ghv_3 : _GEN_9263; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9265 = 8'h4 == new_ptr_66_value ? ghv_4 : _GEN_9264; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9266 = 8'h5 == new_ptr_66_value ? ghv_5 : _GEN_9265; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9267 = 8'h6 == new_ptr_66_value ? ghv_6 : _GEN_9266; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9268 = 8'h7 == new_ptr_66_value ? ghv_7 : _GEN_9267; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9269 = 8'h8 == new_ptr_66_value ? ghv_8 : _GEN_9268; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9270 = 8'h9 == new_ptr_66_value ? ghv_9 : _GEN_9269; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9271 = 8'ha == new_ptr_66_value ? ghv_10 : _GEN_9270; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9272 = 8'hb == new_ptr_66_value ? ghv_11 : _GEN_9271; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9273 = 8'hc == new_ptr_66_value ? ghv_12 : _GEN_9272; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9274 = 8'hd == new_ptr_66_value ? ghv_13 : _GEN_9273; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9275 = 8'he == new_ptr_66_value ? ghv_14 : _GEN_9274; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9276 = 8'hf == new_ptr_66_value ? ghv_15 : _GEN_9275; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9277 = 8'h10 == new_ptr_66_value ? ghv_16 : _GEN_9276; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9278 = 8'h11 == new_ptr_66_value ? ghv_17 : _GEN_9277; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9279 = 8'h12 == new_ptr_66_value ? ghv_18 : _GEN_9278; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9280 = 8'h13 == new_ptr_66_value ? ghv_19 : _GEN_9279; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9281 = 8'h14 == new_ptr_66_value ? ghv_20 : _GEN_9280; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9282 = 8'h15 == new_ptr_66_value ? ghv_21 : _GEN_9281; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9283 = 8'h16 == new_ptr_66_value ? ghv_22 : _GEN_9282; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9284 = 8'h17 == new_ptr_66_value ? ghv_23 : _GEN_9283; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9285 = 8'h18 == new_ptr_66_value ? ghv_24 : _GEN_9284; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9286 = 8'h19 == new_ptr_66_value ? ghv_25 : _GEN_9285; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9287 = 8'h1a == new_ptr_66_value ? ghv_26 : _GEN_9286; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9288 = 8'h1b == new_ptr_66_value ? ghv_27 : _GEN_9287; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9289 = 8'h1c == new_ptr_66_value ? ghv_28 : _GEN_9288; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9290 = 8'h1d == new_ptr_66_value ? ghv_29 : _GEN_9289; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9291 = 8'h1e == new_ptr_66_value ? ghv_30 : _GEN_9290; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9292 = 8'h1f == new_ptr_66_value ? ghv_31 : _GEN_9291; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9293 = 8'h20 == new_ptr_66_value ? ghv_32 : _GEN_9292; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9294 = 8'h21 == new_ptr_66_value ? ghv_33 : _GEN_9293; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9295 = 8'h22 == new_ptr_66_value ? ghv_34 : _GEN_9294; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9296 = 8'h23 == new_ptr_66_value ? ghv_35 : _GEN_9295; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9297 = 8'h24 == new_ptr_66_value ? ghv_36 : _GEN_9296; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9298 = 8'h25 == new_ptr_66_value ? ghv_37 : _GEN_9297; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9299 = 8'h26 == new_ptr_66_value ? ghv_38 : _GEN_9298; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9300 = 8'h27 == new_ptr_66_value ? ghv_39 : _GEN_9299; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9301 = 8'h28 == new_ptr_66_value ? ghv_40 : _GEN_9300; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9302 = 8'h29 == new_ptr_66_value ? ghv_41 : _GEN_9301; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9303 = 8'h2a == new_ptr_66_value ? ghv_42 : _GEN_9302; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9304 = 8'h2b == new_ptr_66_value ? ghv_43 : _GEN_9303; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9305 = 8'h2c == new_ptr_66_value ? ghv_44 : _GEN_9304; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9306 = 8'h2d == new_ptr_66_value ? ghv_45 : _GEN_9305; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9307 = 8'h2e == new_ptr_66_value ? ghv_46 : _GEN_9306; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9308 = 8'h2f == new_ptr_66_value ? ghv_47 : _GEN_9307; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9309 = 8'h30 == new_ptr_66_value ? ghv_48 : _GEN_9308; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9310 = 8'h31 == new_ptr_66_value ? ghv_49 : _GEN_9309; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9311 = 8'h32 == new_ptr_66_value ? ghv_50 : _GEN_9310; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9312 = 8'h33 == new_ptr_66_value ? ghv_51 : _GEN_9311; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9313 = 8'h34 == new_ptr_66_value ? ghv_52 : _GEN_9312; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9314 = 8'h35 == new_ptr_66_value ? ghv_53 : _GEN_9313; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9315 = 8'h36 == new_ptr_66_value ? ghv_54 : _GEN_9314; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9316 = 8'h37 == new_ptr_66_value ? ghv_55 : _GEN_9315; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9317 = 8'h38 == new_ptr_66_value ? ghv_56 : _GEN_9316; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9318 = 8'h39 == new_ptr_66_value ? ghv_57 : _GEN_9317; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9319 = 8'h3a == new_ptr_66_value ? ghv_58 : _GEN_9318; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9320 = 8'h3b == new_ptr_66_value ? ghv_59 : _GEN_9319; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9321 = 8'h3c == new_ptr_66_value ? ghv_60 : _GEN_9320; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9322 = 8'h3d == new_ptr_66_value ? ghv_61 : _GEN_9321; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9323 = 8'h3e == new_ptr_66_value ? ghv_62 : _GEN_9322; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9324 = 8'h3f == new_ptr_66_value ? ghv_63 : _GEN_9323; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9325 = 8'h40 == new_ptr_66_value ? ghv_64 : _GEN_9324; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9326 = 8'h41 == new_ptr_66_value ? ghv_65 : _GEN_9325; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9327 = 8'h42 == new_ptr_66_value ? ghv_66 : _GEN_9326; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9328 = 8'h43 == new_ptr_66_value ? ghv_67 : _GEN_9327; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9329 = 8'h44 == new_ptr_66_value ? ghv_68 : _GEN_9328; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9330 = 8'h45 == new_ptr_66_value ? ghv_69 : _GEN_9329; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9331 = 8'h46 == new_ptr_66_value ? ghv_70 : _GEN_9330; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9332 = 8'h47 == new_ptr_66_value ? ghv_71 : _GEN_9331; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9333 = 8'h48 == new_ptr_66_value ? ghv_72 : _GEN_9332; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9334 = 8'h49 == new_ptr_66_value ? ghv_73 : _GEN_9333; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9335 = 8'h4a == new_ptr_66_value ? ghv_74 : _GEN_9334; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9336 = 8'h4b == new_ptr_66_value ? ghv_75 : _GEN_9335; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9337 = 8'h4c == new_ptr_66_value ? ghv_76 : _GEN_9336; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9338 = 8'h4d == new_ptr_66_value ? ghv_77 : _GEN_9337; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9339 = 8'h4e == new_ptr_66_value ? ghv_78 : _GEN_9338; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9340 = 8'h4f == new_ptr_66_value ? ghv_79 : _GEN_9339; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9341 = 8'h50 == new_ptr_66_value ? ghv_80 : _GEN_9340; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9342 = 8'h51 == new_ptr_66_value ? ghv_81 : _GEN_9341; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9343 = 8'h52 == new_ptr_66_value ? ghv_82 : _GEN_9342; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9344 = 8'h53 == new_ptr_66_value ? ghv_83 : _GEN_9343; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9345 = 8'h54 == new_ptr_66_value ? ghv_84 : _GEN_9344; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9346 = 8'h55 == new_ptr_66_value ? ghv_85 : _GEN_9345; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9347 = 8'h56 == new_ptr_66_value ? ghv_86 : _GEN_9346; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9348 = 8'h57 == new_ptr_66_value ? ghv_87 : _GEN_9347; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9349 = 8'h58 == new_ptr_66_value ? ghv_88 : _GEN_9348; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9350 = 8'h59 == new_ptr_66_value ? ghv_89 : _GEN_9349; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9351 = 8'h5a == new_ptr_66_value ? ghv_90 : _GEN_9350; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9352 = 8'h5b == new_ptr_66_value ? ghv_91 : _GEN_9351; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9353 = 8'h5c == new_ptr_66_value ? ghv_92 : _GEN_9352; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9354 = 8'h5d == new_ptr_66_value ? ghv_93 : _GEN_9353; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9355 = 8'h5e == new_ptr_66_value ? ghv_94 : _GEN_9354; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9356 = 8'h5f == new_ptr_66_value ? ghv_95 : _GEN_9355; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9357 = 8'h60 == new_ptr_66_value ? ghv_96 : _GEN_9356; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9358 = 8'h61 == new_ptr_66_value ? ghv_97 : _GEN_9357; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9359 = 8'h62 == new_ptr_66_value ? ghv_98 : _GEN_9358; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9360 = 8'h63 == new_ptr_66_value ? ghv_99 : _GEN_9359; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9361 = 8'h64 == new_ptr_66_value ? ghv_100 : _GEN_9360; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9362 = 8'h65 == new_ptr_66_value ? ghv_101 : _GEN_9361; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9363 = 8'h66 == new_ptr_66_value ? ghv_102 : _GEN_9362; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9364 = 8'h67 == new_ptr_66_value ? ghv_103 : _GEN_9363; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9365 = 8'h68 == new_ptr_66_value ? ghv_104 : _GEN_9364; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9366 = 8'h69 == new_ptr_66_value ? ghv_105 : _GEN_9365; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9367 = 8'h6a == new_ptr_66_value ? ghv_106 : _GEN_9366; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9368 = 8'h6b == new_ptr_66_value ? ghv_107 : _GEN_9367; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9369 = 8'h6c == new_ptr_66_value ? ghv_108 : _GEN_9368; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9370 = 8'h6d == new_ptr_66_value ? ghv_109 : _GEN_9369; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9371 = 8'h6e == new_ptr_66_value ? ghv_110 : _GEN_9370; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9372 = 8'h6f == new_ptr_66_value ? ghv_111 : _GEN_9371; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9373 = 8'h70 == new_ptr_66_value ? ghv_112 : _GEN_9372; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9374 = 8'h71 == new_ptr_66_value ? ghv_113 : _GEN_9373; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9375 = 8'h72 == new_ptr_66_value ? ghv_114 : _GEN_9374; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9376 = 8'h73 == new_ptr_66_value ? ghv_115 : _GEN_9375; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9377 = 8'h74 == new_ptr_66_value ? ghv_116 : _GEN_9376; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9378 = 8'h75 == new_ptr_66_value ? ghv_117 : _GEN_9377; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9379 = 8'h76 == new_ptr_66_value ? ghv_118 : _GEN_9378; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9380 = 8'h77 == new_ptr_66_value ? ghv_119 : _GEN_9379; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9381 = 8'h78 == new_ptr_66_value ? ghv_120 : _GEN_9380; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9382 = 8'h79 == new_ptr_66_value ? ghv_121 : _GEN_9381; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9383 = 8'h7a == new_ptr_66_value ? ghv_122 : _GEN_9382; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9384 = 8'h7b == new_ptr_66_value ? ghv_123 : _GEN_9383; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9385 = 8'h7c == new_ptr_66_value ? ghv_124 : _GEN_9384; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9386 = 8'h7d == new_ptr_66_value ? ghv_125 : _GEN_9385; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9387 = 8'h7e == new_ptr_66_value ? ghv_126 : _GEN_9386; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9388 = 8'h7f == new_ptr_66_value ? ghv_127 : _GEN_9387; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9389 = 8'h80 == new_ptr_66_value ? ghv_128 : _GEN_9388; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9390 = 8'h81 == new_ptr_66_value ? ghv_129 : _GEN_9389; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9391 = 8'h82 == new_ptr_66_value ? ghv_130 : _GEN_9390; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9392 = 8'h83 == new_ptr_66_value ? ghv_131 : _GEN_9391; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9393 = 8'h84 == new_ptr_66_value ? ghv_132 : _GEN_9392; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9394 = 8'h85 == new_ptr_66_value ? ghv_133 : _GEN_9393; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9395 = 8'h86 == new_ptr_66_value ? ghv_134 : _GEN_9394; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9396 = 8'h87 == new_ptr_66_value ? ghv_135 : _GEN_9395; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9397 = 8'h88 == new_ptr_66_value ? ghv_136 : _GEN_9396; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9398 = 8'h89 == new_ptr_66_value ? ghv_137 : _GEN_9397; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9399 = 8'h8a == new_ptr_66_value ? ghv_138 : _GEN_9398; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9400 = 8'h8b == new_ptr_66_value ? ghv_139 : _GEN_9399; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9401 = 8'h8c == new_ptr_66_value ? ghv_140 : _GEN_9400; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9402 = 8'h8d == new_ptr_66_value ? ghv_141 : _GEN_9401; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9403 = 8'h8e == new_ptr_66_value ? ghv_142 : _GEN_9402; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_72_value = _new_ptr_value_T_145[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_9406 = 8'h1 == new_ptr_72_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9407 = 8'h2 == new_ptr_72_value ? ghv_2 : _GEN_9406; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9408 = 8'h3 == new_ptr_72_value ? ghv_3 : _GEN_9407; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9409 = 8'h4 == new_ptr_72_value ? ghv_4 : _GEN_9408; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9410 = 8'h5 == new_ptr_72_value ? ghv_5 : _GEN_9409; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9411 = 8'h6 == new_ptr_72_value ? ghv_6 : _GEN_9410; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9412 = 8'h7 == new_ptr_72_value ? ghv_7 : _GEN_9411; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9413 = 8'h8 == new_ptr_72_value ? ghv_8 : _GEN_9412; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9414 = 8'h9 == new_ptr_72_value ? ghv_9 : _GEN_9413; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9415 = 8'ha == new_ptr_72_value ? ghv_10 : _GEN_9414; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9416 = 8'hb == new_ptr_72_value ? ghv_11 : _GEN_9415; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9417 = 8'hc == new_ptr_72_value ? ghv_12 : _GEN_9416; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9418 = 8'hd == new_ptr_72_value ? ghv_13 : _GEN_9417; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9419 = 8'he == new_ptr_72_value ? ghv_14 : _GEN_9418; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9420 = 8'hf == new_ptr_72_value ? ghv_15 : _GEN_9419; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9421 = 8'h10 == new_ptr_72_value ? ghv_16 : _GEN_9420; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9422 = 8'h11 == new_ptr_72_value ? ghv_17 : _GEN_9421; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9423 = 8'h12 == new_ptr_72_value ? ghv_18 : _GEN_9422; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9424 = 8'h13 == new_ptr_72_value ? ghv_19 : _GEN_9423; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9425 = 8'h14 == new_ptr_72_value ? ghv_20 : _GEN_9424; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9426 = 8'h15 == new_ptr_72_value ? ghv_21 : _GEN_9425; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9427 = 8'h16 == new_ptr_72_value ? ghv_22 : _GEN_9426; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9428 = 8'h17 == new_ptr_72_value ? ghv_23 : _GEN_9427; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9429 = 8'h18 == new_ptr_72_value ? ghv_24 : _GEN_9428; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9430 = 8'h19 == new_ptr_72_value ? ghv_25 : _GEN_9429; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9431 = 8'h1a == new_ptr_72_value ? ghv_26 : _GEN_9430; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9432 = 8'h1b == new_ptr_72_value ? ghv_27 : _GEN_9431; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9433 = 8'h1c == new_ptr_72_value ? ghv_28 : _GEN_9432; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9434 = 8'h1d == new_ptr_72_value ? ghv_29 : _GEN_9433; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9435 = 8'h1e == new_ptr_72_value ? ghv_30 : _GEN_9434; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9436 = 8'h1f == new_ptr_72_value ? ghv_31 : _GEN_9435; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9437 = 8'h20 == new_ptr_72_value ? ghv_32 : _GEN_9436; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9438 = 8'h21 == new_ptr_72_value ? ghv_33 : _GEN_9437; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9439 = 8'h22 == new_ptr_72_value ? ghv_34 : _GEN_9438; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9440 = 8'h23 == new_ptr_72_value ? ghv_35 : _GEN_9439; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9441 = 8'h24 == new_ptr_72_value ? ghv_36 : _GEN_9440; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9442 = 8'h25 == new_ptr_72_value ? ghv_37 : _GEN_9441; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9443 = 8'h26 == new_ptr_72_value ? ghv_38 : _GEN_9442; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9444 = 8'h27 == new_ptr_72_value ? ghv_39 : _GEN_9443; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9445 = 8'h28 == new_ptr_72_value ? ghv_40 : _GEN_9444; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9446 = 8'h29 == new_ptr_72_value ? ghv_41 : _GEN_9445; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9447 = 8'h2a == new_ptr_72_value ? ghv_42 : _GEN_9446; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9448 = 8'h2b == new_ptr_72_value ? ghv_43 : _GEN_9447; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9449 = 8'h2c == new_ptr_72_value ? ghv_44 : _GEN_9448; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9450 = 8'h2d == new_ptr_72_value ? ghv_45 : _GEN_9449; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9451 = 8'h2e == new_ptr_72_value ? ghv_46 : _GEN_9450; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9452 = 8'h2f == new_ptr_72_value ? ghv_47 : _GEN_9451; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9453 = 8'h30 == new_ptr_72_value ? ghv_48 : _GEN_9452; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9454 = 8'h31 == new_ptr_72_value ? ghv_49 : _GEN_9453; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9455 = 8'h32 == new_ptr_72_value ? ghv_50 : _GEN_9454; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9456 = 8'h33 == new_ptr_72_value ? ghv_51 : _GEN_9455; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9457 = 8'h34 == new_ptr_72_value ? ghv_52 : _GEN_9456; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9458 = 8'h35 == new_ptr_72_value ? ghv_53 : _GEN_9457; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9459 = 8'h36 == new_ptr_72_value ? ghv_54 : _GEN_9458; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9460 = 8'h37 == new_ptr_72_value ? ghv_55 : _GEN_9459; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9461 = 8'h38 == new_ptr_72_value ? ghv_56 : _GEN_9460; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9462 = 8'h39 == new_ptr_72_value ? ghv_57 : _GEN_9461; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9463 = 8'h3a == new_ptr_72_value ? ghv_58 : _GEN_9462; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9464 = 8'h3b == new_ptr_72_value ? ghv_59 : _GEN_9463; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9465 = 8'h3c == new_ptr_72_value ? ghv_60 : _GEN_9464; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9466 = 8'h3d == new_ptr_72_value ? ghv_61 : _GEN_9465; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9467 = 8'h3e == new_ptr_72_value ? ghv_62 : _GEN_9466; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9468 = 8'h3f == new_ptr_72_value ? ghv_63 : _GEN_9467; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9469 = 8'h40 == new_ptr_72_value ? ghv_64 : _GEN_9468; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9470 = 8'h41 == new_ptr_72_value ? ghv_65 : _GEN_9469; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9471 = 8'h42 == new_ptr_72_value ? ghv_66 : _GEN_9470; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9472 = 8'h43 == new_ptr_72_value ? ghv_67 : _GEN_9471; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9473 = 8'h44 == new_ptr_72_value ? ghv_68 : _GEN_9472; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9474 = 8'h45 == new_ptr_72_value ? ghv_69 : _GEN_9473; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9475 = 8'h46 == new_ptr_72_value ? ghv_70 : _GEN_9474; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9476 = 8'h47 == new_ptr_72_value ? ghv_71 : _GEN_9475; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9477 = 8'h48 == new_ptr_72_value ? ghv_72 : _GEN_9476; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9478 = 8'h49 == new_ptr_72_value ? ghv_73 : _GEN_9477; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9479 = 8'h4a == new_ptr_72_value ? ghv_74 : _GEN_9478; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9480 = 8'h4b == new_ptr_72_value ? ghv_75 : _GEN_9479; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9481 = 8'h4c == new_ptr_72_value ? ghv_76 : _GEN_9480; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9482 = 8'h4d == new_ptr_72_value ? ghv_77 : _GEN_9481; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9483 = 8'h4e == new_ptr_72_value ? ghv_78 : _GEN_9482; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9484 = 8'h4f == new_ptr_72_value ? ghv_79 : _GEN_9483; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9485 = 8'h50 == new_ptr_72_value ? ghv_80 : _GEN_9484; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9486 = 8'h51 == new_ptr_72_value ? ghv_81 : _GEN_9485; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9487 = 8'h52 == new_ptr_72_value ? ghv_82 : _GEN_9486; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9488 = 8'h53 == new_ptr_72_value ? ghv_83 : _GEN_9487; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9489 = 8'h54 == new_ptr_72_value ? ghv_84 : _GEN_9488; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9490 = 8'h55 == new_ptr_72_value ? ghv_85 : _GEN_9489; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9491 = 8'h56 == new_ptr_72_value ? ghv_86 : _GEN_9490; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9492 = 8'h57 == new_ptr_72_value ? ghv_87 : _GEN_9491; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9493 = 8'h58 == new_ptr_72_value ? ghv_88 : _GEN_9492; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9494 = 8'h59 == new_ptr_72_value ? ghv_89 : _GEN_9493; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9495 = 8'h5a == new_ptr_72_value ? ghv_90 : _GEN_9494; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9496 = 8'h5b == new_ptr_72_value ? ghv_91 : _GEN_9495; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9497 = 8'h5c == new_ptr_72_value ? ghv_92 : _GEN_9496; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9498 = 8'h5d == new_ptr_72_value ? ghv_93 : _GEN_9497; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9499 = 8'h5e == new_ptr_72_value ? ghv_94 : _GEN_9498; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9500 = 8'h5f == new_ptr_72_value ? ghv_95 : _GEN_9499; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9501 = 8'h60 == new_ptr_72_value ? ghv_96 : _GEN_9500; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9502 = 8'h61 == new_ptr_72_value ? ghv_97 : _GEN_9501; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9503 = 8'h62 == new_ptr_72_value ? ghv_98 : _GEN_9502; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9504 = 8'h63 == new_ptr_72_value ? ghv_99 : _GEN_9503; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9505 = 8'h64 == new_ptr_72_value ? ghv_100 : _GEN_9504; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9506 = 8'h65 == new_ptr_72_value ? ghv_101 : _GEN_9505; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9507 = 8'h66 == new_ptr_72_value ? ghv_102 : _GEN_9506; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9508 = 8'h67 == new_ptr_72_value ? ghv_103 : _GEN_9507; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9509 = 8'h68 == new_ptr_72_value ? ghv_104 : _GEN_9508; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9510 = 8'h69 == new_ptr_72_value ? ghv_105 : _GEN_9509; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9511 = 8'h6a == new_ptr_72_value ? ghv_106 : _GEN_9510; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9512 = 8'h6b == new_ptr_72_value ? ghv_107 : _GEN_9511; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9513 = 8'h6c == new_ptr_72_value ? ghv_108 : _GEN_9512; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9514 = 8'h6d == new_ptr_72_value ? ghv_109 : _GEN_9513; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9515 = 8'h6e == new_ptr_72_value ? ghv_110 : _GEN_9514; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9516 = 8'h6f == new_ptr_72_value ? ghv_111 : _GEN_9515; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9517 = 8'h70 == new_ptr_72_value ? ghv_112 : _GEN_9516; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9518 = 8'h71 == new_ptr_72_value ? ghv_113 : _GEN_9517; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9519 = 8'h72 == new_ptr_72_value ? ghv_114 : _GEN_9518; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9520 = 8'h73 == new_ptr_72_value ? ghv_115 : _GEN_9519; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9521 = 8'h74 == new_ptr_72_value ? ghv_116 : _GEN_9520; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9522 = 8'h75 == new_ptr_72_value ? ghv_117 : _GEN_9521; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9523 = 8'h76 == new_ptr_72_value ? ghv_118 : _GEN_9522; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9524 = 8'h77 == new_ptr_72_value ? ghv_119 : _GEN_9523; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9525 = 8'h78 == new_ptr_72_value ? ghv_120 : _GEN_9524; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9526 = 8'h79 == new_ptr_72_value ? ghv_121 : _GEN_9525; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9527 = 8'h7a == new_ptr_72_value ? ghv_122 : _GEN_9526; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9528 = 8'h7b == new_ptr_72_value ? ghv_123 : _GEN_9527; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9529 = 8'h7c == new_ptr_72_value ? ghv_124 : _GEN_9528; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9530 = 8'h7d == new_ptr_72_value ? ghv_125 : _GEN_9529; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9531 = 8'h7e == new_ptr_72_value ? ghv_126 : _GEN_9530; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9532 = 8'h7f == new_ptr_72_value ? ghv_127 : _GEN_9531; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9533 = 8'h80 == new_ptr_72_value ? ghv_128 : _GEN_9532; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9534 = 8'h81 == new_ptr_72_value ? ghv_129 : _GEN_9533; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9535 = 8'h82 == new_ptr_72_value ? ghv_130 : _GEN_9534; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9536 = 8'h83 == new_ptr_72_value ? ghv_131 : _GEN_9535; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9537 = 8'h84 == new_ptr_72_value ? ghv_132 : _GEN_9536; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9538 = 8'h85 == new_ptr_72_value ? ghv_133 : _GEN_9537; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9539 = 8'h86 == new_ptr_72_value ? ghv_134 : _GEN_9538; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9540 = 8'h87 == new_ptr_72_value ? ghv_135 : _GEN_9539; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9541 = 8'h88 == new_ptr_72_value ? ghv_136 : _GEN_9540; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9542 = 8'h89 == new_ptr_72_value ? ghv_137 : _GEN_9541; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9543 = 8'h8a == new_ptr_72_value ? ghv_138 : _GEN_9542; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9544 = 8'h8b == new_ptr_72_value ? ghv_139 : _GEN_9543; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9545 = 8'h8c == new_ptr_72_value ? ghv_140 : _GEN_9544; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9546 = 8'h8d == new_ptr_72_value ? ghv_141 : _GEN_9545; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9547 = 8'h8e == new_ptr_72_value ? ghv_142 : _GEN_9546; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_75_value = _new_ptr_value_T_151[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_9550 = 8'h1 == new_ptr_75_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9551 = 8'h2 == new_ptr_75_value ? ghv_2 : _GEN_9550; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9552 = 8'h3 == new_ptr_75_value ? ghv_3 : _GEN_9551; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9553 = 8'h4 == new_ptr_75_value ? ghv_4 : _GEN_9552; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9554 = 8'h5 == new_ptr_75_value ? ghv_5 : _GEN_9553; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9555 = 8'h6 == new_ptr_75_value ? ghv_6 : _GEN_9554; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9556 = 8'h7 == new_ptr_75_value ? ghv_7 : _GEN_9555; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9557 = 8'h8 == new_ptr_75_value ? ghv_8 : _GEN_9556; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9558 = 8'h9 == new_ptr_75_value ? ghv_9 : _GEN_9557; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9559 = 8'ha == new_ptr_75_value ? ghv_10 : _GEN_9558; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9560 = 8'hb == new_ptr_75_value ? ghv_11 : _GEN_9559; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9561 = 8'hc == new_ptr_75_value ? ghv_12 : _GEN_9560; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9562 = 8'hd == new_ptr_75_value ? ghv_13 : _GEN_9561; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9563 = 8'he == new_ptr_75_value ? ghv_14 : _GEN_9562; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9564 = 8'hf == new_ptr_75_value ? ghv_15 : _GEN_9563; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9565 = 8'h10 == new_ptr_75_value ? ghv_16 : _GEN_9564; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9566 = 8'h11 == new_ptr_75_value ? ghv_17 : _GEN_9565; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9567 = 8'h12 == new_ptr_75_value ? ghv_18 : _GEN_9566; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9568 = 8'h13 == new_ptr_75_value ? ghv_19 : _GEN_9567; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9569 = 8'h14 == new_ptr_75_value ? ghv_20 : _GEN_9568; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9570 = 8'h15 == new_ptr_75_value ? ghv_21 : _GEN_9569; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9571 = 8'h16 == new_ptr_75_value ? ghv_22 : _GEN_9570; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9572 = 8'h17 == new_ptr_75_value ? ghv_23 : _GEN_9571; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9573 = 8'h18 == new_ptr_75_value ? ghv_24 : _GEN_9572; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9574 = 8'h19 == new_ptr_75_value ? ghv_25 : _GEN_9573; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9575 = 8'h1a == new_ptr_75_value ? ghv_26 : _GEN_9574; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9576 = 8'h1b == new_ptr_75_value ? ghv_27 : _GEN_9575; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9577 = 8'h1c == new_ptr_75_value ? ghv_28 : _GEN_9576; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9578 = 8'h1d == new_ptr_75_value ? ghv_29 : _GEN_9577; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9579 = 8'h1e == new_ptr_75_value ? ghv_30 : _GEN_9578; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9580 = 8'h1f == new_ptr_75_value ? ghv_31 : _GEN_9579; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9581 = 8'h20 == new_ptr_75_value ? ghv_32 : _GEN_9580; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9582 = 8'h21 == new_ptr_75_value ? ghv_33 : _GEN_9581; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9583 = 8'h22 == new_ptr_75_value ? ghv_34 : _GEN_9582; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9584 = 8'h23 == new_ptr_75_value ? ghv_35 : _GEN_9583; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9585 = 8'h24 == new_ptr_75_value ? ghv_36 : _GEN_9584; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9586 = 8'h25 == new_ptr_75_value ? ghv_37 : _GEN_9585; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9587 = 8'h26 == new_ptr_75_value ? ghv_38 : _GEN_9586; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9588 = 8'h27 == new_ptr_75_value ? ghv_39 : _GEN_9587; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9589 = 8'h28 == new_ptr_75_value ? ghv_40 : _GEN_9588; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9590 = 8'h29 == new_ptr_75_value ? ghv_41 : _GEN_9589; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9591 = 8'h2a == new_ptr_75_value ? ghv_42 : _GEN_9590; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9592 = 8'h2b == new_ptr_75_value ? ghv_43 : _GEN_9591; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9593 = 8'h2c == new_ptr_75_value ? ghv_44 : _GEN_9592; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9594 = 8'h2d == new_ptr_75_value ? ghv_45 : _GEN_9593; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9595 = 8'h2e == new_ptr_75_value ? ghv_46 : _GEN_9594; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9596 = 8'h2f == new_ptr_75_value ? ghv_47 : _GEN_9595; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9597 = 8'h30 == new_ptr_75_value ? ghv_48 : _GEN_9596; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9598 = 8'h31 == new_ptr_75_value ? ghv_49 : _GEN_9597; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9599 = 8'h32 == new_ptr_75_value ? ghv_50 : _GEN_9598; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9600 = 8'h33 == new_ptr_75_value ? ghv_51 : _GEN_9599; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9601 = 8'h34 == new_ptr_75_value ? ghv_52 : _GEN_9600; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9602 = 8'h35 == new_ptr_75_value ? ghv_53 : _GEN_9601; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9603 = 8'h36 == new_ptr_75_value ? ghv_54 : _GEN_9602; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9604 = 8'h37 == new_ptr_75_value ? ghv_55 : _GEN_9603; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9605 = 8'h38 == new_ptr_75_value ? ghv_56 : _GEN_9604; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9606 = 8'h39 == new_ptr_75_value ? ghv_57 : _GEN_9605; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9607 = 8'h3a == new_ptr_75_value ? ghv_58 : _GEN_9606; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9608 = 8'h3b == new_ptr_75_value ? ghv_59 : _GEN_9607; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9609 = 8'h3c == new_ptr_75_value ? ghv_60 : _GEN_9608; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9610 = 8'h3d == new_ptr_75_value ? ghv_61 : _GEN_9609; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9611 = 8'h3e == new_ptr_75_value ? ghv_62 : _GEN_9610; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9612 = 8'h3f == new_ptr_75_value ? ghv_63 : _GEN_9611; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9613 = 8'h40 == new_ptr_75_value ? ghv_64 : _GEN_9612; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9614 = 8'h41 == new_ptr_75_value ? ghv_65 : _GEN_9613; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9615 = 8'h42 == new_ptr_75_value ? ghv_66 : _GEN_9614; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9616 = 8'h43 == new_ptr_75_value ? ghv_67 : _GEN_9615; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9617 = 8'h44 == new_ptr_75_value ? ghv_68 : _GEN_9616; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9618 = 8'h45 == new_ptr_75_value ? ghv_69 : _GEN_9617; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9619 = 8'h46 == new_ptr_75_value ? ghv_70 : _GEN_9618; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9620 = 8'h47 == new_ptr_75_value ? ghv_71 : _GEN_9619; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9621 = 8'h48 == new_ptr_75_value ? ghv_72 : _GEN_9620; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9622 = 8'h49 == new_ptr_75_value ? ghv_73 : _GEN_9621; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9623 = 8'h4a == new_ptr_75_value ? ghv_74 : _GEN_9622; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9624 = 8'h4b == new_ptr_75_value ? ghv_75 : _GEN_9623; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9625 = 8'h4c == new_ptr_75_value ? ghv_76 : _GEN_9624; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9626 = 8'h4d == new_ptr_75_value ? ghv_77 : _GEN_9625; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9627 = 8'h4e == new_ptr_75_value ? ghv_78 : _GEN_9626; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9628 = 8'h4f == new_ptr_75_value ? ghv_79 : _GEN_9627; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9629 = 8'h50 == new_ptr_75_value ? ghv_80 : _GEN_9628; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9630 = 8'h51 == new_ptr_75_value ? ghv_81 : _GEN_9629; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9631 = 8'h52 == new_ptr_75_value ? ghv_82 : _GEN_9630; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9632 = 8'h53 == new_ptr_75_value ? ghv_83 : _GEN_9631; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9633 = 8'h54 == new_ptr_75_value ? ghv_84 : _GEN_9632; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9634 = 8'h55 == new_ptr_75_value ? ghv_85 : _GEN_9633; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9635 = 8'h56 == new_ptr_75_value ? ghv_86 : _GEN_9634; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9636 = 8'h57 == new_ptr_75_value ? ghv_87 : _GEN_9635; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9637 = 8'h58 == new_ptr_75_value ? ghv_88 : _GEN_9636; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9638 = 8'h59 == new_ptr_75_value ? ghv_89 : _GEN_9637; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9639 = 8'h5a == new_ptr_75_value ? ghv_90 : _GEN_9638; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9640 = 8'h5b == new_ptr_75_value ? ghv_91 : _GEN_9639; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9641 = 8'h5c == new_ptr_75_value ? ghv_92 : _GEN_9640; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9642 = 8'h5d == new_ptr_75_value ? ghv_93 : _GEN_9641; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9643 = 8'h5e == new_ptr_75_value ? ghv_94 : _GEN_9642; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9644 = 8'h5f == new_ptr_75_value ? ghv_95 : _GEN_9643; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9645 = 8'h60 == new_ptr_75_value ? ghv_96 : _GEN_9644; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9646 = 8'h61 == new_ptr_75_value ? ghv_97 : _GEN_9645; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9647 = 8'h62 == new_ptr_75_value ? ghv_98 : _GEN_9646; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9648 = 8'h63 == new_ptr_75_value ? ghv_99 : _GEN_9647; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9649 = 8'h64 == new_ptr_75_value ? ghv_100 : _GEN_9648; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9650 = 8'h65 == new_ptr_75_value ? ghv_101 : _GEN_9649; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9651 = 8'h66 == new_ptr_75_value ? ghv_102 : _GEN_9650; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9652 = 8'h67 == new_ptr_75_value ? ghv_103 : _GEN_9651; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9653 = 8'h68 == new_ptr_75_value ? ghv_104 : _GEN_9652; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9654 = 8'h69 == new_ptr_75_value ? ghv_105 : _GEN_9653; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9655 = 8'h6a == new_ptr_75_value ? ghv_106 : _GEN_9654; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9656 = 8'h6b == new_ptr_75_value ? ghv_107 : _GEN_9655; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9657 = 8'h6c == new_ptr_75_value ? ghv_108 : _GEN_9656; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9658 = 8'h6d == new_ptr_75_value ? ghv_109 : _GEN_9657; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9659 = 8'h6e == new_ptr_75_value ? ghv_110 : _GEN_9658; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9660 = 8'h6f == new_ptr_75_value ? ghv_111 : _GEN_9659; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9661 = 8'h70 == new_ptr_75_value ? ghv_112 : _GEN_9660; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9662 = 8'h71 == new_ptr_75_value ? ghv_113 : _GEN_9661; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9663 = 8'h72 == new_ptr_75_value ? ghv_114 : _GEN_9662; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9664 = 8'h73 == new_ptr_75_value ? ghv_115 : _GEN_9663; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9665 = 8'h74 == new_ptr_75_value ? ghv_116 : _GEN_9664; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9666 = 8'h75 == new_ptr_75_value ? ghv_117 : _GEN_9665; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9667 = 8'h76 == new_ptr_75_value ? ghv_118 : _GEN_9666; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9668 = 8'h77 == new_ptr_75_value ? ghv_119 : _GEN_9667; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9669 = 8'h78 == new_ptr_75_value ? ghv_120 : _GEN_9668; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9670 = 8'h79 == new_ptr_75_value ? ghv_121 : _GEN_9669; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9671 = 8'h7a == new_ptr_75_value ? ghv_122 : _GEN_9670; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9672 = 8'h7b == new_ptr_75_value ? ghv_123 : _GEN_9671; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9673 = 8'h7c == new_ptr_75_value ? ghv_124 : _GEN_9672; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9674 = 8'h7d == new_ptr_75_value ? ghv_125 : _GEN_9673; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9675 = 8'h7e == new_ptr_75_value ? ghv_126 : _GEN_9674; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9676 = 8'h7f == new_ptr_75_value ? ghv_127 : _GEN_9675; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9677 = 8'h80 == new_ptr_75_value ? ghv_128 : _GEN_9676; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9678 = 8'h81 == new_ptr_75_value ? ghv_129 : _GEN_9677; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9679 = 8'h82 == new_ptr_75_value ? ghv_130 : _GEN_9678; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9680 = 8'h83 == new_ptr_75_value ? ghv_131 : _GEN_9679; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9681 = 8'h84 == new_ptr_75_value ? ghv_132 : _GEN_9680; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9682 = 8'h85 == new_ptr_75_value ? ghv_133 : _GEN_9681; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9683 = 8'h86 == new_ptr_75_value ? ghv_134 : _GEN_9682; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9684 = 8'h87 == new_ptr_75_value ? ghv_135 : _GEN_9683; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9685 = 8'h88 == new_ptr_75_value ? ghv_136 : _GEN_9684; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9686 = 8'h89 == new_ptr_75_value ? ghv_137 : _GEN_9685; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9687 = 8'h8a == new_ptr_75_value ? ghv_138 : _GEN_9686; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9688 = 8'h8b == new_ptr_75_value ? ghv_139 : _GEN_9687; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9689 = 8'h8c == new_ptr_75_value ? ghv_140 : _GEN_9688; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9690 = 8'h8d == new_ptr_75_value ? ghv_141 : _GEN_9689; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9691 = 8'h8e == new_ptr_75_value ? ghv_142 : _GEN_9690; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_62_value = _new_ptr_value_T_125[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_9694 = 8'h1 == new_ptr_62_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9695 = 8'h2 == new_ptr_62_value ? ghv_2 : _GEN_9694; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9696 = 8'h3 == new_ptr_62_value ? ghv_3 : _GEN_9695; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9697 = 8'h4 == new_ptr_62_value ? ghv_4 : _GEN_9696; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9698 = 8'h5 == new_ptr_62_value ? ghv_5 : _GEN_9697; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9699 = 8'h6 == new_ptr_62_value ? ghv_6 : _GEN_9698; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9700 = 8'h7 == new_ptr_62_value ? ghv_7 : _GEN_9699; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9701 = 8'h8 == new_ptr_62_value ? ghv_8 : _GEN_9700; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9702 = 8'h9 == new_ptr_62_value ? ghv_9 : _GEN_9701; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9703 = 8'ha == new_ptr_62_value ? ghv_10 : _GEN_9702; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9704 = 8'hb == new_ptr_62_value ? ghv_11 : _GEN_9703; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9705 = 8'hc == new_ptr_62_value ? ghv_12 : _GEN_9704; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9706 = 8'hd == new_ptr_62_value ? ghv_13 : _GEN_9705; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9707 = 8'he == new_ptr_62_value ? ghv_14 : _GEN_9706; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9708 = 8'hf == new_ptr_62_value ? ghv_15 : _GEN_9707; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9709 = 8'h10 == new_ptr_62_value ? ghv_16 : _GEN_9708; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9710 = 8'h11 == new_ptr_62_value ? ghv_17 : _GEN_9709; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9711 = 8'h12 == new_ptr_62_value ? ghv_18 : _GEN_9710; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9712 = 8'h13 == new_ptr_62_value ? ghv_19 : _GEN_9711; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9713 = 8'h14 == new_ptr_62_value ? ghv_20 : _GEN_9712; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9714 = 8'h15 == new_ptr_62_value ? ghv_21 : _GEN_9713; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9715 = 8'h16 == new_ptr_62_value ? ghv_22 : _GEN_9714; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9716 = 8'h17 == new_ptr_62_value ? ghv_23 : _GEN_9715; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9717 = 8'h18 == new_ptr_62_value ? ghv_24 : _GEN_9716; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9718 = 8'h19 == new_ptr_62_value ? ghv_25 : _GEN_9717; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9719 = 8'h1a == new_ptr_62_value ? ghv_26 : _GEN_9718; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9720 = 8'h1b == new_ptr_62_value ? ghv_27 : _GEN_9719; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9721 = 8'h1c == new_ptr_62_value ? ghv_28 : _GEN_9720; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9722 = 8'h1d == new_ptr_62_value ? ghv_29 : _GEN_9721; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9723 = 8'h1e == new_ptr_62_value ? ghv_30 : _GEN_9722; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9724 = 8'h1f == new_ptr_62_value ? ghv_31 : _GEN_9723; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9725 = 8'h20 == new_ptr_62_value ? ghv_32 : _GEN_9724; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9726 = 8'h21 == new_ptr_62_value ? ghv_33 : _GEN_9725; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9727 = 8'h22 == new_ptr_62_value ? ghv_34 : _GEN_9726; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9728 = 8'h23 == new_ptr_62_value ? ghv_35 : _GEN_9727; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9729 = 8'h24 == new_ptr_62_value ? ghv_36 : _GEN_9728; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9730 = 8'h25 == new_ptr_62_value ? ghv_37 : _GEN_9729; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9731 = 8'h26 == new_ptr_62_value ? ghv_38 : _GEN_9730; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9732 = 8'h27 == new_ptr_62_value ? ghv_39 : _GEN_9731; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9733 = 8'h28 == new_ptr_62_value ? ghv_40 : _GEN_9732; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9734 = 8'h29 == new_ptr_62_value ? ghv_41 : _GEN_9733; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9735 = 8'h2a == new_ptr_62_value ? ghv_42 : _GEN_9734; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9736 = 8'h2b == new_ptr_62_value ? ghv_43 : _GEN_9735; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9737 = 8'h2c == new_ptr_62_value ? ghv_44 : _GEN_9736; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9738 = 8'h2d == new_ptr_62_value ? ghv_45 : _GEN_9737; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9739 = 8'h2e == new_ptr_62_value ? ghv_46 : _GEN_9738; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9740 = 8'h2f == new_ptr_62_value ? ghv_47 : _GEN_9739; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9741 = 8'h30 == new_ptr_62_value ? ghv_48 : _GEN_9740; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9742 = 8'h31 == new_ptr_62_value ? ghv_49 : _GEN_9741; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9743 = 8'h32 == new_ptr_62_value ? ghv_50 : _GEN_9742; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9744 = 8'h33 == new_ptr_62_value ? ghv_51 : _GEN_9743; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9745 = 8'h34 == new_ptr_62_value ? ghv_52 : _GEN_9744; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9746 = 8'h35 == new_ptr_62_value ? ghv_53 : _GEN_9745; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9747 = 8'h36 == new_ptr_62_value ? ghv_54 : _GEN_9746; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9748 = 8'h37 == new_ptr_62_value ? ghv_55 : _GEN_9747; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9749 = 8'h38 == new_ptr_62_value ? ghv_56 : _GEN_9748; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9750 = 8'h39 == new_ptr_62_value ? ghv_57 : _GEN_9749; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9751 = 8'h3a == new_ptr_62_value ? ghv_58 : _GEN_9750; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9752 = 8'h3b == new_ptr_62_value ? ghv_59 : _GEN_9751; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9753 = 8'h3c == new_ptr_62_value ? ghv_60 : _GEN_9752; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9754 = 8'h3d == new_ptr_62_value ? ghv_61 : _GEN_9753; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9755 = 8'h3e == new_ptr_62_value ? ghv_62 : _GEN_9754; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9756 = 8'h3f == new_ptr_62_value ? ghv_63 : _GEN_9755; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9757 = 8'h40 == new_ptr_62_value ? ghv_64 : _GEN_9756; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9758 = 8'h41 == new_ptr_62_value ? ghv_65 : _GEN_9757; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9759 = 8'h42 == new_ptr_62_value ? ghv_66 : _GEN_9758; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9760 = 8'h43 == new_ptr_62_value ? ghv_67 : _GEN_9759; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9761 = 8'h44 == new_ptr_62_value ? ghv_68 : _GEN_9760; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9762 = 8'h45 == new_ptr_62_value ? ghv_69 : _GEN_9761; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9763 = 8'h46 == new_ptr_62_value ? ghv_70 : _GEN_9762; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9764 = 8'h47 == new_ptr_62_value ? ghv_71 : _GEN_9763; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9765 = 8'h48 == new_ptr_62_value ? ghv_72 : _GEN_9764; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9766 = 8'h49 == new_ptr_62_value ? ghv_73 : _GEN_9765; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9767 = 8'h4a == new_ptr_62_value ? ghv_74 : _GEN_9766; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9768 = 8'h4b == new_ptr_62_value ? ghv_75 : _GEN_9767; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9769 = 8'h4c == new_ptr_62_value ? ghv_76 : _GEN_9768; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9770 = 8'h4d == new_ptr_62_value ? ghv_77 : _GEN_9769; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9771 = 8'h4e == new_ptr_62_value ? ghv_78 : _GEN_9770; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9772 = 8'h4f == new_ptr_62_value ? ghv_79 : _GEN_9771; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9773 = 8'h50 == new_ptr_62_value ? ghv_80 : _GEN_9772; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9774 = 8'h51 == new_ptr_62_value ? ghv_81 : _GEN_9773; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9775 = 8'h52 == new_ptr_62_value ? ghv_82 : _GEN_9774; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9776 = 8'h53 == new_ptr_62_value ? ghv_83 : _GEN_9775; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9777 = 8'h54 == new_ptr_62_value ? ghv_84 : _GEN_9776; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9778 = 8'h55 == new_ptr_62_value ? ghv_85 : _GEN_9777; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9779 = 8'h56 == new_ptr_62_value ? ghv_86 : _GEN_9778; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9780 = 8'h57 == new_ptr_62_value ? ghv_87 : _GEN_9779; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9781 = 8'h58 == new_ptr_62_value ? ghv_88 : _GEN_9780; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9782 = 8'h59 == new_ptr_62_value ? ghv_89 : _GEN_9781; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9783 = 8'h5a == new_ptr_62_value ? ghv_90 : _GEN_9782; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9784 = 8'h5b == new_ptr_62_value ? ghv_91 : _GEN_9783; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9785 = 8'h5c == new_ptr_62_value ? ghv_92 : _GEN_9784; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9786 = 8'h5d == new_ptr_62_value ? ghv_93 : _GEN_9785; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9787 = 8'h5e == new_ptr_62_value ? ghv_94 : _GEN_9786; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9788 = 8'h5f == new_ptr_62_value ? ghv_95 : _GEN_9787; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9789 = 8'h60 == new_ptr_62_value ? ghv_96 : _GEN_9788; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9790 = 8'h61 == new_ptr_62_value ? ghv_97 : _GEN_9789; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9791 = 8'h62 == new_ptr_62_value ? ghv_98 : _GEN_9790; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9792 = 8'h63 == new_ptr_62_value ? ghv_99 : _GEN_9791; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9793 = 8'h64 == new_ptr_62_value ? ghv_100 : _GEN_9792; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9794 = 8'h65 == new_ptr_62_value ? ghv_101 : _GEN_9793; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9795 = 8'h66 == new_ptr_62_value ? ghv_102 : _GEN_9794; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9796 = 8'h67 == new_ptr_62_value ? ghv_103 : _GEN_9795; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9797 = 8'h68 == new_ptr_62_value ? ghv_104 : _GEN_9796; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9798 = 8'h69 == new_ptr_62_value ? ghv_105 : _GEN_9797; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9799 = 8'h6a == new_ptr_62_value ? ghv_106 : _GEN_9798; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9800 = 8'h6b == new_ptr_62_value ? ghv_107 : _GEN_9799; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9801 = 8'h6c == new_ptr_62_value ? ghv_108 : _GEN_9800; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9802 = 8'h6d == new_ptr_62_value ? ghv_109 : _GEN_9801; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9803 = 8'h6e == new_ptr_62_value ? ghv_110 : _GEN_9802; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9804 = 8'h6f == new_ptr_62_value ? ghv_111 : _GEN_9803; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9805 = 8'h70 == new_ptr_62_value ? ghv_112 : _GEN_9804; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9806 = 8'h71 == new_ptr_62_value ? ghv_113 : _GEN_9805; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9807 = 8'h72 == new_ptr_62_value ? ghv_114 : _GEN_9806; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9808 = 8'h73 == new_ptr_62_value ? ghv_115 : _GEN_9807; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9809 = 8'h74 == new_ptr_62_value ? ghv_116 : _GEN_9808; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9810 = 8'h75 == new_ptr_62_value ? ghv_117 : _GEN_9809; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9811 = 8'h76 == new_ptr_62_value ? ghv_118 : _GEN_9810; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9812 = 8'h77 == new_ptr_62_value ? ghv_119 : _GEN_9811; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9813 = 8'h78 == new_ptr_62_value ? ghv_120 : _GEN_9812; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9814 = 8'h79 == new_ptr_62_value ? ghv_121 : _GEN_9813; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9815 = 8'h7a == new_ptr_62_value ? ghv_122 : _GEN_9814; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9816 = 8'h7b == new_ptr_62_value ? ghv_123 : _GEN_9815; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9817 = 8'h7c == new_ptr_62_value ? ghv_124 : _GEN_9816; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9818 = 8'h7d == new_ptr_62_value ? ghv_125 : _GEN_9817; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9819 = 8'h7e == new_ptr_62_value ? ghv_126 : _GEN_9818; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9820 = 8'h7f == new_ptr_62_value ? ghv_127 : _GEN_9819; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9821 = 8'h80 == new_ptr_62_value ? ghv_128 : _GEN_9820; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9822 = 8'h81 == new_ptr_62_value ? ghv_129 : _GEN_9821; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9823 = 8'h82 == new_ptr_62_value ? ghv_130 : _GEN_9822; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9824 = 8'h83 == new_ptr_62_value ? ghv_131 : _GEN_9823; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9825 = 8'h84 == new_ptr_62_value ? ghv_132 : _GEN_9824; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9826 = 8'h85 == new_ptr_62_value ? ghv_133 : _GEN_9825; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9827 = 8'h86 == new_ptr_62_value ? ghv_134 : _GEN_9826; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9828 = 8'h87 == new_ptr_62_value ? ghv_135 : _GEN_9827; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9829 = 8'h88 == new_ptr_62_value ? ghv_136 : _GEN_9828; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9830 = 8'h89 == new_ptr_62_value ? ghv_137 : _GEN_9829; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9831 = 8'h8a == new_ptr_62_value ? ghv_138 : _GEN_9830; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9832 = 8'h8b == new_ptr_62_value ? ghv_139 : _GEN_9831; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9833 = 8'h8c == new_ptr_62_value ? ghv_140 : _GEN_9832; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9834 = 8'h8d == new_ptr_62_value ? ghv_141 : _GEN_9833; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9835 = 8'h8e == new_ptr_62_value ? ghv_142 : _GEN_9834; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_74_value = _new_ptr_value_T_149[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_9838 = 8'h1 == new_ptr_74_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9839 = 8'h2 == new_ptr_74_value ? ghv_2 : _GEN_9838; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9840 = 8'h3 == new_ptr_74_value ? ghv_3 : _GEN_9839; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9841 = 8'h4 == new_ptr_74_value ? ghv_4 : _GEN_9840; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9842 = 8'h5 == new_ptr_74_value ? ghv_5 : _GEN_9841; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9843 = 8'h6 == new_ptr_74_value ? ghv_6 : _GEN_9842; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9844 = 8'h7 == new_ptr_74_value ? ghv_7 : _GEN_9843; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9845 = 8'h8 == new_ptr_74_value ? ghv_8 : _GEN_9844; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9846 = 8'h9 == new_ptr_74_value ? ghv_9 : _GEN_9845; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9847 = 8'ha == new_ptr_74_value ? ghv_10 : _GEN_9846; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9848 = 8'hb == new_ptr_74_value ? ghv_11 : _GEN_9847; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9849 = 8'hc == new_ptr_74_value ? ghv_12 : _GEN_9848; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9850 = 8'hd == new_ptr_74_value ? ghv_13 : _GEN_9849; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9851 = 8'he == new_ptr_74_value ? ghv_14 : _GEN_9850; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9852 = 8'hf == new_ptr_74_value ? ghv_15 : _GEN_9851; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9853 = 8'h10 == new_ptr_74_value ? ghv_16 : _GEN_9852; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9854 = 8'h11 == new_ptr_74_value ? ghv_17 : _GEN_9853; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9855 = 8'h12 == new_ptr_74_value ? ghv_18 : _GEN_9854; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9856 = 8'h13 == new_ptr_74_value ? ghv_19 : _GEN_9855; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9857 = 8'h14 == new_ptr_74_value ? ghv_20 : _GEN_9856; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9858 = 8'h15 == new_ptr_74_value ? ghv_21 : _GEN_9857; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9859 = 8'h16 == new_ptr_74_value ? ghv_22 : _GEN_9858; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9860 = 8'h17 == new_ptr_74_value ? ghv_23 : _GEN_9859; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9861 = 8'h18 == new_ptr_74_value ? ghv_24 : _GEN_9860; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9862 = 8'h19 == new_ptr_74_value ? ghv_25 : _GEN_9861; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9863 = 8'h1a == new_ptr_74_value ? ghv_26 : _GEN_9862; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9864 = 8'h1b == new_ptr_74_value ? ghv_27 : _GEN_9863; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9865 = 8'h1c == new_ptr_74_value ? ghv_28 : _GEN_9864; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9866 = 8'h1d == new_ptr_74_value ? ghv_29 : _GEN_9865; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9867 = 8'h1e == new_ptr_74_value ? ghv_30 : _GEN_9866; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9868 = 8'h1f == new_ptr_74_value ? ghv_31 : _GEN_9867; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9869 = 8'h20 == new_ptr_74_value ? ghv_32 : _GEN_9868; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9870 = 8'h21 == new_ptr_74_value ? ghv_33 : _GEN_9869; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9871 = 8'h22 == new_ptr_74_value ? ghv_34 : _GEN_9870; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9872 = 8'h23 == new_ptr_74_value ? ghv_35 : _GEN_9871; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9873 = 8'h24 == new_ptr_74_value ? ghv_36 : _GEN_9872; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9874 = 8'h25 == new_ptr_74_value ? ghv_37 : _GEN_9873; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9875 = 8'h26 == new_ptr_74_value ? ghv_38 : _GEN_9874; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9876 = 8'h27 == new_ptr_74_value ? ghv_39 : _GEN_9875; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9877 = 8'h28 == new_ptr_74_value ? ghv_40 : _GEN_9876; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9878 = 8'h29 == new_ptr_74_value ? ghv_41 : _GEN_9877; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9879 = 8'h2a == new_ptr_74_value ? ghv_42 : _GEN_9878; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9880 = 8'h2b == new_ptr_74_value ? ghv_43 : _GEN_9879; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9881 = 8'h2c == new_ptr_74_value ? ghv_44 : _GEN_9880; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9882 = 8'h2d == new_ptr_74_value ? ghv_45 : _GEN_9881; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9883 = 8'h2e == new_ptr_74_value ? ghv_46 : _GEN_9882; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9884 = 8'h2f == new_ptr_74_value ? ghv_47 : _GEN_9883; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9885 = 8'h30 == new_ptr_74_value ? ghv_48 : _GEN_9884; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9886 = 8'h31 == new_ptr_74_value ? ghv_49 : _GEN_9885; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9887 = 8'h32 == new_ptr_74_value ? ghv_50 : _GEN_9886; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9888 = 8'h33 == new_ptr_74_value ? ghv_51 : _GEN_9887; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9889 = 8'h34 == new_ptr_74_value ? ghv_52 : _GEN_9888; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9890 = 8'h35 == new_ptr_74_value ? ghv_53 : _GEN_9889; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9891 = 8'h36 == new_ptr_74_value ? ghv_54 : _GEN_9890; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9892 = 8'h37 == new_ptr_74_value ? ghv_55 : _GEN_9891; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9893 = 8'h38 == new_ptr_74_value ? ghv_56 : _GEN_9892; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9894 = 8'h39 == new_ptr_74_value ? ghv_57 : _GEN_9893; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9895 = 8'h3a == new_ptr_74_value ? ghv_58 : _GEN_9894; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9896 = 8'h3b == new_ptr_74_value ? ghv_59 : _GEN_9895; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9897 = 8'h3c == new_ptr_74_value ? ghv_60 : _GEN_9896; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9898 = 8'h3d == new_ptr_74_value ? ghv_61 : _GEN_9897; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9899 = 8'h3e == new_ptr_74_value ? ghv_62 : _GEN_9898; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9900 = 8'h3f == new_ptr_74_value ? ghv_63 : _GEN_9899; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9901 = 8'h40 == new_ptr_74_value ? ghv_64 : _GEN_9900; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9902 = 8'h41 == new_ptr_74_value ? ghv_65 : _GEN_9901; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9903 = 8'h42 == new_ptr_74_value ? ghv_66 : _GEN_9902; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9904 = 8'h43 == new_ptr_74_value ? ghv_67 : _GEN_9903; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9905 = 8'h44 == new_ptr_74_value ? ghv_68 : _GEN_9904; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9906 = 8'h45 == new_ptr_74_value ? ghv_69 : _GEN_9905; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9907 = 8'h46 == new_ptr_74_value ? ghv_70 : _GEN_9906; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9908 = 8'h47 == new_ptr_74_value ? ghv_71 : _GEN_9907; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9909 = 8'h48 == new_ptr_74_value ? ghv_72 : _GEN_9908; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9910 = 8'h49 == new_ptr_74_value ? ghv_73 : _GEN_9909; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9911 = 8'h4a == new_ptr_74_value ? ghv_74 : _GEN_9910; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9912 = 8'h4b == new_ptr_74_value ? ghv_75 : _GEN_9911; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9913 = 8'h4c == new_ptr_74_value ? ghv_76 : _GEN_9912; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9914 = 8'h4d == new_ptr_74_value ? ghv_77 : _GEN_9913; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9915 = 8'h4e == new_ptr_74_value ? ghv_78 : _GEN_9914; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9916 = 8'h4f == new_ptr_74_value ? ghv_79 : _GEN_9915; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9917 = 8'h50 == new_ptr_74_value ? ghv_80 : _GEN_9916; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9918 = 8'h51 == new_ptr_74_value ? ghv_81 : _GEN_9917; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9919 = 8'h52 == new_ptr_74_value ? ghv_82 : _GEN_9918; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9920 = 8'h53 == new_ptr_74_value ? ghv_83 : _GEN_9919; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9921 = 8'h54 == new_ptr_74_value ? ghv_84 : _GEN_9920; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9922 = 8'h55 == new_ptr_74_value ? ghv_85 : _GEN_9921; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9923 = 8'h56 == new_ptr_74_value ? ghv_86 : _GEN_9922; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9924 = 8'h57 == new_ptr_74_value ? ghv_87 : _GEN_9923; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9925 = 8'h58 == new_ptr_74_value ? ghv_88 : _GEN_9924; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9926 = 8'h59 == new_ptr_74_value ? ghv_89 : _GEN_9925; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9927 = 8'h5a == new_ptr_74_value ? ghv_90 : _GEN_9926; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9928 = 8'h5b == new_ptr_74_value ? ghv_91 : _GEN_9927; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9929 = 8'h5c == new_ptr_74_value ? ghv_92 : _GEN_9928; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9930 = 8'h5d == new_ptr_74_value ? ghv_93 : _GEN_9929; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9931 = 8'h5e == new_ptr_74_value ? ghv_94 : _GEN_9930; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9932 = 8'h5f == new_ptr_74_value ? ghv_95 : _GEN_9931; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9933 = 8'h60 == new_ptr_74_value ? ghv_96 : _GEN_9932; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9934 = 8'h61 == new_ptr_74_value ? ghv_97 : _GEN_9933; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9935 = 8'h62 == new_ptr_74_value ? ghv_98 : _GEN_9934; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9936 = 8'h63 == new_ptr_74_value ? ghv_99 : _GEN_9935; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9937 = 8'h64 == new_ptr_74_value ? ghv_100 : _GEN_9936; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9938 = 8'h65 == new_ptr_74_value ? ghv_101 : _GEN_9937; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9939 = 8'h66 == new_ptr_74_value ? ghv_102 : _GEN_9938; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9940 = 8'h67 == new_ptr_74_value ? ghv_103 : _GEN_9939; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9941 = 8'h68 == new_ptr_74_value ? ghv_104 : _GEN_9940; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9942 = 8'h69 == new_ptr_74_value ? ghv_105 : _GEN_9941; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9943 = 8'h6a == new_ptr_74_value ? ghv_106 : _GEN_9942; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9944 = 8'h6b == new_ptr_74_value ? ghv_107 : _GEN_9943; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9945 = 8'h6c == new_ptr_74_value ? ghv_108 : _GEN_9944; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9946 = 8'h6d == new_ptr_74_value ? ghv_109 : _GEN_9945; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9947 = 8'h6e == new_ptr_74_value ? ghv_110 : _GEN_9946; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9948 = 8'h6f == new_ptr_74_value ? ghv_111 : _GEN_9947; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9949 = 8'h70 == new_ptr_74_value ? ghv_112 : _GEN_9948; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9950 = 8'h71 == new_ptr_74_value ? ghv_113 : _GEN_9949; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9951 = 8'h72 == new_ptr_74_value ? ghv_114 : _GEN_9950; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9952 = 8'h73 == new_ptr_74_value ? ghv_115 : _GEN_9951; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9953 = 8'h74 == new_ptr_74_value ? ghv_116 : _GEN_9952; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9954 = 8'h75 == new_ptr_74_value ? ghv_117 : _GEN_9953; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9955 = 8'h76 == new_ptr_74_value ? ghv_118 : _GEN_9954; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9956 = 8'h77 == new_ptr_74_value ? ghv_119 : _GEN_9955; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9957 = 8'h78 == new_ptr_74_value ? ghv_120 : _GEN_9956; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9958 = 8'h79 == new_ptr_74_value ? ghv_121 : _GEN_9957; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9959 = 8'h7a == new_ptr_74_value ? ghv_122 : _GEN_9958; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9960 = 8'h7b == new_ptr_74_value ? ghv_123 : _GEN_9959; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9961 = 8'h7c == new_ptr_74_value ? ghv_124 : _GEN_9960; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9962 = 8'h7d == new_ptr_74_value ? ghv_125 : _GEN_9961; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9963 = 8'h7e == new_ptr_74_value ? ghv_126 : _GEN_9962; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9964 = 8'h7f == new_ptr_74_value ? ghv_127 : _GEN_9963; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9965 = 8'h80 == new_ptr_74_value ? ghv_128 : _GEN_9964; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9966 = 8'h81 == new_ptr_74_value ? ghv_129 : _GEN_9965; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9967 = 8'h82 == new_ptr_74_value ? ghv_130 : _GEN_9966; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9968 = 8'h83 == new_ptr_74_value ? ghv_131 : _GEN_9967; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9969 = 8'h84 == new_ptr_74_value ? ghv_132 : _GEN_9968; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9970 = 8'h85 == new_ptr_74_value ? ghv_133 : _GEN_9969; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9971 = 8'h86 == new_ptr_74_value ? ghv_134 : _GEN_9970; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9972 = 8'h87 == new_ptr_74_value ? ghv_135 : _GEN_9971; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9973 = 8'h88 == new_ptr_74_value ? ghv_136 : _GEN_9972; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9974 = 8'h89 == new_ptr_74_value ? ghv_137 : _GEN_9973; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9975 = 8'h8a == new_ptr_74_value ? ghv_138 : _GEN_9974; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9976 = 8'h8b == new_ptr_74_value ? ghv_139 : _GEN_9975; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9977 = 8'h8c == new_ptr_74_value ? ghv_140 : _GEN_9976; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9978 = 8'h8d == new_ptr_74_value ? ghv_141 : _GEN_9977; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9979 = 8'h8e == new_ptr_74_value ? ghv_142 : _GEN_9978; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_77_value = _new_ptr_value_T_155[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_9982 = 8'h1 == new_ptr_77_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9983 = 8'h2 == new_ptr_77_value ? ghv_2 : _GEN_9982; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9984 = 8'h3 == new_ptr_77_value ? ghv_3 : _GEN_9983; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9985 = 8'h4 == new_ptr_77_value ? ghv_4 : _GEN_9984; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9986 = 8'h5 == new_ptr_77_value ? ghv_5 : _GEN_9985; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9987 = 8'h6 == new_ptr_77_value ? ghv_6 : _GEN_9986; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9988 = 8'h7 == new_ptr_77_value ? ghv_7 : _GEN_9987; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9989 = 8'h8 == new_ptr_77_value ? ghv_8 : _GEN_9988; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9990 = 8'h9 == new_ptr_77_value ? ghv_9 : _GEN_9989; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9991 = 8'ha == new_ptr_77_value ? ghv_10 : _GEN_9990; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9992 = 8'hb == new_ptr_77_value ? ghv_11 : _GEN_9991; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9993 = 8'hc == new_ptr_77_value ? ghv_12 : _GEN_9992; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9994 = 8'hd == new_ptr_77_value ? ghv_13 : _GEN_9993; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9995 = 8'he == new_ptr_77_value ? ghv_14 : _GEN_9994; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9996 = 8'hf == new_ptr_77_value ? ghv_15 : _GEN_9995; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9997 = 8'h10 == new_ptr_77_value ? ghv_16 : _GEN_9996; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9998 = 8'h11 == new_ptr_77_value ? ghv_17 : _GEN_9997; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_9999 = 8'h12 == new_ptr_77_value ? ghv_18 : _GEN_9998; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10000 = 8'h13 == new_ptr_77_value ? ghv_19 : _GEN_9999; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10001 = 8'h14 == new_ptr_77_value ? ghv_20 : _GEN_10000; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10002 = 8'h15 == new_ptr_77_value ? ghv_21 : _GEN_10001; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10003 = 8'h16 == new_ptr_77_value ? ghv_22 : _GEN_10002; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10004 = 8'h17 == new_ptr_77_value ? ghv_23 : _GEN_10003; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10005 = 8'h18 == new_ptr_77_value ? ghv_24 : _GEN_10004; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10006 = 8'h19 == new_ptr_77_value ? ghv_25 : _GEN_10005; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10007 = 8'h1a == new_ptr_77_value ? ghv_26 : _GEN_10006; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10008 = 8'h1b == new_ptr_77_value ? ghv_27 : _GEN_10007; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10009 = 8'h1c == new_ptr_77_value ? ghv_28 : _GEN_10008; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10010 = 8'h1d == new_ptr_77_value ? ghv_29 : _GEN_10009; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10011 = 8'h1e == new_ptr_77_value ? ghv_30 : _GEN_10010; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10012 = 8'h1f == new_ptr_77_value ? ghv_31 : _GEN_10011; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10013 = 8'h20 == new_ptr_77_value ? ghv_32 : _GEN_10012; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10014 = 8'h21 == new_ptr_77_value ? ghv_33 : _GEN_10013; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10015 = 8'h22 == new_ptr_77_value ? ghv_34 : _GEN_10014; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10016 = 8'h23 == new_ptr_77_value ? ghv_35 : _GEN_10015; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10017 = 8'h24 == new_ptr_77_value ? ghv_36 : _GEN_10016; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10018 = 8'h25 == new_ptr_77_value ? ghv_37 : _GEN_10017; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10019 = 8'h26 == new_ptr_77_value ? ghv_38 : _GEN_10018; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10020 = 8'h27 == new_ptr_77_value ? ghv_39 : _GEN_10019; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10021 = 8'h28 == new_ptr_77_value ? ghv_40 : _GEN_10020; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10022 = 8'h29 == new_ptr_77_value ? ghv_41 : _GEN_10021; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10023 = 8'h2a == new_ptr_77_value ? ghv_42 : _GEN_10022; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10024 = 8'h2b == new_ptr_77_value ? ghv_43 : _GEN_10023; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10025 = 8'h2c == new_ptr_77_value ? ghv_44 : _GEN_10024; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10026 = 8'h2d == new_ptr_77_value ? ghv_45 : _GEN_10025; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10027 = 8'h2e == new_ptr_77_value ? ghv_46 : _GEN_10026; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10028 = 8'h2f == new_ptr_77_value ? ghv_47 : _GEN_10027; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10029 = 8'h30 == new_ptr_77_value ? ghv_48 : _GEN_10028; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10030 = 8'h31 == new_ptr_77_value ? ghv_49 : _GEN_10029; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10031 = 8'h32 == new_ptr_77_value ? ghv_50 : _GEN_10030; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10032 = 8'h33 == new_ptr_77_value ? ghv_51 : _GEN_10031; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10033 = 8'h34 == new_ptr_77_value ? ghv_52 : _GEN_10032; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10034 = 8'h35 == new_ptr_77_value ? ghv_53 : _GEN_10033; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10035 = 8'h36 == new_ptr_77_value ? ghv_54 : _GEN_10034; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10036 = 8'h37 == new_ptr_77_value ? ghv_55 : _GEN_10035; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10037 = 8'h38 == new_ptr_77_value ? ghv_56 : _GEN_10036; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10038 = 8'h39 == new_ptr_77_value ? ghv_57 : _GEN_10037; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10039 = 8'h3a == new_ptr_77_value ? ghv_58 : _GEN_10038; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10040 = 8'h3b == new_ptr_77_value ? ghv_59 : _GEN_10039; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10041 = 8'h3c == new_ptr_77_value ? ghv_60 : _GEN_10040; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10042 = 8'h3d == new_ptr_77_value ? ghv_61 : _GEN_10041; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10043 = 8'h3e == new_ptr_77_value ? ghv_62 : _GEN_10042; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10044 = 8'h3f == new_ptr_77_value ? ghv_63 : _GEN_10043; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10045 = 8'h40 == new_ptr_77_value ? ghv_64 : _GEN_10044; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10046 = 8'h41 == new_ptr_77_value ? ghv_65 : _GEN_10045; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10047 = 8'h42 == new_ptr_77_value ? ghv_66 : _GEN_10046; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10048 = 8'h43 == new_ptr_77_value ? ghv_67 : _GEN_10047; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10049 = 8'h44 == new_ptr_77_value ? ghv_68 : _GEN_10048; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10050 = 8'h45 == new_ptr_77_value ? ghv_69 : _GEN_10049; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10051 = 8'h46 == new_ptr_77_value ? ghv_70 : _GEN_10050; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10052 = 8'h47 == new_ptr_77_value ? ghv_71 : _GEN_10051; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10053 = 8'h48 == new_ptr_77_value ? ghv_72 : _GEN_10052; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10054 = 8'h49 == new_ptr_77_value ? ghv_73 : _GEN_10053; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10055 = 8'h4a == new_ptr_77_value ? ghv_74 : _GEN_10054; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10056 = 8'h4b == new_ptr_77_value ? ghv_75 : _GEN_10055; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10057 = 8'h4c == new_ptr_77_value ? ghv_76 : _GEN_10056; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10058 = 8'h4d == new_ptr_77_value ? ghv_77 : _GEN_10057; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10059 = 8'h4e == new_ptr_77_value ? ghv_78 : _GEN_10058; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10060 = 8'h4f == new_ptr_77_value ? ghv_79 : _GEN_10059; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10061 = 8'h50 == new_ptr_77_value ? ghv_80 : _GEN_10060; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10062 = 8'h51 == new_ptr_77_value ? ghv_81 : _GEN_10061; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10063 = 8'h52 == new_ptr_77_value ? ghv_82 : _GEN_10062; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10064 = 8'h53 == new_ptr_77_value ? ghv_83 : _GEN_10063; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10065 = 8'h54 == new_ptr_77_value ? ghv_84 : _GEN_10064; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10066 = 8'h55 == new_ptr_77_value ? ghv_85 : _GEN_10065; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10067 = 8'h56 == new_ptr_77_value ? ghv_86 : _GEN_10066; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10068 = 8'h57 == new_ptr_77_value ? ghv_87 : _GEN_10067; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10069 = 8'h58 == new_ptr_77_value ? ghv_88 : _GEN_10068; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10070 = 8'h59 == new_ptr_77_value ? ghv_89 : _GEN_10069; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10071 = 8'h5a == new_ptr_77_value ? ghv_90 : _GEN_10070; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10072 = 8'h5b == new_ptr_77_value ? ghv_91 : _GEN_10071; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10073 = 8'h5c == new_ptr_77_value ? ghv_92 : _GEN_10072; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10074 = 8'h5d == new_ptr_77_value ? ghv_93 : _GEN_10073; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10075 = 8'h5e == new_ptr_77_value ? ghv_94 : _GEN_10074; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10076 = 8'h5f == new_ptr_77_value ? ghv_95 : _GEN_10075; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10077 = 8'h60 == new_ptr_77_value ? ghv_96 : _GEN_10076; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10078 = 8'h61 == new_ptr_77_value ? ghv_97 : _GEN_10077; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10079 = 8'h62 == new_ptr_77_value ? ghv_98 : _GEN_10078; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10080 = 8'h63 == new_ptr_77_value ? ghv_99 : _GEN_10079; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10081 = 8'h64 == new_ptr_77_value ? ghv_100 : _GEN_10080; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10082 = 8'h65 == new_ptr_77_value ? ghv_101 : _GEN_10081; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10083 = 8'h66 == new_ptr_77_value ? ghv_102 : _GEN_10082; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10084 = 8'h67 == new_ptr_77_value ? ghv_103 : _GEN_10083; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10085 = 8'h68 == new_ptr_77_value ? ghv_104 : _GEN_10084; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10086 = 8'h69 == new_ptr_77_value ? ghv_105 : _GEN_10085; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10087 = 8'h6a == new_ptr_77_value ? ghv_106 : _GEN_10086; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10088 = 8'h6b == new_ptr_77_value ? ghv_107 : _GEN_10087; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10089 = 8'h6c == new_ptr_77_value ? ghv_108 : _GEN_10088; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10090 = 8'h6d == new_ptr_77_value ? ghv_109 : _GEN_10089; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10091 = 8'h6e == new_ptr_77_value ? ghv_110 : _GEN_10090; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10092 = 8'h6f == new_ptr_77_value ? ghv_111 : _GEN_10091; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10093 = 8'h70 == new_ptr_77_value ? ghv_112 : _GEN_10092; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10094 = 8'h71 == new_ptr_77_value ? ghv_113 : _GEN_10093; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10095 = 8'h72 == new_ptr_77_value ? ghv_114 : _GEN_10094; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10096 = 8'h73 == new_ptr_77_value ? ghv_115 : _GEN_10095; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10097 = 8'h74 == new_ptr_77_value ? ghv_116 : _GEN_10096; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10098 = 8'h75 == new_ptr_77_value ? ghv_117 : _GEN_10097; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10099 = 8'h76 == new_ptr_77_value ? ghv_118 : _GEN_10098; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10100 = 8'h77 == new_ptr_77_value ? ghv_119 : _GEN_10099; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10101 = 8'h78 == new_ptr_77_value ? ghv_120 : _GEN_10100; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10102 = 8'h79 == new_ptr_77_value ? ghv_121 : _GEN_10101; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10103 = 8'h7a == new_ptr_77_value ? ghv_122 : _GEN_10102; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10104 = 8'h7b == new_ptr_77_value ? ghv_123 : _GEN_10103; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10105 = 8'h7c == new_ptr_77_value ? ghv_124 : _GEN_10104; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10106 = 8'h7d == new_ptr_77_value ? ghv_125 : _GEN_10105; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10107 = 8'h7e == new_ptr_77_value ? ghv_126 : _GEN_10106; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10108 = 8'h7f == new_ptr_77_value ? ghv_127 : _GEN_10107; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10109 = 8'h80 == new_ptr_77_value ? ghv_128 : _GEN_10108; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10110 = 8'h81 == new_ptr_77_value ? ghv_129 : _GEN_10109; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10111 = 8'h82 == new_ptr_77_value ? ghv_130 : _GEN_10110; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10112 = 8'h83 == new_ptr_77_value ? ghv_131 : _GEN_10111; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10113 = 8'h84 == new_ptr_77_value ? ghv_132 : _GEN_10112; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10114 = 8'h85 == new_ptr_77_value ? ghv_133 : _GEN_10113; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10115 = 8'h86 == new_ptr_77_value ? ghv_134 : _GEN_10114; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10116 = 8'h87 == new_ptr_77_value ? ghv_135 : _GEN_10115; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10117 = 8'h88 == new_ptr_77_value ? ghv_136 : _GEN_10116; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10118 = 8'h89 == new_ptr_77_value ? ghv_137 : _GEN_10117; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10119 = 8'h8a == new_ptr_77_value ? ghv_138 : _GEN_10118; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10120 = 8'h8b == new_ptr_77_value ? ghv_139 : _GEN_10119; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10121 = 8'h8c == new_ptr_77_value ? ghv_140 : _GEN_10120; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10122 = 8'h8d == new_ptr_77_value ? ghv_141 : _GEN_10121; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10123 = 8'h8e == new_ptr_77_value ? ghv_142 : _GEN_10122; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_64_value = _new_ptr_value_T_129[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_10126 = 8'h1 == new_ptr_64_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10127 = 8'h2 == new_ptr_64_value ? ghv_2 : _GEN_10126; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10128 = 8'h3 == new_ptr_64_value ? ghv_3 : _GEN_10127; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10129 = 8'h4 == new_ptr_64_value ? ghv_4 : _GEN_10128; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10130 = 8'h5 == new_ptr_64_value ? ghv_5 : _GEN_10129; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10131 = 8'h6 == new_ptr_64_value ? ghv_6 : _GEN_10130; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10132 = 8'h7 == new_ptr_64_value ? ghv_7 : _GEN_10131; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10133 = 8'h8 == new_ptr_64_value ? ghv_8 : _GEN_10132; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10134 = 8'h9 == new_ptr_64_value ? ghv_9 : _GEN_10133; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10135 = 8'ha == new_ptr_64_value ? ghv_10 : _GEN_10134; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10136 = 8'hb == new_ptr_64_value ? ghv_11 : _GEN_10135; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10137 = 8'hc == new_ptr_64_value ? ghv_12 : _GEN_10136; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10138 = 8'hd == new_ptr_64_value ? ghv_13 : _GEN_10137; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10139 = 8'he == new_ptr_64_value ? ghv_14 : _GEN_10138; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10140 = 8'hf == new_ptr_64_value ? ghv_15 : _GEN_10139; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10141 = 8'h10 == new_ptr_64_value ? ghv_16 : _GEN_10140; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10142 = 8'h11 == new_ptr_64_value ? ghv_17 : _GEN_10141; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10143 = 8'h12 == new_ptr_64_value ? ghv_18 : _GEN_10142; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10144 = 8'h13 == new_ptr_64_value ? ghv_19 : _GEN_10143; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10145 = 8'h14 == new_ptr_64_value ? ghv_20 : _GEN_10144; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10146 = 8'h15 == new_ptr_64_value ? ghv_21 : _GEN_10145; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10147 = 8'h16 == new_ptr_64_value ? ghv_22 : _GEN_10146; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10148 = 8'h17 == new_ptr_64_value ? ghv_23 : _GEN_10147; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10149 = 8'h18 == new_ptr_64_value ? ghv_24 : _GEN_10148; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10150 = 8'h19 == new_ptr_64_value ? ghv_25 : _GEN_10149; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10151 = 8'h1a == new_ptr_64_value ? ghv_26 : _GEN_10150; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10152 = 8'h1b == new_ptr_64_value ? ghv_27 : _GEN_10151; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10153 = 8'h1c == new_ptr_64_value ? ghv_28 : _GEN_10152; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10154 = 8'h1d == new_ptr_64_value ? ghv_29 : _GEN_10153; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10155 = 8'h1e == new_ptr_64_value ? ghv_30 : _GEN_10154; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10156 = 8'h1f == new_ptr_64_value ? ghv_31 : _GEN_10155; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10157 = 8'h20 == new_ptr_64_value ? ghv_32 : _GEN_10156; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10158 = 8'h21 == new_ptr_64_value ? ghv_33 : _GEN_10157; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10159 = 8'h22 == new_ptr_64_value ? ghv_34 : _GEN_10158; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10160 = 8'h23 == new_ptr_64_value ? ghv_35 : _GEN_10159; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10161 = 8'h24 == new_ptr_64_value ? ghv_36 : _GEN_10160; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10162 = 8'h25 == new_ptr_64_value ? ghv_37 : _GEN_10161; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10163 = 8'h26 == new_ptr_64_value ? ghv_38 : _GEN_10162; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10164 = 8'h27 == new_ptr_64_value ? ghv_39 : _GEN_10163; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10165 = 8'h28 == new_ptr_64_value ? ghv_40 : _GEN_10164; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10166 = 8'h29 == new_ptr_64_value ? ghv_41 : _GEN_10165; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10167 = 8'h2a == new_ptr_64_value ? ghv_42 : _GEN_10166; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10168 = 8'h2b == new_ptr_64_value ? ghv_43 : _GEN_10167; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10169 = 8'h2c == new_ptr_64_value ? ghv_44 : _GEN_10168; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10170 = 8'h2d == new_ptr_64_value ? ghv_45 : _GEN_10169; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10171 = 8'h2e == new_ptr_64_value ? ghv_46 : _GEN_10170; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10172 = 8'h2f == new_ptr_64_value ? ghv_47 : _GEN_10171; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10173 = 8'h30 == new_ptr_64_value ? ghv_48 : _GEN_10172; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10174 = 8'h31 == new_ptr_64_value ? ghv_49 : _GEN_10173; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10175 = 8'h32 == new_ptr_64_value ? ghv_50 : _GEN_10174; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10176 = 8'h33 == new_ptr_64_value ? ghv_51 : _GEN_10175; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10177 = 8'h34 == new_ptr_64_value ? ghv_52 : _GEN_10176; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10178 = 8'h35 == new_ptr_64_value ? ghv_53 : _GEN_10177; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10179 = 8'h36 == new_ptr_64_value ? ghv_54 : _GEN_10178; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10180 = 8'h37 == new_ptr_64_value ? ghv_55 : _GEN_10179; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10181 = 8'h38 == new_ptr_64_value ? ghv_56 : _GEN_10180; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10182 = 8'h39 == new_ptr_64_value ? ghv_57 : _GEN_10181; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10183 = 8'h3a == new_ptr_64_value ? ghv_58 : _GEN_10182; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10184 = 8'h3b == new_ptr_64_value ? ghv_59 : _GEN_10183; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10185 = 8'h3c == new_ptr_64_value ? ghv_60 : _GEN_10184; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10186 = 8'h3d == new_ptr_64_value ? ghv_61 : _GEN_10185; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10187 = 8'h3e == new_ptr_64_value ? ghv_62 : _GEN_10186; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10188 = 8'h3f == new_ptr_64_value ? ghv_63 : _GEN_10187; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10189 = 8'h40 == new_ptr_64_value ? ghv_64 : _GEN_10188; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10190 = 8'h41 == new_ptr_64_value ? ghv_65 : _GEN_10189; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10191 = 8'h42 == new_ptr_64_value ? ghv_66 : _GEN_10190; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10192 = 8'h43 == new_ptr_64_value ? ghv_67 : _GEN_10191; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10193 = 8'h44 == new_ptr_64_value ? ghv_68 : _GEN_10192; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10194 = 8'h45 == new_ptr_64_value ? ghv_69 : _GEN_10193; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10195 = 8'h46 == new_ptr_64_value ? ghv_70 : _GEN_10194; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10196 = 8'h47 == new_ptr_64_value ? ghv_71 : _GEN_10195; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10197 = 8'h48 == new_ptr_64_value ? ghv_72 : _GEN_10196; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10198 = 8'h49 == new_ptr_64_value ? ghv_73 : _GEN_10197; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10199 = 8'h4a == new_ptr_64_value ? ghv_74 : _GEN_10198; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10200 = 8'h4b == new_ptr_64_value ? ghv_75 : _GEN_10199; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10201 = 8'h4c == new_ptr_64_value ? ghv_76 : _GEN_10200; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10202 = 8'h4d == new_ptr_64_value ? ghv_77 : _GEN_10201; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10203 = 8'h4e == new_ptr_64_value ? ghv_78 : _GEN_10202; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10204 = 8'h4f == new_ptr_64_value ? ghv_79 : _GEN_10203; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10205 = 8'h50 == new_ptr_64_value ? ghv_80 : _GEN_10204; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10206 = 8'h51 == new_ptr_64_value ? ghv_81 : _GEN_10205; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10207 = 8'h52 == new_ptr_64_value ? ghv_82 : _GEN_10206; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10208 = 8'h53 == new_ptr_64_value ? ghv_83 : _GEN_10207; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10209 = 8'h54 == new_ptr_64_value ? ghv_84 : _GEN_10208; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10210 = 8'h55 == new_ptr_64_value ? ghv_85 : _GEN_10209; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10211 = 8'h56 == new_ptr_64_value ? ghv_86 : _GEN_10210; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10212 = 8'h57 == new_ptr_64_value ? ghv_87 : _GEN_10211; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10213 = 8'h58 == new_ptr_64_value ? ghv_88 : _GEN_10212; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10214 = 8'h59 == new_ptr_64_value ? ghv_89 : _GEN_10213; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10215 = 8'h5a == new_ptr_64_value ? ghv_90 : _GEN_10214; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10216 = 8'h5b == new_ptr_64_value ? ghv_91 : _GEN_10215; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10217 = 8'h5c == new_ptr_64_value ? ghv_92 : _GEN_10216; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10218 = 8'h5d == new_ptr_64_value ? ghv_93 : _GEN_10217; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10219 = 8'h5e == new_ptr_64_value ? ghv_94 : _GEN_10218; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10220 = 8'h5f == new_ptr_64_value ? ghv_95 : _GEN_10219; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10221 = 8'h60 == new_ptr_64_value ? ghv_96 : _GEN_10220; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10222 = 8'h61 == new_ptr_64_value ? ghv_97 : _GEN_10221; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10223 = 8'h62 == new_ptr_64_value ? ghv_98 : _GEN_10222; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10224 = 8'h63 == new_ptr_64_value ? ghv_99 : _GEN_10223; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10225 = 8'h64 == new_ptr_64_value ? ghv_100 : _GEN_10224; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10226 = 8'h65 == new_ptr_64_value ? ghv_101 : _GEN_10225; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10227 = 8'h66 == new_ptr_64_value ? ghv_102 : _GEN_10226; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10228 = 8'h67 == new_ptr_64_value ? ghv_103 : _GEN_10227; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10229 = 8'h68 == new_ptr_64_value ? ghv_104 : _GEN_10228; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10230 = 8'h69 == new_ptr_64_value ? ghv_105 : _GEN_10229; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10231 = 8'h6a == new_ptr_64_value ? ghv_106 : _GEN_10230; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10232 = 8'h6b == new_ptr_64_value ? ghv_107 : _GEN_10231; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10233 = 8'h6c == new_ptr_64_value ? ghv_108 : _GEN_10232; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10234 = 8'h6d == new_ptr_64_value ? ghv_109 : _GEN_10233; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10235 = 8'h6e == new_ptr_64_value ? ghv_110 : _GEN_10234; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10236 = 8'h6f == new_ptr_64_value ? ghv_111 : _GEN_10235; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10237 = 8'h70 == new_ptr_64_value ? ghv_112 : _GEN_10236; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10238 = 8'h71 == new_ptr_64_value ? ghv_113 : _GEN_10237; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10239 = 8'h72 == new_ptr_64_value ? ghv_114 : _GEN_10238; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10240 = 8'h73 == new_ptr_64_value ? ghv_115 : _GEN_10239; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10241 = 8'h74 == new_ptr_64_value ? ghv_116 : _GEN_10240; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10242 = 8'h75 == new_ptr_64_value ? ghv_117 : _GEN_10241; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10243 = 8'h76 == new_ptr_64_value ? ghv_118 : _GEN_10242; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10244 = 8'h77 == new_ptr_64_value ? ghv_119 : _GEN_10243; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10245 = 8'h78 == new_ptr_64_value ? ghv_120 : _GEN_10244; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10246 = 8'h79 == new_ptr_64_value ? ghv_121 : _GEN_10245; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10247 = 8'h7a == new_ptr_64_value ? ghv_122 : _GEN_10246; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10248 = 8'h7b == new_ptr_64_value ? ghv_123 : _GEN_10247; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10249 = 8'h7c == new_ptr_64_value ? ghv_124 : _GEN_10248; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10250 = 8'h7d == new_ptr_64_value ? ghv_125 : _GEN_10249; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10251 = 8'h7e == new_ptr_64_value ? ghv_126 : _GEN_10250; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10252 = 8'h7f == new_ptr_64_value ? ghv_127 : _GEN_10251; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10253 = 8'h80 == new_ptr_64_value ? ghv_128 : _GEN_10252; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10254 = 8'h81 == new_ptr_64_value ? ghv_129 : _GEN_10253; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10255 = 8'h82 == new_ptr_64_value ? ghv_130 : _GEN_10254; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10256 = 8'h83 == new_ptr_64_value ? ghv_131 : _GEN_10255; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10257 = 8'h84 == new_ptr_64_value ? ghv_132 : _GEN_10256; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10258 = 8'h85 == new_ptr_64_value ? ghv_133 : _GEN_10257; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10259 = 8'h86 == new_ptr_64_value ? ghv_134 : _GEN_10258; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10260 = 8'h87 == new_ptr_64_value ? ghv_135 : _GEN_10259; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10261 = 8'h88 == new_ptr_64_value ? ghv_136 : _GEN_10260; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10262 = 8'h89 == new_ptr_64_value ? ghv_137 : _GEN_10261; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10263 = 8'h8a == new_ptr_64_value ? ghv_138 : _GEN_10262; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10264 = 8'h8b == new_ptr_64_value ? ghv_139 : _GEN_10263; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10265 = 8'h8c == new_ptr_64_value ? ghv_140 : _GEN_10264; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10266 = 8'h8d == new_ptr_64_value ? ghv_141 : _GEN_10265; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10267 = 8'h8e == new_ptr_64_value ? ghv_142 : _GEN_10266; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_68_value = _new_ptr_value_T_137[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_10270 = 8'h1 == new_ptr_68_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10271 = 8'h2 == new_ptr_68_value ? ghv_2 : _GEN_10270; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10272 = 8'h3 == new_ptr_68_value ? ghv_3 : _GEN_10271; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10273 = 8'h4 == new_ptr_68_value ? ghv_4 : _GEN_10272; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10274 = 8'h5 == new_ptr_68_value ? ghv_5 : _GEN_10273; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10275 = 8'h6 == new_ptr_68_value ? ghv_6 : _GEN_10274; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10276 = 8'h7 == new_ptr_68_value ? ghv_7 : _GEN_10275; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10277 = 8'h8 == new_ptr_68_value ? ghv_8 : _GEN_10276; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10278 = 8'h9 == new_ptr_68_value ? ghv_9 : _GEN_10277; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10279 = 8'ha == new_ptr_68_value ? ghv_10 : _GEN_10278; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10280 = 8'hb == new_ptr_68_value ? ghv_11 : _GEN_10279; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10281 = 8'hc == new_ptr_68_value ? ghv_12 : _GEN_10280; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10282 = 8'hd == new_ptr_68_value ? ghv_13 : _GEN_10281; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10283 = 8'he == new_ptr_68_value ? ghv_14 : _GEN_10282; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10284 = 8'hf == new_ptr_68_value ? ghv_15 : _GEN_10283; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10285 = 8'h10 == new_ptr_68_value ? ghv_16 : _GEN_10284; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10286 = 8'h11 == new_ptr_68_value ? ghv_17 : _GEN_10285; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10287 = 8'h12 == new_ptr_68_value ? ghv_18 : _GEN_10286; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10288 = 8'h13 == new_ptr_68_value ? ghv_19 : _GEN_10287; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10289 = 8'h14 == new_ptr_68_value ? ghv_20 : _GEN_10288; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10290 = 8'h15 == new_ptr_68_value ? ghv_21 : _GEN_10289; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10291 = 8'h16 == new_ptr_68_value ? ghv_22 : _GEN_10290; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10292 = 8'h17 == new_ptr_68_value ? ghv_23 : _GEN_10291; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10293 = 8'h18 == new_ptr_68_value ? ghv_24 : _GEN_10292; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10294 = 8'h19 == new_ptr_68_value ? ghv_25 : _GEN_10293; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10295 = 8'h1a == new_ptr_68_value ? ghv_26 : _GEN_10294; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10296 = 8'h1b == new_ptr_68_value ? ghv_27 : _GEN_10295; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10297 = 8'h1c == new_ptr_68_value ? ghv_28 : _GEN_10296; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10298 = 8'h1d == new_ptr_68_value ? ghv_29 : _GEN_10297; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10299 = 8'h1e == new_ptr_68_value ? ghv_30 : _GEN_10298; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10300 = 8'h1f == new_ptr_68_value ? ghv_31 : _GEN_10299; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10301 = 8'h20 == new_ptr_68_value ? ghv_32 : _GEN_10300; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10302 = 8'h21 == new_ptr_68_value ? ghv_33 : _GEN_10301; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10303 = 8'h22 == new_ptr_68_value ? ghv_34 : _GEN_10302; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10304 = 8'h23 == new_ptr_68_value ? ghv_35 : _GEN_10303; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10305 = 8'h24 == new_ptr_68_value ? ghv_36 : _GEN_10304; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10306 = 8'h25 == new_ptr_68_value ? ghv_37 : _GEN_10305; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10307 = 8'h26 == new_ptr_68_value ? ghv_38 : _GEN_10306; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10308 = 8'h27 == new_ptr_68_value ? ghv_39 : _GEN_10307; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10309 = 8'h28 == new_ptr_68_value ? ghv_40 : _GEN_10308; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10310 = 8'h29 == new_ptr_68_value ? ghv_41 : _GEN_10309; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10311 = 8'h2a == new_ptr_68_value ? ghv_42 : _GEN_10310; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10312 = 8'h2b == new_ptr_68_value ? ghv_43 : _GEN_10311; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10313 = 8'h2c == new_ptr_68_value ? ghv_44 : _GEN_10312; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10314 = 8'h2d == new_ptr_68_value ? ghv_45 : _GEN_10313; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10315 = 8'h2e == new_ptr_68_value ? ghv_46 : _GEN_10314; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10316 = 8'h2f == new_ptr_68_value ? ghv_47 : _GEN_10315; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10317 = 8'h30 == new_ptr_68_value ? ghv_48 : _GEN_10316; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10318 = 8'h31 == new_ptr_68_value ? ghv_49 : _GEN_10317; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10319 = 8'h32 == new_ptr_68_value ? ghv_50 : _GEN_10318; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10320 = 8'h33 == new_ptr_68_value ? ghv_51 : _GEN_10319; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10321 = 8'h34 == new_ptr_68_value ? ghv_52 : _GEN_10320; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10322 = 8'h35 == new_ptr_68_value ? ghv_53 : _GEN_10321; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10323 = 8'h36 == new_ptr_68_value ? ghv_54 : _GEN_10322; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10324 = 8'h37 == new_ptr_68_value ? ghv_55 : _GEN_10323; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10325 = 8'h38 == new_ptr_68_value ? ghv_56 : _GEN_10324; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10326 = 8'h39 == new_ptr_68_value ? ghv_57 : _GEN_10325; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10327 = 8'h3a == new_ptr_68_value ? ghv_58 : _GEN_10326; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10328 = 8'h3b == new_ptr_68_value ? ghv_59 : _GEN_10327; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10329 = 8'h3c == new_ptr_68_value ? ghv_60 : _GEN_10328; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10330 = 8'h3d == new_ptr_68_value ? ghv_61 : _GEN_10329; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10331 = 8'h3e == new_ptr_68_value ? ghv_62 : _GEN_10330; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10332 = 8'h3f == new_ptr_68_value ? ghv_63 : _GEN_10331; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10333 = 8'h40 == new_ptr_68_value ? ghv_64 : _GEN_10332; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10334 = 8'h41 == new_ptr_68_value ? ghv_65 : _GEN_10333; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10335 = 8'h42 == new_ptr_68_value ? ghv_66 : _GEN_10334; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10336 = 8'h43 == new_ptr_68_value ? ghv_67 : _GEN_10335; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10337 = 8'h44 == new_ptr_68_value ? ghv_68 : _GEN_10336; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10338 = 8'h45 == new_ptr_68_value ? ghv_69 : _GEN_10337; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10339 = 8'h46 == new_ptr_68_value ? ghv_70 : _GEN_10338; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10340 = 8'h47 == new_ptr_68_value ? ghv_71 : _GEN_10339; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10341 = 8'h48 == new_ptr_68_value ? ghv_72 : _GEN_10340; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10342 = 8'h49 == new_ptr_68_value ? ghv_73 : _GEN_10341; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10343 = 8'h4a == new_ptr_68_value ? ghv_74 : _GEN_10342; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10344 = 8'h4b == new_ptr_68_value ? ghv_75 : _GEN_10343; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10345 = 8'h4c == new_ptr_68_value ? ghv_76 : _GEN_10344; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10346 = 8'h4d == new_ptr_68_value ? ghv_77 : _GEN_10345; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10347 = 8'h4e == new_ptr_68_value ? ghv_78 : _GEN_10346; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10348 = 8'h4f == new_ptr_68_value ? ghv_79 : _GEN_10347; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10349 = 8'h50 == new_ptr_68_value ? ghv_80 : _GEN_10348; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10350 = 8'h51 == new_ptr_68_value ? ghv_81 : _GEN_10349; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10351 = 8'h52 == new_ptr_68_value ? ghv_82 : _GEN_10350; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10352 = 8'h53 == new_ptr_68_value ? ghv_83 : _GEN_10351; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10353 = 8'h54 == new_ptr_68_value ? ghv_84 : _GEN_10352; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10354 = 8'h55 == new_ptr_68_value ? ghv_85 : _GEN_10353; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10355 = 8'h56 == new_ptr_68_value ? ghv_86 : _GEN_10354; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10356 = 8'h57 == new_ptr_68_value ? ghv_87 : _GEN_10355; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10357 = 8'h58 == new_ptr_68_value ? ghv_88 : _GEN_10356; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10358 = 8'h59 == new_ptr_68_value ? ghv_89 : _GEN_10357; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10359 = 8'h5a == new_ptr_68_value ? ghv_90 : _GEN_10358; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10360 = 8'h5b == new_ptr_68_value ? ghv_91 : _GEN_10359; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10361 = 8'h5c == new_ptr_68_value ? ghv_92 : _GEN_10360; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10362 = 8'h5d == new_ptr_68_value ? ghv_93 : _GEN_10361; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10363 = 8'h5e == new_ptr_68_value ? ghv_94 : _GEN_10362; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10364 = 8'h5f == new_ptr_68_value ? ghv_95 : _GEN_10363; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10365 = 8'h60 == new_ptr_68_value ? ghv_96 : _GEN_10364; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10366 = 8'h61 == new_ptr_68_value ? ghv_97 : _GEN_10365; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10367 = 8'h62 == new_ptr_68_value ? ghv_98 : _GEN_10366; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10368 = 8'h63 == new_ptr_68_value ? ghv_99 : _GEN_10367; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10369 = 8'h64 == new_ptr_68_value ? ghv_100 : _GEN_10368; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10370 = 8'h65 == new_ptr_68_value ? ghv_101 : _GEN_10369; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10371 = 8'h66 == new_ptr_68_value ? ghv_102 : _GEN_10370; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10372 = 8'h67 == new_ptr_68_value ? ghv_103 : _GEN_10371; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10373 = 8'h68 == new_ptr_68_value ? ghv_104 : _GEN_10372; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10374 = 8'h69 == new_ptr_68_value ? ghv_105 : _GEN_10373; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10375 = 8'h6a == new_ptr_68_value ? ghv_106 : _GEN_10374; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10376 = 8'h6b == new_ptr_68_value ? ghv_107 : _GEN_10375; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10377 = 8'h6c == new_ptr_68_value ? ghv_108 : _GEN_10376; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10378 = 8'h6d == new_ptr_68_value ? ghv_109 : _GEN_10377; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10379 = 8'h6e == new_ptr_68_value ? ghv_110 : _GEN_10378; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10380 = 8'h6f == new_ptr_68_value ? ghv_111 : _GEN_10379; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10381 = 8'h70 == new_ptr_68_value ? ghv_112 : _GEN_10380; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10382 = 8'h71 == new_ptr_68_value ? ghv_113 : _GEN_10381; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10383 = 8'h72 == new_ptr_68_value ? ghv_114 : _GEN_10382; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10384 = 8'h73 == new_ptr_68_value ? ghv_115 : _GEN_10383; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10385 = 8'h74 == new_ptr_68_value ? ghv_116 : _GEN_10384; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10386 = 8'h75 == new_ptr_68_value ? ghv_117 : _GEN_10385; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10387 = 8'h76 == new_ptr_68_value ? ghv_118 : _GEN_10386; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10388 = 8'h77 == new_ptr_68_value ? ghv_119 : _GEN_10387; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10389 = 8'h78 == new_ptr_68_value ? ghv_120 : _GEN_10388; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10390 = 8'h79 == new_ptr_68_value ? ghv_121 : _GEN_10389; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10391 = 8'h7a == new_ptr_68_value ? ghv_122 : _GEN_10390; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10392 = 8'h7b == new_ptr_68_value ? ghv_123 : _GEN_10391; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10393 = 8'h7c == new_ptr_68_value ? ghv_124 : _GEN_10392; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10394 = 8'h7d == new_ptr_68_value ? ghv_125 : _GEN_10393; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10395 = 8'h7e == new_ptr_68_value ? ghv_126 : _GEN_10394; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10396 = 8'h7f == new_ptr_68_value ? ghv_127 : _GEN_10395; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10397 = 8'h80 == new_ptr_68_value ? ghv_128 : _GEN_10396; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10398 = 8'h81 == new_ptr_68_value ? ghv_129 : _GEN_10397; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10399 = 8'h82 == new_ptr_68_value ? ghv_130 : _GEN_10398; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10400 = 8'h83 == new_ptr_68_value ? ghv_131 : _GEN_10399; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10401 = 8'h84 == new_ptr_68_value ? ghv_132 : _GEN_10400; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10402 = 8'h85 == new_ptr_68_value ? ghv_133 : _GEN_10401; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10403 = 8'h86 == new_ptr_68_value ? ghv_134 : _GEN_10402; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10404 = 8'h87 == new_ptr_68_value ? ghv_135 : _GEN_10403; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10405 = 8'h88 == new_ptr_68_value ? ghv_136 : _GEN_10404; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10406 = 8'h89 == new_ptr_68_value ? ghv_137 : _GEN_10405; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10407 = 8'h8a == new_ptr_68_value ? ghv_138 : _GEN_10406; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10408 = 8'h8b == new_ptr_68_value ? ghv_139 : _GEN_10407; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10409 = 8'h8c == new_ptr_68_value ? ghv_140 : _GEN_10408; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10410 = 8'h8d == new_ptr_68_value ? ghv_141 : _GEN_10409; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10411 = 8'h8e == new_ptr_68_value ? ghv_142 : _GEN_10410; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_79_value = _new_ptr_value_T_159[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_10414 = 8'h1 == new_ptr_79_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10415 = 8'h2 == new_ptr_79_value ? ghv_2 : _GEN_10414; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10416 = 8'h3 == new_ptr_79_value ? ghv_3 : _GEN_10415; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10417 = 8'h4 == new_ptr_79_value ? ghv_4 : _GEN_10416; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10418 = 8'h5 == new_ptr_79_value ? ghv_5 : _GEN_10417; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10419 = 8'h6 == new_ptr_79_value ? ghv_6 : _GEN_10418; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10420 = 8'h7 == new_ptr_79_value ? ghv_7 : _GEN_10419; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10421 = 8'h8 == new_ptr_79_value ? ghv_8 : _GEN_10420; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10422 = 8'h9 == new_ptr_79_value ? ghv_9 : _GEN_10421; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10423 = 8'ha == new_ptr_79_value ? ghv_10 : _GEN_10422; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10424 = 8'hb == new_ptr_79_value ? ghv_11 : _GEN_10423; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10425 = 8'hc == new_ptr_79_value ? ghv_12 : _GEN_10424; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10426 = 8'hd == new_ptr_79_value ? ghv_13 : _GEN_10425; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10427 = 8'he == new_ptr_79_value ? ghv_14 : _GEN_10426; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10428 = 8'hf == new_ptr_79_value ? ghv_15 : _GEN_10427; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10429 = 8'h10 == new_ptr_79_value ? ghv_16 : _GEN_10428; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10430 = 8'h11 == new_ptr_79_value ? ghv_17 : _GEN_10429; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10431 = 8'h12 == new_ptr_79_value ? ghv_18 : _GEN_10430; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10432 = 8'h13 == new_ptr_79_value ? ghv_19 : _GEN_10431; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10433 = 8'h14 == new_ptr_79_value ? ghv_20 : _GEN_10432; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10434 = 8'h15 == new_ptr_79_value ? ghv_21 : _GEN_10433; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10435 = 8'h16 == new_ptr_79_value ? ghv_22 : _GEN_10434; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10436 = 8'h17 == new_ptr_79_value ? ghv_23 : _GEN_10435; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10437 = 8'h18 == new_ptr_79_value ? ghv_24 : _GEN_10436; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10438 = 8'h19 == new_ptr_79_value ? ghv_25 : _GEN_10437; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10439 = 8'h1a == new_ptr_79_value ? ghv_26 : _GEN_10438; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10440 = 8'h1b == new_ptr_79_value ? ghv_27 : _GEN_10439; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10441 = 8'h1c == new_ptr_79_value ? ghv_28 : _GEN_10440; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10442 = 8'h1d == new_ptr_79_value ? ghv_29 : _GEN_10441; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10443 = 8'h1e == new_ptr_79_value ? ghv_30 : _GEN_10442; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10444 = 8'h1f == new_ptr_79_value ? ghv_31 : _GEN_10443; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10445 = 8'h20 == new_ptr_79_value ? ghv_32 : _GEN_10444; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10446 = 8'h21 == new_ptr_79_value ? ghv_33 : _GEN_10445; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10447 = 8'h22 == new_ptr_79_value ? ghv_34 : _GEN_10446; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10448 = 8'h23 == new_ptr_79_value ? ghv_35 : _GEN_10447; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10449 = 8'h24 == new_ptr_79_value ? ghv_36 : _GEN_10448; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10450 = 8'h25 == new_ptr_79_value ? ghv_37 : _GEN_10449; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10451 = 8'h26 == new_ptr_79_value ? ghv_38 : _GEN_10450; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10452 = 8'h27 == new_ptr_79_value ? ghv_39 : _GEN_10451; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10453 = 8'h28 == new_ptr_79_value ? ghv_40 : _GEN_10452; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10454 = 8'h29 == new_ptr_79_value ? ghv_41 : _GEN_10453; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10455 = 8'h2a == new_ptr_79_value ? ghv_42 : _GEN_10454; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10456 = 8'h2b == new_ptr_79_value ? ghv_43 : _GEN_10455; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10457 = 8'h2c == new_ptr_79_value ? ghv_44 : _GEN_10456; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10458 = 8'h2d == new_ptr_79_value ? ghv_45 : _GEN_10457; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10459 = 8'h2e == new_ptr_79_value ? ghv_46 : _GEN_10458; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10460 = 8'h2f == new_ptr_79_value ? ghv_47 : _GEN_10459; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10461 = 8'h30 == new_ptr_79_value ? ghv_48 : _GEN_10460; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10462 = 8'h31 == new_ptr_79_value ? ghv_49 : _GEN_10461; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10463 = 8'h32 == new_ptr_79_value ? ghv_50 : _GEN_10462; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10464 = 8'h33 == new_ptr_79_value ? ghv_51 : _GEN_10463; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10465 = 8'h34 == new_ptr_79_value ? ghv_52 : _GEN_10464; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10466 = 8'h35 == new_ptr_79_value ? ghv_53 : _GEN_10465; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10467 = 8'h36 == new_ptr_79_value ? ghv_54 : _GEN_10466; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10468 = 8'h37 == new_ptr_79_value ? ghv_55 : _GEN_10467; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10469 = 8'h38 == new_ptr_79_value ? ghv_56 : _GEN_10468; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10470 = 8'h39 == new_ptr_79_value ? ghv_57 : _GEN_10469; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10471 = 8'h3a == new_ptr_79_value ? ghv_58 : _GEN_10470; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10472 = 8'h3b == new_ptr_79_value ? ghv_59 : _GEN_10471; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10473 = 8'h3c == new_ptr_79_value ? ghv_60 : _GEN_10472; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10474 = 8'h3d == new_ptr_79_value ? ghv_61 : _GEN_10473; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10475 = 8'h3e == new_ptr_79_value ? ghv_62 : _GEN_10474; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10476 = 8'h3f == new_ptr_79_value ? ghv_63 : _GEN_10475; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10477 = 8'h40 == new_ptr_79_value ? ghv_64 : _GEN_10476; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10478 = 8'h41 == new_ptr_79_value ? ghv_65 : _GEN_10477; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10479 = 8'h42 == new_ptr_79_value ? ghv_66 : _GEN_10478; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10480 = 8'h43 == new_ptr_79_value ? ghv_67 : _GEN_10479; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10481 = 8'h44 == new_ptr_79_value ? ghv_68 : _GEN_10480; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10482 = 8'h45 == new_ptr_79_value ? ghv_69 : _GEN_10481; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10483 = 8'h46 == new_ptr_79_value ? ghv_70 : _GEN_10482; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10484 = 8'h47 == new_ptr_79_value ? ghv_71 : _GEN_10483; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10485 = 8'h48 == new_ptr_79_value ? ghv_72 : _GEN_10484; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10486 = 8'h49 == new_ptr_79_value ? ghv_73 : _GEN_10485; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10487 = 8'h4a == new_ptr_79_value ? ghv_74 : _GEN_10486; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10488 = 8'h4b == new_ptr_79_value ? ghv_75 : _GEN_10487; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10489 = 8'h4c == new_ptr_79_value ? ghv_76 : _GEN_10488; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10490 = 8'h4d == new_ptr_79_value ? ghv_77 : _GEN_10489; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10491 = 8'h4e == new_ptr_79_value ? ghv_78 : _GEN_10490; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10492 = 8'h4f == new_ptr_79_value ? ghv_79 : _GEN_10491; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10493 = 8'h50 == new_ptr_79_value ? ghv_80 : _GEN_10492; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10494 = 8'h51 == new_ptr_79_value ? ghv_81 : _GEN_10493; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10495 = 8'h52 == new_ptr_79_value ? ghv_82 : _GEN_10494; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10496 = 8'h53 == new_ptr_79_value ? ghv_83 : _GEN_10495; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10497 = 8'h54 == new_ptr_79_value ? ghv_84 : _GEN_10496; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10498 = 8'h55 == new_ptr_79_value ? ghv_85 : _GEN_10497; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10499 = 8'h56 == new_ptr_79_value ? ghv_86 : _GEN_10498; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10500 = 8'h57 == new_ptr_79_value ? ghv_87 : _GEN_10499; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10501 = 8'h58 == new_ptr_79_value ? ghv_88 : _GEN_10500; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10502 = 8'h59 == new_ptr_79_value ? ghv_89 : _GEN_10501; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10503 = 8'h5a == new_ptr_79_value ? ghv_90 : _GEN_10502; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10504 = 8'h5b == new_ptr_79_value ? ghv_91 : _GEN_10503; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10505 = 8'h5c == new_ptr_79_value ? ghv_92 : _GEN_10504; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10506 = 8'h5d == new_ptr_79_value ? ghv_93 : _GEN_10505; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10507 = 8'h5e == new_ptr_79_value ? ghv_94 : _GEN_10506; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10508 = 8'h5f == new_ptr_79_value ? ghv_95 : _GEN_10507; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10509 = 8'h60 == new_ptr_79_value ? ghv_96 : _GEN_10508; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10510 = 8'h61 == new_ptr_79_value ? ghv_97 : _GEN_10509; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10511 = 8'h62 == new_ptr_79_value ? ghv_98 : _GEN_10510; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10512 = 8'h63 == new_ptr_79_value ? ghv_99 : _GEN_10511; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10513 = 8'h64 == new_ptr_79_value ? ghv_100 : _GEN_10512; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10514 = 8'h65 == new_ptr_79_value ? ghv_101 : _GEN_10513; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10515 = 8'h66 == new_ptr_79_value ? ghv_102 : _GEN_10514; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10516 = 8'h67 == new_ptr_79_value ? ghv_103 : _GEN_10515; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10517 = 8'h68 == new_ptr_79_value ? ghv_104 : _GEN_10516; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10518 = 8'h69 == new_ptr_79_value ? ghv_105 : _GEN_10517; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10519 = 8'h6a == new_ptr_79_value ? ghv_106 : _GEN_10518; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10520 = 8'h6b == new_ptr_79_value ? ghv_107 : _GEN_10519; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10521 = 8'h6c == new_ptr_79_value ? ghv_108 : _GEN_10520; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10522 = 8'h6d == new_ptr_79_value ? ghv_109 : _GEN_10521; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10523 = 8'h6e == new_ptr_79_value ? ghv_110 : _GEN_10522; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10524 = 8'h6f == new_ptr_79_value ? ghv_111 : _GEN_10523; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10525 = 8'h70 == new_ptr_79_value ? ghv_112 : _GEN_10524; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10526 = 8'h71 == new_ptr_79_value ? ghv_113 : _GEN_10525; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10527 = 8'h72 == new_ptr_79_value ? ghv_114 : _GEN_10526; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10528 = 8'h73 == new_ptr_79_value ? ghv_115 : _GEN_10527; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10529 = 8'h74 == new_ptr_79_value ? ghv_116 : _GEN_10528; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10530 = 8'h75 == new_ptr_79_value ? ghv_117 : _GEN_10529; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10531 = 8'h76 == new_ptr_79_value ? ghv_118 : _GEN_10530; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10532 = 8'h77 == new_ptr_79_value ? ghv_119 : _GEN_10531; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10533 = 8'h78 == new_ptr_79_value ? ghv_120 : _GEN_10532; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10534 = 8'h79 == new_ptr_79_value ? ghv_121 : _GEN_10533; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10535 = 8'h7a == new_ptr_79_value ? ghv_122 : _GEN_10534; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10536 = 8'h7b == new_ptr_79_value ? ghv_123 : _GEN_10535; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10537 = 8'h7c == new_ptr_79_value ? ghv_124 : _GEN_10536; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10538 = 8'h7d == new_ptr_79_value ? ghv_125 : _GEN_10537; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10539 = 8'h7e == new_ptr_79_value ? ghv_126 : _GEN_10538; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10540 = 8'h7f == new_ptr_79_value ? ghv_127 : _GEN_10539; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10541 = 8'h80 == new_ptr_79_value ? ghv_128 : _GEN_10540; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10542 = 8'h81 == new_ptr_79_value ? ghv_129 : _GEN_10541; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10543 = 8'h82 == new_ptr_79_value ? ghv_130 : _GEN_10542; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10544 = 8'h83 == new_ptr_79_value ? ghv_131 : _GEN_10543; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10545 = 8'h84 == new_ptr_79_value ? ghv_132 : _GEN_10544; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10546 = 8'h85 == new_ptr_79_value ? ghv_133 : _GEN_10545; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10547 = 8'h86 == new_ptr_79_value ? ghv_134 : _GEN_10546; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10548 = 8'h87 == new_ptr_79_value ? ghv_135 : _GEN_10547; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10549 = 8'h88 == new_ptr_79_value ? ghv_136 : _GEN_10548; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10550 = 8'h89 == new_ptr_79_value ? ghv_137 : _GEN_10549; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10551 = 8'h8a == new_ptr_79_value ? ghv_138 : _GEN_10550; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10552 = 8'h8b == new_ptr_79_value ? ghv_139 : _GEN_10551; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10553 = 8'h8c == new_ptr_79_value ? ghv_140 : _GEN_10552; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10554 = 8'h8d == new_ptr_79_value ? ghv_141 : _GEN_10553; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10555 = 8'h8e == new_ptr_79_value ? ghv_142 : _GEN_10554; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_63_value = _new_ptr_value_T_127[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_10558 = 8'h1 == new_ptr_63_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10559 = 8'h2 == new_ptr_63_value ? ghv_2 : _GEN_10558; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10560 = 8'h3 == new_ptr_63_value ? ghv_3 : _GEN_10559; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10561 = 8'h4 == new_ptr_63_value ? ghv_4 : _GEN_10560; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10562 = 8'h5 == new_ptr_63_value ? ghv_5 : _GEN_10561; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10563 = 8'h6 == new_ptr_63_value ? ghv_6 : _GEN_10562; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10564 = 8'h7 == new_ptr_63_value ? ghv_7 : _GEN_10563; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10565 = 8'h8 == new_ptr_63_value ? ghv_8 : _GEN_10564; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10566 = 8'h9 == new_ptr_63_value ? ghv_9 : _GEN_10565; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10567 = 8'ha == new_ptr_63_value ? ghv_10 : _GEN_10566; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10568 = 8'hb == new_ptr_63_value ? ghv_11 : _GEN_10567; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10569 = 8'hc == new_ptr_63_value ? ghv_12 : _GEN_10568; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10570 = 8'hd == new_ptr_63_value ? ghv_13 : _GEN_10569; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10571 = 8'he == new_ptr_63_value ? ghv_14 : _GEN_10570; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10572 = 8'hf == new_ptr_63_value ? ghv_15 : _GEN_10571; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10573 = 8'h10 == new_ptr_63_value ? ghv_16 : _GEN_10572; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10574 = 8'h11 == new_ptr_63_value ? ghv_17 : _GEN_10573; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10575 = 8'h12 == new_ptr_63_value ? ghv_18 : _GEN_10574; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10576 = 8'h13 == new_ptr_63_value ? ghv_19 : _GEN_10575; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10577 = 8'h14 == new_ptr_63_value ? ghv_20 : _GEN_10576; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10578 = 8'h15 == new_ptr_63_value ? ghv_21 : _GEN_10577; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10579 = 8'h16 == new_ptr_63_value ? ghv_22 : _GEN_10578; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10580 = 8'h17 == new_ptr_63_value ? ghv_23 : _GEN_10579; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10581 = 8'h18 == new_ptr_63_value ? ghv_24 : _GEN_10580; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10582 = 8'h19 == new_ptr_63_value ? ghv_25 : _GEN_10581; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10583 = 8'h1a == new_ptr_63_value ? ghv_26 : _GEN_10582; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10584 = 8'h1b == new_ptr_63_value ? ghv_27 : _GEN_10583; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10585 = 8'h1c == new_ptr_63_value ? ghv_28 : _GEN_10584; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10586 = 8'h1d == new_ptr_63_value ? ghv_29 : _GEN_10585; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10587 = 8'h1e == new_ptr_63_value ? ghv_30 : _GEN_10586; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10588 = 8'h1f == new_ptr_63_value ? ghv_31 : _GEN_10587; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10589 = 8'h20 == new_ptr_63_value ? ghv_32 : _GEN_10588; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10590 = 8'h21 == new_ptr_63_value ? ghv_33 : _GEN_10589; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10591 = 8'h22 == new_ptr_63_value ? ghv_34 : _GEN_10590; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10592 = 8'h23 == new_ptr_63_value ? ghv_35 : _GEN_10591; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10593 = 8'h24 == new_ptr_63_value ? ghv_36 : _GEN_10592; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10594 = 8'h25 == new_ptr_63_value ? ghv_37 : _GEN_10593; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10595 = 8'h26 == new_ptr_63_value ? ghv_38 : _GEN_10594; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10596 = 8'h27 == new_ptr_63_value ? ghv_39 : _GEN_10595; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10597 = 8'h28 == new_ptr_63_value ? ghv_40 : _GEN_10596; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10598 = 8'h29 == new_ptr_63_value ? ghv_41 : _GEN_10597; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10599 = 8'h2a == new_ptr_63_value ? ghv_42 : _GEN_10598; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10600 = 8'h2b == new_ptr_63_value ? ghv_43 : _GEN_10599; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10601 = 8'h2c == new_ptr_63_value ? ghv_44 : _GEN_10600; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10602 = 8'h2d == new_ptr_63_value ? ghv_45 : _GEN_10601; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10603 = 8'h2e == new_ptr_63_value ? ghv_46 : _GEN_10602; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10604 = 8'h2f == new_ptr_63_value ? ghv_47 : _GEN_10603; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10605 = 8'h30 == new_ptr_63_value ? ghv_48 : _GEN_10604; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10606 = 8'h31 == new_ptr_63_value ? ghv_49 : _GEN_10605; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10607 = 8'h32 == new_ptr_63_value ? ghv_50 : _GEN_10606; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10608 = 8'h33 == new_ptr_63_value ? ghv_51 : _GEN_10607; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10609 = 8'h34 == new_ptr_63_value ? ghv_52 : _GEN_10608; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10610 = 8'h35 == new_ptr_63_value ? ghv_53 : _GEN_10609; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10611 = 8'h36 == new_ptr_63_value ? ghv_54 : _GEN_10610; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10612 = 8'h37 == new_ptr_63_value ? ghv_55 : _GEN_10611; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10613 = 8'h38 == new_ptr_63_value ? ghv_56 : _GEN_10612; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10614 = 8'h39 == new_ptr_63_value ? ghv_57 : _GEN_10613; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10615 = 8'h3a == new_ptr_63_value ? ghv_58 : _GEN_10614; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10616 = 8'h3b == new_ptr_63_value ? ghv_59 : _GEN_10615; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10617 = 8'h3c == new_ptr_63_value ? ghv_60 : _GEN_10616; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10618 = 8'h3d == new_ptr_63_value ? ghv_61 : _GEN_10617; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10619 = 8'h3e == new_ptr_63_value ? ghv_62 : _GEN_10618; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10620 = 8'h3f == new_ptr_63_value ? ghv_63 : _GEN_10619; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10621 = 8'h40 == new_ptr_63_value ? ghv_64 : _GEN_10620; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10622 = 8'h41 == new_ptr_63_value ? ghv_65 : _GEN_10621; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10623 = 8'h42 == new_ptr_63_value ? ghv_66 : _GEN_10622; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10624 = 8'h43 == new_ptr_63_value ? ghv_67 : _GEN_10623; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10625 = 8'h44 == new_ptr_63_value ? ghv_68 : _GEN_10624; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10626 = 8'h45 == new_ptr_63_value ? ghv_69 : _GEN_10625; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10627 = 8'h46 == new_ptr_63_value ? ghv_70 : _GEN_10626; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10628 = 8'h47 == new_ptr_63_value ? ghv_71 : _GEN_10627; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10629 = 8'h48 == new_ptr_63_value ? ghv_72 : _GEN_10628; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10630 = 8'h49 == new_ptr_63_value ? ghv_73 : _GEN_10629; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10631 = 8'h4a == new_ptr_63_value ? ghv_74 : _GEN_10630; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10632 = 8'h4b == new_ptr_63_value ? ghv_75 : _GEN_10631; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10633 = 8'h4c == new_ptr_63_value ? ghv_76 : _GEN_10632; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10634 = 8'h4d == new_ptr_63_value ? ghv_77 : _GEN_10633; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10635 = 8'h4e == new_ptr_63_value ? ghv_78 : _GEN_10634; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10636 = 8'h4f == new_ptr_63_value ? ghv_79 : _GEN_10635; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10637 = 8'h50 == new_ptr_63_value ? ghv_80 : _GEN_10636; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10638 = 8'h51 == new_ptr_63_value ? ghv_81 : _GEN_10637; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10639 = 8'h52 == new_ptr_63_value ? ghv_82 : _GEN_10638; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10640 = 8'h53 == new_ptr_63_value ? ghv_83 : _GEN_10639; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10641 = 8'h54 == new_ptr_63_value ? ghv_84 : _GEN_10640; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10642 = 8'h55 == new_ptr_63_value ? ghv_85 : _GEN_10641; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10643 = 8'h56 == new_ptr_63_value ? ghv_86 : _GEN_10642; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10644 = 8'h57 == new_ptr_63_value ? ghv_87 : _GEN_10643; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10645 = 8'h58 == new_ptr_63_value ? ghv_88 : _GEN_10644; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10646 = 8'h59 == new_ptr_63_value ? ghv_89 : _GEN_10645; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10647 = 8'h5a == new_ptr_63_value ? ghv_90 : _GEN_10646; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10648 = 8'h5b == new_ptr_63_value ? ghv_91 : _GEN_10647; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10649 = 8'h5c == new_ptr_63_value ? ghv_92 : _GEN_10648; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10650 = 8'h5d == new_ptr_63_value ? ghv_93 : _GEN_10649; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10651 = 8'h5e == new_ptr_63_value ? ghv_94 : _GEN_10650; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10652 = 8'h5f == new_ptr_63_value ? ghv_95 : _GEN_10651; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10653 = 8'h60 == new_ptr_63_value ? ghv_96 : _GEN_10652; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10654 = 8'h61 == new_ptr_63_value ? ghv_97 : _GEN_10653; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10655 = 8'h62 == new_ptr_63_value ? ghv_98 : _GEN_10654; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10656 = 8'h63 == new_ptr_63_value ? ghv_99 : _GEN_10655; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10657 = 8'h64 == new_ptr_63_value ? ghv_100 : _GEN_10656; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10658 = 8'h65 == new_ptr_63_value ? ghv_101 : _GEN_10657; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10659 = 8'h66 == new_ptr_63_value ? ghv_102 : _GEN_10658; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10660 = 8'h67 == new_ptr_63_value ? ghv_103 : _GEN_10659; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10661 = 8'h68 == new_ptr_63_value ? ghv_104 : _GEN_10660; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10662 = 8'h69 == new_ptr_63_value ? ghv_105 : _GEN_10661; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10663 = 8'h6a == new_ptr_63_value ? ghv_106 : _GEN_10662; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10664 = 8'h6b == new_ptr_63_value ? ghv_107 : _GEN_10663; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10665 = 8'h6c == new_ptr_63_value ? ghv_108 : _GEN_10664; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10666 = 8'h6d == new_ptr_63_value ? ghv_109 : _GEN_10665; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10667 = 8'h6e == new_ptr_63_value ? ghv_110 : _GEN_10666; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10668 = 8'h6f == new_ptr_63_value ? ghv_111 : _GEN_10667; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10669 = 8'h70 == new_ptr_63_value ? ghv_112 : _GEN_10668; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10670 = 8'h71 == new_ptr_63_value ? ghv_113 : _GEN_10669; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10671 = 8'h72 == new_ptr_63_value ? ghv_114 : _GEN_10670; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10672 = 8'h73 == new_ptr_63_value ? ghv_115 : _GEN_10671; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10673 = 8'h74 == new_ptr_63_value ? ghv_116 : _GEN_10672; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10674 = 8'h75 == new_ptr_63_value ? ghv_117 : _GEN_10673; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10675 = 8'h76 == new_ptr_63_value ? ghv_118 : _GEN_10674; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10676 = 8'h77 == new_ptr_63_value ? ghv_119 : _GEN_10675; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10677 = 8'h78 == new_ptr_63_value ? ghv_120 : _GEN_10676; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10678 = 8'h79 == new_ptr_63_value ? ghv_121 : _GEN_10677; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10679 = 8'h7a == new_ptr_63_value ? ghv_122 : _GEN_10678; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10680 = 8'h7b == new_ptr_63_value ? ghv_123 : _GEN_10679; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10681 = 8'h7c == new_ptr_63_value ? ghv_124 : _GEN_10680; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10682 = 8'h7d == new_ptr_63_value ? ghv_125 : _GEN_10681; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10683 = 8'h7e == new_ptr_63_value ? ghv_126 : _GEN_10682; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10684 = 8'h7f == new_ptr_63_value ? ghv_127 : _GEN_10683; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10685 = 8'h80 == new_ptr_63_value ? ghv_128 : _GEN_10684; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10686 = 8'h81 == new_ptr_63_value ? ghv_129 : _GEN_10685; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10687 = 8'h82 == new_ptr_63_value ? ghv_130 : _GEN_10686; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10688 = 8'h83 == new_ptr_63_value ? ghv_131 : _GEN_10687; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10689 = 8'h84 == new_ptr_63_value ? ghv_132 : _GEN_10688; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10690 = 8'h85 == new_ptr_63_value ? ghv_133 : _GEN_10689; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10691 = 8'h86 == new_ptr_63_value ? ghv_134 : _GEN_10690; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10692 = 8'h87 == new_ptr_63_value ? ghv_135 : _GEN_10691; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10693 = 8'h88 == new_ptr_63_value ? ghv_136 : _GEN_10692; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10694 = 8'h89 == new_ptr_63_value ? ghv_137 : _GEN_10693; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10695 = 8'h8a == new_ptr_63_value ? ghv_138 : _GEN_10694; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10696 = 8'h8b == new_ptr_63_value ? ghv_139 : _GEN_10695; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10697 = 8'h8c == new_ptr_63_value ? ghv_140 : _GEN_10696; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10698 = 8'h8d == new_ptr_63_value ? ghv_141 : _GEN_10697; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10699 = 8'h8e == new_ptr_63_value ? ghv_142 : _GEN_10698; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_70_value = _new_ptr_value_T_141[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_10702 = 8'h1 == new_ptr_70_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10703 = 8'h2 == new_ptr_70_value ? ghv_2 : _GEN_10702; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10704 = 8'h3 == new_ptr_70_value ? ghv_3 : _GEN_10703; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10705 = 8'h4 == new_ptr_70_value ? ghv_4 : _GEN_10704; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10706 = 8'h5 == new_ptr_70_value ? ghv_5 : _GEN_10705; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10707 = 8'h6 == new_ptr_70_value ? ghv_6 : _GEN_10706; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10708 = 8'h7 == new_ptr_70_value ? ghv_7 : _GEN_10707; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10709 = 8'h8 == new_ptr_70_value ? ghv_8 : _GEN_10708; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10710 = 8'h9 == new_ptr_70_value ? ghv_9 : _GEN_10709; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10711 = 8'ha == new_ptr_70_value ? ghv_10 : _GEN_10710; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10712 = 8'hb == new_ptr_70_value ? ghv_11 : _GEN_10711; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10713 = 8'hc == new_ptr_70_value ? ghv_12 : _GEN_10712; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10714 = 8'hd == new_ptr_70_value ? ghv_13 : _GEN_10713; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10715 = 8'he == new_ptr_70_value ? ghv_14 : _GEN_10714; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10716 = 8'hf == new_ptr_70_value ? ghv_15 : _GEN_10715; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10717 = 8'h10 == new_ptr_70_value ? ghv_16 : _GEN_10716; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10718 = 8'h11 == new_ptr_70_value ? ghv_17 : _GEN_10717; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10719 = 8'h12 == new_ptr_70_value ? ghv_18 : _GEN_10718; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10720 = 8'h13 == new_ptr_70_value ? ghv_19 : _GEN_10719; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10721 = 8'h14 == new_ptr_70_value ? ghv_20 : _GEN_10720; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10722 = 8'h15 == new_ptr_70_value ? ghv_21 : _GEN_10721; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10723 = 8'h16 == new_ptr_70_value ? ghv_22 : _GEN_10722; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10724 = 8'h17 == new_ptr_70_value ? ghv_23 : _GEN_10723; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10725 = 8'h18 == new_ptr_70_value ? ghv_24 : _GEN_10724; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10726 = 8'h19 == new_ptr_70_value ? ghv_25 : _GEN_10725; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10727 = 8'h1a == new_ptr_70_value ? ghv_26 : _GEN_10726; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10728 = 8'h1b == new_ptr_70_value ? ghv_27 : _GEN_10727; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10729 = 8'h1c == new_ptr_70_value ? ghv_28 : _GEN_10728; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10730 = 8'h1d == new_ptr_70_value ? ghv_29 : _GEN_10729; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10731 = 8'h1e == new_ptr_70_value ? ghv_30 : _GEN_10730; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10732 = 8'h1f == new_ptr_70_value ? ghv_31 : _GEN_10731; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10733 = 8'h20 == new_ptr_70_value ? ghv_32 : _GEN_10732; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10734 = 8'h21 == new_ptr_70_value ? ghv_33 : _GEN_10733; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10735 = 8'h22 == new_ptr_70_value ? ghv_34 : _GEN_10734; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10736 = 8'h23 == new_ptr_70_value ? ghv_35 : _GEN_10735; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10737 = 8'h24 == new_ptr_70_value ? ghv_36 : _GEN_10736; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10738 = 8'h25 == new_ptr_70_value ? ghv_37 : _GEN_10737; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10739 = 8'h26 == new_ptr_70_value ? ghv_38 : _GEN_10738; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10740 = 8'h27 == new_ptr_70_value ? ghv_39 : _GEN_10739; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10741 = 8'h28 == new_ptr_70_value ? ghv_40 : _GEN_10740; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10742 = 8'h29 == new_ptr_70_value ? ghv_41 : _GEN_10741; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10743 = 8'h2a == new_ptr_70_value ? ghv_42 : _GEN_10742; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10744 = 8'h2b == new_ptr_70_value ? ghv_43 : _GEN_10743; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10745 = 8'h2c == new_ptr_70_value ? ghv_44 : _GEN_10744; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10746 = 8'h2d == new_ptr_70_value ? ghv_45 : _GEN_10745; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10747 = 8'h2e == new_ptr_70_value ? ghv_46 : _GEN_10746; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10748 = 8'h2f == new_ptr_70_value ? ghv_47 : _GEN_10747; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10749 = 8'h30 == new_ptr_70_value ? ghv_48 : _GEN_10748; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10750 = 8'h31 == new_ptr_70_value ? ghv_49 : _GEN_10749; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10751 = 8'h32 == new_ptr_70_value ? ghv_50 : _GEN_10750; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10752 = 8'h33 == new_ptr_70_value ? ghv_51 : _GEN_10751; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10753 = 8'h34 == new_ptr_70_value ? ghv_52 : _GEN_10752; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10754 = 8'h35 == new_ptr_70_value ? ghv_53 : _GEN_10753; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10755 = 8'h36 == new_ptr_70_value ? ghv_54 : _GEN_10754; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10756 = 8'h37 == new_ptr_70_value ? ghv_55 : _GEN_10755; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10757 = 8'h38 == new_ptr_70_value ? ghv_56 : _GEN_10756; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10758 = 8'h39 == new_ptr_70_value ? ghv_57 : _GEN_10757; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10759 = 8'h3a == new_ptr_70_value ? ghv_58 : _GEN_10758; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10760 = 8'h3b == new_ptr_70_value ? ghv_59 : _GEN_10759; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10761 = 8'h3c == new_ptr_70_value ? ghv_60 : _GEN_10760; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10762 = 8'h3d == new_ptr_70_value ? ghv_61 : _GEN_10761; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10763 = 8'h3e == new_ptr_70_value ? ghv_62 : _GEN_10762; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10764 = 8'h3f == new_ptr_70_value ? ghv_63 : _GEN_10763; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10765 = 8'h40 == new_ptr_70_value ? ghv_64 : _GEN_10764; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10766 = 8'h41 == new_ptr_70_value ? ghv_65 : _GEN_10765; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10767 = 8'h42 == new_ptr_70_value ? ghv_66 : _GEN_10766; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10768 = 8'h43 == new_ptr_70_value ? ghv_67 : _GEN_10767; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10769 = 8'h44 == new_ptr_70_value ? ghv_68 : _GEN_10768; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10770 = 8'h45 == new_ptr_70_value ? ghv_69 : _GEN_10769; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10771 = 8'h46 == new_ptr_70_value ? ghv_70 : _GEN_10770; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10772 = 8'h47 == new_ptr_70_value ? ghv_71 : _GEN_10771; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10773 = 8'h48 == new_ptr_70_value ? ghv_72 : _GEN_10772; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10774 = 8'h49 == new_ptr_70_value ? ghv_73 : _GEN_10773; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10775 = 8'h4a == new_ptr_70_value ? ghv_74 : _GEN_10774; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10776 = 8'h4b == new_ptr_70_value ? ghv_75 : _GEN_10775; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10777 = 8'h4c == new_ptr_70_value ? ghv_76 : _GEN_10776; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10778 = 8'h4d == new_ptr_70_value ? ghv_77 : _GEN_10777; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10779 = 8'h4e == new_ptr_70_value ? ghv_78 : _GEN_10778; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10780 = 8'h4f == new_ptr_70_value ? ghv_79 : _GEN_10779; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10781 = 8'h50 == new_ptr_70_value ? ghv_80 : _GEN_10780; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10782 = 8'h51 == new_ptr_70_value ? ghv_81 : _GEN_10781; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10783 = 8'h52 == new_ptr_70_value ? ghv_82 : _GEN_10782; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10784 = 8'h53 == new_ptr_70_value ? ghv_83 : _GEN_10783; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10785 = 8'h54 == new_ptr_70_value ? ghv_84 : _GEN_10784; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10786 = 8'h55 == new_ptr_70_value ? ghv_85 : _GEN_10785; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10787 = 8'h56 == new_ptr_70_value ? ghv_86 : _GEN_10786; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10788 = 8'h57 == new_ptr_70_value ? ghv_87 : _GEN_10787; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10789 = 8'h58 == new_ptr_70_value ? ghv_88 : _GEN_10788; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10790 = 8'h59 == new_ptr_70_value ? ghv_89 : _GEN_10789; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10791 = 8'h5a == new_ptr_70_value ? ghv_90 : _GEN_10790; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10792 = 8'h5b == new_ptr_70_value ? ghv_91 : _GEN_10791; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10793 = 8'h5c == new_ptr_70_value ? ghv_92 : _GEN_10792; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10794 = 8'h5d == new_ptr_70_value ? ghv_93 : _GEN_10793; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10795 = 8'h5e == new_ptr_70_value ? ghv_94 : _GEN_10794; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10796 = 8'h5f == new_ptr_70_value ? ghv_95 : _GEN_10795; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10797 = 8'h60 == new_ptr_70_value ? ghv_96 : _GEN_10796; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10798 = 8'h61 == new_ptr_70_value ? ghv_97 : _GEN_10797; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10799 = 8'h62 == new_ptr_70_value ? ghv_98 : _GEN_10798; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10800 = 8'h63 == new_ptr_70_value ? ghv_99 : _GEN_10799; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10801 = 8'h64 == new_ptr_70_value ? ghv_100 : _GEN_10800; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10802 = 8'h65 == new_ptr_70_value ? ghv_101 : _GEN_10801; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10803 = 8'h66 == new_ptr_70_value ? ghv_102 : _GEN_10802; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10804 = 8'h67 == new_ptr_70_value ? ghv_103 : _GEN_10803; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10805 = 8'h68 == new_ptr_70_value ? ghv_104 : _GEN_10804; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10806 = 8'h69 == new_ptr_70_value ? ghv_105 : _GEN_10805; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10807 = 8'h6a == new_ptr_70_value ? ghv_106 : _GEN_10806; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10808 = 8'h6b == new_ptr_70_value ? ghv_107 : _GEN_10807; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10809 = 8'h6c == new_ptr_70_value ? ghv_108 : _GEN_10808; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10810 = 8'h6d == new_ptr_70_value ? ghv_109 : _GEN_10809; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10811 = 8'h6e == new_ptr_70_value ? ghv_110 : _GEN_10810; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10812 = 8'h6f == new_ptr_70_value ? ghv_111 : _GEN_10811; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10813 = 8'h70 == new_ptr_70_value ? ghv_112 : _GEN_10812; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10814 = 8'h71 == new_ptr_70_value ? ghv_113 : _GEN_10813; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10815 = 8'h72 == new_ptr_70_value ? ghv_114 : _GEN_10814; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10816 = 8'h73 == new_ptr_70_value ? ghv_115 : _GEN_10815; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10817 = 8'h74 == new_ptr_70_value ? ghv_116 : _GEN_10816; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10818 = 8'h75 == new_ptr_70_value ? ghv_117 : _GEN_10817; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10819 = 8'h76 == new_ptr_70_value ? ghv_118 : _GEN_10818; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10820 = 8'h77 == new_ptr_70_value ? ghv_119 : _GEN_10819; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10821 = 8'h78 == new_ptr_70_value ? ghv_120 : _GEN_10820; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10822 = 8'h79 == new_ptr_70_value ? ghv_121 : _GEN_10821; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10823 = 8'h7a == new_ptr_70_value ? ghv_122 : _GEN_10822; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10824 = 8'h7b == new_ptr_70_value ? ghv_123 : _GEN_10823; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10825 = 8'h7c == new_ptr_70_value ? ghv_124 : _GEN_10824; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10826 = 8'h7d == new_ptr_70_value ? ghv_125 : _GEN_10825; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10827 = 8'h7e == new_ptr_70_value ? ghv_126 : _GEN_10826; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10828 = 8'h7f == new_ptr_70_value ? ghv_127 : _GEN_10827; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10829 = 8'h80 == new_ptr_70_value ? ghv_128 : _GEN_10828; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10830 = 8'h81 == new_ptr_70_value ? ghv_129 : _GEN_10829; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10831 = 8'h82 == new_ptr_70_value ? ghv_130 : _GEN_10830; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10832 = 8'h83 == new_ptr_70_value ? ghv_131 : _GEN_10831; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10833 = 8'h84 == new_ptr_70_value ? ghv_132 : _GEN_10832; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10834 = 8'h85 == new_ptr_70_value ? ghv_133 : _GEN_10833; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10835 = 8'h86 == new_ptr_70_value ? ghv_134 : _GEN_10834; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10836 = 8'h87 == new_ptr_70_value ? ghv_135 : _GEN_10835; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10837 = 8'h88 == new_ptr_70_value ? ghv_136 : _GEN_10836; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10838 = 8'h89 == new_ptr_70_value ? ghv_137 : _GEN_10837; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10839 = 8'h8a == new_ptr_70_value ? ghv_138 : _GEN_10838; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10840 = 8'h8b == new_ptr_70_value ? ghv_139 : _GEN_10839; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10841 = 8'h8c == new_ptr_70_value ? ghv_140 : _GEN_10840; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10842 = 8'h8d == new_ptr_70_value ? ghv_141 : _GEN_10841; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10843 = 8'h8e == new_ptr_70_value ? ghv_142 : _GEN_10842; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_61_value = _new_ptr_value_T_123[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_10846 = 8'h1 == new_ptr_61_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10847 = 8'h2 == new_ptr_61_value ? ghv_2 : _GEN_10846; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10848 = 8'h3 == new_ptr_61_value ? ghv_3 : _GEN_10847; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10849 = 8'h4 == new_ptr_61_value ? ghv_4 : _GEN_10848; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10850 = 8'h5 == new_ptr_61_value ? ghv_5 : _GEN_10849; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10851 = 8'h6 == new_ptr_61_value ? ghv_6 : _GEN_10850; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10852 = 8'h7 == new_ptr_61_value ? ghv_7 : _GEN_10851; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10853 = 8'h8 == new_ptr_61_value ? ghv_8 : _GEN_10852; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10854 = 8'h9 == new_ptr_61_value ? ghv_9 : _GEN_10853; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10855 = 8'ha == new_ptr_61_value ? ghv_10 : _GEN_10854; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10856 = 8'hb == new_ptr_61_value ? ghv_11 : _GEN_10855; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10857 = 8'hc == new_ptr_61_value ? ghv_12 : _GEN_10856; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10858 = 8'hd == new_ptr_61_value ? ghv_13 : _GEN_10857; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10859 = 8'he == new_ptr_61_value ? ghv_14 : _GEN_10858; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10860 = 8'hf == new_ptr_61_value ? ghv_15 : _GEN_10859; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10861 = 8'h10 == new_ptr_61_value ? ghv_16 : _GEN_10860; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10862 = 8'h11 == new_ptr_61_value ? ghv_17 : _GEN_10861; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10863 = 8'h12 == new_ptr_61_value ? ghv_18 : _GEN_10862; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10864 = 8'h13 == new_ptr_61_value ? ghv_19 : _GEN_10863; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10865 = 8'h14 == new_ptr_61_value ? ghv_20 : _GEN_10864; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10866 = 8'h15 == new_ptr_61_value ? ghv_21 : _GEN_10865; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10867 = 8'h16 == new_ptr_61_value ? ghv_22 : _GEN_10866; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10868 = 8'h17 == new_ptr_61_value ? ghv_23 : _GEN_10867; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10869 = 8'h18 == new_ptr_61_value ? ghv_24 : _GEN_10868; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10870 = 8'h19 == new_ptr_61_value ? ghv_25 : _GEN_10869; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10871 = 8'h1a == new_ptr_61_value ? ghv_26 : _GEN_10870; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10872 = 8'h1b == new_ptr_61_value ? ghv_27 : _GEN_10871; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10873 = 8'h1c == new_ptr_61_value ? ghv_28 : _GEN_10872; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10874 = 8'h1d == new_ptr_61_value ? ghv_29 : _GEN_10873; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10875 = 8'h1e == new_ptr_61_value ? ghv_30 : _GEN_10874; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10876 = 8'h1f == new_ptr_61_value ? ghv_31 : _GEN_10875; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10877 = 8'h20 == new_ptr_61_value ? ghv_32 : _GEN_10876; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10878 = 8'h21 == new_ptr_61_value ? ghv_33 : _GEN_10877; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10879 = 8'h22 == new_ptr_61_value ? ghv_34 : _GEN_10878; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10880 = 8'h23 == new_ptr_61_value ? ghv_35 : _GEN_10879; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10881 = 8'h24 == new_ptr_61_value ? ghv_36 : _GEN_10880; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10882 = 8'h25 == new_ptr_61_value ? ghv_37 : _GEN_10881; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10883 = 8'h26 == new_ptr_61_value ? ghv_38 : _GEN_10882; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10884 = 8'h27 == new_ptr_61_value ? ghv_39 : _GEN_10883; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10885 = 8'h28 == new_ptr_61_value ? ghv_40 : _GEN_10884; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10886 = 8'h29 == new_ptr_61_value ? ghv_41 : _GEN_10885; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10887 = 8'h2a == new_ptr_61_value ? ghv_42 : _GEN_10886; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10888 = 8'h2b == new_ptr_61_value ? ghv_43 : _GEN_10887; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10889 = 8'h2c == new_ptr_61_value ? ghv_44 : _GEN_10888; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10890 = 8'h2d == new_ptr_61_value ? ghv_45 : _GEN_10889; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10891 = 8'h2e == new_ptr_61_value ? ghv_46 : _GEN_10890; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10892 = 8'h2f == new_ptr_61_value ? ghv_47 : _GEN_10891; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10893 = 8'h30 == new_ptr_61_value ? ghv_48 : _GEN_10892; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10894 = 8'h31 == new_ptr_61_value ? ghv_49 : _GEN_10893; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10895 = 8'h32 == new_ptr_61_value ? ghv_50 : _GEN_10894; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10896 = 8'h33 == new_ptr_61_value ? ghv_51 : _GEN_10895; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10897 = 8'h34 == new_ptr_61_value ? ghv_52 : _GEN_10896; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10898 = 8'h35 == new_ptr_61_value ? ghv_53 : _GEN_10897; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10899 = 8'h36 == new_ptr_61_value ? ghv_54 : _GEN_10898; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10900 = 8'h37 == new_ptr_61_value ? ghv_55 : _GEN_10899; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10901 = 8'h38 == new_ptr_61_value ? ghv_56 : _GEN_10900; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10902 = 8'h39 == new_ptr_61_value ? ghv_57 : _GEN_10901; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10903 = 8'h3a == new_ptr_61_value ? ghv_58 : _GEN_10902; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10904 = 8'h3b == new_ptr_61_value ? ghv_59 : _GEN_10903; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10905 = 8'h3c == new_ptr_61_value ? ghv_60 : _GEN_10904; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10906 = 8'h3d == new_ptr_61_value ? ghv_61 : _GEN_10905; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10907 = 8'h3e == new_ptr_61_value ? ghv_62 : _GEN_10906; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10908 = 8'h3f == new_ptr_61_value ? ghv_63 : _GEN_10907; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10909 = 8'h40 == new_ptr_61_value ? ghv_64 : _GEN_10908; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10910 = 8'h41 == new_ptr_61_value ? ghv_65 : _GEN_10909; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10911 = 8'h42 == new_ptr_61_value ? ghv_66 : _GEN_10910; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10912 = 8'h43 == new_ptr_61_value ? ghv_67 : _GEN_10911; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10913 = 8'h44 == new_ptr_61_value ? ghv_68 : _GEN_10912; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10914 = 8'h45 == new_ptr_61_value ? ghv_69 : _GEN_10913; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10915 = 8'h46 == new_ptr_61_value ? ghv_70 : _GEN_10914; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10916 = 8'h47 == new_ptr_61_value ? ghv_71 : _GEN_10915; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10917 = 8'h48 == new_ptr_61_value ? ghv_72 : _GEN_10916; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10918 = 8'h49 == new_ptr_61_value ? ghv_73 : _GEN_10917; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10919 = 8'h4a == new_ptr_61_value ? ghv_74 : _GEN_10918; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10920 = 8'h4b == new_ptr_61_value ? ghv_75 : _GEN_10919; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10921 = 8'h4c == new_ptr_61_value ? ghv_76 : _GEN_10920; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10922 = 8'h4d == new_ptr_61_value ? ghv_77 : _GEN_10921; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10923 = 8'h4e == new_ptr_61_value ? ghv_78 : _GEN_10922; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10924 = 8'h4f == new_ptr_61_value ? ghv_79 : _GEN_10923; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10925 = 8'h50 == new_ptr_61_value ? ghv_80 : _GEN_10924; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10926 = 8'h51 == new_ptr_61_value ? ghv_81 : _GEN_10925; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10927 = 8'h52 == new_ptr_61_value ? ghv_82 : _GEN_10926; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10928 = 8'h53 == new_ptr_61_value ? ghv_83 : _GEN_10927; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10929 = 8'h54 == new_ptr_61_value ? ghv_84 : _GEN_10928; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10930 = 8'h55 == new_ptr_61_value ? ghv_85 : _GEN_10929; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10931 = 8'h56 == new_ptr_61_value ? ghv_86 : _GEN_10930; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10932 = 8'h57 == new_ptr_61_value ? ghv_87 : _GEN_10931; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10933 = 8'h58 == new_ptr_61_value ? ghv_88 : _GEN_10932; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10934 = 8'h59 == new_ptr_61_value ? ghv_89 : _GEN_10933; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10935 = 8'h5a == new_ptr_61_value ? ghv_90 : _GEN_10934; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10936 = 8'h5b == new_ptr_61_value ? ghv_91 : _GEN_10935; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10937 = 8'h5c == new_ptr_61_value ? ghv_92 : _GEN_10936; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10938 = 8'h5d == new_ptr_61_value ? ghv_93 : _GEN_10937; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10939 = 8'h5e == new_ptr_61_value ? ghv_94 : _GEN_10938; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10940 = 8'h5f == new_ptr_61_value ? ghv_95 : _GEN_10939; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10941 = 8'h60 == new_ptr_61_value ? ghv_96 : _GEN_10940; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10942 = 8'h61 == new_ptr_61_value ? ghv_97 : _GEN_10941; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10943 = 8'h62 == new_ptr_61_value ? ghv_98 : _GEN_10942; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10944 = 8'h63 == new_ptr_61_value ? ghv_99 : _GEN_10943; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10945 = 8'h64 == new_ptr_61_value ? ghv_100 : _GEN_10944; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10946 = 8'h65 == new_ptr_61_value ? ghv_101 : _GEN_10945; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10947 = 8'h66 == new_ptr_61_value ? ghv_102 : _GEN_10946; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10948 = 8'h67 == new_ptr_61_value ? ghv_103 : _GEN_10947; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10949 = 8'h68 == new_ptr_61_value ? ghv_104 : _GEN_10948; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10950 = 8'h69 == new_ptr_61_value ? ghv_105 : _GEN_10949; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10951 = 8'h6a == new_ptr_61_value ? ghv_106 : _GEN_10950; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10952 = 8'h6b == new_ptr_61_value ? ghv_107 : _GEN_10951; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10953 = 8'h6c == new_ptr_61_value ? ghv_108 : _GEN_10952; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10954 = 8'h6d == new_ptr_61_value ? ghv_109 : _GEN_10953; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10955 = 8'h6e == new_ptr_61_value ? ghv_110 : _GEN_10954; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10956 = 8'h6f == new_ptr_61_value ? ghv_111 : _GEN_10955; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10957 = 8'h70 == new_ptr_61_value ? ghv_112 : _GEN_10956; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10958 = 8'h71 == new_ptr_61_value ? ghv_113 : _GEN_10957; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10959 = 8'h72 == new_ptr_61_value ? ghv_114 : _GEN_10958; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10960 = 8'h73 == new_ptr_61_value ? ghv_115 : _GEN_10959; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10961 = 8'h74 == new_ptr_61_value ? ghv_116 : _GEN_10960; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10962 = 8'h75 == new_ptr_61_value ? ghv_117 : _GEN_10961; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10963 = 8'h76 == new_ptr_61_value ? ghv_118 : _GEN_10962; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10964 = 8'h77 == new_ptr_61_value ? ghv_119 : _GEN_10963; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10965 = 8'h78 == new_ptr_61_value ? ghv_120 : _GEN_10964; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10966 = 8'h79 == new_ptr_61_value ? ghv_121 : _GEN_10965; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10967 = 8'h7a == new_ptr_61_value ? ghv_122 : _GEN_10966; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10968 = 8'h7b == new_ptr_61_value ? ghv_123 : _GEN_10967; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10969 = 8'h7c == new_ptr_61_value ? ghv_124 : _GEN_10968; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10970 = 8'h7d == new_ptr_61_value ? ghv_125 : _GEN_10969; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10971 = 8'h7e == new_ptr_61_value ? ghv_126 : _GEN_10970; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10972 = 8'h7f == new_ptr_61_value ? ghv_127 : _GEN_10971; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10973 = 8'h80 == new_ptr_61_value ? ghv_128 : _GEN_10972; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10974 = 8'h81 == new_ptr_61_value ? ghv_129 : _GEN_10973; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10975 = 8'h82 == new_ptr_61_value ? ghv_130 : _GEN_10974; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10976 = 8'h83 == new_ptr_61_value ? ghv_131 : _GEN_10975; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10977 = 8'h84 == new_ptr_61_value ? ghv_132 : _GEN_10976; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10978 = 8'h85 == new_ptr_61_value ? ghv_133 : _GEN_10977; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10979 = 8'h86 == new_ptr_61_value ? ghv_134 : _GEN_10978; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10980 = 8'h87 == new_ptr_61_value ? ghv_135 : _GEN_10979; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10981 = 8'h88 == new_ptr_61_value ? ghv_136 : _GEN_10980; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10982 = 8'h89 == new_ptr_61_value ? ghv_137 : _GEN_10981; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10983 = 8'h8a == new_ptr_61_value ? ghv_138 : _GEN_10982; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10984 = 8'h8b == new_ptr_61_value ? ghv_139 : _GEN_10983; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10985 = 8'h8c == new_ptr_61_value ? ghv_140 : _GEN_10984; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10986 = 8'h8d == new_ptr_61_value ? ghv_141 : _GEN_10985; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10987 = 8'h8e == new_ptr_61_value ? ghv_142 : _GEN_10986; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_78_value = _new_ptr_value_T_157[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_10990 = 8'h1 == new_ptr_78_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10991 = 8'h2 == new_ptr_78_value ? ghv_2 : _GEN_10990; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10992 = 8'h3 == new_ptr_78_value ? ghv_3 : _GEN_10991; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10993 = 8'h4 == new_ptr_78_value ? ghv_4 : _GEN_10992; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10994 = 8'h5 == new_ptr_78_value ? ghv_5 : _GEN_10993; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10995 = 8'h6 == new_ptr_78_value ? ghv_6 : _GEN_10994; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10996 = 8'h7 == new_ptr_78_value ? ghv_7 : _GEN_10995; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10997 = 8'h8 == new_ptr_78_value ? ghv_8 : _GEN_10996; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10998 = 8'h9 == new_ptr_78_value ? ghv_9 : _GEN_10997; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_10999 = 8'ha == new_ptr_78_value ? ghv_10 : _GEN_10998; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11000 = 8'hb == new_ptr_78_value ? ghv_11 : _GEN_10999; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11001 = 8'hc == new_ptr_78_value ? ghv_12 : _GEN_11000; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11002 = 8'hd == new_ptr_78_value ? ghv_13 : _GEN_11001; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11003 = 8'he == new_ptr_78_value ? ghv_14 : _GEN_11002; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11004 = 8'hf == new_ptr_78_value ? ghv_15 : _GEN_11003; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11005 = 8'h10 == new_ptr_78_value ? ghv_16 : _GEN_11004; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11006 = 8'h11 == new_ptr_78_value ? ghv_17 : _GEN_11005; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11007 = 8'h12 == new_ptr_78_value ? ghv_18 : _GEN_11006; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11008 = 8'h13 == new_ptr_78_value ? ghv_19 : _GEN_11007; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11009 = 8'h14 == new_ptr_78_value ? ghv_20 : _GEN_11008; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11010 = 8'h15 == new_ptr_78_value ? ghv_21 : _GEN_11009; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11011 = 8'h16 == new_ptr_78_value ? ghv_22 : _GEN_11010; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11012 = 8'h17 == new_ptr_78_value ? ghv_23 : _GEN_11011; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11013 = 8'h18 == new_ptr_78_value ? ghv_24 : _GEN_11012; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11014 = 8'h19 == new_ptr_78_value ? ghv_25 : _GEN_11013; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11015 = 8'h1a == new_ptr_78_value ? ghv_26 : _GEN_11014; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11016 = 8'h1b == new_ptr_78_value ? ghv_27 : _GEN_11015; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11017 = 8'h1c == new_ptr_78_value ? ghv_28 : _GEN_11016; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11018 = 8'h1d == new_ptr_78_value ? ghv_29 : _GEN_11017; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11019 = 8'h1e == new_ptr_78_value ? ghv_30 : _GEN_11018; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11020 = 8'h1f == new_ptr_78_value ? ghv_31 : _GEN_11019; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11021 = 8'h20 == new_ptr_78_value ? ghv_32 : _GEN_11020; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11022 = 8'h21 == new_ptr_78_value ? ghv_33 : _GEN_11021; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11023 = 8'h22 == new_ptr_78_value ? ghv_34 : _GEN_11022; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11024 = 8'h23 == new_ptr_78_value ? ghv_35 : _GEN_11023; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11025 = 8'h24 == new_ptr_78_value ? ghv_36 : _GEN_11024; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11026 = 8'h25 == new_ptr_78_value ? ghv_37 : _GEN_11025; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11027 = 8'h26 == new_ptr_78_value ? ghv_38 : _GEN_11026; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11028 = 8'h27 == new_ptr_78_value ? ghv_39 : _GEN_11027; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11029 = 8'h28 == new_ptr_78_value ? ghv_40 : _GEN_11028; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11030 = 8'h29 == new_ptr_78_value ? ghv_41 : _GEN_11029; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11031 = 8'h2a == new_ptr_78_value ? ghv_42 : _GEN_11030; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11032 = 8'h2b == new_ptr_78_value ? ghv_43 : _GEN_11031; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11033 = 8'h2c == new_ptr_78_value ? ghv_44 : _GEN_11032; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11034 = 8'h2d == new_ptr_78_value ? ghv_45 : _GEN_11033; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11035 = 8'h2e == new_ptr_78_value ? ghv_46 : _GEN_11034; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11036 = 8'h2f == new_ptr_78_value ? ghv_47 : _GEN_11035; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11037 = 8'h30 == new_ptr_78_value ? ghv_48 : _GEN_11036; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11038 = 8'h31 == new_ptr_78_value ? ghv_49 : _GEN_11037; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11039 = 8'h32 == new_ptr_78_value ? ghv_50 : _GEN_11038; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11040 = 8'h33 == new_ptr_78_value ? ghv_51 : _GEN_11039; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11041 = 8'h34 == new_ptr_78_value ? ghv_52 : _GEN_11040; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11042 = 8'h35 == new_ptr_78_value ? ghv_53 : _GEN_11041; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11043 = 8'h36 == new_ptr_78_value ? ghv_54 : _GEN_11042; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11044 = 8'h37 == new_ptr_78_value ? ghv_55 : _GEN_11043; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11045 = 8'h38 == new_ptr_78_value ? ghv_56 : _GEN_11044; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11046 = 8'h39 == new_ptr_78_value ? ghv_57 : _GEN_11045; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11047 = 8'h3a == new_ptr_78_value ? ghv_58 : _GEN_11046; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11048 = 8'h3b == new_ptr_78_value ? ghv_59 : _GEN_11047; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11049 = 8'h3c == new_ptr_78_value ? ghv_60 : _GEN_11048; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11050 = 8'h3d == new_ptr_78_value ? ghv_61 : _GEN_11049; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11051 = 8'h3e == new_ptr_78_value ? ghv_62 : _GEN_11050; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11052 = 8'h3f == new_ptr_78_value ? ghv_63 : _GEN_11051; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11053 = 8'h40 == new_ptr_78_value ? ghv_64 : _GEN_11052; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11054 = 8'h41 == new_ptr_78_value ? ghv_65 : _GEN_11053; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11055 = 8'h42 == new_ptr_78_value ? ghv_66 : _GEN_11054; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11056 = 8'h43 == new_ptr_78_value ? ghv_67 : _GEN_11055; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11057 = 8'h44 == new_ptr_78_value ? ghv_68 : _GEN_11056; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11058 = 8'h45 == new_ptr_78_value ? ghv_69 : _GEN_11057; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11059 = 8'h46 == new_ptr_78_value ? ghv_70 : _GEN_11058; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11060 = 8'h47 == new_ptr_78_value ? ghv_71 : _GEN_11059; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11061 = 8'h48 == new_ptr_78_value ? ghv_72 : _GEN_11060; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11062 = 8'h49 == new_ptr_78_value ? ghv_73 : _GEN_11061; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11063 = 8'h4a == new_ptr_78_value ? ghv_74 : _GEN_11062; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11064 = 8'h4b == new_ptr_78_value ? ghv_75 : _GEN_11063; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11065 = 8'h4c == new_ptr_78_value ? ghv_76 : _GEN_11064; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11066 = 8'h4d == new_ptr_78_value ? ghv_77 : _GEN_11065; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11067 = 8'h4e == new_ptr_78_value ? ghv_78 : _GEN_11066; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11068 = 8'h4f == new_ptr_78_value ? ghv_79 : _GEN_11067; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11069 = 8'h50 == new_ptr_78_value ? ghv_80 : _GEN_11068; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11070 = 8'h51 == new_ptr_78_value ? ghv_81 : _GEN_11069; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11071 = 8'h52 == new_ptr_78_value ? ghv_82 : _GEN_11070; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11072 = 8'h53 == new_ptr_78_value ? ghv_83 : _GEN_11071; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11073 = 8'h54 == new_ptr_78_value ? ghv_84 : _GEN_11072; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11074 = 8'h55 == new_ptr_78_value ? ghv_85 : _GEN_11073; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11075 = 8'h56 == new_ptr_78_value ? ghv_86 : _GEN_11074; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11076 = 8'h57 == new_ptr_78_value ? ghv_87 : _GEN_11075; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11077 = 8'h58 == new_ptr_78_value ? ghv_88 : _GEN_11076; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11078 = 8'h59 == new_ptr_78_value ? ghv_89 : _GEN_11077; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11079 = 8'h5a == new_ptr_78_value ? ghv_90 : _GEN_11078; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11080 = 8'h5b == new_ptr_78_value ? ghv_91 : _GEN_11079; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11081 = 8'h5c == new_ptr_78_value ? ghv_92 : _GEN_11080; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11082 = 8'h5d == new_ptr_78_value ? ghv_93 : _GEN_11081; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11083 = 8'h5e == new_ptr_78_value ? ghv_94 : _GEN_11082; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11084 = 8'h5f == new_ptr_78_value ? ghv_95 : _GEN_11083; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11085 = 8'h60 == new_ptr_78_value ? ghv_96 : _GEN_11084; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11086 = 8'h61 == new_ptr_78_value ? ghv_97 : _GEN_11085; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11087 = 8'h62 == new_ptr_78_value ? ghv_98 : _GEN_11086; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11088 = 8'h63 == new_ptr_78_value ? ghv_99 : _GEN_11087; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11089 = 8'h64 == new_ptr_78_value ? ghv_100 : _GEN_11088; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11090 = 8'h65 == new_ptr_78_value ? ghv_101 : _GEN_11089; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11091 = 8'h66 == new_ptr_78_value ? ghv_102 : _GEN_11090; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11092 = 8'h67 == new_ptr_78_value ? ghv_103 : _GEN_11091; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11093 = 8'h68 == new_ptr_78_value ? ghv_104 : _GEN_11092; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11094 = 8'h69 == new_ptr_78_value ? ghv_105 : _GEN_11093; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11095 = 8'h6a == new_ptr_78_value ? ghv_106 : _GEN_11094; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11096 = 8'h6b == new_ptr_78_value ? ghv_107 : _GEN_11095; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11097 = 8'h6c == new_ptr_78_value ? ghv_108 : _GEN_11096; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11098 = 8'h6d == new_ptr_78_value ? ghv_109 : _GEN_11097; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11099 = 8'h6e == new_ptr_78_value ? ghv_110 : _GEN_11098; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11100 = 8'h6f == new_ptr_78_value ? ghv_111 : _GEN_11099; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11101 = 8'h70 == new_ptr_78_value ? ghv_112 : _GEN_11100; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11102 = 8'h71 == new_ptr_78_value ? ghv_113 : _GEN_11101; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11103 = 8'h72 == new_ptr_78_value ? ghv_114 : _GEN_11102; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11104 = 8'h73 == new_ptr_78_value ? ghv_115 : _GEN_11103; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11105 = 8'h74 == new_ptr_78_value ? ghv_116 : _GEN_11104; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11106 = 8'h75 == new_ptr_78_value ? ghv_117 : _GEN_11105; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11107 = 8'h76 == new_ptr_78_value ? ghv_118 : _GEN_11106; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11108 = 8'h77 == new_ptr_78_value ? ghv_119 : _GEN_11107; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11109 = 8'h78 == new_ptr_78_value ? ghv_120 : _GEN_11108; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11110 = 8'h79 == new_ptr_78_value ? ghv_121 : _GEN_11109; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11111 = 8'h7a == new_ptr_78_value ? ghv_122 : _GEN_11110; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11112 = 8'h7b == new_ptr_78_value ? ghv_123 : _GEN_11111; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11113 = 8'h7c == new_ptr_78_value ? ghv_124 : _GEN_11112; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11114 = 8'h7d == new_ptr_78_value ? ghv_125 : _GEN_11113; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11115 = 8'h7e == new_ptr_78_value ? ghv_126 : _GEN_11114; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11116 = 8'h7f == new_ptr_78_value ? ghv_127 : _GEN_11115; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11117 = 8'h80 == new_ptr_78_value ? ghv_128 : _GEN_11116; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11118 = 8'h81 == new_ptr_78_value ? ghv_129 : _GEN_11117; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11119 = 8'h82 == new_ptr_78_value ? ghv_130 : _GEN_11118; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11120 = 8'h83 == new_ptr_78_value ? ghv_131 : _GEN_11119; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11121 = 8'h84 == new_ptr_78_value ? ghv_132 : _GEN_11120; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11122 = 8'h85 == new_ptr_78_value ? ghv_133 : _GEN_11121; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11123 = 8'h86 == new_ptr_78_value ? ghv_134 : _GEN_11122; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11124 = 8'h87 == new_ptr_78_value ? ghv_135 : _GEN_11123; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11125 = 8'h88 == new_ptr_78_value ? ghv_136 : _GEN_11124; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11126 = 8'h89 == new_ptr_78_value ? ghv_137 : _GEN_11125; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11127 = 8'h8a == new_ptr_78_value ? ghv_138 : _GEN_11126; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11128 = 8'h8b == new_ptr_78_value ? ghv_139 : _GEN_11127; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11129 = 8'h8c == new_ptr_78_value ? ghv_140 : _GEN_11128; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11130 = 8'h8d == new_ptr_78_value ? ghv_141 : _GEN_11129; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11131 = 8'h8e == new_ptr_78_value ? ghv_142 : _GEN_11130; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_71_value = _new_ptr_value_T_143[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_11134 = 8'h1 == new_ptr_71_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11135 = 8'h2 == new_ptr_71_value ? ghv_2 : _GEN_11134; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11136 = 8'h3 == new_ptr_71_value ? ghv_3 : _GEN_11135; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11137 = 8'h4 == new_ptr_71_value ? ghv_4 : _GEN_11136; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11138 = 8'h5 == new_ptr_71_value ? ghv_5 : _GEN_11137; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11139 = 8'h6 == new_ptr_71_value ? ghv_6 : _GEN_11138; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11140 = 8'h7 == new_ptr_71_value ? ghv_7 : _GEN_11139; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11141 = 8'h8 == new_ptr_71_value ? ghv_8 : _GEN_11140; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11142 = 8'h9 == new_ptr_71_value ? ghv_9 : _GEN_11141; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11143 = 8'ha == new_ptr_71_value ? ghv_10 : _GEN_11142; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11144 = 8'hb == new_ptr_71_value ? ghv_11 : _GEN_11143; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11145 = 8'hc == new_ptr_71_value ? ghv_12 : _GEN_11144; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11146 = 8'hd == new_ptr_71_value ? ghv_13 : _GEN_11145; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11147 = 8'he == new_ptr_71_value ? ghv_14 : _GEN_11146; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11148 = 8'hf == new_ptr_71_value ? ghv_15 : _GEN_11147; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11149 = 8'h10 == new_ptr_71_value ? ghv_16 : _GEN_11148; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11150 = 8'h11 == new_ptr_71_value ? ghv_17 : _GEN_11149; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11151 = 8'h12 == new_ptr_71_value ? ghv_18 : _GEN_11150; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11152 = 8'h13 == new_ptr_71_value ? ghv_19 : _GEN_11151; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11153 = 8'h14 == new_ptr_71_value ? ghv_20 : _GEN_11152; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11154 = 8'h15 == new_ptr_71_value ? ghv_21 : _GEN_11153; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11155 = 8'h16 == new_ptr_71_value ? ghv_22 : _GEN_11154; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11156 = 8'h17 == new_ptr_71_value ? ghv_23 : _GEN_11155; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11157 = 8'h18 == new_ptr_71_value ? ghv_24 : _GEN_11156; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11158 = 8'h19 == new_ptr_71_value ? ghv_25 : _GEN_11157; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11159 = 8'h1a == new_ptr_71_value ? ghv_26 : _GEN_11158; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11160 = 8'h1b == new_ptr_71_value ? ghv_27 : _GEN_11159; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11161 = 8'h1c == new_ptr_71_value ? ghv_28 : _GEN_11160; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11162 = 8'h1d == new_ptr_71_value ? ghv_29 : _GEN_11161; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11163 = 8'h1e == new_ptr_71_value ? ghv_30 : _GEN_11162; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11164 = 8'h1f == new_ptr_71_value ? ghv_31 : _GEN_11163; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11165 = 8'h20 == new_ptr_71_value ? ghv_32 : _GEN_11164; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11166 = 8'h21 == new_ptr_71_value ? ghv_33 : _GEN_11165; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11167 = 8'h22 == new_ptr_71_value ? ghv_34 : _GEN_11166; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11168 = 8'h23 == new_ptr_71_value ? ghv_35 : _GEN_11167; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11169 = 8'h24 == new_ptr_71_value ? ghv_36 : _GEN_11168; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11170 = 8'h25 == new_ptr_71_value ? ghv_37 : _GEN_11169; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11171 = 8'h26 == new_ptr_71_value ? ghv_38 : _GEN_11170; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11172 = 8'h27 == new_ptr_71_value ? ghv_39 : _GEN_11171; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11173 = 8'h28 == new_ptr_71_value ? ghv_40 : _GEN_11172; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11174 = 8'h29 == new_ptr_71_value ? ghv_41 : _GEN_11173; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11175 = 8'h2a == new_ptr_71_value ? ghv_42 : _GEN_11174; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11176 = 8'h2b == new_ptr_71_value ? ghv_43 : _GEN_11175; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11177 = 8'h2c == new_ptr_71_value ? ghv_44 : _GEN_11176; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11178 = 8'h2d == new_ptr_71_value ? ghv_45 : _GEN_11177; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11179 = 8'h2e == new_ptr_71_value ? ghv_46 : _GEN_11178; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11180 = 8'h2f == new_ptr_71_value ? ghv_47 : _GEN_11179; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11181 = 8'h30 == new_ptr_71_value ? ghv_48 : _GEN_11180; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11182 = 8'h31 == new_ptr_71_value ? ghv_49 : _GEN_11181; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11183 = 8'h32 == new_ptr_71_value ? ghv_50 : _GEN_11182; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11184 = 8'h33 == new_ptr_71_value ? ghv_51 : _GEN_11183; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11185 = 8'h34 == new_ptr_71_value ? ghv_52 : _GEN_11184; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11186 = 8'h35 == new_ptr_71_value ? ghv_53 : _GEN_11185; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11187 = 8'h36 == new_ptr_71_value ? ghv_54 : _GEN_11186; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11188 = 8'h37 == new_ptr_71_value ? ghv_55 : _GEN_11187; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11189 = 8'h38 == new_ptr_71_value ? ghv_56 : _GEN_11188; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11190 = 8'h39 == new_ptr_71_value ? ghv_57 : _GEN_11189; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11191 = 8'h3a == new_ptr_71_value ? ghv_58 : _GEN_11190; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11192 = 8'h3b == new_ptr_71_value ? ghv_59 : _GEN_11191; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11193 = 8'h3c == new_ptr_71_value ? ghv_60 : _GEN_11192; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11194 = 8'h3d == new_ptr_71_value ? ghv_61 : _GEN_11193; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11195 = 8'h3e == new_ptr_71_value ? ghv_62 : _GEN_11194; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11196 = 8'h3f == new_ptr_71_value ? ghv_63 : _GEN_11195; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11197 = 8'h40 == new_ptr_71_value ? ghv_64 : _GEN_11196; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11198 = 8'h41 == new_ptr_71_value ? ghv_65 : _GEN_11197; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11199 = 8'h42 == new_ptr_71_value ? ghv_66 : _GEN_11198; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11200 = 8'h43 == new_ptr_71_value ? ghv_67 : _GEN_11199; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11201 = 8'h44 == new_ptr_71_value ? ghv_68 : _GEN_11200; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11202 = 8'h45 == new_ptr_71_value ? ghv_69 : _GEN_11201; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11203 = 8'h46 == new_ptr_71_value ? ghv_70 : _GEN_11202; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11204 = 8'h47 == new_ptr_71_value ? ghv_71 : _GEN_11203; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11205 = 8'h48 == new_ptr_71_value ? ghv_72 : _GEN_11204; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11206 = 8'h49 == new_ptr_71_value ? ghv_73 : _GEN_11205; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11207 = 8'h4a == new_ptr_71_value ? ghv_74 : _GEN_11206; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11208 = 8'h4b == new_ptr_71_value ? ghv_75 : _GEN_11207; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11209 = 8'h4c == new_ptr_71_value ? ghv_76 : _GEN_11208; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11210 = 8'h4d == new_ptr_71_value ? ghv_77 : _GEN_11209; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11211 = 8'h4e == new_ptr_71_value ? ghv_78 : _GEN_11210; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11212 = 8'h4f == new_ptr_71_value ? ghv_79 : _GEN_11211; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11213 = 8'h50 == new_ptr_71_value ? ghv_80 : _GEN_11212; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11214 = 8'h51 == new_ptr_71_value ? ghv_81 : _GEN_11213; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11215 = 8'h52 == new_ptr_71_value ? ghv_82 : _GEN_11214; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11216 = 8'h53 == new_ptr_71_value ? ghv_83 : _GEN_11215; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11217 = 8'h54 == new_ptr_71_value ? ghv_84 : _GEN_11216; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11218 = 8'h55 == new_ptr_71_value ? ghv_85 : _GEN_11217; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11219 = 8'h56 == new_ptr_71_value ? ghv_86 : _GEN_11218; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11220 = 8'h57 == new_ptr_71_value ? ghv_87 : _GEN_11219; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11221 = 8'h58 == new_ptr_71_value ? ghv_88 : _GEN_11220; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11222 = 8'h59 == new_ptr_71_value ? ghv_89 : _GEN_11221; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11223 = 8'h5a == new_ptr_71_value ? ghv_90 : _GEN_11222; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11224 = 8'h5b == new_ptr_71_value ? ghv_91 : _GEN_11223; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11225 = 8'h5c == new_ptr_71_value ? ghv_92 : _GEN_11224; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11226 = 8'h5d == new_ptr_71_value ? ghv_93 : _GEN_11225; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11227 = 8'h5e == new_ptr_71_value ? ghv_94 : _GEN_11226; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11228 = 8'h5f == new_ptr_71_value ? ghv_95 : _GEN_11227; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11229 = 8'h60 == new_ptr_71_value ? ghv_96 : _GEN_11228; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11230 = 8'h61 == new_ptr_71_value ? ghv_97 : _GEN_11229; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11231 = 8'h62 == new_ptr_71_value ? ghv_98 : _GEN_11230; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11232 = 8'h63 == new_ptr_71_value ? ghv_99 : _GEN_11231; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11233 = 8'h64 == new_ptr_71_value ? ghv_100 : _GEN_11232; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11234 = 8'h65 == new_ptr_71_value ? ghv_101 : _GEN_11233; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11235 = 8'h66 == new_ptr_71_value ? ghv_102 : _GEN_11234; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11236 = 8'h67 == new_ptr_71_value ? ghv_103 : _GEN_11235; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11237 = 8'h68 == new_ptr_71_value ? ghv_104 : _GEN_11236; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11238 = 8'h69 == new_ptr_71_value ? ghv_105 : _GEN_11237; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11239 = 8'h6a == new_ptr_71_value ? ghv_106 : _GEN_11238; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11240 = 8'h6b == new_ptr_71_value ? ghv_107 : _GEN_11239; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11241 = 8'h6c == new_ptr_71_value ? ghv_108 : _GEN_11240; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11242 = 8'h6d == new_ptr_71_value ? ghv_109 : _GEN_11241; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11243 = 8'h6e == new_ptr_71_value ? ghv_110 : _GEN_11242; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11244 = 8'h6f == new_ptr_71_value ? ghv_111 : _GEN_11243; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11245 = 8'h70 == new_ptr_71_value ? ghv_112 : _GEN_11244; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11246 = 8'h71 == new_ptr_71_value ? ghv_113 : _GEN_11245; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11247 = 8'h72 == new_ptr_71_value ? ghv_114 : _GEN_11246; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11248 = 8'h73 == new_ptr_71_value ? ghv_115 : _GEN_11247; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11249 = 8'h74 == new_ptr_71_value ? ghv_116 : _GEN_11248; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11250 = 8'h75 == new_ptr_71_value ? ghv_117 : _GEN_11249; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11251 = 8'h76 == new_ptr_71_value ? ghv_118 : _GEN_11250; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11252 = 8'h77 == new_ptr_71_value ? ghv_119 : _GEN_11251; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11253 = 8'h78 == new_ptr_71_value ? ghv_120 : _GEN_11252; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11254 = 8'h79 == new_ptr_71_value ? ghv_121 : _GEN_11253; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11255 = 8'h7a == new_ptr_71_value ? ghv_122 : _GEN_11254; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11256 = 8'h7b == new_ptr_71_value ? ghv_123 : _GEN_11255; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11257 = 8'h7c == new_ptr_71_value ? ghv_124 : _GEN_11256; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11258 = 8'h7d == new_ptr_71_value ? ghv_125 : _GEN_11257; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11259 = 8'h7e == new_ptr_71_value ? ghv_126 : _GEN_11258; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11260 = 8'h7f == new_ptr_71_value ? ghv_127 : _GEN_11259; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11261 = 8'h80 == new_ptr_71_value ? ghv_128 : _GEN_11260; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11262 = 8'h81 == new_ptr_71_value ? ghv_129 : _GEN_11261; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11263 = 8'h82 == new_ptr_71_value ? ghv_130 : _GEN_11262; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11264 = 8'h83 == new_ptr_71_value ? ghv_131 : _GEN_11263; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11265 = 8'h84 == new_ptr_71_value ? ghv_132 : _GEN_11264; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11266 = 8'h85 == new_ptr_71_value ? ghv_133 : _GEN_11265; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11267 = 8'h86 == new_ptr_71_value ? ghv_134 : _GEN_11266; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11268 = 8'h87 == new_ptr_71_value ? ghv_135 : _GEN_11267; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11269 = 8'h88 == new_ptr_71_value ? ghv_136 : _GEN_11268; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11270 = 8'h89 == new_ptr_71_value ? ghv_137 : _GEN_11269; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11271 = 8'h8a == new_ptr_71_value ? ghv_138 : _GEN_11270; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11272 = 8'h8b == new_ptr_71_value ? ghv_139 : _GEN_11271; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11273 = 8'h8c == new_ptr_71_value ? ghv_140 : _GEN_11272; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11274 = 8'h8d == new_ptr_71_value ? ghv_141 : _GEN_11273; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11275 = 8'h8e == new_ptr_71_value ? ghv_142 : _GEN_11274; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_67_value = _new_ptr_value_T_135[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_11278 = 8'h1 == new_ptr_67_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11279 = 8'h2 == new_ptr_67_value ? ghv_2 : _GEN_11278; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11280 = 8'h3 == new_ptr_67_value ? ghv_3 : _GEN_11279; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11281 = 8'h4 == new_ptr_67_value ? ghv_4 : _GEN_11280; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11282 = 8'h5 == new_ptr_67_value ? ghv_5 : _GEN_11281; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11283 = 8'h6 == new_ptr_67_value ? ghv_6 : _GEN_11282; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11284 = 8'h7 == new_ptr_67_value ? ghv_7 : _GEN_11283; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11285 = 8'h8 == new_ptr_67_value ? ghv_8 : _GEN_11284; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11286 = 8'h9 == new_ptr_67_value ? ghv_9 : _GEN_11285; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11287 = 8'ha == new_ptr_67_value ? ghv_10 : _GEN_11286; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11288 = 8'hb == new_ptr_67_value ? ghv_11 : _GEN_11287; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11289 = 8'hc == new_ptr_67_value ? ghv_12 : _GEN_11288; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11290 = 8'hd == new_ptr_67_value ? ghv_13 : _GEN_11289; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11291 = 8'he == new_ptr_67_value ? ghv_14 : _GEN_11290; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11292 = 8'hf == new_ptr_67_value ? ghv_15 : _GEN_11291; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11293 = 8'h10 == new_ptr_67_value ? ghv_16 : _GEN_11292; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11294 = 8'h11 == new_ptr_67_value ? ghv_17 : _GEN_11293; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11295 = 8'h12 == new_ptr_67_value ? ghv_18 : _GEN_11294; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11296 = 8'h13 == new_ptr_67_value ? ghv_19 : _GEN_11295; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11297 = 8'h14 == new_ptr_67_value ? ghv_20 : _GEN_11296; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11298 = 8'h15 == new_ptr_67_value ? ghv_21 : _GEN_11297; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11299 = 8'h16 == new_ptr_67_value ? ghv_22 : _GEN_11298; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11300 = 8'h17 == new_ptr_67_value ? ghv_23 : _GEN_11299; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11301 = 8'h18 == new_ptr_67_value ? ghv_24 : _GEN_11300; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11302 = 8'h19 == new_ptr_67_value ? ghv_25 : _GEN_11301; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11303 = 8'h1a == new_ptr_67_value ? ghv_26 : _GEN_11302; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11304 = 8'h1b == new_ptr_67_value ? ghv_27 : _GEN_11303; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11305 = 8'h1c == new_ptr_67_value ? ghv_28 : _GEN_11304; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11306 = 8'h1d == new_ptr_67_value ? ghv_29 : _GEN_11305; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11307 = 8'h1e == new_ptr_67_value ? ghv_30 : _GEN_11306; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11308 = 8'h1f == new_ptr_67_value ? ghv_31 : _GEN_11307; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11309 = 8'h20 == new_ptr_67_value ? ghv_32 : _GEN_11308; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11310 = 8'h21 == new_ptr_67_value ? ghv_33 : _GEN_11309; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11311 = 8'h22 == new_ptr_67_value ? ghv_34 : _GEN_11310; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11312 = 8'h23 == new_ptr_67_value ? ghv_35 : _GEN_11311; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11313 = 8'h24 == new_ptr_67_value ? ghv_36 : _GEN_11312; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11314 = 8'h25 == new_ptr_67_value ? ghv_37 : _GEN_11313; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11315 = 8'h26 == new_ptr_67_value ? ghv_38 : _GEN_11314; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11316 = 8'h27 == new_ptr_67_value ? ghv_39 : _GEN_11315; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11317 = 8'h28 == new_ptr_67_value ? ghv_40 : _GEN_11316; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11318 = 8'h29 == new_ptr_67_value ? ghv_41 : _GEN_11317; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11319 = 8'h2a == new_ptr_67_value ? ghv_42 : _GEN_11318; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11320 = 8'h2b == new_ptr_67_value ? ghv_43 : _GEN_11319; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11321 = 8'h2c == new_ptr_67_value ? ghv_44 : _GEN_11320; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11322 = 8'h2d == new_ptr_67_value ? ghv_45 : _GEN_11321; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11323 = 8'h2e == new_ptr_67_value ? ghv_46 : _GEN_11322; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11324 = 8'h2f == new_ptr_67_value ? ghv_47 : _GEN_11323; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11325 = 8'h30 == new_ptr_67_value ? ghv_48 : _GEN_11324; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11326 = 8'h31 == new_ptr_67_value ? ghv_49 : _GEN_11325; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11327 = 8'h32 == new_ptr_67_value ? ghv_50 : _GEN_11326; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11328 = 8'h33 == new_ptr_67_value ? ghv_51 : _GEN_11327; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11329 = 8'h34 == new_ptr_67_value ? ghv_52 : _GEN_11328; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11330 = 8'h35 == new_ptr_67_value ? ghv_53 : _GEN_11329; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11331 = 8'h36 == new_ptr_67_value ? ghv_54 : _GEN_11330; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11332 = 8'h37 == new_ptr_67_value ? ghv_55 : _GEN_11331; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11333 = 8'h38 == new_ptr_67_value ? ghv_56 : _GEN_11332; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11334 = 8'h39 == new_ptr_67_value ? ghv_57 : _GEN_11333; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11335 = 8'h3a == new_ptr_67_value ? ghv_58 : _GEN_11334; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11336 = 8'h3b == new_ptr_67_value ? ghv_59 : _GEN_11335; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11337 = 8'h3c == new_ptr_67_value ? ghv_60 : _GEN_11336; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11338 = 8'h3d == new_ptr_67_value ? ghv_61 : _GEN_11337; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11339 = 8'h3e == new_ptr_67_value ? ghv_62 : _GEN_11338; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11340 = 8'h3f == new_ptr_67_value ? ghv_63 : _GEN_11339; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11341 = 8'h40 == new_ptr_67_value ? ghv_64 : _GEN_11340; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11342 = 8'h41 == new_ptr_67_value ? ghv_65 : _GEN_11341; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11343 = 8'h42 == new_ptr_67_value ? ghv_66 : _GEN_11342; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11344 = 8'h43 == new_ptr_67_value ? ghv_67 : _GEN_11343; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11345 = 8'h44 == new_ptr_67_value ? ghv_68 : _GEN_11344; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11346 = 8'h45 == new_ptr_67_value ? ghv_69 : _GEN_11345; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11347 = 8'h46 == new_ptr_67_value ? ghv_70 : _GEN_11346; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11348 = 8'h47 == new_ptr_67_value ? ghv_71 : _GEN_11347; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11349 = 8'h48 == new_ptr_67_value ? ghv_72 : _GEN_11348; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11350 = 8'h49 == new_ptr_67_value ? ghv_73 : _GEN_11349; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11351 = 8'h4a == new_ptr_67_value ? ghv_74 : _GEN_11350; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11352 = 8'h4b == new_ptr_67_value ? ghv_75 : _GEN_11351; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11353 = 8'h4c == new_ptr_67_value ? ghv_76 : _GEN_11352; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11354 = 8'h4d == new_ptr_67_value ? ghv_77 : _GEN_11353; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11355 = 8'h4e == new_ptr_67_value ? ghv_78 : _GEN_11354; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11356 = 8'h4f == new_ptr_67_value ? ghv_79 : _GEN_11355; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11357 = 8'h50 == new_ptr_67_value ? ghv_80 : _GEN_11356; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11358 = 8'h51 == new_ptr_67_value ? ghv_81 : _GEN_11357; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11359 = 8'h52 == new_ptr_67_value ? ghv_82 : _GEN_11358; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11360 = 8'h53 == new_ptr_67_value ? ghv_83 : _GEN_11359; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11361 = 8'h54 == new_ptr_67_value ? ghv_84 : _GEN_11360; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11362 = 8'h55 == new_ptr_67_value ? ghv_85 : _GEN_11361; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11363 = 8'h56 == new_ptr_67_value ? ghv_86 : _GEN_11362; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11364 = 8'h57 == new_ptr_67_value ? ghv_87 : _GEN_11363; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11365 = 8'h58 == new_ptr_67_value ? ghv_88 : _GEN_11364; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11366 = 8'h59 == new_ptr_67_value ? ghv_89 : _GEN_11365; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11367 = 8'h5a == new_ptr_67_value ? ghv_90 : _GEN_11366; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11368 = 8'h5b == new_ptr_67_value ? ghv_91 : _GEN_11367; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11369 = 8'h5c == new_ptr_67_value ? ghv_92 : _GEN_11368; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11370 = 8'h5d == new_ptr_67_value ? ghv_93 : _GEN_11369; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11371 = 8'h5e == new_ptr_67_value ? ghv_94 : _GEN_11370; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11372 = 8'h5f == new_ptr_67_value ? ghv_95 : _GEN_11371; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11373 = 8'h60 == new_ptr_67_value ? ghv_96 : _GEN_11372; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11374 = 8'h61 == new_ptr_67_value ? ghv_97 : _GEN_11373; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11375 = 8'h62 == new_ptr_67_value ? ghv_98 : _GEN_11374; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11376 = 8'h63 == new_ptr_67_value ? ghv_99 : _GEN_11375; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11377 = 8'h64 == new_ptr_67_value ? ghv_100 : _GEN_11376; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11378 = 8'h65 == new_ptr_67_value ? ghv_101 : _GEN_11377; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11379 = 8'h66 == new_ptr_67_value ? ghv_102 : _GEN_11378; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11380 = 8'h67 == new_ptr_67_value ? ghv_103 : _GEN_11379; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11381 = 8'h68 == new_ptr_67_value ? ghv_104 : _GEN_11380; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11382 = 8'h69 == new_ptr_67_value ? ghv_105 : _GEN_11381; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11383 = 8'h6a == new_ptr_67_value ? ghv_106 : _GEN_11382; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11384 = 8'h6b == new_ptr_67_value ? ghv_107 : _GEN_11383; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11385 = 8'h6c == new_ptr_67_value ? ghv_108 : _GEN_11384; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11386 = 8'h6d == new_ptr_67_value ? ghv_109 : _GEN_11385; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11387 = 8'h6e == new_ptr_67_value ? ghv_110 : _GEN_11386; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11388 = 8'h6f == new_ptr_67_value ? ghv_111 : _GEN_11387; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11389 = 8'h70 == new_ptr_67_value ? ghv_112 : _GEN_11388; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11390 = 8'h71 == new_ptr_67_value ? ghv_113 : _GEN_11389; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11391 = 8'h72 == new_ptr_67_value ? ghv_114 : _GEN_11390; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11392 = 8'h73 == new_ptr_67_value ? ghv_115 : _GEN_11391; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11393 = 8'h74 == new_ptr_67_value ? ghv_116 : _GEN_11392; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11394 = 8'h75 == new_ptr_67_value ? ghv_117 : _GEN_11393; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11395 = 8'h76 == new_ptr_67_value ? ghv_118 : _GEN_11394; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11396 = 8'h77 == new_ptr_67_value ? ghv_119 : _GEN_11395; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11397 = 8'h78 == new_ptr_67_value ? ghv_120 : _GEN_11396; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11398 = 8'h79 == new_ptr_67_value ? ghv_121 : _GEN_11397; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11399 = 8'h7a == new_ptr_67_value ? ghv_122 : _GEN_11398; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11400 = 8'h7b == new_ptr_67_value ? ghv_123 : _GEN_11399; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11401 = 8'h7c == new_ptr_67_value ? ghv_124 : _GEN_11400; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11402 = 8'h7d == new_ptr_67_value ? ghv_125 : _GEN_11401; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11403 = 8'h7e == new_ptr_67_value ? ghv_126 : _GEN_11402; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11404 = 8'h7f == new_ptr_67_value ? ghv_127 : _GEN_11403; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11405 = 8'h80 == new_ptr_67_value ? ghv_128 : _GEN_11404; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11406 = 8'h81 == new_ptr_67_value ? ghv_129 : _GEN_11405; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11407 = 8'h82 == new_ptr_67_value ? ghv_130 : _GEN_11406; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11408 = 8'h83 == new_ptr_67_value ? ghv_131 : _GEN_11407; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11409 = 8'h84 == new_ptr_67_value ? ghv_132 : _GEN_11408; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11410 = 8'h85 == new_ptr_67_value ? ghv_133 : _GEN_11409; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11411 = 8'h86 == new_ptr_67_value ? ghv_134 : _GEN_11410; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11412 = 8'h87 == new_ptr_67_value ? ghv_135 : _GEN_11411; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11413 = 8'h88 == new_ptr_67_value ? ghv_136 : _GEN_11412; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11414 = 8'h89 == new_ptr_67_value ? ghv_137 : _GEN_11413; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11415 = 8'h8a == new_ptr_67_value ? ghv_138 : _GEN_11414; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11416 = 8'h8b == new_ptr_67_value ? ghv_139 : _GEN_11415; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11417 = 8'h8c == new_ptr_67_value ? ghv_140 : _GEN_11416; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11418 = 8'h8d == new_ptr_67_value ? ghv_141 : _GEN_11417; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11419 = 8'h8e == new_ptr_67_value ? ghv_142 : _GEN_11418; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_65_value = _new_ptr_value_T_131[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_11422 = 8'h1 == new_ptr_65_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11423 = 8'h2 == new_ptr_65_value ? ghv_2 : _GEN_11422; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11424 = 8'h3 == new_ptr_65_value ? ghv_3 : _GEN_11423; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11425 = 8'h4 == new_ptr_65_value ? ghv_4 : _GEN_11424; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11426 = 8'h5 == new_ptr_65_value ? ghv_5 : _GEN_11425; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11427 = 8'h6 == new_ptr_65_value ? ghv_6 : _GEN_11426; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11428 = 8'h7 == new_ptr_65_value ? ghv_7 : _GEN_11427; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11429 = 8'h8 == new_ptr_65_value ? ghv_8 : _GEN_11428; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11430 = 8'h9 == new_ptr_65_value ? ghv_9 : _GEN_11429; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11431 = 8'ha == new_ptr_65_value ? ghv_10 : _GEN_11430; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11432 = 8'hb == new_ptr_65_value ? ghv_11 : _GEN_11431; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11433 = 8'hc == new_ptr_65_value ? ghv_12 : _GEN_11432; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11434 = 8'hd == new_ptr_65_value ? ghv_13 : _GEN_11433; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11435 = 8'he == new_ptr_65_value ? ghv_14 : _GEN_11434; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11436 = 8'hf == new_ptr_65_value ? ghv_15 : _GEN_11435; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11437 = 8'h10 == new_ptr_65_value ? ghv_16 : _GEN_11436; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11438 = 8'h11 == new_ptr_65_value ? ghv_17 : _GEN_11437; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11439 = 8'h12 == new_ptr_65_value ? ghv_18 : _GEN_11438; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11440 = 8'h13 == new_ptr_65_value ? ghv_19 : _GEN_11439; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11441 = 8'h14 == new_ptr_65_value ? ghv_20 : _GEN_11440; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11442 = 8'h15 == new_ptr_65_value ? ghv_21 : _GEN_11441; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11443 = 8'h16 == new_ptr_65_value ? ghv_22 : _GEN_11442; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11444 = 8'h17 == new_ptr_65_value ? ghv_23 : _GEN_11443; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11445 = 8'h18 == new_ptr_65_value ? ghv_24 : _GEN_11444; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11446 = 8'h19 == new_ptr_65_value ? ghv_25 : _GEN_11445; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11447 = 8'h1a == new_ptr_65_value ? ghv_26 : _GEN_11446; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11448 = 8'h1b == new_ptr_65_value ? ghv_27 : _GEN_11447; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11449 = 8'h1c == new_ptr_65_value ? ghv_28 : _GEN_11448; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11450 = 8'h1d == new_ptr_65_value ? ghv_29 : _GEN_11449; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11451 = 8'h1e == new_ptr_65_value ? ghv_30 : _GEN_11450; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11452 = 8'h1f == new_ptr_65_value ? ghv_31 : _GEN_11451; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11453 = 8'h20 == new_ptr_65_value ? ghv_32 : _GEN_11452; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11454 = 8'h21 == new_ptr_65_value ? ghv_33 : _GEN_11453; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11455 = 8'h22 == new_ptr_65_value ? ghv_34 : _GEN_11454; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11456 = 8'h23 == new_ptr_65_value ? ghv_35 : _GEN_11455; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11457 = 8'h24 == new_ptr_65_value ? ghv_36 : _GEN_11456; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11458 = 8'h25 == new_ptr_65_value ? ghv_37 : _GEN_11457; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11459 = 8'h26 == new_ptr_65_value ? ghv_38 : _GEN_11458; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11460 = 8'h27 == new_ptr_65_value ? ghv_39 : _GEN_11459; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11461 = 8'h28 == new_ptr_65_value ? ghv_40 : _GEN_11460; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11462 = 8'h29 == new_ptr_65_value ? ghv_41 : _GEN_11461; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11463 = 8'h2a == new_ptr_65_value ? ghv_42 : _GEN_11462; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11464 = 8'h2b == new_ptr_65_value ? ghv_43 : _GEN_11463; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11465 = 8'h2c == new_ptr_65_value ? ghv_44 : _GEN_11464; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11466 = 8'h2d == new_ptr_65_value ? ghv_45 : _GEN_11465; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11467 = 8'h2e == new_ptr_65_value ? ghv_46 : _GEN_11466; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11468 = 8'h2f == new_ptr_65_value ? ghv_47 : _GEN_11467; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11469 = 8'h30 == new_ptr_65_value ? ghv_48 : _GEN_11468; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11470 = 8'h31 == new_ptr_65_value ? ghv_49 : _GEN_11469; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11471 = 8'h32 == new_ptr_65_value ? ghv_50 : _GEN_11470; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11472 = 8'h33 == new_ptr_65_value ? ghv_51 : _GEN_11471; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11473 = 8'h34 == new_ptr_65_value ? ghv_52 : _GEN_11472; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11474 = 8'h35 == new_ptr_65_value ? ghv_53 : _GEN_11473; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11475 = 8'h36 == new_ptr_65_value ? ghv_54 : _GEN_11474; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11476 = 8'h37 == new_ptr_65_value ? ghv_55 : _GEN_11475; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11477 = 8'h38 == new_ptr_65_value ? ghv_56 : _GEN_11476; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11478 = 8'h39 == new_ptr_65_value ? ghv_57 : _GEN_11477; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11479 = 8'h3a == new_ptr_65_value ? ghv_58 : _GEN_11478; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11480 = 8'h3b == new_ptr_65_value ? ghv_59 : _GEN_11479; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11481 = 8'h3c == new_ptr_65_value ? ghv_60 : _GEN_11480; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11482 = 8'h3d == new_ptr_65_value ? ghv_61 : _GEN_11481; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11483 = 8'h3e == new_ptr_65_value ? ghv_62 : _GEN_11482; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11484 = 8'h3f == new_ptr_65_value ? ghv_63 : _GEN_11483; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11485 = 8'h40 == new_ptr_65_value ? ghv_64 : _GEN_11484; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11486 = 8'h41 == new_ptr_65_value ? ghv_65 : _GEN_11485; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11487 = 8'h42 == new_ptr_65_value ? ghv_66 : _GEN_11486; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11488 = 8'h43 == new_ptr_65_value ? ghv_67 : _GEN_11487; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11489 = 8'h44 == new_ptr_65_value ? ghv_68 : _GEN_11488; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11490 = 8'h45 == new_ptr_65_value ? ghv_69 : _GEN_11489; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11491 = 8'h46 == new_ptr_65_value ? ghv_70 : _GEN_11490; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11492 = 8'h47 == new_ptr_65_value ? ghv_71 : _GEN_11491; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11493 = 8'h48 == new_ptr_65_value ? ghv_72 : _GEN_11492; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11494 = 8'h49 == new_ptr_65_value ? ghv_73 : _GEN_11493; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11495 = 8'h4a == new_ptr_65_value ? ghv_74 : _GEN_11494; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11496 = 8'h4b == new_ptr_65_value ? ghv_75 : _GEN_11495; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11497 = 8'h4c == new_ptr_65_value ? ghv_76 : _GEN_11496; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11498 = 8'h4d == new_ptr_65_value ? ghv_77 : _GEN_11497; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11499 = 8'h4e == new_ptr_65_value ? ghv_78 : _GEN_11498; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11500 = 8'h4f == new_ptr_65_value ? ghv_79 : _GEN_11499; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11501 = 8'h50 == new_ptr_65_value ? ghv_80 : _GEN_11500; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11502 = 8'h51 == new_ptr_65_value ? ghv_81 : _GEN_11501; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11503 = 8'h52 == new_ptr_65_value ? ghv_82 : _GEN_11502; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11504 = 8'h53 == new_ptr_65_value ? ghv_83 : _GEN_11503; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11505 = 8'h54 == new_ptr_65_value ? ghv_84 : _GEN_11504; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11506 = 8'h55 == new_ptr_65_value ? ghv_85 : _GEN_11505; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11507 = 8'h56 == new_ptr_65_value ? ghv_86 : _GEN_11506; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11508 = 8'h57 == new_ptr_65_value ? ghv_87 : _GEN_11507; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11509 = 8'h58 == new_ptr_65_value ? ghv_88 : _GEN_11508; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11510 = 8'h59 == new_ptr_65_value ? ghv_89 : _GEN_11509; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11511 = 8'h5a == new_ptr_65_value ? ghv_90 : _GEN_11510; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11512 = 8'h5b == new_ptr_65_value ? ghv_91 : _GEN_11511; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11513 = 8'h5c == new_ptr_65_value ? ghv_92 : _GEN_11512; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11514 = 8'h5d == new_ptr_65_value ? ghv_93 : _GEN_11513; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11515 = 8'h5e == new_ptr_65_value ? ghv_94 : _GEN_11514; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11516 = 8'h5f == new_ptr_65_value ? ghv_95 : _GEN_11515; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11517 = 8'h60 == new_ptr_65_value ? ghv_96 : _GEN_11516; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11518 = 8'h61 == new_ptr_65_value ? ghv_97 : _GEN_11517; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11519 = 8'h62 == new_ptr_65_value ? ghv_98 : _GEN_11518; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11520 = 8'h63 == new_ptr_65_value ? ghv_99 : _GEN_11519; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11521 = 8'h64 == new_ptr_65_value ? ghv_100 : _GEN_11520; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11522 = 8'h65 == new_ptr_65_value ? ghv_101 : _GEN_11521; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11523 = 8'h66 == new_ptr_65_value ? ghv_102 : _GEN_11522; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11524 = 8'h67 == new_ptr_65_value ? ghv_103 : _GEN_11523; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11525 = 8'h68 == new_ptr_65_value ? ghv_104 : _GEN_11524; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11526 = 8'h69 == new_ptr_65_value ? ghv_105 : _GEN_11525; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11527 = 8'h6a == new_ptr_65_value ? ghv_106 : _GEN_11526; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11528 = 8'h6b == new_ptr_65_value ? ghv_107 : _GEN_11527; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11529 = 8'h6c == new_ptr_65_value ? ghv_108 : _GEN_11528; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11530 = 8'h6d == new_ptr_65_value ? ghv_109 : _GEN_11529; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11531 = 8'h6e == new_ptr_65_value ? ghv_110 : _GEN_11530; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11532 = 8'h6f == new_ptr_65_value ? ghv_111 : _GEN_11531; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11533 = 8'h70 == new_ptr_65_value ? ghv_112 : _GEN_11532; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11534 = 8'h71 == new_ptr_65_value ? ghv_113 : _GEN_11533; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11535 = 8'h72 == new_ptr_65_value ? ghv_114 : _GEN_11534; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11536 = 8'h73 == new_ptr_65_value ? ghv_115 : _GEN_11535; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11537 = 8'h74 == new_ptr_65_value ? ghv_116 : _GEN_11536; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11538 = 8'h75 == new_ptr_65_value ? ghv_117 : _GEN_11537; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11539 = 8'h76 == new_ptr_65_value ? ghv_118 : _GEN_11538; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11540 = 8'h77 == new_ptr_65_value ? ghv_119 : _GEN_11539; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11541 = 8'h78 == new_ptr_65_value ? ghv_120 : _GEN_11540; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11542 = 8'h79 == new_ptr_65_value ? ghv_121 : _GEN_11541; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11543 = 8'h7a == new_ptr_65_value ? ghv_122 : _GEN_11542; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11544 = 8'h7b == new_ptr_65_value ? ghv_123 : _GEN_11543; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11545 = 8'h7c == new_ptr_65_value ? ghv_124 : _GEN_11544; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11546 = 8'h7d == new_ptr_65_value ? ghv_125 : _GEN_11545; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11547 = 8'h7e == new_ptr_65_value ? ghv_126 : _GEN_11546; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11548 = 8'h7f == new_ptr_65_value ? ghv_127 : _GEN_11547; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11549 = 8'h80 == new_ptr_65_value ? ghv_128 : _GEN_11548; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11550 = 8'h81 == new_ptr_65_value ? ghv_129 : _GEN_11549; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11551 = 8'h82 == new_ptr_65_value ? ghv_130 : _GEN_11550; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11552 = 8'h83 == new_ptr_65_value ? ghv_131 : _GEN_11551; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11553 = 8'h84 == new_ptr_65_value ? ghv_132 : _GEN_11552; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11554 = 8'h85 == new_ptr_65_value ? ghv_133 : _GEN_11553; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11555 = 8'h86 == new_ptr_65_value ? ghv_134 : _GEN_11554; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11556 = 8'h87 == new_ptr_65_value ? ghv_135 : _GEN_11555; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11557 = 8'h88 == new_ptr_65_value ? ghv_136 : _GEN_11556; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11558 = 8'h89 == new_ptr_65_value ? ghv_137 : _GEN_11557; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11559 = 8'h8a == new_ptr_65_value ? ghv_138 : _GEN_11558; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11560 = 8'h8b == new_ptr_65_value ? ghv_139 : _GEN_11559; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11561 = 8'h8c == new_ptr_65_value ? ghv_140 : _GEN_11560; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11562 = 8'h8d == new_ptr_65_value ? ghv_141 : _GEN_11561; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11563 = 8'h8e == new_ptr_65_value ? ghv_142 : _GEN_11562; // @[FrontendBundle.scala 329:{20,20}]
  wire [7:0] new_ptr_60_value = _new_ptr_value_T_121[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  wire  _GEN_11566 = 8'h1 == new_ptr_60_value ? ghv_1 : ghv_0; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11567 = 8'h2 == new_ptr_60_value ? ghv_2 : _GEN_11566; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11568 = 8'h3 == new_ptr_60_value ? ghv_3 : _GEN_11567; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11569 = 8'h4 == new_ptr_60_value ? ghv_4 : _GEN_11568; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11570 = 8'h5 == new_ptr_60_value ? ghv_5 : _GEN_11569; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11571 = 8'h6 == new_ptr_60_value ? ghv_6 : _GEN_11570; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11572 = 8'h7 == new_ptr_60_value ? ghv_7 : _GEN_11571; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11573 = 8'h8 == new_ptr_60_value ? ghv_8 : _GEN_11572; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11574 = 8'h9 == new_ptr_60_value ? ghv_9 : _GEN_11573; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11575 = 8'ha == new_ptr_60_value ? ghv_10 : _GEN_11574; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11576 = 8'hb == new_ptr_60_value ? ghv_11 : _GEN_11575; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11577 = 8'hc == new_ptr_60_value ? ghv_12 : _GEN_11576; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11578 = 8'hd == new_ptr_60_value ? ghv_13 : _GEN_11577; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11579 = 8'he == new_ptr_60_value ? ghv_14 : _GEN_11578; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11580 = 8'hf == new_ptr_60_value ? ghv_15 : _GEN_11579; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11581 = 8'h10 == new_ptr_60_value ? ghv_16 : _GEN_11580; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11582 = 8'h11 == new_ptr_60_value ? ghv_17 : _GEN_11581; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11583 = 8'h12 == new_ptr_60_value ? ghv_18 : _GEN_11582; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11584 = 8'h13 == new_ptr_60_value ? ghv_19 : _GEN_11583; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11585 = 8'h14 == new_ptr_60_value ? ghv_20 : _GEN_11584; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11586 = 8'h15 == new_ptr_60_value ? ghv_21 : _GEN_11585; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11587 = 8'h16 == new_ptr_60_value ? ghv_22 : _GEN_11586; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11588 = 8'h17 == new_ptr_60_value ? ghv_23 : _GEN_11587; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11589 = 8'h18 == new_ptr_60_value ? ghv_24 : _GEN_11588; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11590 = 8'h19 == new_ptr_60_value ? ghv_25 : _GEN_11589; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11591 = 8'h1a == new_ptr_60_value ? ghv_26 : _GEN_11590; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11592 = 8'h1b == new_ptr_60_value ? ghv_27 : _GEN_11591; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11593 = 8'h1c == new_ptr_60_value ? ghv_28 : _GEN_11592; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11594 = 8'h1d == new_ptr_60_value ? ghv_29 : _GEN_11593; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11595 = 8'h1e == new_ptr_60_value ? ghv_30 : _GEN_11594; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11596 = 8'h1f == new_ptr_60_value ? ghv_31 : _GEN_11595; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11597 = 8'h20 == new_ptr_60_value ? ghv_32 : _GEN_11596; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11598 = 8'h21 == new_ptr_60_value ? ghv_33 : _GEN_11597; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11599 = 8'h22 == new_ptr_60_value ? ghv_34 : _GEN_11598; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11600 = 8'h23 == new_ptr_60_value ? ghv_35 : _GEN_11599; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11601 = 8'h24 == new_ptr_60_value ? ghv_36 : _GEN_11600; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11602 = 8'h25 == new_ptr_60_value ? ghv_37 : _GEN_11601; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11603 = 8'h26 == new_ptr_60_value ? ghv_38 : _GEN_11602; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11604 = 8'h27 == new_ptr_60_value ? ghv_39 : _GEN_11603; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11605 = 8'h28 == new_ptr_60_value ? ghv_40 : _GEN_11604; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11606 = 8'h29 == new_ptr_60_value ? ghv_41 : _GEN_11605; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11607 = 8'h2a == new_ptr_60_value ? ghv_42 : _GEN_11606; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11608 = 8'h2b == new_ptr_60_value ? ghv_43 : _GEN_11607; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11609 = 8'h2c == new_ptr_60_value ? ghv_44 : _GEN_11608; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11610 = 8'h2d == new_ptr_60_value ? ghv_45 : _GEN_11609; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11611 = 8'h2e == new_ptr_60_value ? ghv_46 : _GEN_11610; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11612 = 8'h2f == new_ptr_60_value ? ghv_47 : _GEN_11611; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11613 = 8'h30 == new_ptr_60_value ? ghv_48 : _GEN_11612; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11614 = 8'h31 == new_ptr_60_value ? ghv_49 : _GEN_11613; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11615 = 8'h32 == new_ptr_60_value ? ghv_50 : _GEN_11614; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11616 = 8'h33 == new_ptr_60_value ? ghv_51 : _GEN_11615; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11617 = 8'h34 == new_ptr_60_value ? ghv_52 : _GEN_11616; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11618 = 8'h35 == new_ptr_60_value ? ghv_53 : _GEN_11617; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11619 = 8'h36 == new_ptr_60_value ? ghv_54 : _GEN_11618; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11620 = 8'h37 == new_ptr_60_value ? ghv_55 : _GEN_11619; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11621 = 8'h38 == new_ptr_60_value ? ghv_56 : _GEN_11620; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11622 = 8'h39 == new_ptr_60_value ? ghv_57 : _GEN_11621; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11623 = 8'h3a == new_ptr_60_value ? ghv_58 : _GEN_11622; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11624 = 8'h3b == new_ptr_60_value ? ghv_59 : _GEN_11623; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11625 = 8'h3c == new_ptr_60_value ? ghv_60 : _GEN_11624; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11626 = 8'h3d == new_ptr_60_value ? ghv_61 : _GEN_11625; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11627 = 8'h3e == new_ptr_60_value ? ghv_62 : _GEN_11626; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11628 = 8'h3f == new_ptr_60_value ? ghv_63 : _GEN_11627; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11629 = 8'h40 == new_ptr_60_value ? ghv_64 : _GEN_11628; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11630 = 8'h41 == new_ptr_60_value ? ghv_65 : _GEN_11629; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11631 = 8'h42 == new_ptr_60_value ? ghv_66 : _GEN_11630; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11632 = 8'h43 == new_ptr_60_value ? ghv_67 : _GEN_11631; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11633 = 8'h44 == new_ptr_60_value ? ghv_68 : _GEN_11632; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11634 = 8'h45 == new_ptr_60_value ? ghv_69 : _GEN_11633; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11635 = 8'h46 == new_ptr_60_value ? ghv_70 : _GEN_11634; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11636 = 8'h47 == new_ptr_60_value ? ghv_71 : _GEN_11635; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11637 = 8'h48 == new_ptr_60_value ? ghv_72 : _GEN_11636; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11638 = 8'h49 == new_ptr_60_value ? ghv_73 : _GEN_11637; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11639 = 8'h4a == new_ptr_60_value ? ghv_74 : _GEN_11638; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11640 = 8'h4b == new_ptr_60_value ? ghv_75 : _GEN_11639; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11641 = 8'h4c == new_ptr_60_value ? ghv_76 : _GEN_11640; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11642 = 8'h4d == new_ptr_60_value ? ghv_77 : _GEN_11641; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11643 = 8'h4e == new_ptr_60_value ? ghv_78 : _GEN_11642; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11644 = 8'h4f == new_ptr_60_value ? ghv_79 : _GEN_11643; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11645 = 8'h50 == new_ptr_60_value ? ghv_80 : _GEN_11644; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11646 = 8'h51 == new_ptr_60_value ? ghv_81 : _GEN_11645; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11647 = 8'h52 == new_ptr_60_value ? ghv_82 : _GEN_11646; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11648 = 8'h53 == new_ptr_60_value ? ghv_83 : _GEN_11647; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11649 = 8'h54 == new_ptr_60_value ? ghv_84 : _GEN_11648; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11650 = 8'h55 == new_ptr_60_value ? ghv_85 : _GEN_11649; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11651 = 8'h56 == new_ptr_60_value ? ghv_86 : _GEN_11650; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11652 = 8'h57 == new_ptr_60_value ? ghv_87 : _GEN_11651; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11653 = 8'h58 == new_ptr_60_value ? ghv_88 : _GEN_11652; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11654 = 8'h59 == new_ptr_60_value ? ghv_89 : _GEN_11653; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11655 = 8'h5a == new_ptr_60_value ? ghv_90 : _GEN_11654; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11656 = 8'h5b == new_ptr_60_value ? ghv_91 : _GEN_11655; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11657 = 8'h5c == new_ptr_60_value ? ghv_92 : _GEN_11656; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11658 = 8'h5d == new_ptr_60_value ? ghv_93 : _GEN_11657; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11659 = 8'h5e == new_ptr_60_value ? ghv_94 : _GEN_11658; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11660 = 8'h5f == new_ptr_60_value ? ghv_95 : _GEN_11659; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11661 = 8'h60 == new_ptr_60_value ? ghv_96 : _GEN_11660; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11662 = 8'h61 == new_ptr_60_value ? ghv_97 : _GEN_11661; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11663 = 8'h62 == new_ptr_60_value ? ghv_98 : _GEN_11662; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11664 = 8'h63 == new_ptr_60_value ? ghv_99 : _GEN_11663; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11665 = 8'h64 == new_ptr_60_value ? ghv_100 : _GEN_11664; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11666 = 8'h65 == new_ptr_60_value ? ghv_101 : _GEN_11665; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11667 = 8'h66 == new_ptr_60_value ? ghv_102 : _GEN_11666; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11668 = 8'h67 == new_ptr_60_value ? ghv_103 : _GEN_11667; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11669 = 8'h68 == new_ptr_60_value ? ghv_104 : _GEN_11668; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11670 = 8'h69 == new_ptr_60_value ? ghv_105 : _GEN_11669; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11671 = 8'h6a == new_ptr_60_value ? ghv_106 : _GEN_11670; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11672 = 8'h6b == new_ptr_60_value ? ghv_107 : _GEN_11671; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11673 = 8'h6c == new_ptr_60_value ? ghv_108 : _GEN_11672; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11674 = 8'h6d == new_ptr_60_value ? ghv_109 : _GEN_11673; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11675 = 8'h6e == new_ptr_60_value ? ghv_110 : _GEN_11674; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11676 = 8'h6f == new_ptr_60_value ? ghv_111 : _GEN_11675; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11677 = 8'h70 == new_ptr_60_value ? ghv_112 : _GEN_11676; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11678 = 8'h71 == new_ptr_60_value ? ghv_113 : _GEN_11677; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11679 = 8'h72 == new_ptr_60_value ? ghv_114 : _GEN_11678; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11680 = 8'h73 == new_ptr_60_value ? ghv_115 : _GEN_11679; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11681 = 8'h74 == new_ptr_60_value ? ghv_116 : _GEN_11680; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11682 = 8'h75 == new_ptr_60_value ? ghv_117 : _GEN_11681; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11683 = 8'h76 == new_ptr_60_value ? ghv_118 : _GEN_11682; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11684 = 8'h77 == new_ptr_60_value ? ghv_119 : _GEN_11683; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11685 = 8'h78 == new_ptr_60_value ? ghv_120 : _GEN_11684; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11686 = 8'h79 == new_ptr_60_value ? ghv_121 : _GEN_11685; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11687 = 8'h7a == new_ptr_60_value ? ghv_122 : _GEN_11686; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11688 = 8'h7b == new_ptr_60_value ? ghv_123 : _GEN_11687; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11689 = 8'h7c == new_ptr_60_value ? ghv_124 : _GEN_11688; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11690 = 8'h7d == new_ptr_60_value ? ghv_125 : _GEN_11689; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11691 = 8'h7e == new_ptr_60_value ? ghv_126 : _GEN_11690; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11692 = 8'h7f == new_ptr_60_value ? ghv_127 : _GEN_11691; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11693 = 8'h80 == new_ptr_60_value ? ghv_128 : _GEN_11692; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11694 = 8'h81 == new_ptr_60_value ? ghv_129 : _GEN_11693; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11695 = 8'h82 == new_ptr_60_value ? ghv_130 : _GEN_11694; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11696 = 8'h83 == new_ptr_60_value ? ghv_131 : _GEN_11695; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11697 = 8'h84 == new_ptr_60_value ? ghv_132 : _GEN_11696; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11698 = 8'h85 == new_ptr_60_value ? ghv_133 : _GEN_11697; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11699 = 8'h86 == new_ptr_60_value ? ghv_134 : _GEN_11698; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11700 = 8'h87 == new_ptr_60_value ? ghv_135 : _GEN_11699; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11701 = 8'h88 == new_ptr_60_value ? ghv_136 : _GEN_11700; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11702 = 8'h89 == new_ptr_60_value ? ghv_137 : _GEN_11701; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11703 = 8'h8a == new_ptr_60_value ? ghv_138 : _GEN_11702; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11704 = 8'h8b == new_ptr_60_value ? ghv_139 : _GEN_11703; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11705 = 8'h8c == new_ptr_60_value ? ghv_140 : _GEN_11704; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11706 = 8'h8d == new_ptr_60_value ? ghv_141 : _GEN_11705; // @[FrontendBundle.scala 329:{20,20}]
  wire  _GEN_11707 = 8'h8e == new_ptr_60_value ? ghv_142 : _GEN_11706; // @[FrontendBundle.scala 329:{20,20}]
  wire  _redirect_ghv_wens_T_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_0_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_value & shouldShiftVec_0
     & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_3 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_1_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_0_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_1_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_5 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_1_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_1_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_1_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_7 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_3_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_1_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_3_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_9 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_3_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_2_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_3_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_11 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_5_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_2_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_5_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_13 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_5_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_3_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_5_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_15 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_7_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_3_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_7_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_17 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_7_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_4_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_7_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_19 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_9_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_4_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_9_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_21 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_9_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_5_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_9_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_23 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_11_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_5_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_11_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_25 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_11_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_6_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_11_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_27 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_13_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_6_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_13_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_29 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_13_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_7_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_13_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_31 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_15_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_7_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_15_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_33 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_15_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_8_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_15_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_35 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_17_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_8_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_17_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_37 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_17_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_9_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_17_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_39 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_19_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_9_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_19_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_41 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_19_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_10_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_19_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_43 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_21_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_10_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_21_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_45 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_21_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_11_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_21_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_47 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_23_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_11_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_23_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_49 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_23_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_12_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_23_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_51 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_25_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_12_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_25_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_53 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_25_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_13_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_25_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_55 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_27_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_13_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_27_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_57 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_27_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_14_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_27_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_59 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_29_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_14_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_29_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_61 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_29_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_15_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_29_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_63 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_31_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_15_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_31_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_65 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_31_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_16_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_31_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_67 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_33_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_16_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_33_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_69 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_33_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_17_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_33_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_71 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_35_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_17_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_35_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_73 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_35_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_18_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_35_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_75 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_37_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_18_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_37_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_77 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_37_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_19_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_37_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_79 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_39_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_19_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_39_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_81 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_39_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_20_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_39_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_83 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_41_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_20_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_41_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_85 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_41_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_21_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_41_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_87 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_43_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_21_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_43_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_89 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_43_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_22_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_43_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_91 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_45_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_22_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_45_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_93 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_45_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_23_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_45_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_95 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_47_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_23_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_47_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_97 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_47_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_24_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_47_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_99 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_49_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_24_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_49_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_101 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_49_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_25_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_49_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_103 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_51_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_25_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_51_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_105 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_51_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_26_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_51_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_107 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_53_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_26_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_53_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_109 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_53_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_27_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_53_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_111 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_55_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_27_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_55_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_113 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_55_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_28_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_55_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_115 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_57_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_28_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_57_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_117 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_57_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_29_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_57_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_119 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_59_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_29_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_59_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_121 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_59_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_30_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_59_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_123 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_61_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_30_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_61_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_125 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_61_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_31_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_61_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_127 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_63_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_31_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_63_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_129 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_63_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_32_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_63_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_131 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_65_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_32_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_65_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_133 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_65_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_33_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_65_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_135 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_67_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_33_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_67_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_137 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_67_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_34_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_67_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_139 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_69_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_34_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_69_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_141 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_69_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_35_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_69_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_143 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_71_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_35_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_71_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_145 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_71_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_36_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_71_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_147 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_73_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_36_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_73_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_149 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_73_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_37_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_73_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_151 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_75_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_37_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_75_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_153 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_75_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_38_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_75_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_155 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_77_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_38_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_77_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_157 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_77_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_39_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_77_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_159 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_79_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_39_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_79_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_161 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_79_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_40_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_79_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_163 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_81_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_40_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_81_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_165 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_81_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_41_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_81_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_167 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_83_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_41_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_83_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_169 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_83_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_42_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_83_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_171 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_85_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_42_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_85_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_173 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_85_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_43_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_85_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_175 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_87_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_43_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_87_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_177 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_87_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_44_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_87_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_179 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_89_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_44_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_89_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_181 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_89_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_45_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_89_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_183 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_91_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_45_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_91_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_185 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_91_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_46_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_91_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_187 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_93_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_46_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_93_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_189 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_93_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_47_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_93_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_191 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_95_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_47_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_95_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_193 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_95_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_48_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_95_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_195 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_97_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_48_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_97_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_197 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_97_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_49_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_97_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_199 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_99_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_49_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_99_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_201 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_99_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_50_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_99_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_203 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_101_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_50_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_101_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_205 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_101_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_51_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_101_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_207 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_103_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_51_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_103_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_209 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_103_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_52_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_103_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_211 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_105_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_52_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_105_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_213 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_105_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_53_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_105_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_215 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_107_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_53_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_107_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_217 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_107_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_54_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_107_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_219 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_109_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_54_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_109_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_221 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_109_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_55_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_109_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_223 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_111_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_55_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_111_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_225 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_111_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_56_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_111_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_227 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_113_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_56_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_113_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_229 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_113_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_57_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_113_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_231 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_115_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_57_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_115_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_233 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_115_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_58_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_115_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_235 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_117_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_58_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_117_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_237 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_117_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_59_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_117_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_239 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_119_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_59_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_119_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_241 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_119_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_60_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_119_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_243 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_121_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_60_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_121_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_245 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_121_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_61_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_121_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_247 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_123_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_61_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_123_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_249 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_123_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_62_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_123_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_251 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_125_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_62_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_125_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_253 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_125_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_63_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_125_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_255 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_127_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_63_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_127_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_257 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_127_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_64_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_127_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_259 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_129_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_64_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_129_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_261 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_129_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_65_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_129_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_263 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_131_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_65_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_131_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_265 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_131_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_66_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_131_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_267 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_133_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_66_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_133_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_269 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_133_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_67_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_133_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_271 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_135_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_67_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_135_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_273 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_135_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_68_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_135_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_275 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_137_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_68_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_137_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_277 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_137_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_69_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_137_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_279 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_139_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_69_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_139_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_281 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_139_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_70_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_139_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_283 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_141_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_70_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_141_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_285 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_141_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_71_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_141_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_287 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_143_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_71_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_143_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_289 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_143_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_72_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_143_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_291 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_145_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_72_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_145_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_293 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_145_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_73_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_145_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_295 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_147_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_73_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_147_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_297 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_147_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_74_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_147_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_299 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_149_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_74_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_149_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_301 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_149_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_75_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_149_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_303 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_151_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_75_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_151_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_305 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_151_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_76_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_151_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_307 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_153_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_76_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_153_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_309 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_153_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_77_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_153_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_311 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_155_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_77_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_155_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_313 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_155_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_78_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_155_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_315 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_157_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_78_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_157_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_317 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_157_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_79_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_157_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_319 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_159_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_79_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_159_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_321 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_159_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_80_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_159_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_323 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_161_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_80_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_161_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_325 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_161_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_81_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_161_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_327 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_163_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_81_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_163_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_329 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_163_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_82_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_163_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_331 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_165_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_82_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_165_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_333 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_165_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_83_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_165_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_335 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_167_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_83_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_167_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_337 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_167_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_84_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_167_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_339 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_169_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_84_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_169_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_341 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_169_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_85_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_169_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_343 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_171_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_85_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_171_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_345 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_171_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_86_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_171_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_347 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_173_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_86_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_173_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_349 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_173_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_87_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_173_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_351 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_175_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_87_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_175_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_353 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_175_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_88_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_175_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_355 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_177_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_88_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_177_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_357 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_177_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_89_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_177_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_359 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_179_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_89_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_179_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_361 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_179_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_90_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_179_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_363 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_181_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_90_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_181_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_365 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_181_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_91_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_181_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_367 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_183_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_91_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_183_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_369 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_183_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_92_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_183_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_371 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_185_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_92_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_185_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_373 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_185_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_93_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_185_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_375 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_187_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_93_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_187_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_377 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_187_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_94_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_187_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_379 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_189_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_94_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_189_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_381 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_189_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_95_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_189_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_383 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_191_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_95_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_191_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_385 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_191_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_96_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_191_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_387 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_193_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_96_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_193_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_389 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_193_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_97_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_193_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_391 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_195_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_97_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_195_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_393 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_195_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_98_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_195_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_395 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_197_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_98_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_197_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_397 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_197_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_99_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_197_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_399 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_199_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_99_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_199_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_401 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_199_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_100_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_199_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_403 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_201_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_100_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_201_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_405 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_201_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_101_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_201_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_407 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_203_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_101_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_203_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_409 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_203_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_102_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_203_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_411 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_205_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_102_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_205_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_413 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_205_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_103_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_205_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_415 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_207_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_103_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_207_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_417 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_207_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_104_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_207_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_419 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_209_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_104_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_209_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_421 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_209_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_105_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_209_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_423 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_211_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_105_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_211_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_425 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_211_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_106_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_211_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_427 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_213_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_106_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_213_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_429 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_213_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_107_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_213_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_431 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_215_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_107_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_215_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_433 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_215_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_108_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_215_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_435 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_217_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_108_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_217_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_437 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_217_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_109_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_217_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_439 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_219_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_109_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_219_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_441 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_219_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_110_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_219_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_443 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_221_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_110_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_221_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_445 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_221_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_111_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_221_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_447 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_223_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_111_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_223_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_449 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_223_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_112_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_223_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_451 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_225_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_112_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_225_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_453 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_225_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_113_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_225_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_455 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_227_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_113_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_227_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_457 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_227_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_114_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_227_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_459 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_229_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_114_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_229_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_461 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_229_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_115_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_229_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_463 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_231_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_115_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_231_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_465 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_231_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_116_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_231_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_467 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_233_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_116_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_233_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_469 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_233_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_117_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_233_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_471 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_235_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_117_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_235_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_473 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_235_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_118_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_235_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_475 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_237_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_118_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_237_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_477 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_237_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_119_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_237_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_479 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_239_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_119_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_239_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_481 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_239_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_120_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_239_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_483 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_241_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_120_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_241_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_485 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_241_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_121_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_241_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_487 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_243_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_121_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_243_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_489 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_243_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_122_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_243_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_491 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_245_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_122_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_245_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_493 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_245_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_123_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_245_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_495 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_247_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_123_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_247_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_497 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_247_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_124_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_247_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_499 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_249_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_124_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_249_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_501 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_249_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_125_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_249_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_503 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_251_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_125_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_251_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_505 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_251_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_126_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_251_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_507 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_253_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_126_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_253_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_509 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_253_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_127_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_253_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_511 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_255_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_127_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_255_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_513 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_255_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_128_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_255_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_515 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_257_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_128_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_257_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_517 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_257_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_129_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_257_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_519 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_259_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_129_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_259_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_521 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_259_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_130_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_259_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_523 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_261_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_130_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_261_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_525 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_261_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_131_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_261_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_527 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_263_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_131_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_263_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_529 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_263_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_132_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_263_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_531 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_265_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_132_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_265_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_533 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_265_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_133_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_265_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_535 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_267_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_133_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_267_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_537 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_267_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_134_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_267_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_539 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_269_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_134_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_269_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_541 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_269_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_135_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_269_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_543 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_271_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_135_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_271_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_545 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_271_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_136_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_271_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_547 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_273_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_136_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_273_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_549 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_273_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_137_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_273_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_551 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_275_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_137_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_275_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_553 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_275_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_138_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_275_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_555 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_277_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_138_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_277_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_557 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_277_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_139_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_277_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_559 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_279_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_139_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_279_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_561 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_279_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_140_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_279_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_563 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_281_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_140_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_281_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_565 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_281_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_141_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_281_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_567 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_283_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_141_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_283_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_569 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_283_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_142_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_283_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_571 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_285_value &
    shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_142_1 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_285_value &
    shouldShiftVec_1 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_573 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_285_value &
    shouldShiftVec_0; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_143_0 = do_redirect_bits_cfiUpdate_histPtr_value == s1_ghv_wens_new_ptr_285_value &
    shouldShiftVec_0 & do_redirect_valid; // @[BPU.scala 627:103]
  wire  _redirect_ghv_wens_T_575 = do_redirect_bits_cfiUpdate_histPtr_value == 8'h0 & shouldShiftVec_1; // @[BPU.scala 627:82]
  wire  redirect_ghv_wens_143_1 = do_redirect_bits_cfiUpdate_histPtr_value == 8'h0 & shouldShiftVec_1 &
    do_redirect_valid; // @[BPU.scala 627:103]
  wire  _T_812 = redirect_ghv_wens_0_0 | redirect_ghv_wens_0_1; // @[BPU.scala 656:26]
  wire  _T_813 = redirect_ghv_wens_1_0 | redirect_ghv_wens_1_1; // @[BPU.scala 656:26]
  wire  _T_814 = redirect_ghv_wens_2_0 | redirect_ghv_wens_2_1; // @[BPU.scala 656:26]
  wire  _T_815 = redirect_ghv_wens_3_0 | redirect_ghv_wens_3_1; // @[BPU.scala 656:26]
  wire  _T_816 = redirect_ghv_wens_4_0 | redirect_ghv_wens_4_1; // @[BPU.scala 656:26]
  wire  _T_817 = redirect_ghv_wens_5_0 | redirect_ghv_wens_5_1; // @[BPU.scala 656:26]
  wire  _T_818 = redirect_ghv_wens_6_0 | redirect_ghv_wens_6_1; // @[BPU.scala 656:26]
  wire  _T_819 = redirect_ghv_wens_7_0 | redirect_ghv_wens_7_1; // @[BPU.scala 656:26]
  wire  _T_820 = redirect_ghv_wens_8_0 | redirect_ghv_wens_8_1; // @[BPU.scala 656:26]
  wire  _T_821 = redirect_ghv_wens_9_0 | redirect_ghv_wens_9_1; // @[BPU.scala 656:26]
  wire  _T_822 = redirect_ghv_wens_10_0 | redirect_ghv_wens_10_1; // @[BPU.scala 656:26]
  wire  _T_823 = redirect_ghv_wens_11_0 | redirect_ghv_wens_11_1; // @[BPU.scala 656:26]
  wire  _T_824 = redirect_ghv_wens_12_0 | redirect_ghv_wens_12_1; // @[BPU.scala 656:26]
  wire  _T_825 = redirect_ghv_wens_13_0 | redirect_ghv_wens_13_1; // @[BPU.scala 656:26]
  wire  _T_826 = redirect_ghv_wens_14_0 | redirect_ghv_wens_14_1; // @[BPU.scala 656:26]
  wire  _T_827 = redirect_ghv_wens_15_0 | redirect_ghv_wens_15_1; // @[BPU.scala 656:26]
  wire  _T_828 = redirect_ghv_wens_16_0 | redirect_ghv_wens_16_1; // @[BPU.scala 656:26]
  wire  _T_829 = redirect_ghv_wens_17_0 | redirect_ghv_wens_17_1; // @[BPU.scala 656:26]
  wire  _T_830 = redirect_ghv_wens_18_0 | redirect_ghv_wens_18_1; // @[BPU.scala 656:26]
  wire  _T_831 = redirect_ghv_wens_19_0 | redirect_ghv_wens_19_1; // @[BPU.scala 656:26]
  wire  _T_832 = redirect_ghv_wens_20_0 | redirect_ghv_wens_20_1; // @[BPU.scala 656:26]
  wire  _T_833 = redirect_ghv_wens_21_0 | redirect_ghv_wens_21_1; // @[BPU.scala 656:26]
  wire  _T_834 = redirect_ghv_wens_22_0 | redirect_ghv_wens_22_1; // @[BPU.scala 656:26]
  wire  _T_835 = redirect_ghv_wens_23_0 | redirect_ghv_wens_23_1; // @[BPU.scala 656:26]
  wire  _T_836 = redirect_ghv_wens_24_0 | redirect_ghv_wens_24_1; // @[BPU.scala 656:26]
  wire  _T_837 = redirect_ghv_wens_25_0 | redirect_ghv_wens_25_1; // @[BPU.scala 656:26]
  wire  _T_838 = redirect_ghv_wens_26_0 | redirect_ghv_wens_26_1; // @[BPU.scala 656:26]
  wire  _T_839 = redirect_ghv_wens_27_0 | redirect_ghv_wens_27_1; // @[BPU.scala 656:26]
  wire  _T_840 = redirect_ghv_wens_28_0 | redirect_ghv_wens_28_1; // @[BPU.scala 656:26]
  wire  _T_841 = redirect_ghv_wens_29_0 | redirect_ghv_wens_29_1; // @[BPU.scala 656:26]
  wire  _T_842 = redirect_ghv_wens_30_0 | redirect_ghv_wens_30_1; // @[BPU.scala 656:26]
  wire  _T_843 = redirect_ghv_wens_31_0 | redirect_ghv_wens_31_1; // @[BPU.scala 656:26]
  wire  _T_844 = redirect_ghv_wens_32_0 | redirect_ghv_wens_32_1; // @[BPU.scala 656:26]
  wire  _T_845 = redirect_ghv_wens_33_0 | redirect_ghv_wens_33_1; // @[BPU.scala 656:26]
  wire  _T_846 = redirect_ghv_wens_34_0 | redirect_ghv_wens_34_1; // @[BPU.scala 656:26]
  wire  _T_847 = redirect_ghv_wens_35_0 | redirect_ghv_wens_35_1; // @[BPU.scala 656:26]
  wire  _T_848 = redirect_ghv_wens_36_0 | redirect_ghv_wens_36_1; // @[BPU.scala 656:26]
  wire  _T_849 = redirect_ghv_wens_37_0 | redirect_ghv_wens_37_1; // @[BPU.scala 656:26]
  wire  _T_850 = redirect_ghv_wens_38_0 | redirect_ghv_wens_38_1; // @[BPU.scala 656:26]
  wire  _T_851 = redirect_ghv_wens_39_0 | redirect_ghv_wens_39_1; // @[BPU.scala 656:26]
  wire  _T_852 = redirect_ghv_wens_40_0 | redirect_ghv_wens_40_1; // @[BPU.scala 656:26]
  wire  _T_853 = redirect_ghv_wens_41_0 | redirect_ghv_wens_41_1; // @[BPU.scala 656:26]
  wire  _T_854 = redirect_ghv_wens_42_0 | redirect_ghv_wens_42_1; // @[BPU.scala 656:26]
  wire  _T_855 = redirect_ghv_wens_43_0 | redirect_ghv_wens_43_1; // @[BPU.scala 656:26]
  wire  _T_856 = redirect_ghv_wens_44_0 | redirect_ghv_wens_44_1; // @[BPU.scala 656:26]
  wire  _T_857 = redirect_ghv_wens_45_0 | redirect_ghv_wens_45_1; // @[BPU.scala 656:26]
  wire  _T_858 = redirect_ghv_wens_46_0 | redirect_ghv_wens_46_1; // @[BPU.scala 656:26]
  wire  _T_859 = redirect_ghv_wens_47_0 | redirect_ghv_wens_47_1; // @[BPU.scala 656:26]
  wire  _T_860 = redirect_ghv_wens_48_0 | redirect_ghv_wens_48_1; // @[BPU.scala 656:26]
  wire  _T_861 = redirect_ghv_wens_49_0 | redirect_ghv_wens_49_1; // @[BPU.scala 656:26]
  wire  _T_862 = redirect_ghv_wens_50_0 | redirect_ghv_wens_50_1; // @[BPU.scala 656:26]
  wire  _T_863 = redirect_ghv_wens_51_0 | redirect_ghv_wens_51_1; // @[BPU.scala 656:26]
  wire  _T_864 = redirect_ghv_wens_52_0 | redirect_ghv_wens_52_1; // @[BPU.scala 656:26]
  wire  _T_865 = redirect_ghv_wens_53_0 | redirect_ghv_wens_53_1; // @[BPU.scala 656:26]
  wire  _T_866 = redirect_ghv_wens_54_0 | redirect_ghv_wens_54_1; // @[BPU.scala 656:26]
  wire  _T_867 = redirect_ghv_wens_55_0 | redirect_ghv_wens_55_1; // @[BPU.scala 656:26]
  wire  _T_868 = redirect_ghv_wens_56_0 | redirect_ghv_wens_56_1; // @[BPU.scala 656:26]
  wire  _T_869 = redirect_ghv_wens_57_0 | redirect_ghv_wens_57_1; // @[BPU.scala 656:26]
  wire  _T_870 = redirect_ghv_wens_58_0 | redirect_ghv_wens_58_1; // @[BPU.scala 656:26]
  wire  _T_871 = redirect_ghv_wens_59_0 | redirect_ghv_wens_59_1; // @[BPU.scala 656:26]
  wire  _T_872 = redirect_ghv_wens_60_0 | redirect_ghv_wens_60_1; // @[BPU.scala 656:26]
  wire  _T_873 = redirect_ghv_wens_61_0 | redirect_ghv_wens_61_1; // @[BPU.scala 656:26]
  wire  _T_874 = redirect_ghv_wens_62_0 | redirect_ghv_wens_62_1; // @[BPU.scala 656:26]
  wire  _T_875 = redirect_ghv_wens_63_0 | redirect_ghv_wens_63_1; // @[BPU.scala 656:26]
  wire  _T_876 = redirect_ghv_wens_64_0 | redirect_ghv_wens_64_1; // @[BPU.scala 656:26]
  wire  _T_877 = redirect_ghv_wens_65_0 | redirect_ghv_wens_65_1; // @[BPU.scala 656:26]
  wire  _T_878 = redirect_ghv_wens_66_0 | redirect_ghv_wens_66_1; // @[BPU.scala 656:26]
  wire  _T_879 = redirect_ghv_wens_67_0 | redirect_ghv_wens_67_1; // @[BPU.scala 656:26]
  wire  _T_880 = redirect_ghv_wens_68_0 | redirect_ghv_wens_68_1; // @[BPU.scala 656:26]
  wire  _T_881 = redirect_ghv_wens_69_0 | redirect_ghv_wens_69_1; // @[BPU.scala 656:26]
  wire  _T_882 = redirect_ghv_wens_70_0 | redirect_ghv_wens_70_1; // @[BPU.scala 656:26]
  wire  _T_883 = redirect_ghv_wens_71_0 | redirect_ghv_wens_71_1; // @[BPU.scala 656:26]
  wire  _T_884 = redirect_ghv_wens_72_0 | redirect_ghv_wens_72_1; // @[BPU.scala 656:26]
  wire  _T_885 = redirect_ghv_wens_73_0 | redirect_ghv_wens_73_1; // @[BPU.scala 656:26]
  wire  _T_886 = redirect_ghv_wens_74_0 | redirect_ghv_wens_74_1; // @[BPU.scala 656:26]
  wire  _T_887 = redirect_ghv_wens_75_0 | redirect_ghv_wens_75_1; // @[BPU.scala 656:26]
  wire  _T_888 = redirect_ghv_wens_76_0 | redirect_ghv_wens_76_1; // @[BPU.scala 656:26]
  wire  _T_889 = redirect_ghv_wens_77_0 | redirect_ghv_wens_77_1; // @[BPU.scala 656:26]
  wire  _T_890 = redirect_ghv_wens_78_0 | redirect_ghv_wens_78_1; // @[BPU.scala 656:26]
  wire  _T_891 = redirect_ghv_wens_79_0 | redirect_ghv_wens_79_1; // @[BPU.scala 656:26]
  wire  _T_892 = redirect_ghv_wens_80_0 | redirect_ghv_wens_80_1; // @[BPU.scala 656:26]
  wire  _T_893 = redirect_ghv_wens_81_0 | redirect_ghv_wens_81_1; // @[BPU.scala 656:26]
  wire  _T_894 = redirect_ghv_wens_82_0 | redirect_ghv_wens_82_1; // @[BPU.scala 656:26]
  wire  _T_895 = redirect_ghv_wens_83_0 | redirect_ghv_wens_83_1; // @[BPU.scala 656:26]
  wire  _T_896 = redirect_ghv_wens_84_0 | redirect_ghv_wens_84_1; // @[BPU.scala 656:26]
  wire  _T_897 = redirect_ghv_wens_85_0 | redirect_ghv_wens_85_1; // @[BPU.scala 656:26]
  wire  _T_898 = redirect_ghv_wens_86_0 | redirect_ghv_wens_86_1; // @[BPU.scala 656:26]
  wire  _T_899 = redirect_ghv_wens_87_0 | redirect_ghv_wens_87_1; // @[BPU.scala 656:26]
  wire  _T_900 = redirect_ghv_wens_88_0 | redirect_ghv_wens_88_1; // @[BPU.scala 656:26]
  wire  _T_901 = redirect_ghv_wens_89_0 | redirect_ghv_wens_89_1; // @[BPU.scala 656:26]
  wire  _T_902 = redirect_ghv_wens_90_0 | redirect_ghv_wens_90_1; // @[BPU.scala 656:26]
  wire  _T_903 = redirect_ghv_wens_91_0 | redirect_ghv_wens_91_1; // @[BPU.scala 656:26]
  wire  _T_904 = redirect_ghv_wens_92_0 | redirect_ghv_wens_92_1; // @[BPU.scala 656:26]
  wire  _T_905 = redirect_ghv_wens_93_0 | redirect_ghv_wens_93_1; // @[BPU.scala 656:26]
  wire  _T_906 = redirect_ghv_wens_94_0 | redirect_ghv_wens_94_1; // @[BPU.scala 656:26]
  wire  _T_907 = redirect_ghv_wens_95_0 | redirect_ghv_wens_95_1; // @[BPU.scala 656:26]
  wire  _T_908 = redirect_ghv_wens_96_0 | redirect_ghv_wens_96_1; // @[BPU.scala 656:26]
  wire  _T_909 = redirect_ghv_wens_97_0 | redirect_ghv_wens_97_1; // @[BPU.scala 656:26]
  wire  _T_910 = redirect_ghv_wens_98_0 | redirect_ghv_wens_98_1; // @[BPU.scala 656:26]
  wire  _T_911 = redirect_ghv_wens_99_0 | redirect_ghv_wens_99_1; // @[BPU.scala 656:26]
  wire  _T_912 = redirect_ghv_wens_100_0 | redirect_ghv_wens_100_1; // @[BPU.scala 656:26]
  wire  _T_913 = redirect_ghv_wens_101_0 | redirect_ghv_wens_101_1; // @[BPU.scala 656:26]
  wire  _T_914 = redirect_ghv_wens_102_0 | redirect_ghv_wens_102_1; // @[BPU.scala 656:26]
  wire  _T_915 = redirect_ghv_wens_103_0 | redirect_ghv_wens_103_1; // @[BPU.scala 656:26]
  wire  _T_916 = redirect_ghv_wens_104_0 | redirect_ghv_wens_104_1; // @[BPU.scala 656:26]
  wire  _T_917 = redirect_ghv_wens_105_0 | redirect_ghv_wens_105_1; // @[BPU.scala 656:26]
  wire  _T_918 = redirect_ghv_wens_106_0 | redirect_ghv_wens_106_1; // @[BPU.scala 656:26]
  wire  _T_919 = redirect_ghv_wens_107_0 | redirect_ghv_wens_107_1; // @[BPU.scala 656:26]
  wire  _T_920 = redirect_ghv_wens_108_0 | redirect_ghv_wens_108_1; // @[BPU.scala 656:26]
  wire  _T_921 = redirect_ghv_wens_109_0 | redirect_ghv_wens_109_1; // @[BPU.scala 656:26]
  wire  _T_922 = redirect_ghv_wens_110_0 | redirect_ghv_wens_110_1; // @[BPU.scala 656:26]
  wire  _T_923 = redirect_ghv_wens_111_0 | redirect_ghv_wens_111_1; // @[BPU.scala 656:26]
  wire  _T_924 = redirect_ghv_wens_112_0 | redirect_ghv_wens_112_1; // @[BPU.scala 656:26]
  wire  _T_925 = redirect_ghv_wens_113_0 | redirect_ghv_wens_113_1; // @[BPU.scala 656:26]
  wire  _T_926 = redirect_ghv_wens_114_0 | redirect_ghv_wens_114_1; // @[BPU.scala 656:26]
  wire  _T_927 = redirect_ghv_wens_115_0 | redirect_ghv_wens_115_1; // @[BPU.scala 656:26]
  wire  _T_928 = redirect_ghv_wens_116_0 | redirect_ghv_wens_116_1; // @[BPU.scala 656:26]
  wire  _T_929 = redirect_ghv_wens_117_0 | redirect_ghv_wens_117_1; // @[BPU.scala 656:26]
  wire  _T_930 = redirect_ghv_wens_118_0 | redirect_ghv_wens_118_1; // @[BPU.scala 656:26]
  wire  _T_931 = redirect_ghv_wens_119_0 | redirect_ghv_wens_119_1; // @[BPU.scala 656:26]
  wire  _T_932 = redirect_ghv_wens_120_0 | redirect_ghv_wens_120_1; // @[BPU.scala 656:26]
  wire  _T_933 = redirect_ghv_wens_121_0 | redirect_ghv_wens_121_1; // @[BPU.scala 656:26]
  wire  _T_934 = redirect_ghv_wens_122_0 | redirect_ghv_wens_122_1; // @[BPU.scala 656:26]
  wire  _T_935 = redirect_ghv_wens_123_0 | redirect_ghv_wens_123_1; // @[BPU.scala 656:26]
  wire  _T_936 = redirect_ghv_wens_124_0 | redirect_ghv_wens_124_1; // @[BPU.scala 656:26]
  wire  _T_937 = redirect_ghv_wens_125_0 | redirect_ghv_wens_125_1; // @[BPU.scala 656:26]
  wire  _T_938 = redirect_ghv_wens_126_0 | redirect_ghv_wens_126_1; // @[BPU.scala 656:26]
  wire  _T_939 = redirect_ghv_wens_127_0 | redirect_ghv_wens_127_1; // @[BPU.scala 656:26]
  wire  _T_940 = redirect_ghv_wens_128_0 | redirect_ghv_wens_128_1; // @[BPU.scala 656:26]
  wire  _T_941 = redirect_ghv_wens_129_0 | redirect_ghv_wens_129_1; // @[BPU.scala 656:26]
  wire  _T_942 = redirect_ghv_wens_130_0 | redirect_ghv_wens_130_1; // @[BPU.scala 656:26]
  wire  _T_943 = redirect_ghv_wens_131_0 | redirect_ghv_wens_131_1; // @[BPU.scala 656:26]
  wire  _T_944 = redirect_ghv_wens_132_0 | redirect_ghv_wens_132_1; // @[BPU.scala 656:26]
  wire  _T_945 = redirect_ghv_wens_133_0 | redirect_ghv_wens_133_1; // @[BPU.scala 656:26]
  wire  _T_946 = redirect_ghv_wens_134_0 | redirect_ghv_wens_134_1; // @[BPU.scala 656:26]
  wire  _T_947 = redirect_ghv_wens_135_0 | redirect_ghv_wens_135_1; // @[BPU.scala 656:26]
  wire  _T_948 = redirect_ghv_wens_136_0 | redirect_ghv_wens_136_1; // @[BPU.scala 656:26]
  wire  _T_949 = redirect_ghv_wens_137_0 | redirect_ghv_wens_137_1; // @[BPU.scala 656:26]
  wire  _T_950 = redirect_ghv_wens_138_0 | redirect_ghv_wens_138_1; // @[BPU.scala 656:26]
  wire  _T_951 = redirect_ghv_wens_139_0 | redirect_ghv_wens_139_1; // @[BPU.scala 656:26]
  wire  _T_952 = redirect_ghv_wens_140_0 | redirect_ghv_wens_140_1; // @[BPU.scala 656:26]
  wire  _T_953 = redirect_ghv_wens_141_0 | redirect_ghv_wens_141_1; // @[BPU.scala 656:26]
  wire  _T_954 = redirect_ghv_wens_142_0 | redirect_ghv_wens_142_1; // @[BPU.scala 656:26]
  wire  _T_955 = redirect_ghv_wens_143_0 | redirect_ghv_wens_143_1; // @[BPU.scala 656:26]
  wire [7:0] _GEN_11713 = 2'h1 == do_redirect_bits_cfiUpdate_shift ? updated_fh_res_hist_0_new_folded_hist_1 :
    updated_fh_res_hist_0_new_folded_hist; // @[PriorityMuxGen.scala 140:{24,24}]
  wire [7:0] _GEN_11716 = 2'h1 == do_redirect_bits_cfiUpdate_shift ? updated_fh_res_hist_1_new_folded_hist_1 :
    updated_fh_res_hist_1_new_folded_hist; // @[PriorityMuxGen.scala 140:{24,24}]
  wire [7:0] _GEN_11719 = 2'h1 == do_redirect_bits_cfiUpdate_shift ? updated_fh_res_hist_2_new_folded_hist_1 :
    updated_fh_res_hist_2_new_folded_hist; // @[PriorityMuxGen.scala 140:{24,24}]
  wire [10:0] _GEN_11722 = 2'h1 == do_redirect_bits_cfiUpdate_shift ? updated_fh_res_hist_3_new_folded_hist_1 :
    updated_fh_res_hist_3_new_folded_hist; // @[PriorityMuxGen.scala 140:{24,24}]
  wire [3:0] _GEN_11725 = 2'h1 == do_redirect_bits_cfiUpdate_shift ? updated_fh_res_hist_4_new_folded_hist_1 :
    updated_fh_res_hist_4_new_folded_hist; // @[PriorityMuxGen.scala 140:{24,24}]
  wire [10:0] _GEN_11728 = 2'h1 == do_redirect_bits_cfiUpdate_shift ? updated_fh_res_hist_5_new_folded_hist_1 :
    updated_fh_res_hist_5_new_folded_hist; // @[PriorityMuxGen.scala 140:{24,24}]
  wire [8:0] _GEN_11731 = 2'h1 == do_redirect_bits_cfiUpdate_shift ? updated_fh_res_hist_6_new_folded_hist_1 :
    updated_fh_res_hist_6_new_folded_hist; // @[PriorityMuxGen.scala 140:{24,24}]
  wire [8:0] _GEN_11734 = 2'h1 == do_redirect_bits_cfiUpdate_shift ? updated_fh_res_hist_7_new_folded_hist_1 :
    updated_fh_res_hist_7_new_folded_hist; // @[PriorityMuxGen.scala 140:{24,24}]
  wire [7:0] _GEN_11737 = 2'h1 == do_redirect_bits_cfiUpdate_shift ? updated_fh_res_hist_8_new_folded_hist_1 :
    updated_fh_res_hist_8_new_folded_hist; // @[PriorityMuxGen.scala 140:{24,24}]
  wire [6:0] _GEN_11740 = 2'h1 == do_redirect_bits_cfiUpdate_shift ? updated_fh_res_hist_9_new_folded_hist_1 :
    updated_fh_res_hist_9_new_folded_hist; // @[PriorityMuxGen.scala 140:{24,24}]
  wire [8:0] _GEN_11743 = 2'h1 == do_redirect_bits_cfiUpdate_shift ? updated_fh_res_hist_10_new_folded_hist_1 :
    updated_fh_res_hist_10_new_folded_hist; // @[PriorityMuxGen.scala 140:{24,24}]
  wire [7:0] _GEN_11746 = 2'h1 == do_redirect_bits_cfiUpdate_shift ? updated_fh_res_hist_11_new_folded_hist_1 :
    updated_fh_res_hist_11_new_folded_hist; // @[PriorityMuxGen.scala 140:{24,24}]
  wire [6:0] _GEN_11749 = 2'h1 == do_redirect_bits_cfiUpdate_shift ? updated_fh_res_hist_12_new_folded_hist_1 :
    updated_fh_res_hist_12_new_folded_hist; // @[PriorityMuxGen.scala 140:{24,24}]
  wire [6:0] _GEN_11752 = 2'h1 == do_redirect_bits_cfiUpdate_shift ? updated_fh_res_hist_13_new_folded_hist_1 :
    updated_fh_res_hist_13_new_folded_hist; // @[PriorityMuxGen.scala 140:{24,24}]
  wire [6:0] _GEN_11755 = 2'h1 == do_redirect_bits_cfiUpdate_shift ? updated_fh_res_hist_14_new_folded_hist_1 :
    updated_fh_res_hist_14_new_folded_hist; // @[PriorityMuxGen.scala 140:{24,24}]
  wire [10:0] _GEN_11758 = 2'h1 == do_redirect_bits_cfiUpdate_shift ? updated_fh_res_hist_15_new_folded_hist_1 :
    updated_fh_res_hist_15_new_folded_hist; // @[PriorityMuxGen.scala 140:{24,24}]
  wire [7:0] _GEN_11761 = 2'h1 == do_redirect_bits_cfiUpdate_shift ? updated_fh_res_hist_16_new_folded_hist_1 :
    updated_fh_res_hist_16_new_folded_hist; // @[PriorityMuxGen.scala 140:{24,24}]
  wire [7:0] _GEN_11764 = 2'h1 == do_redirect_bits_cfiUpdate_shift ? updated_fh_res_hist_17_new_folded_hist_1 :
    updated_fh_res_hist_17_new_folded_hist; // @[PriorityMuxGen.scala 140:{24,24}]
  wire  ghv_wens_0 = _T_123 | _T_385 | _T_666 | _T_812; // @[BPU.scala 674:113]
  wire  ghv_write_datas_0 = ghv_write_datas_0_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_1 = _T_124 | _T_386 | _T_667 | _T_813; // @[BPU.scala 674:113]
  wire  ghv_write_datas_1 = ghv_write_datas_1_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_2 = _T_125 | _T_387 | _T_668 | _T_814; // @[BPU.scala 674:113]
  wire  ghv_write_datas_2 = ghv_write_datas_2_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_3 = _T_126 | _T_388 | _T_669 | _T_815; // @[BPU.scala 674:113]
  wire  ghv_write_datas_3 = ghv_write_datas_3_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_4 = _T_127 | _T_389 | _T_670 | _T_816; // @[BPU.scala 674:113]
  wire  ghv_write_datas_4 = ghv_write_datas_4_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_5 = _T_128 | _T_390 | _T_671 | _T_817; // @[BPU.scala 674:113]
  wire  ghv_write_datas_5 = ghv_write_datas_5_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_6 = _T_129 | _T_391 | _T_672 | _T_818; // @[BPU.scala 674:113]
  wire  ghv_write_datas_6 = ghv_write_datas_6_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_7 = _T_130 | _T_392 | _T_673 | _T_819; // @[BPU.scala 674:113]
  wire  ghv_write_datas_7 = ghv_write_datas_7_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_8 = _T_131 | _T_393 | _T_674 | _T_820; // @[BPU.scala 674:113]
  wire  ghv_write_datas_8 = ghv_write_datas_8_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_9 = _T_132 | _T_394 | _T_675 | _T_821; // @[BPU.scala 674:113]
  wire  ghv_write_datas_9 = ghv_write_datas_9_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_10 = _T_133 | _T_395 | _T_676 | _T_822; // @[BPU.scala 674:113]
  wire  ghv_write_datas_10 = ghv_write_datas_10_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_11 = _T_134 | _T_396 | _T_677 | _T_823; // @[BPU.scala 674:113]
  wire  ghv_write_datas_11 = ghv_write_datas_11_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_12 = _T_135 | _T_397 | _T_678 | _T_824; // @[BPU.scala 674:113]
  wire  ghv_write_datas_12 = ghv_write_datas_12_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_13 = _T_136 | _T_398 | _T_679 | _T_825; // @[BPU.scala 674:113]
  wire  ghv_write_datas_13 = ghv_write_datas_13_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_14 = _T_137 | _T_399 | _T_680 | _T_826; // @[BPU.scala 674:113]
  wire  ghv_write_datas_14 = ghv_write_datas_14_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_15 = _T_138 | _T_400 | _T_681 | _T_827; // @[BPU.scala 674:113]
  wire  ghv_write_datas_15 = ghv_write_datas_15_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_16 = _T_139 | _T_401 | _T_682 | _T_828; // @[BPU.scala 674:113]
  wire  ghv_write_datas_16 = ghv_write_datas_16_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_17 = _T_140 | _T_402 | _T_683 | _T_829; // @[BPU.scala 674:113]
  wire  ghv_write_datas_17 = ghv_write_datas_17_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_18 = _T_141 | _T_403 | _T_684 | _T_830; // @[BPU.scala 674:113]
  wire  ghv_write_datas_18 = ghv_write_datas_18_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_19 = _T_142 | _T_404 | _T_685 | _T_831; // @[BPU.scala 674:113]
  wire  ghv_write_datas_19 = ghv_write_datas_19_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_20 = _T_143 | _T_405 | _T_686 | _T_832; // @[BPU.scala 674:113]
  wire  ghv_write_datas_20 = ghv_write_datas_20_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_21 = _T_144 | _T_406 | _T_687 | _T_833; // @[BPU.scala 674:113]
  wire  ghv_write_datas_21 = ghv_write_datas_21_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_22 = _T_145 | _T_407 | _T_688 | _T_834; // @[BPU.scala 674:113]
  wire  ghv_write_datas_22 = ghv_write_datas_22_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_23 = _T_146 | _T_408 | _T_689 | _T_835; // @[BPU.scala 674:113]
  wire  ghv_write_datas_23 = ghv_write_datas_23_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_24 = _T_147 | _T_409 | _T_690 | _T_836; // @[BPU.scala 674:113]
  wire  ghv_write_datas_24 = ghv_write_datas_24_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_25 = _T_148 | _T_410 | _T_691 | _T_837; // @[BPU.scala 674:113]
  wire  ghv_write_datas_25 = ghv_write_datas_25_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_26 = _T_149 | _T_411 | _T_692 | _T_838; // @[BPU.scala 674:113]
  wire  ghv_write_datas_26 = ghv_write_datas_26_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_27 = _T_150 | _T_412 | _T_693 | _T_839; // @[BPU.scala 674:113]
  wire  ghv_write_datas_27 = ghv_write_datas_27_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_28 = _T_151 | _T_413 | _T_694 | _T_840; // @[BPU.scala 674:113]
  wire  ghv_write_datas_28 = ghv_write_datas_28_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_29 = _T_152 | _T_414 | _T_695 | _T_841; // @[BPU.scala 674:113]
  wire  ghv_write_datas_29 = ghv_write_datas_29_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_30 = _T_153 | _T_415 | _T_696 | _T_842; // @[BPU.scala 674:113]
  wire  ghv_write_datas_30 = ghv_write_datas_30_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_31 = _T_154 | _T_416 | _T_697 | _T_843; // @[BPU.scala 674:113]
  wire  ghv_write_datas_31 = ghv_write_datas_31_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_32 = _T_155 | _T_417 | _T_698 | _T_844; // @[BPU.scala 674:113]
  wire  ghv_write_datas_32 = ghv_write_datas_32_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_33 = _T_156 | _T_418 | _T_699 | _T_845; // @[BPU.scala 674:113]
  wire  ghv_write_datas_33 = ghv_write_datas_33_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_34 = _T_157 | _T_419 | _T_700 | _T_846; // @[BPU.scala 674:113]
  wire  ghv_write_datas_34 = ghv_write_datas_34_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_35 = _T_158 | _T_420 | _T_701 | _T_847; // @[BPU.scala 674:113]
  wire  ghv_write_datas_35 = ghv_write_datas_35_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_36 = _T_159 | _T_421 | _T_702 | _T_848; // @[BPU.scala 674:113]
  wire  ghv_write_datas_36 = ghv_write_datas_36_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_37 = _T_160 | _T_422 | _T_703 | _T_849; // @[BPU.scala 674:113]
  wire  ghv_write_datas_37 = ghv_write_datas_37_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_38 = _T_161 | _T_423 | _T_704 | _T_850; // @[BPU.scala 674:113]
  wire  ghv_write_datas_38 = ghv_write_datas_38_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_39 = _T_162 | _T_424 | _T_705 | _T_851; // @[BPU.scala 674:113]
  wire  ghv_write_datas_39 = ghv_write_datas_39_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_40 = _T_163 | _T_425 | _T_706 | _T_852; // @[BPU.scala 674:113]
  wire  ghv_write_datas_40 = ghv_write_datas_40_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_41 = _T_164 | _T_426 | _T_707 | _T_853; // @[BPU.scala 674:113]
  wire  ghv_write_datas_41 = ghv_write_datas_41_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_42 = _T_165 | _T_427 | _T_708 | _T_854; // @[BPU.scala 674:113]
  wire  ghv_write_datas_42 = ghv_write_datas_42_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_43 = _T_166 | _T_428 | _T_709 | _T_855; // @[BPU.scala 674:113]
  wire  ghv_write_datas_43 = ghv_write_datas_43_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_44 = _T_167 | _T_429 | _T_710 | _T_856; // @[BPU.scala 674:113]
  wire  ghv_write_datas_44 = ghv_write_datas_44_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_45 = _T_168 | _T_430 | _T_711 | _T_857; // @[BPU.scala 674:113]
  wire  ghv_write_datas_45 = ghv_write_datas_45_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_46 = _T_169 | _T_431 | _T_712 | _T_858; // @[BPU.scala 674:113]
  wire  ghv_write_datas_46 = ghv_write_datas_46_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_47 = _T_170 | _T_432 | _T_713 | _T_859; // @[BPU.scala 674:113]
  wire  ghv_write_datas_47 = ghv_write_datas_47_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_48 = _T_171 | _T_433 | _T_714 | _T_860; // @[BPU.scala 674:113]
  wire  ghv_write_datas_48 = ghv_write_datas_48_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_49 = _T_172 | _T_434 | _T_715 | _T_861; // @[BPU.scala 674:113]
  wire  ghv_write_datas_49 = ghv_write_datas_49_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_50 = _T_173 | _T_435 | _T_716 | _T_862; // @[BPU.scala 674:113]
  wire  ghv_write_datas_50 = ghv_write_datas_50_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_51 = _T_174 | _T_436 | _T_717 | _T_863; // @[BPU.scala 674:113]
  wire  ghv_write_datas_51 = ghv_write_datas_51_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_52 = _T_175 | _T_437 | _T_718 | _T_864; // @[BPU.scala 674:113]
  wire  ghv_write_datas_52 = ghv_write_datas_52_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_53 = _T_176 | _T_438 | _T_719 | _T_865; // @[BPU.scala 674:113]
  wire  ghv_write_datas_53 = ghv_write_datas_53_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_54 = _T_177 | _T_439 | _T_720 | _T_866; // @[BPU.scala 674:113]
  wire  ghv_write_datas_54 = ghv_write_datas_54_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_55 = _T_178 | _T_440 | _T_721 | _T_867; // @[BPU.scala 674:113]
  wire  ghv_write_datas_55 = ghv_write_datas_55_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_56 = _T_179 | _T_441 | _T_722 | _T_868; // @[BPU.scala 674:113]
  wire  ghv_write_datas_56 = ghv_write_datas_56_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_57 = _T_180 | _T_442 | _T_723 | _T_869; // @[BPU.scala 674:113]
  wire  ghv_write_datas_57 = ghv_write_datas_57_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_58 = _T_181 | _T_443 | _T_724 | _T_870; // @[BPU.scala 674:113]
  wire  ghv_write_datas_58 = ghv_write_datas_58_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_59 = _T_182 | _T_444 | _T_725 | _T_871; // @[BPU.scala 674:113]
  wire  ghv_write_datas_59 = ghv_write_datas_59_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_60 = _T_183 | _T_445 | _T_726 | _T_872; // @[BPU.scala 674:113]
  wire  ghv_write_datas_60 = ghv_write_datas_60_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_61 = _T_184 | _T_446 | _T_727 | _T_873; // @[BPU.scala 674:113]
  wire  ghv_write_datas_61 = ghv_write_datas_61_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_62 = _T_185 | _T_447 | _T_728 | _T_874; // @[BPU.scala 674:113]
  wire  ghv_write_datas_62 = ghv_write_datas_62_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_63 = _T_186 | _T_448 | _T_729 | _T_875; // @[BPU.scala 674:113]
  wire  ghv_write_datas_63 = ghv_write_datas_63_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_64 = _T_187 | _T_449 | _T_730 | _T_876; // @[BPU.scala 674:113]
  wire  ghv_write_datas_64 = ghv_write_datas_64_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_65 = _T_188 | _T_450 | _T_731 | _T_877; // @[BPU.scala 674:113]
  wire  ghv_write_datas_65 = ghv_write_datas_65_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_66 = _T_189 | _T_451 | _T_732 | _T_878; // @[BPU.scala 674:113]
  wire  ghv_write_datas_66 = ghv_write_datas_66_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_67 = _T_190 | _T_452 | _T_733 | _T_879; // @[BPU.scala 674:113]
  wire  ghv_write_datas_67 = ghv_write_datas_67_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_68 = _T_191 | _T_453 | _T_734 | _T_880; // @[BPU.scala 674:113]
  wire  ghv_write_datas_68 = ghv_write_datas_68_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_69 = _T_192 | _T_454 | _T_735 | _T_881; // @[BPU.scala 674:113]
  wire  ghv_write_datas_69 = ghv_write_datas_69_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_70 = _T_193 | _T_455 | _T_736 | _T_882; // @[BPU.scala 674:113]
  wire  ghv_write_datas_70 = ghv_write_datas_70_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_71 = _T_194 | _T_456 | _T_737 | _T_883; // @[BPU.scala 674:113]
  wire  ghv_write_datas_71 = ghv_write_datas_71_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_72 = _T_195 | _T_457 | _T_738 | _T_884; // @[BPU.scala 674:113]
  wire  ghv_write_datas_72 = ghv_write_datas_72_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_73 = _T_196 | _T_458 | _T_739 | _T_885; // @[BPU.scala 674:113]
  wire  ghv_write_datas_73 = ghv_write_datas_73_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_74 = _T_197 | _T_459 | _T_740 | _T_886; // @[BPU.scala 674:113]
  wire  ghv_write_datas_74 = ghv_write_datas_74_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_75 = _T_198 | _T_460 | _T_741 | _T_887; // @[BPU.scala 674:113]
  wire  ghv_write_datas_75 = ghv_write_datas_75_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_76 = _T_199 | _T_461 | _T_742 | _T_888; // @[BPU.scala 674:113]
  wire  ghv_write_datas_76 = ghv_write_datas_76_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_77 = _T_200 | _T_462 | _T_743 | _T_889; // @[BPU.scala 674:113]
  wire  ghv_write_datas_77 = ghv_write_datas_77_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_78 = _T_201 | _T_463 | _T_744 | _T_890; // @[BPU.scala 674:113]
  wire  ghv_write_datas_78 = ghv_write_datas_78_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_79 = _T_202 | _T_464 | _T_745 | _T_891; // @[BPU.scala 674:113]
  wire  ghv_write_datas_79 = ghv_write_datas_79_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_80 = _T_203 | _T_465 | _T_746 | _T_892; // @[BPU.scala 674:113]
  wire  ghv_write_datas_80 = ghv_write_datas_80_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_81 = _T_204 | _T_466 | _T_747 | _T_893; // @[BPU.scala 674:113]
  wire  ghv_write_datas_81 = ghv_write_datas_81_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_82 = _T_205 | _T_467 | _T_748 | _T_894; // @[BPU.scala 674:113]
  wire  ghv_write_datas_82 = ghv_write_datas_82_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_83 = _T_206 | _T_468 | _T_749 | _T_895; // @[BPU.scala 674:113]
  wire  ghv_write_datas_83 = ghv_write_datas_83_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_84 = _T_207 | _T_469 | _T_750 | _T_896; // @[BPU.scala 674:113]
  wire  ghv_write_datas_84 = ghv_write_datas_84_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_85 = _T_208 | _T_470 | _T_751 | _T_897; // @[BPU.scala 674:113]
  wire  ghv_write_datas_85 = ghv_write_datas_85_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_86 = _T_209 | _T_471 | _T_752 | _T_898; // @[BPU.scala 674:113]
  wire  ghv_write_datas_86 = ghv_write_datas_86_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_87 = _T_210 | _T_472 | _T_753 | _T_899; // @[BPU.scala 674:113]
  wire  ghv_write_datas_87 = ghv_write_datas_87_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_88 = _T_211 | _T_473 | _T_754 | _T_900; // @[BPU.scala 674:113]
  wire  ghv_write_datas_88 = ghv_write_datas_88_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_89 = _T_212 | _T_474 | _T_755 | _T_901; // @[BPU.scala 674:113]
  wire  ghv_write_datas_89 = ghv_write_datas_89_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_90 = _T_213 | _T_475 | _T_756 | _T_902; // @[BPU.scala 674:113]
  wire  ghv_write_datas_90 = ghv_write_datas_90_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_91 = _T_214 | _T_476 | _T_757 | _T_903; // @[BPU.scala 674:113]
  wire  ghv_write_datas_91 = ghv_write_datas_91_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_92 = _T_215 | _T_477 | _T_758 | _T_904; // @[BPU.scala 674:113]
  wire  ghv_write_datas_92 = ghv_write_datas_92_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_93 = _T_216 | _T_478 | _T_759 | _T_905; // @[BPU.scala 674:113]
  wire  ghv_write_datas_93 = ghv_write_datas_93_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_94 = _T_217 | _T_479 | _T_760 | _T_906; // @[BPU.scala 674:113]
  wire  ghv_write_datas_94 = ghv_write_datas_94_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_95 = _T_218 | _T_480 | _T_761 | _T_907; // @[BPU.scala 674:113]
  wire  ghv_write_datas_95 = ghv_write_datas_95_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_96 = _T_219 | _T_481 | _T_762 | _T_908; // @[BPU.scala 674:113]
  wire  ghv_write_datas_96 = ghv_write_datas_96_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_97 = _T_220 | _T_482 | _T_763 | _T_909; // @[BPU.scala 674:113]
  wire  ghv_write_datas_97 = ghv_write_datas_97_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_98 = _T_221 | _T_483 | _T_764 | _T_910; // @[BPU.scala 674:113]
  wire  ghv_write_datas_98 = ghv_write_datas_98_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_99 = _T_222 | _T_484 | _T_765 | _T_911; // @[BPU.scala 674:113]
  wire  ghv_write_datas_99 = ghv_write_datas_99_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_100 = _T_223 | _T_485 | _T_766 | _T_912; // @[BPU.scala 674:113]
  wire  ghv_write_datas_100 = ghv_write_datas_100_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_101 = _T_224 | _T_486 | _T_767 | _T_913; // @[BPU.scala 674:113]
  wire  ghv_write_datas_101 = ghv_write_datas_101_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_102 = _T_225 | _T_487 | _T_768 | _T_914; // @[BPU.scala 674:113]
  wire  ghv_write_datas_102 = ghv_write_datas_102_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_103 = _T_226 | _T_488 | _T_769 | _T_915; // @[BPU.scala 674:113]
  wire  ghv_write_datas_103 = ghv_write_datas_103_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_104 = _T_227 | _T_489 | _T_770 | _T_916; // @[BPU.scala 674:113]
  wire  ghv_write_datas_104 = ghv_write_datas_104_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_105 = _T_228 | _T_490 | _T_771 | _T_917; // @[BPU.scala 674:113]
  wire  ghv_write_datas_105 = ghv_write_datas_105_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_106 = _T_229 | _T_491 | _T_772 | _T_918; // @[BPU.scala 674:113]
  wire  ghv_write_datas_106 = ghv_write_datas_106_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_107 = _T_230 | _T_492 | _T_773 | _T_919; // @[BPU.scala 674:113]
  wire  ghv_write_datas_107 = ghv_write_datas_107_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_108 = _T_231 | _T_493 | _T_774 | _T_920; // @[BPU.scala 674:113]
  wire  ghv_write_datas_108 = ghv_write_datas_108_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_109 = _T_232 | _T_494 | _T_775 | _T_921; // @[BPU.scala 674:113]
  wire  ghv_write_datas_109 = ghv_write_datas_109_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_110 = _T_233 | _T_495 | _T_776 | _T_922; // @[BPU.scala 674:113]
  wire  ghv_write_datas_110 = ghv_write_datas_110_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_111 = _T_234 | _T_496 | _T_777 | _T_923; // @[BPU.scala 674:113]
  wire  ghv_write_datas_111 = ghv_write_datas_111_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_112 = _T_235 | _T_497 | _T_778 | _T_924; // @[BPU.scala 674:113]
  wire  ghv_write_datas_112 = ghv_write_datas_112_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_113 = _T_236 | _T_498 | _T_779 | _T_925; // @[BPU.scala 674:113]
  wire  ghv_write_datas_113 = ghv_write_datas_113_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_114 = _T_237 | _T_499 | _T_780 | _T_926; // @[BPU.scala 674:113]
  wire  ghv_write_datas_114 = ghv_write_datas_114_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_115 = _T_238 | _T_500 | _T_781 | _T_927; // @[BPU.scala 674:113]
  wire  ghv_write_datas_115 = ghv_write_datas_115_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_116 = _T_239 | _T_501 | _T_782 | _T_928; // @[BPU.scala 674:113]
  wire  ghv_write_datas_116 = ghv_write_datas_116_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_117 = _T_240 | _T_502 | _T_783 | _T_929; // @[BPU.scala 674:113]
  wire  ghv_write_datas_117 = ghv_write_datas_117_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_118 = _T_241 | _T_503 | _T_784 | _T_930; // @[BPU.scala 674:113]
  wire  ghv_write_datas_118 = ghv_write_datas_118_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_119 = _T_242 | _T_504 | _T_785 | _T_931; // @[BPU.scala 674:113]
  wire  ghv_write_datas_119 = ghv_write_datas_119_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_120 = _T_243 | _T_505 | _T_786 | _T_932; // @[BPU.scala 674:113]
  wire  ghv_write_datas_120 = ghv_write_datas_120_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_121 = _T_244 | _T_506 | _T_787 | _T_933; // @[BPU.scala 674:113]
  wire  ghv_write_datas_121 = ghv_write_datas_121_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_122 = _T_245 | _T_507 | _T_788 | _T_934; // @[BPU.scala 674:113]
  wire  ghv_write_datas_122 = ghv_write_datas_122_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_123 = _T_246 | _T_508 | _T_789 | _T_935; // @[BPU.scala 674:113]
  wire  ghv_write_datas_123 = ghv_write_datas_123_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_124 = _T_247 | _T_509 | _T_790 | _T_936; // @[BPU.scala 674:113]
  wire  ghv_write_datas_124 = ghv_write_datas_124_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_125 = _T_248 | _T_510 | _T_791 | _T_937; // @[BPU.scala 674:113]
  wire  ghv_write_datas_125 = ghv_write_datas_125_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_126 = _T_249 | _T_511 | _T_792 | _T_938; // @[BPU.scala 674:113]
  wire  ghv_write_datas_126 = ghv_write_datas_126_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_127 = _T_250 | _T_512 | _T_793 | _T_939; // @[BPU.scala 674:113]
  wire  ghv_write_datas_127 = ghv_write_datas_127_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_128 = _T_251 | _T_513 | _T_794 | _T_940; // @[BPU.scala 674:113]
  wire  ghv_write_datas_128 = ghv_write_datas_128_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_129 = _T_252 | _T_514 | _T_795 | _T_941; // @[BPU.scala 674:113]
  wire  ghv_write_datas_129 = ghv_write_datas_129_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_130 = _T_253 | _T_515 | _T_796 | _T_942; // @[BPU.scala 674:113]
  wire  ghv_write_datas_130 = ghv_write_datas_130_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_131 = _T_254 | _T_516 | _T_797 | _T_943; // @[BPU.scala 674:113]
  wire  ghv_write_datas_131 = ghv_write_datas_131_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_132 = _T_255 | _T_517 | _T_798 | _T_944; // @[BPU.scala 674:113]
  wire  ghv_write_datas_132 = ghv_write_datas_132_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_133 = _T_256 | _T_518 | _T_799 | _T_945; // @[BPU.scala 674:113]
  wire  ghv_write_datas_133 = ghv_write_datas_133_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_134 = _T_257 | _T_519 | _T_800 | _T_946; // @[BPU.scala 674:113]
  wire  ghv_write_datas_134 = ghv_write_datas_134_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_135 = _T_258 | _T_520 | _T_801 | _T_947; // @[BPU.scala 674:113]
  wire  ghv_write_datas_135 = ghv_write_datas_135_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_136 = _T_259 | _T_521 | _T_802 | _T_948; // @[BPU.scala 674:113]
  wire  ghv_write_datas_136 = ghv_write_datas_136_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_137 = _T_260 | _T_522 | _T_803 | _T_949; // @[BPU.scala 674:113]
  wire  ghv_write_datas_137 = ghv_write_datas_137_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_138 = _T_261 | _T_523 | _T_804 | _T_950; // @[BPU.scala 674:113]
  wire  ghv_write_datas_138 = ghv_write_datas_138_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_139 = _T_262 | _T_524 | _T_805 | _T_951; // @[BPU.scala 674:113]
  wire  ghv_write_datas_139 = ghv_write_datas_139_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_140 = _T_263 | _T_525 | _T_806 | _T_952; // @[BPU.scala 674:113]
  wire  ghv_write_datas_140 = ghv_write_datas_140_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_141 = _T_264 | _T_526 | _T_807 | _T_953; // @[BPU.scala 674:113]
  wire  ghv_write_datas_141 = ghv_write_datas_141_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_142 = _T_265 | _T_527 | _T_808 | _T_954; // @[BPU.scala 674:113]
  wire  ghv_write_datas_142 = ghv_write_datas_142_ppm_out_res; // @[BPU.scala 300:29 672:64]
  wire  ghv_wens_143 = _T_266 | _T_528 | _T_809 | _T_955; // @[BPU.scala 674:113]
  wire  ghv_write_datas_143 = ghv_write_datas_143_ppm_out_res; // @[BPU.scala 300:29 672:64]
  reg [5:0] io_perf_0_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg [5:0] io_perf_0_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg [5:0] io_perf_1_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg [5:0] io_perf_1_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg [5:0] io_perf_2_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg [5:0] io_perf_2_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg [5:0] io_perf_3_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg [5:0] io_perf_3_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg [5:0] io_perf_4_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg [5:0] io_perf_4_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg [5:0] io_perf_5_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg [5:0] io_perf_5_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg [5:0] io_perf_6_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg [5:0] io_perf_6_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  DelayN_1 ctrl_delay ( // @[Hold.scala 97:23]
    .clock(ctrl_delay_clock),
    .io_in_ubtb_enable(ctrl_delay_io_in_ubtb_enable),
    .io_in_btb_enable(ctrl_delay_io_in_btb_enable),
    .io_in_tage_enable(ctrl_delay_io_in_tage_enable),
    .io_in_sc_enable(ctrl_delay_io_in_sc_enable),
    .io_in_ras_enable(ctrl_delay_io_in_ras_enable),
    .io_out_ubtb_enable(ctrl_delay_io_out_ubtb_enable),
    .io_out_btb_enable(ctrl_delay_io_out_btb_enable),
    .io_out_tage_enable(ctrl_delay_io_out_tage_enable),
    .io_out_sc_enable(ctrl_delay_io_out_sc_enable),
    .io_out_ras_enable(ctrl_delay_io_out_ras_enable)
  );
  Composer predictors ( // @[BPU.scala 245:26]
    .clock(predictors_clock),
    .reset(predictors_reset),
    .io_reset_vector(predictors_io_reset_vector),
    .io_in_bits_s0_pc(predictors_io_in_bits_s0_pc),
    .io_in_bits_folded_hist_hist_17_folded_hist(predictors_io_in_bits_folded_hist_hist_17_folded_hist),
    .io_in_bits_folded_hist_hist_16_folded_hist(predictors_io_in_bits_folded_hist_hist_16_folded_hist),
    .io_in_bits_folded_hist_hist_15_folded_hist(predictors_io_in_bits_folded_hist_hist_15_folded_hist),
    .io_in_bits_folded_hist_hist_14_folded_hist(predictors_io_in_bits_folded_hist_hist_14_folded_hist),
    .io_in_bits_folded_hist_hist_13_folded_hist(predictors_io_in_bits_folded_hist_hist_13_folded_hist),
    .io_in_bits_folded_hist_hist_12_folded_hist(predictors_io_in_bits_folded_hist_hist_12_folded_hist),
    .io_in_bits_folded_hist_hist_10_folded_hist(predictors_io_in_bits_folded_hist_hist_10_folded_hist),
    .io_in_bits_folded_hist_hist_9_folded_hist(predictors_io_in_bits_folded_hist_hist_9_folded_hist),
    .io_in_bits_folded_hist_hist_8_folded_hist(predictors_io_in_bits_folded_hist_hist_8_folded_hist),
    .io_in_bits_folded_hist_hist_7_folded_hist(predictors_io_in_bits_folded_hist_hist_7_folded_hist),
    .io_in_bits_folded_hist_hist_6_folded_hist(predictors_io_in_bits_folded_hist_hist_6_folded_hist),
    .io_in_bits_folded_hist_hist_5_folded_hist(predictors_io_in_bits_folded_hist_hist_5_folded_hist),
    .io_in_bits_folded_hist_hist_4_folded_hist(predictors_io_in_bits_folded_hist_hist_4_folded_hist),
    .io_in_bits_folded_hist_hist_3_folded_hist(predictors_io_in_bits_folded_hist_hist_3_folded_hist),
    .io_in_bits_folded_hist_hist_2_folded_hist(predictors_io_in_bits_folded_hist_hist_2_folded_hist),
    .io_in_bits_folded_hist_hist_1_folded_hist(predictors_io_in_bits_folded_hist_hist_1_folded_hist),
    .io_in_bits_folded_hist_hist_0_folded_hist(predictors_io_in_bits_folded_hist_hist_0_folded_hist),
    .io_out_s1_pc(predictors_io_out_s1_pc),
    .io_out_s1_full_pred_br_taken_mask_0(predictors_io_out_s1_full_pred_br_taken_mask_0),
    .io_out_s1_full_pred_br_taken_mask_1(predictors_io_out_s1_full_pred_br_taken_mask_1),
    .io_out_s1_full_pred_slot_valids_0(predictors_io_out_s1_full_pred_slot_valids_0),
    .io_out_s1_full_pred_slot_valids_1(predictors_io_out_s1_full_pred_slot_valids_1),
    .io_out_s1_full_pred_targets_0(predictors_io_out_s1_full_pred_targets_0),
    .io_out_s1_full_pred_targets_1(predictors_io_out_s1_full_pred_targets_1),
    .io_out_s1_full_pred_offsets_0(predictors_io_out_s1_full_pred_offsets_0),
    .io_out_s1_full_pred_offsets_1(predictors_io_out_s1_full_pred_offsets_1),
    .io_out_s1_full_pred_fallThroughAddr(predictors_io_out_s1_full_pred_fallThroughAddr),
    .io_out_s1_full_pred_fallThroughErr(predictors_io_out_s1_full_pred_fallThroughErr),
    .io_out_s1_full_pred_is_br_sharing(predictors_io_out_s1_full_pred_is_br_sharing),
    .io_out_s1_full_pred_hit(predictors_io_out_s1_full_pred_hit),
    .io_out_s2_pc(predictors_io_out_s2_pc),
    .io_out_s2_full_pred_br_taken_mask_0(predictors_io_out_s2_full_pred_br_taken_mask_0),
    .io_out_s2_full_pred_br_taken_mask_1(predictors_io_out_s2_full_pred_br_taken_mask_1),
    .io_out_s2_full_pred_slot_valids_0(predictors_io_out_s2_full_pred_slot_valids_0),
    .io_out_s2_full_pred_slot_valids_1(predictors_io_out_s2_full_pred_slot_valids_1),
    .io_out_s2_full_pred_targets_0(predictors_io_out_s2_full_pred_targets_0),
    .io_out_s2_full_pred_targets_1(predictors_io_out_s2_full_pred_targets_1),
    .io_out_s2_full_pred_offsets_0(predictors_io_out_s2_full_pred_offsets_0),
    .io_out_s2_full_pred_offsets_1(predictors_io_out_s2_full_pred_offsets_1),
    .io_out_s2_full_pred_fallThroughAddr(predictors_io_out_s2_full_pred_fallThroughAddr),
    .io_out_s2_full_pred_fallThroughErr(predictors_io_out_s2_full_pred_fallThroughErr),
    .io_out_s2_full_pred_is_br_sharing(predictors_io_out_s2_full_pred_is_br_sharing),
    .io_out_s2_full_pred_hit(predictors_io_out_s2_full_pred_hit),
    .io_out_s3_pc(predictors_io_out_s3_pc),
    .io_out_s3_full_pred_br_taken_mask_0(predictors_io_out_s3_full_pred_br_taken_mask_0),
    .io_out_s3_full_pred_br_taken_mask_1(predictors_io_out_s3_full_pred_br_taken_mask_1),
    .io_out_s3_full_pred_slot_valids_0(predictors_io_out_s3_full_pred_slot_valids_0),
    .io_out_s3_full_pred_slot_valids_1(predictors_io_out_s3_full_pred_slot_valids_1),
    .io_out_s3_full_pred_targets_0(predictors_io_out_s3_full_pred_targets_0),
    .io_out_s3_full_pred_targets_1(predictors_io_out_s3_full_pred_targets_1),
    .io_out_s3_full_pred_offsets_0(predictors_io_out_s3_full_pred_offsets_0),
    .io_out_s3_full_pred_offsets_1(predictors_io_out_s3_full_pred_offsets_1),
    .io_out_s3_full_pred_fallThroughAddr(predictors_io_out_s3_full_pred_fallThroughAddr),
    .io_out_s3_full_pred_fallThroughErr(predictors_io_out_s3_full_pred_fallThroughErr),
    .io_out_s3_full_pred_is_br_sharing(predictors_io_out_s3_full_pred_is_br_sharing),
    .io_out_s3_full_pred_hit(predictors_io_out_s3_full_pred_hit),
    .io_out_last_stage_meta(predictors_io_out_last_stage_meta),
    .io_out_last_stage_spec_info_rasSp(predictors_io_out_last_stage_spec_info_rasSp),
    .io_out_last_stage_spec_info_rasTop_retAddr(predictors_io_out_last_stage_spec_info_rasTop_retAddr),
    .io_out_last_stage_spec_info_rasTop_ctr(predictors_io_out_last_stage_spec_info_rasTop_ctr),
    .io_out_last_stage_ftb_entry_valid(predictors_io_out_last_stage_ftb_entry_valid),
    .io_out_last_stage_ftb_entry_brSlots_0_offset(predictors_io_out_last_stage_ftb_entry_brSlots_0_offset),
    .io_out_last_stage_ftb_entry_brSlots_0_lower(predictors_io_out_last_stage_ftb_entry_brSlots_0_lower),
    .io_out_last_stage_ftb_entry_brSlots_0_tarStat(predictors_io_out_last_stage_ftb_entry_brSlots_0_tarStat),
    .io_out_last_stage_ftb_entry_brSlots_0_sharing(predictors_io_out_last_stage_ftb_entry_brSlots_0_sharing),
    .io_out_last_stage_ftb_entry_brSlots_0_valid(predictors_io_out_last_stage_ftb_entry_brSlots_0_valid),
    .io_out_last_stage_ftb_entry_tailSlot_offset(predictors_io_out_last_stage_ftb_entry_tailSlot_offset),
    .io_out_last_stage_ftb_entry_tailSlot_lower(predictors_io_out_last_stage_ftb_entry_tailSlot_lower),
    .io_out_last_stage_ftb_entry_tailSlot_tarStat(predictors_io_out_last_stage_ftb_entry_tailSlot_tarStat),
    .io_out_last_stage_ftb_entry_tailSlot_sharing(predictors_io_out_last_stage_ftb_entry_tailSlot_sharing),
    .io_out_last_stage_ftb_entry_tailSlot_valid(predictors_io_out_last_stage_ftb_entry_tailSlot_valid),
    .io_out_last_stage_ftb_entry_pftAddr(predictors_io_out_last_stage_ftb_entry_pftAddr),
    .io_out_last_stage_ftb_entry_carry(predictors_io_out_last_stage_ftb_entry_carry),
    .io_out_last_stage_ftb_entry_isCall(predictors_io_out_last_stage_ftb_entry_isCall),
    .io_out_last_stage_ftb_entry_isRet(predictors_io_out_last_stage_ftb_entry_isRet),
    .io_out_last_stage_ftb_entry_isJalr(predictors_io_out_last_stage_ftb_entry_isJalr),
    .io_out_last_stage_ftb_entry_last_may_be_rvi_call(predictors_io_out_last_stage_ftb_entry_last_may_be_rvi_call),
    .io_out_last_stage_ftb_entry_always_taken_0(predictors_io_out_last_stage_ftb_entry_always_taken_0),
    .io_out_last_stage_ftb_entry_always_taken_1(predictors_io_out_last_stage_ftb_entry_always_taken_1),
    .io_ctrl_ubtb_enable(predictors_io_ctrl_ubtb_enable),
    .io_ctrl_btb_enable(predictors_io_ctrl_btb_enable),
    .io_ctrl_tage_enable(predictors_io_ctrl_tage_enable),
    .io_ctrl_sc_enable(predictors_io_ctrl_sc_enable),
    .io_ctrl_ras_enable(predictors_io_ctrl_ras_enable),
    .io_s0_fire(predictors_io_s0_fire),
    .io_s1_fire(predictors_io_s1_fire),
    .io_s2_fire(predictors_io_s2_fire),
    .io_s3_fire(predictors_io_s3_fire),
    .io_s3_redirect(predictors_io_s3_redirect),
    .io_s1_ready(predictors_io_s1_ready),
    .io_update_valid(predictors_io_update_valid),
    .io_update_bits_pc(predictors_io_update_bits_pc),
    .io_update_bits_spec_info_folded_hist_hist_17_folded_hist(
      predictors_io_update_bits_spec_info_folded_hist_hist_17_folded_hist),
    .io_update_bits_spec_info_folded_hist_hist_16_folded_hist(
      predictors_io_update_bits_spec_info_folded_hist_hist_16_folded_hist),
    .io_update_bits_spec_info_folded_hist_hist_15_folded_hist(
      predictors_io_update_bits_spec_info_folded_hist_hist_15_folded_hist),
    .io_update_bits_spec_info_folded_hist_hist_14_folded_hist(
      predictors_io_update_bits_spec_info_folded_hist_hist_14_folded_hist),
    .io_update_bits_spec_info_folded_hist_hist_13_folded_hist(
      predictors_io_update_bits_spec_info_folded_hist_hist_13_folded_hist),
    .io_update_bits_spec_info_folded_hist_hist_12_folded_hist(
      predictors_io_update_bits_spec_info_folded_hist_hist_12_folded_hist),
    .io_update_bits_spec_info_folded_hist_hist_10_folded_hist(
      predictors_io_update_bits_spec_info_folded_hist_hist_10_folded_hist),
    .io_update_bits_spec_info_folded_hist_hist_9_folded_hist(
      predictors_io_update_bits_spec_info_folded_hist_hist_9_folded_hist),
    .io_update_bits_spec_info_folded_hist_hist_8_folded_hist(
      predictors_io_update_bits_spec_info_folded_hist_hist_8_folded_hist),
    .io_update_bits_spec_info_folded_hist_hist_7_folded_hist(
      predictors_io_update_bits_spec_info_folded_hist_hist_7_folded_hist),
    .io_update_bits_spec_info_folded_hist_hist_6_folded_hist(
      predictors_io_update_bits_spec_info_folded_hist_hist_6_folded_hist),
    .io_update_bits_spec_info_folded_hist_hist_5_folded_hist(
      predictors_io_update_bits_spec_info_folded_hist_hist_5_folded_hist),
    .io_update_bits_spec_info_folded_hist_hist_4_folded_hist(
      predictors_io_update_bits_spec_info_folded_hist_hist_4_folded_hist),
    .io_update_bits_spec_info_folded_hist_hist_3_folded_hist(
      predictors_io_update_bits_spec_info_folded_hist_hist_3_folded_hist),
    .io_update_bits_spec_info_folded_hist_hist_2_folded_hist(
      predictors_io_update_bits_spec_info_folded_hist_hist_2_folded_hist),
    .io_update_bits_spec_info_folded_hist_hist_1_folded_hist(
      predictors_io_update_bits_spec_info_folded_hist_hist_1_folded_hist),
    .io_update_bits_spec_info_folded_hist_hist_0_folded_hist(
      predictors_io_update_bits_spec_info_folded_hist_hist_0_folded_hist),
    .io_update_bits_ftb_entry_valid(predictors_io_update_bits_ftb_entry_valid),
    .io_update_bits_ftb_entry_brSlots_0_offset(predictors_io_update_bits_ftb_entry_brSlots_0_offset),
    .io_update_bits_ftb_entry_brSlots_0_lower(predictors_io_update_bits_ftb_entry_brSlots_0_lower),
    .io_update_bits_ftb_entry_brSlots_0_tarStat(predictors_io_update_bits_ftb_entry_brSlots_0_tarStat),
    .io_update_bits_ftb_entry_brSlots_0_sharing(predictors_io_update_bits_ftb_entry_brSlots_0_sharing),
    .io_update_bits_ftb_entry_brSlots_0_valid(predictors_io_update_bits_ftb_entry_brSlots_0_valid),
    .io_update_bits_ftb_entry_tailSlot_offset(predictors_io_update_bits_ftb_entry_tailSlot_offset),
    .io_update_bits_ftb_entry_tailSlot_lower(predictors_io_update_bits_ftb_entry_tailSlot_lower),
    .io_update_bits_ftb_entry_tailSlot_tarStat(predictors_io_update_bits_ftb_entry_tailSlot_tarStat),
    .io_update_bits_ftb_entry_tailSlot_sharing(predictors_io_update_bits_ftb_entry_tailSlot_sharing),
    .io_update_bits_ftb_entry_tailSlot_valid(predictors_io_update_bits_ftb_entry_tailSlot_valid),
    .io_update_bits_ftb_entry_pftAddr(predictors_io_update_bits_ftb_entry_pftAddr),
    .io_update_bits_ftb_entry_carry(predictors_io_update_bits_ftb_entry_carry),
    .io_update_bits_ftb_entry_isCall(predictors_io_update_bits_ftb_entry_isCall),
    .io_update_bits_ftb_entry_isRet(predictors_io_update_bits_ftb_entry_isRet),
    .io_update_bits_ftb_entry_isJalr(predictors_io_update_bits_ftb_entry_isJalr),
    .io_update_bits_ftb_entry_last_may_be_rvi_call(predictors_io_update_bits_ftb_entry_last_may_be_rvi_call),
    .io_update_bits_ftb_entry_always_taken_0(predictors_io_update_bits_ftb_entry_always_taken_0),
    .io_update_bits_ftb_entry_always_taken_1(predictors_io_update_bits_ftb_entry_always_taken_1),
    .io_update_bits_br_taken_mask_0(predictors_io_update_bits_br_taken_mask_0),
    .io_update_bits_br_taken_mask_1(predictors_io_update_bits_br_taken_mask_1),
    .io_update_bits_jmp_taken(predictors_io_update_bits_jmp_taken),
    .io_update_bits_mispred_mask_0(predictors_io_update_bits_mispred_mask_0),
    .io_update_bits_mispred_mask_1(predictors_io_update_bits_mispred_mask_1),
    .io_update_bits_mispred_mask_2(predictors_io_update_bits_mispred_mask_2),
    .io_update_bits_old_entry(predictors_io_update_bits_old_entry),
    .io_update_bits_meta(predictors_io_update_bits_meta),
    .io_update_bits_full_target(predictors_io_update_bits_full_target),
    .io_redirect_valid(predictors_io_redirect_valid),
    .io_redirect_bits_level(predictors_io_redirect_bits_level),
    .io_redirect_bits_cfiUpdate_pc(predictors_io_redirect_bits_cfiUpdate_pc),
    .io_redirect_bits_cfiUpdate_pd_isRVC(predictors_io_redirect_bits_cfiUpdate_pd_isRVC),
    .io_redirect_bits_cfiUpdate_pd_isCall(predictors_io_redirect_bits_cfiUpdate_pd_isCall),
    .io_redirect_bits_cfiUpdate_pd_isRet(predictors_io_redirect_bits_cfiUpdate_pd_isRet),
    .io_redirect_bits_cfiUpdate_rasSp(predictors_io_redirect_bits_cfiUpdate_rasSp),
    .io_redirect_bits_cfiUpdate_rasEntry_retAddr(predictors_io_redirect_bits_cfiUpdate_rasEntry_retAddr),
    .io_redirect_bits_cfiUpdate_rasEntry_ctr(predictors_io_redirect_bits_cfiUpdate_rasEntry_ctr),
    .io_perf_0_value(predictors_io_perf_0_value),
    .io_perf_1_value(predictors_io_perf_1_value),
    .io_perf_2_value(predictors_io_perf_2_value),
    .io_perf_3_value(predictors_io_perf_3_value),
    .io_perf_4_value(predictors_io_perf_4_value),
    .io_perf_5_value(predictors_io_perf_5_value),
    .io_perf_6_value(predictors_io_perf_6_value)
  );
  DelayN_2 reset_vector_delay ( // @[Hold.scala 97:23]
    .clock(reset_vector_delay_clock),
    .io_in(reset_vector_delay_io_in),
    .io_out(reset_vector_delay_io_out)
  );
  PriorityMuxModule s0_pc_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_target_sel(s0_pc_ppm_s2_target_sel),
    .s2_target_src(s0_pc_ppm_s2_target_src),
    .s1_target_sel(s0_pc_ppm_s1_target_sel),
    .s1_target_src(s0_pc_ppm_s1_target_src),
    .s3_target_sel(s0_pc_ppm_s3_target_sel),
    .s3_target_src(s0_pc_ppm_s3_target_src),
    .redirect_target_sel(s0_pc_ppm_redirect_target_sel),
    .redirect_target_src(s0_pc_ppm_redirect_target_src),
    .stallPC_src(s0_pc_ppm_stallPC_src),
    .out_res(s0_pc_ppm_out_res)
  );
  PriorityMuxModule_1 s0_folded_gh_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_FGH_sel(s0_folded_gh_ppm_s2_FGH_sel),
    .s2_FGH_src_hist_17_folded_hist(s0_folded_gh_ppm_s2_FGH_src_hist_17_folded_hist),
    .s2_FGH_src_hist_16_folded_hist(s0_folded_gh_ppm_s2_FGH_src_hist_16_folded_hist),
    .s2_FGH_src_hist_15_folded_hist(s0_folded_gh_ppm_s2_FGH_src_hist_15_folded_hist),
    .s2_FGH_src_hist_14_folded_hist(s0_folded_gh_ppm_s2_FGH_src_hist_14_folded_hist),
    .s2_FGH_src_hist_13_folded_hist(s0_folded_gh_ppm_s2_FGH_src_hist_13_folded_hist),
    .s2_FGH_src_hist_12_folded_hist(s0_folded_gh_ppm_s2_FGH_src_hist_12_folded_hist),
    .s2_FGH_src_hist_11_folded_hist(s0_folded_gh_ppm_s2_FGH_src_hist_11_folded_hist),
    .s2_FGH_src_hist_10_folded_hist(s0_folded_gh_ppm_s2_FGH_src_hist_10_folded_hist),
    .s2_FGH_src_hist_9_folded_hist(s0_folded_gh_ppm_s2_FGH_src_hist_9_folded_hist),
    .s2_FGH_src_hist_8_folded_hist(s0_folded_gh_ppm_s2_FGH_src_hist_8_folded_hist),
    .s2_FGH_src_hist_7_folded_hist(s0_folded_gh_ppm_s2_FGH_src_hist_7_folded_hist),
    .s2_FGH_src_hist_6_folded_hist(s0_folded_gh_ppm_s2_FGH_src_hist_6_folded_hist),
    .s2_FGH_src_hist_5_folded_hist(s0_folded_gh_ppm_s2_FGH_src_hist_5_folded_hist),
    .s2_FGH_src_hist_4_folded_hist(s0_folded_gh_ppm_s2_FGH_src_hist_4_folded_hist),
    .s2_FGH_src_hist_3_folded_hist(s0_folded_gh_ppm_s2_FGH_src_hist_3_folded_hist),
    .s2_FGH_src_hist_2_folded_hist(s0_folded_gh_ppm_s2_FGH_src_hist_2_folded_hist),
    .s2_FGH_src_hist_1_folded_hist(s0_folded_gh_ppm_s2_FGH_src_hist_1_folded_hist),
    .s2_FGH_src_hist_0_folded_hist(s0_folded_gh_ppm_s2_FGH_src_hist_0_folded_hist),
    .s1_FGH_sel(s0_folded_gh_ppm_s1_FGH_sel),
    .s1_FGH_src_hist_17_folded_hist(s0_folded_gh_ppm_s1_FGH_src_hist_17_folded_hist),
    .s1_FGH_src_hist_16_folded_hist(s0_folded_gh_ppm_s1_FGH_src_hist_16_folded_hist),
    .s1_FGH_src_hist_15_folded_hist(s0_folded_gh_ppm_s1_FGH_src_hist_15_folded_hist),
    .s1_FGH_src_hist_14_folded_hist(s0_folded_gh_ppm_s1_FGH_src_hist_14_folded_hist),
    .s1_FGH_src_hist_13_folded_hist(s0_folded_gh_ppm_s1_FGH_src_hist_13_folded_hist),
    .s1_FGH_src_hist_12_folded_hist(s0_folded_gh_ppm_s1_FGH_src_hist_12_folded_hist),
    .s1_FGH_src_hist_11_folded_hist(s0_folded_gh_ppm_s1_FGH_src_hist_11_folded_hist),
    .s1_FGH_src_hist_10_folded_hist(s0_folded_gh_ppm_s1_FGH_src_hist_10_folded_hist),
    .s1_FGH_src_hist_9_folded_hist(s0_folded_gh_ppm_s1_FGH_src_hist_9_folded_hist),
    .s1_FGH_src_hist_8_folded_hist(s0_folded_gh_ppm_s1_FGH_src_hist_8_folded_hist),
    .s1_FGH_src_hist_7_folded_hist(s0_folded_gh_ppm_s1_FGH_src_hist_7_folded_hist),
    .s1_FGH_src_hist_6_folded_hist(s0_folded_gh_ppm_s1_FGH_src_hist_6_folded_hist),
    .s1_FGH_src_hist_5_folded_hist(s0_folded_gh_ppm_s1_FGH_src_hist_5_folded_hist),
    .s1_FGH_src_hist_4_folded_hist(s0_folded_gh_ppm_s1_FGH_src_hist_4_folded_hist),
    .s1_FGH_src_hist_3_folded_hist(s0_folded_gh_ppm_s1_FGH_src_hist_3_folded_hist),
    .s1_FGH_src_hist_2_folded_hist(s0_folded_gh_ppm_s1_FGH_src_hist_2_folded_hist),
    .s1_FGH_src_hist_1_folded_hist(s0_folded_gh_ppm_s1_FGH_src_hist_1_folded_hist),
    .s1_FGH_src_hist_0_folded_hist(s0_folded_gh_ppm_s1_FGH_src_hist_0_folded_hist),
    .s3_FGH_sel(s0_folded_gh_ppm_s3_FGH_sel),
    .s3_FGH_src_hist_17_folded_hist(s0_folded_gh_ppm_s3_FGH_src_hist_17_folded_hist),
    .s3_FGH_src_hist_16_folded_hist(s0_folded_gh_ppm_s3_FGH_src_hist_16_folded_hist),
    .s3_FGH_src_hist_15_folded_hist(s0_folded_gh_ppm_s3_FGH_src_hist_15_folded_hist),
    .s3_FGH_src_hist_14_folded_hist(s0_folded_gh_ppm_s3_FGH_src_hist_14_folded_hist),
    .s3_FGH_src_hist_13_folded_hist(s0_folded_gh_ppm_s3_FGH_src_hist_13_folded_hist),
    .s3_FGH_src_hist_12_folded_hist(s0_folded_gh_ppm_s3_FGH_src_hist_12_folded_hist),
    .s3_FGH_src_hist_11_folded_hist(s0_folded_gh_ppm_s3_FGH_src_hist_11_folded_hist),
    .s3_FGH_src_hist_10_folded_hist(s0_folded_gh_ppm_s3_FGH_src_hist_10_folded_hist),
    .s3_FGH_src_hist_9_folded_hist(s0_folded_gh_ppm_s3_FGH_src_hist_9_folded_hist),
    .s3_FGH_src_hist_8_folded_hist(s0_folded_gh_ppm_s3_FGH_src_hist_8_folded_hist),
    .s3_FGH_src_hist_7_folded_hist(s0_folded_gh_ppm_s3_FGH_src_hist_7_folded_hist),
    .s3_FGH_src_hist_6_folded_hist(s0_folded_gh_ppm_s3_FGH_src_hist_6_folded_hist),
    .s3_FGH_src_hist_5_folded_hist(s0_folded_gh_ppm_s3_FGH_src_hist_5_folded_hist),
    .s3_FGH_src_hist_4_folded_hist(s0_folded_gh_ppm_s3_FGH_src_hist_4_folded_hist),
    .s3_FGH_src_hist_3_folded_hist(s0_folded_gh_ppm_s3_FGH_src_hist_3_folded_hist),
    .s3_FGH_src_hist_2_folded_hist(s0_folded_gh_ppm_s3_FGH_src_hist_2_folded_hist),
    .s3_FGH_src_hist_1_folded_hist(s0_folded_gh_ppm_s3_FGH_src_hist_1_folded_hist),
    .s3_FGH_src_hist_0_folded_hist(s0_folded_gh_ppm_s3_FGH_src_hist_0_folded_hist),
    .redirect_FGHT_sel(s0_folded_gh_ppm_redirect_FGHT_sel),
    .redirect_FGHT_src_hist_17_folded_hist(s0_folded_gh_ppm_redirect_FGHT_src_hist_17_folded_hist),
    .redirect_FGHT_src_hist_16_folded_hist(s0_folded_gh_ppm_redirect_FGHT_src_hist_16_folded_hist),
    .redirect_FGHT_src_hist_15_folded_hist(s0_folded_gh_ppm_redirect_FGHT_src_hist_15_folded_hist),
    .redirect_FGHT_src_hist_14_folded_hist(s0_folded_gh_ppm_redirect_FGHT_src_hist_14_folded_hist),
    .redirect_FGHT_src_hist_13_folded_hist(s0_folded_gh_ppm_redirect_FGHT_src_hist_13_folded_hist),
    .redirect_FGHT_src_hist_12_folded_hist(s0_folded_gh_ppm_redirect_FGHT_src_hist_12_folded_hist),
    .redirect_FGHT_src_hist_11_folded_hist(s0_folded_gh_ppm_redirect_FGHT_src_hist_11_folded_hist),
    .redirect_FGHT_src_hist_10_folded_hist(s0_folded_gh_ppm_redirect_FGHT_src_hist_10_folded_hist),
    .redirect_FGHT_src_hist_9_folded_hist(s0_folded_gh_ppm_redirect_FGHT_src_hist_9_folded_hist),
    .redirect_FGHT_src_hist_8_folded_hist(s0_folded_gh_ppm_redirect_FGHT_src_hist_8_folded_hist),
    .redirect_FGHT_src_hist_7_folded_hist(s0_folded_gh_ppm_redirect_FGHT_src_hist_7_folded_hist),
    .redirect_FGHT_src_hist_6_folded_hist(s0_folded_gh_ppm_redirect_FGHT_src_hist_6_folded_hist),
    .redirect_FGHT_src_hist_5_folded_hist(s0_folded_gh_ppm_redirect_FGHT_src_hist_5_folded_hist),
    .redirect_FGHT_src_hist_4_folded_hist(s0_folded_gh_ppm_redirect_FGHT_src_hist_4_folded_hist),
    .redirect_FGHT_src_hist_3_folded_hist(s0_folded_gh_ppm_redirect_FGHT_src_hist_3_folded_hist),
    .redirect_FGHT_src_hist_2_folded_hist(s0_folded_gh_ppm_redirect_FGHT_src_hist_2_folded_hist),
    .redirect_FGHT_src_hist_1_folded_hist(s0_folded_gh_ppm_redirect_FGHT_src_hist_1_folded_hist),
    .redirect_FGHT_src_hist_0_folded_hist(s0_folded_gh_ppm_redirect_FGHT_src_hist_0_folded_hist),
    .stallFGH_src_hist_17_folded_hist(s0_folded_gh_ppm_stallFGH_src_hist_17_folded_hist),
    .stallFGH_src_hist_16_folded_hist(s0_folded_gh_ppm_stallFGH_src_hist_16_folded_hist),
    .stallFGH_src_hist_15_folded_hist(s0_folded_gh_ppm_stallFGH_src_hist_15_folded_hist),
    .stallFGH_src_hist_14_folded_hist(s0_folded_gh_ppm_stallFGH_src_hist_14_folded_hist),
    .stallFGH_src_hist_13_folded_hist(s0_folded_gh_ppm_stallFGH_src_hist_13_folded_hist),
    .stallFGH_src_hist_12_folded_hist(s0_folded_gh_ppm_stallFGH_src_hist_12_folded_hist),
    .stallFGH_src_hist_11_folded_hist(s0_folded_gh_ppm_stallFGH_src_hist_11_folded_hist),
    .stallFGH_src_hist_10_folded_hist(s0_folded_gh_ppm_stallFGH_src_hist_10_folded_hist),
    .stallFGH_src_hist_9_folded_hist(s0_folded_gh_ppm_stallFGH_src_hist_9_folded_hist),
    .stallFGH_src_hist_8_folded_hist(s0_folded_gh_ppm_stallFGH_src_hist_8_folded_hist),
    .stallFGH_src_hist_7_folded_hist(s0_folded_gh_ppm_stallFGH_src_hist_7_folded_hist),
    .stallFGH_src_hist_6_folded_hist(s0_folded_gh_ppm_stallFGH_src_hist_6_folded_hist),
    .stallFGH_src_hist_5_folded_hist(s0_folded_gh_ppm_stallFGH_src_hist_5_folded_hist),
    .stallFGH_src_hist_4_folded_hist(s0_folded_gh_ppm_stallFGH_src_hist_4_folded_hist),
    .stallFGH_src_hist_3_folded_hist(s0_folded_gh_ppm_stallFGH_src_hist_3_folded_hist),
    .stallFGH_src_hist_2_folded_hist(s0_folded_gh_ppm_stallFGH_src_hist_2_folded_hist),
    .stallFGH_src_hist_1_folded_hist(s0_folded_gh_ppm_stallFGH_src_hist_1_folded_hist),
    .stallFGH_src_hist_0_folded_hist(s0_folded_gh_ppm_stallFGH_src_hist_0_folded_hist),
    .out_res_hist_17_folded_hist(s0_folded_gh_ppm_out_res_hist_17_folded_hist),
    .out_res_hist_16_folded_hist(s0_folded_gh_ppm_out_res_hist_16_folded_hist),
    .out_res_hist_15_folded_hist(s0_folded_gh_ppm_out_res_hist_15_folded_hist),
    .out_res_hist_14_folded_hist(s0_folded_gh_ppm_out_res_hist_14_folded_hist),
    .out_res_hist_13_folded_hist(s0_folded_gh_ppm_out_res_hist_13_folded_hist),
    .out_res_hist_12_folded_hist(s0_folded_gh_ppm_out_res_hist_12_folded_hist),
    .out_res_hist_11_folded_hist(s0_folded_gh_ppm_out_res_hist_11_folded_hist),
    .out_res_hist_10_folded_hist(s0_folded_gh_ppm_out_res_hist_10_folded_hist),
    .out_res_hist_9_folded_hist(s0_folded_gh_ppm_out_res_hist_9_folded_hist),
    .out_res_hist_8_folded_hist(s0_folded_gh_ppm_out_res_hist_8_folded_hist),
    .out_res_hist_7_folded_hist(s0_folded_gh_ppm_out_res_hist_7_folded_hist),
    .out_res_hist_6_folded_hist(s0_folded_gh_ppm_out_res_hist_6_folded_hist),
    .out_res_hist_5_folded_hist(s0_folded_gh_ppm_out_res_hist_5_folded_hist),
    .out_res_hist_4_folded_hist(s0_folded_gh_ppm_out_res_hist_4_folded_hist),
    .out_res_hist_3_folded_hist(s0_folded_gh_ppm_out_res_hist_3_folded_hist),
    .out_res_hist_2_folded_hist(s0_folded_gh_ppm_out_res_hist_2_folded_hist),
    .out_res_hist_1_folded_hist(s0_folded_gh_ppm_out_res_hist_1_folded_hist),
    .out_res_hist_0_folded_hist(s0_folded_gh_ppm_out_res_hist_0_folded_hist)
  );
  PriorityMuxModule_2 s0_ghist_ptr_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_GHPtr_sel(s0_ghist_ptr_ppm_s2_GHPtr_sel),
    .s2_GHPtr_src_flag(s0_ghist_ptr_ppm_s2_GHPtr_src_flag),
    .s2_GHPtr_src_value(s0_ghist_ptr_ppm_s2_GHPtr_src_value),
    .s1_GHPtr_sel(s0_ghist_ptr_ppm_s1_GHPtr_sel),
    .s1_GHPtr_src_flag(s0_ghist_ptr_ppm_s1_GHPtr_src_flag),
    .s1_GHPtr_src_value(s0_ghist_ptr_ppm_s1_GHPtr_src_value),
    .s3_GHPtr_sel(s0_ghist_ptr_ppm_s3_GHPtr_sel),
    .s3_GHPtr_src_flag(s0_ghist_ptr_ppm_s3_GHPtr_src_flag),
    .s3_GHPtr_src_value(s0_ghist_ptr_ppm_s3_GHPtr_src_value),
    .redirect_GHPtr_sel(s0_ghist_ptr_ppm_redirect_GHPtr_sel),
    .redirect_GHPtr_src_flag(s0_ghist_ptr_ppm_redirect_GHPtr_src_flag),
    .redirect_GHPtr_src_value(s0_ghist_ptr_ppm_redirect_GHPtr_src_value),
    .stallGHPtr_src_flag(s0_ghist_ptr_ppm_stallGHPtr_src_flag),
    .stallGHPtr_src_value(s0_ghist_ptr_ppm_stallGHPtr_src_value),
    .out_res_flag(s0_ghist_ptr_ppm_out_res_flag),
    .out_res_value(s0_ghist_ptr_ppm_out_res_value)
  );
  PriorityMuxModule_3 s0_ahead_fh_oldest_bits_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_AFHOB_sel(s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_sel),
    .s2_AFHOB_src_afhob_5_bits_0(s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_src_afhob_5_bits_0),
    .s2_AFHOB_src_afhob_5_bits_1(s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_src_afhob_5_bits_1),
    .s2_AFHOB_src_afhob_5_bits_2(s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_src_afhob_5_bits_2),
    .s2_AFHOB_src_afhob_5_bits_3(s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_src_afhob_5_bits_3),
    .s2_AFHOB_src_afhob_4_bits_0(s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_src_afhob_4_bits_0),
    .s2_AFHOB_src_afhob_4_bits_1(s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_src_afhob_4_bits_1),
    .s2_AFHOB_src_afhob_4_bits_2(s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_src_afhob_4_bits_2),
    .s2_AFHOB_src_afhob_4_bits_3(s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_src_afhob_4_bits_3),
    .s2_AFHOB_src_afhob_3_bits_0(s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_src_afhob_3_bits_0),
    .s2_AFHOB_src_afhob_3_bits_1(s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_src_afhob_3_bits_1),
    .s2_AFHOB_src_afhob_3_bits_2(s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_src_afhob_3_bits_2),
    .s2_AFHOB_src_afhob_3_bits_3(s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_src_afhob_3_bits_3),
    .s2_AFHOB_src_afhob_2_bits_0(s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_src_afhob_2_bits_0),
    .s2_AFHOB_src_afhob_2_bits_1(s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_src_afhob_2_bits_1),
    .s2_AFHOB_src_afhob_2_bits_2(s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_src_afhob_2_bits_2),
    .s2_AFHOB_src_afhob_2_bits_3(s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_src_afhob_2_bits_3),
    .s2_AFHOB_src_afhob_1_bits_0(s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_src_afhob_1_bits_0),
    .s2_AFHOB_src_afhob_1_bits_1(s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_src_afhob_1_bits_1),
    .s2_AFHOB_src_afhob_1_bits_2(s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_src_afhob_1_bits_2),
    .s2_AFHOB_src_afhob_1_bits_3(s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_src_afhob_1_bits_3),
    .s2_AFHOB_src_afhob_0_bits_0(s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_src_afhob_0_bits_0),
    .s2_AFHOB_src_afhob_0_bits_1(s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_src_afhob_0_bits_1),
    .s2_AFHOB_src_afhob_0_bits_2(s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_src_afhob_0_bits_2),
    .s2_AFHOB_src_afhob_0_bits_3(s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_src_afhob_0_bits_3),
    .s1_AFHOB_sel(s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_sel),
    .s1_AFHOB_src_afhob_5_bits_0(s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_src_afhob_5_bits_0),
    .s1_AFHOB_src_afhob_5_bits_1(s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_src_afhob_5_bits_1),
    .s1_AFHOB_src_afhob_5_bits_2(s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_src_afhob_5_bits_2),
    .s1_AFHOB_src_afhob_5_bits_3(s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_src_afhob_5_bits_3),
    .s1_AFHOB_src_afhob_4_bits_0(s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_src_afhob_4_bits_0),
    .s1_AFHOB_src_afhob_4_bits_1(s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_src_afhob_4_bits_1),
    .s1_AFHOB_src_afhob_4_bits_2(s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_src_afhob_4_bits_2),
    .s1_AFHOB_src_afhob_4_bits_3(s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_src_afhob_4_bits_3),
    .s1_AFHOB_src_afhob_3_bits_0(s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_src_afhob_3_bits_0),
    .s1_AFHOB_src_afhob_3_bits_1(s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_src_afhob_3_bits_1),
    .s1_AFHOB_src_afhob_3_bits_2(s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_src_afhob_3_bits_2),
    .s1_AFHOB_src_afhob_3_bits_3(s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_src_afhob_3_bits_3),
    .s1_AFHOB_src_afhob_2_bits_0(s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_src_afhob_2_bits_0),
    .s1_AFHOB_src_afhob_2_bits_1(s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_src_afhob_2_bits_1),
    .s1_AFHOB_src_afhob_2_bits_2(s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_src_afhob_2_bits_2),
    .s1_AFHOB_src_afhob_2_bits_3(s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_src_afhob_2_bits_3),
    .s1_AFHOB_src_afhob_1_bits_0(s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_src_afhob_1_bits_0),
    .s1_AFHOB_src_afhob_1_bits_1(s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_src_afhob_1_bits_1),
    .s1_AFHOB_src_afhob_1_bits_2(s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_src_afhob_1_bits_2),
    .s1_AFHOB_src_afhob_1_bits_3(s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_src_afhob_1_bits_3),
    .s1_AFHOB_src_afhob_0_bits_0(s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_src_afhob_0_bits_0),
    .s1_AFHOB_src_afhob_0_bits_1(s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_src_afhob_0_bits_1),
    .s1_AFHOB_src_afhob_0_bits_2(s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_src_afhob_0_bits_2),
    .s1_AFHOB_src_afhob_0_bits_3(s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_src_afhob_0_bits_3),
    .s3_AFHOB_sel(s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_sel),
    .s3_AFHOB_src_afhob_5_bits_0(s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_src_afhob_5_bits_0),
    .s3_AFHOB_src_afhob_5_bits_1(s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_src_afhob_5_bits_1),
    .s3_AFHOB_src_afhob_5_bits_2(s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_src_afhob_5_bits_2),
    .s3_AFHOB_src_afhob_5_bits_3(s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_src_afhob_5_bits_3),
    .s3_AFHOB_src_afhob_4_bits_0(s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_src_afhob_4_bits_0),
    .s3_AFHOB_src_afhob_4_bits_1(s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_src_afhob_4_bits_1),
    .s3_AFHOB_src_afhob_4_bits_2(s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_src_afhob_4_bits_2),
    .s3_AFHOB_src_afhob_4_bits_3(s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_src_afhob_4_bits_3),
    .s3_AFHOB_src_afhob_3_bits_0(s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_src_afhob_3_bits_0),
    .s3_AFHOB_src_afhob_3_bits_1(s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_src_afhob_3_bits_1),
    .s3_AFHOB_src_afhob_3_bits_2(s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_src_afhob_3_bits_2),
    .s3_AFHOB_src_afhob_3_bits_3(s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_src_afhob_3_bits_3),
    .s3_AFHOB_src_afhob_2_bits_0(s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_src_afhob_2_bits_0),
    .s3_AFHOB_src_afhob_2_bits_1(s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_src_afhob_2_bits_1),
    .s3_AFHOB_src_afhob_2_bits_2(s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_src_afhob_2_bits_2),
    .s3_AFHOB_src_afhob_2_bits_3(s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_src_afhob_2_bits_3),
    .s3_AFHOB_src_afhob_1_bits_0(s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_src_afhob_1_bits_0),
    .s3_AFHOB_src_afhob_1_bits_1(s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_src_afhob_1_bits_1),
    .s3_AFHOB_src_afhob_1_bits_2(s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_src_afhob_1_bits_2),
    .s3_AFHOB_src_afhob_1_bits_3(s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_src_afhob_1_bits_3),
    .s3_AFHOB_src_afhob_0_bits_0(s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_src_afhob_0_bits_0),
    .s3_AFHOB_src_afhob_0_bits_1(s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_src_afhob_0_bits_1),
    .s3_AFHOB_src_afhob_0_bits_2(s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_src_afhob_0_bits_2),
    .s3_AFHOB_src_afhob_0_bits_3(s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_src_afhob_0_bits_3),
    .redirect_AFHOB_sel(s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_sel),
    .redirect_AFHOB_src_afhob_5_bits_0(s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_src_afhob_5_bits_0),
    .redirect_AFHOB_src_afhob_5_bits_1(s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_src_afhob_5_bits_1),
    .redirect_AFHOB_src_afhob_5_bits_2(s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_src_afhob_5_bits_2),
    .redirect_AFHOB_src_afhob_5_bits_3(s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_src_afhob_5_bits_3),
    .redirect_AFHOB_src_afhob_4_bits_0(s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_src_afhob_4_bits_0),
    .redirect_AFHOB_src_afhob_4_bits_1(s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_src_afhob_4_bits_1),
    .redirect_AFHOB_src_afhob_4_bits_2(s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_src_afhob_4_bits_2),
    .redirect_AFHOB_src_afhob_4_bits_3(s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_src_afhob_4_bits_3),
    .redirect_AFHOB_src_afhob_3_bits_0(s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_src_afhob_3_bits_0),
    .redirect_AFHOB_src_afhob_3_bits_1(s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_src_afhob_3_bits_1),
    .redirect_AFHOB_src_afhob_3_bits_2(s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_src_afhob_3_bits_2),
    .redirect_AFHOB_src_afhob_3_bits_3(s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_src_afhob_3_bits_3),
    .redirect_AFHOB_src_afhob_2_bits_0(s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_src_afhob_2_bits_0),
    .redirect_AFHOB_src_afhob_2_bits_1(s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_src_afhob_2_bits_1),
    .redirect_AFHOB_src_afhob_2_bits_2(s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_src_afhob_2_bits_2),
    .redirect_AFHOB_src_afhob_2_bits_3(s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_src_afhob_2_bits_3),
    .redirect_AFHOB_src_afhob_1_bits_0(s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_src_afhob_1_bits_0),
    .redirect_AFHOB_src_afhob_1_bits_1(s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_src_afhob_1_bits_1),
    .redirect_AFHOB_src_afhob_1_bits_2(s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_src_afhob_1_bits_2),
    .redirect_AFHOB_src_afhob_1_bits_3(s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_src_afhob_1_bits_3),
    .redirect_AFHOB_src_afhob_0_bits_0(s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_src_afhob_0_bits_0),
    .redirect_AFHOB_src_afhob_0_bits_1(s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_src_afhob_0_bits_1),
    .redirect_AFHOB_src_afhob_0_bits_2(s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_src_afhob_0_bits_2),
    .redirect_AFHOB_src_afhob_0_bits_3(s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_src_afhob_0_bits_3),
    .stallAFHOB_src_afhob_5_bits_0(s0_ahead_fh_oldest_bits_ppm_stallAFHOB_src_afhob_5_bits_0),
    .stallAFHOB_src_afhob_5_bits_1(s0_ahead_fh_oldest_bits_ppm_stallAFHOB_src_afhob_5_bits_1),
    .stallAFHOB_src_afhob_5_bits_2(s0_ahead_fh_oldest_bits_ppm_stallAFHOB_src_afhob_5_bits_2),
    .stallAFHOB_src_afhob_5_bits_3(s0_ahead_fh_oldest_bits_ppm_stallAFHOB_src_afhob_5_bits_3),
    .stallAFHOB_src_afhob_4_bits_0(s0_ahead_fh_oldest_bits_ppm_stallAFHOB_src_afhob_4_bits_0),
    .stallAFHOB_src_afhob_4_bits_1(s0_ahead_fh_oldest_bits_ppm_stallAFHOB_src_afhob_4_bits_1),
    .stallAFHOB_src_afhob_4_bits_2(s0_ahead_fh_oldest_bits_ppm_stallAFHOB_src_afhob_4_bits_2),
    .stallAFHOB_src_afhob_4_bits_3(s0_ahead_fh_oldest_bits_ppm_stallAFHOB_src_afhob_4_bits_3),
    .stallAFHOB_src_afhob_3_bits_0(s0_ahead_fh_oldest_bits_ppm_stallAFHOB_src_afhob_3_bits_0),
    .stallAFHOB_src_afhob_3_bits_1(s0_ahead_fh_oldest_bits_ppm_stallAFHOB_src_afhob_3_bits_1),
    .stallAFHOB_src_afhob_3_bits_2(s0_ahead_fh_oldest_bits_ppm_stallAFHOB_src_afhob_3_bits_2),
    .stallAFHOB_src_afhob_3_bits_3(s0_ahead_fh_oldest_bits_ppm_stallAFHOB_src_afhob_3_bits_3),
    .stallAFHOB_src_afhob_2_bits_0(s0_ahead_fh_oldest_bits_ppm_stallAFHOB_src_afhob_2_bits_0),
    .stallAFHOB_src_afhob_2_bits_1(s0_ahead_fh_oldest_bits_ppm_stallAFHOB_src_afhob_2_bits_1),
    .stallAFHOB_src_afhob_2_bits_2(s0_ahead_fh_oldest_bits_ppm_stallAFHOB_src_afhob_2_bits_2),
    .stallAFHOB_src_afhob_2_bits_3(s0_ahead_fh_oldest_bits_ppm_stallAFHOB_src_afhob_2_bits_3),
    .stallAFHOB_src_afhob_1_bits_0(s0_ahead_fh_oldest_bits_ppm_stallAFHOB_src_afhob_1_bits_0),
    .stallAFHOB_src_afhob_1_bits_1(s0_ahead_fh_oldest_bits_ppm_stallAFHOB_src_afhob_1_bits_1),
    .stallAFHOB_src_afhob_1_bits_2(s0_ahead_fh_oldest_bits_ppm_stallAFHOB_src_afhob_1_bits_2),
    .stallAFHOB_src_afhob_1_bits_3(s0_ahead_fh_oldest_bits_ppm_stallAFHOB_src_afhob_1_bits_3),
    .stallAFHOB_src_afhob_0_bits_0(s0_ahead_fh_oldest_bits_ppm_stallAFHOB_src_afhob_0_bits_0),
    .stallAFHOB_src_afhob_0_bits_1(s0_ahead_fh_oldest_bits_ppm_stallAFHOB_src_afhob_0_bits_1),
    .stallAFHOB_src_afhob_0_bits_2(s0_ahead_fh_oldest_bits_ppm_stallAFHOB_src_afhob_0_bits_2),
    .stallAFHOB_src_afhob_0_bits_3(s0_ahead_fh_oldest_bits_ppm_stallAFHOB_src_afhob_0_bits_3),
    .out_res_afhob_5_bits_0(s0_ahead_fh_oldest_bits_ppm_out_res_afhob_5_bits_0),
    .out_res_afhob_5_bits_1(s0_ahead_fh_oldest_bits_ppm_out_res_afhob_5_bits_1),
    .out_res_afhob_5_bits_2(s0_ahead_fh_oldest_bits_ppm_out_res_afhob_5_bits_2),
    .out_res_afhob_5_bits_3(s0_ahead_fh_oldest_bits_ppm_out_res_afhob_5_bits_3),
    .out_res_afhob_4_bits_0(s0_ahead_fh_oldest_bits_ppm_out_res_afhob_4_bits_0),
    .out_res_afhob_4_bits_1(s0_ahead_fh_oldest_bits_ppm_out_res_afhob_4_bits_1),
    .out_res_afhob_4_bits_2(s0_ahead_fh_oldest_bits_ppm_out_res_afhob_4_bits_2),
    .out_res_afhob_4_bits_3(s0_ahead_fh_oldest_bits_ppm_out_res_afhob_4_bits_3),
    .out_res_afhob_3_bits_0(s0_ahead_fh_oldest_bits_ppm_out_res_afhob_3_bits_0),
    .out_res_afhob_3_bits_1(s0_ahead_fh_oldest_bits_ppm_out_res_afhob_3_bits_1),
    .out_res_afhob_3_bits_2(s0_ahead_fh_oldest_bits_ppm_out_res_afhob_3_bits_2),
    .out_res_afhob_3_bits_3(s0_ahead_fh_oldest_bits_ppm_out_res_afhob_3_bits_3),
    .out_res_afhob_2_bits_0(s0_ahead_fh_oldest_bits_ppm_out_res_afhob_2_bits_0),
    .out_res_afhob_2_bits_1(s0_ahead_fh_oldest_bits_ppm_out_res_afhob_2_bits_1),
    .out_res_afhob_2_bits_2(s0_ahead_fh_oldest_bits_ppm_out_res_afhob_2_bits_2),
    .out_res_afhob_2_bits_3(s0_ahead_fh_oldest_bits_ppm_out_res_afhob_2_bits_3),
    .out_res_afhob_1_bits_0(s0_ahead_fh_oldest_bits_ppm_out_res_afhob_1_bits_0),
    .out_res_afhob_1_bits_1(s0_ahead_fh_oldest_bits_ppm_out_res_afhob_1_bits_1),
    .out_res_afhob_1_bits_2(s0_ahead_fh_oldest_bits_ppm_out_res_afhob_1_bits_2),
    .out_res_afhob_1_bits_3(s0_ahead_fh_oldest_bits_ppm_out_res_afhob_1_bits_3),
    .out_res_afhob_0_bits_0(s0_ahead_fh_oldest_bits_ppm_out_res_afhob_0_bits_0),
    .out_res_afhob_0_bits_1(s0_ahead_fh_oldest_bits_ppm_out_res_afhob_0_bits_1),
    .out_res_afhob_0_bits_2(s0_ahead_fh_oldest_bits_ppm_out_res_afhob_0_bits_2),
    .out_res_afhob_0_bits_3(s0_ahead_fh_oldest_bits_ppm_out_res_afhob_0_bits_3)
  );
  PriorityMuxModule_4 s0_last_br_num_oh_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_BrNumOH_sel(s0_last_br_num_oh_ppm_s2_BrNumOH_sel),
    .s2_BrNumOH_src(s0_last_br_num_oh_ppm_s2_BrNumOH_src),
    .s1_BrNumOH_sel(s0_last_br_num_oh_ppm_s1_BrNumOH_sel),
    .s1_BrNumOH_src(s0_last_br_num_oh_ppm_s1_BrNumOH_src),
    .s3_BrNumOH_sel(s0_last_br_num_oh_ppm_s3_BrNumOH_sel),
    .s3_BrNumOH_src(s0_last_br_num_oh_ppm_s3_BrNumOH_src),
    .redirect_BrNumOH_sel(s0_last_br_num_oh_ppm_redirect_BrNumOH_sel),
    .redirect_BrNumOH_src(s0_last_br_num_oh_ppm_redirect_BrNumOH_src),
    .stallBrNumOH_src(s0_last_br_num_oh_ppm_stallBrNumOH_src),
    .out_res(s0_last_br_num_oh_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_0_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_0_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_0_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_0_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_0_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_0_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_0_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_0_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_0_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_1_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_1_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_1_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_1_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_1_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_1_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_1_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_1_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_1_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_2_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_2_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_2_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_2_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_2_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_2_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_2_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_2_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_2_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_3_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_3_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_3_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_3_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_3_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_3_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_3_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_3_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_3_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_4_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_4_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_4_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_4_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_4_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_4_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_4_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_4_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_4_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_5_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_5_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_5_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_5_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_5_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_5_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_5_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_5_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_5_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_6_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_6_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_6_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_6_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_6_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_6_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_6_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_6_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_6_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_7_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_7_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_7_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_7_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_7_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_7_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_7_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_7_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_7_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_8_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_8_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_8_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_8_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_8_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_8_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_8_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_8_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_8_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_9_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_9_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_9_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_9_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_9_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_9_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_9_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_9_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_9_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_10_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_10_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_10_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_10_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_10_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_10_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_10_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_10_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_10_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_11_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_11_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_11_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_11_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_11_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_11_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_11_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_11_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_11_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_12_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_12_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_12_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_12_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_12_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_12_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_12_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_12_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_12_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_13_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_13_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_13_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_13_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_13_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_13_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_13_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_13_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_13_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_14_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_14_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_14_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_14_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_14_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_14_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_14_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_14_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_14_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_15_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_15_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_15_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_15_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_15_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_15_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_15_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_15_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_15_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_16_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_16_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_16_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_16_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_16_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_16_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_16_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_16_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_16_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_17_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_17_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_17_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_17_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_17_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_17_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_17_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_17_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_17_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_18_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_18_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_18_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_18_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_18_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_18_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_18_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_18_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_18_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_19_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_19_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_19_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_19_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_19_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_19_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_19_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_19_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_19_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_20_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_20_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_20_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_20_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_20_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_20_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_20_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_20_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_20_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_21_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_21_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_21_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_21_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_21_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_21_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_21_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_21_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_21_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_22_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_22_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_22_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_22_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_22_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_22_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_22_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_22_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_22_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_23_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_23_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_23_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_23_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_23_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_23_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_23_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_23_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_23_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_24_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_24_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_24_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_24_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_24_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_24_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_24_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_24_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_24_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_25_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_25_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_25_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_25_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_25_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_25_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_25_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_25_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_25_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_26_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_26_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_26_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_26_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_26_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_26_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_26_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_26_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_26_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_27_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_27_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_27_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_27_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_27_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_27_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_27_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_27_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_27_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_28_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_28_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_28_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_28_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_28_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_28_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_28_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_28_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_28_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_29_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_29_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_29_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_29_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_29_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_29_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_29_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_29_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_29_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_30_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_30_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_30_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_30_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_30_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_30_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_30_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_30_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_30_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_31_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_31_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_31_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_31_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_31_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_31_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_31_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_31_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_31_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_32_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_32_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_32_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_32_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_32_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_32_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_32_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_32_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_32_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_33_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_33_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_33_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_33_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_33_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_33_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_33_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_33_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_33_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_34_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_34_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_34_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_34_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_34_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_34_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_34_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_34_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_34_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_35_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_35_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_35_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_35_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_35_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_35_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_35_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_35_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_35_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_36_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_36_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_36_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_36_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_36_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_36_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_36_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_36_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_36_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_37_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_37_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_37_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_37_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_37_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_37_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_37_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_37_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_37_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_38_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_38_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_38_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_38_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_38_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_38_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_38_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_38_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_38_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_39_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_39_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_39_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_39_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_39_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_39_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_39_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_39_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_39_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_40_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_40_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_40_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_40_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_40_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_40_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_40_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_40_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_40_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_41_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_41_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_41_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_41_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_41_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_41_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_41_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_41_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_41_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_42_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_42_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_42_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_42_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_42_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_42_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_42_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_42_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_42_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_43_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_43_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_43_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_43_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_43_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_43_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_43_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_43_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_43_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_44_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_44_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_44_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_44_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_44_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_44_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_44_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_44_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_44_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_45_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_45_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_45_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_45_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_45_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_45_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_45_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_45_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_45_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_46_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_46_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_46_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_46_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_46_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_46_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_46_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_46_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_46_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_47_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_47_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_47_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_47_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_47_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_47_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_47_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_47_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_47_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_48_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_48_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_48_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_48_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_48_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_48_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_48_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_48_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_48_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_49_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_49_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_49_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_49_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_49_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_49_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_49_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_49_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_49_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_50_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_50_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_50_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_50_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_50_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_50_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_50_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_50_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_50_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_51_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_51_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_51_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_51_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_51_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_51_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_51_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_51_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_51_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_52_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_52_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_52_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_52_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_52_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_52_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_52_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_52_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_52_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_53_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_53_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_53_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_53_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_53_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_53_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_53_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_53_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_53_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_54_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_54_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_54_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_54_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_54_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_54_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_54_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_54_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_54_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_55_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_55_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_55_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_55_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_55_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_55_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_55_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_55_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_55_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_56_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_56_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_56_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_56_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_56_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_56_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_56_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_56_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_56_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_57_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_57_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_57_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_57_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_57_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_57_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_57_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_57_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_57_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_58_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_58_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_58_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_58_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_58_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_58_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_58_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_58_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_58_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_59_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_59_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_59_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_59_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_59_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_59_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_59_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_59_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_59_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_60_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_60_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_60_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_60_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_60_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_60_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_60_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_60_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_60_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_61_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_61_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_61_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_61_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_61_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_61_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_61_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_61_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_61_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_62_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_62_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_62_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_62_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_62_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_62_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_62_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_62_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_62_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_63_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_63_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_63_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_63_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_63_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_63_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_63_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_63_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_63_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_64_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_64_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_64_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_64_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_64_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_64_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_64_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_64_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_64_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_65_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_65_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_65_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_65_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_65_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_65_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_65_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_65_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_65_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_66_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_66_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_66_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_66_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_66_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_66_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_66_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_66_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_66_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_67_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_67_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_67_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_67_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_67_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_67_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_67_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_67_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_67_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_68_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_68_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_68_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_68_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_68_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_68_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_68_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_68_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_68_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_69_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_69_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_69_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_69_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_69_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_69_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_69_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_69_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_69_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_70_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_70_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_70_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_70_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_70_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_70_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_70_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_70_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_70_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_71_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_71_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_71_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_71_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_71_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_71_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_71_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_71_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_71_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_72_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_72_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_72_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_72_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_72_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_72_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_72_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_72_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_72_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_73_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_73_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_73_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_73_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_73_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_73_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_73_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_73_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_73_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_74_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_74_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_74_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_74_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_74_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_74_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_74_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_74_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_74_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_75_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_75_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_75_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_75_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_75_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_75_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_75_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_75_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_75_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_76_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_76_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_76_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_76_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_76_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_76_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_76_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_76_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_76_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_77_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_77_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_77_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_77_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_77_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_77_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_77_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_77_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_77_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_78_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_78_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_78_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_78_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_78_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_78_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_78_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_78_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_78_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_79_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_79_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_79_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_79_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_79_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_79_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_79_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_79_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_79_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_80_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_80_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_80_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_80_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_80_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_80_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_80_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_80_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_80_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_81_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_81_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_81_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_81_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_81_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_81_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_81_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_81_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_81_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_82_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_82_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_82_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_82_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_82_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_82_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_82_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_82_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_82_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_83_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_83_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_83_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_83_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_83_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_83_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_83_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_83_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_83_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_84_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_84_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_84_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_84_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_84_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_84_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_84_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_84_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_84_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_85_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_85_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_85_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_85_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_85_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_85_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_85_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_85_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_85_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_86_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_86_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_86_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_86_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_86_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_86_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_86_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_86_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_86_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_87_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_87_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_87_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_87_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_87_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_87_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_87_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_87_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_87_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_88_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_88_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_88_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_88_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_88_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_88_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_88_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_88_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_88_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_89_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_89_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_89_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_89_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_89_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_89_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_89_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_89_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_89_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_90_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_90_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_90_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_90_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_90_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_90_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_90_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_90_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_90_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_91_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_91_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_91_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_91_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_91_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_91_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_91_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_91_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_91_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_92_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_92_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_92_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_92_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_92_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_92_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_92_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_92_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_92_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_93_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_93_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_93_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_93_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_93_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_93_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_93_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_93_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_93_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_94_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_94_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_94_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_94_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_94_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_94_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_94_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_94_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_94_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_95_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_95_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_95_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_95_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_95_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_95_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_95_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_95_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_95_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_96_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_96_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_96_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_96_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_96_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_96_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_96_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_96_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_96_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_97_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_97_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_97_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_97_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_97_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_97_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_97_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_97_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_97_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_98_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_98_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_98_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_98_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_98_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_98_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_98_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_98_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_98_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_99_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_99_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_99_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_99_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_99_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_99_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_99_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_99_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_99_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_100_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_100_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_100_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_100_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_100_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_100_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_100_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_100_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_100_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_101_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_101_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_101_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_101_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_101_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_101_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_101_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_101_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_101_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_102_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_102_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_102_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_102_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_102_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_102_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_102_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_102_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_102_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_103_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_103_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_103_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_103_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_103_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_103_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_103_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_103_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_103_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_104_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_104_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_104_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_104_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_104_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_104_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_104_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_104_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_104_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_105_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_105_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_105_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_105_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_105_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_105_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_105_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_105_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_105_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_106_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_106_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_106_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_106_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_106_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_106_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_106_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_106_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_106_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_107_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_107_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_107_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_107_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_107_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_107_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_107_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_107_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_107_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_108_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_108_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_108_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_108_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_108_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_108_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_108_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_108_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_108_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_109_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_109_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_109_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_109_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_109_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_109_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_109_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_109_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_109_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_110_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_110_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_110_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_110_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_110_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_110_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_110_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_110_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_110_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_111_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_111_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_111_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_111_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_111_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_111_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_111_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_111_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_111_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_112_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_112_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_112_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_112_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_112_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_112_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_112_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_112_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_112_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_113_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_113_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_113_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_113_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_113_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_113_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_113_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_113_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_113_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_114_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_114_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_114_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_114_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_114_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_114_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_114_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_114_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_114_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_115_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_115_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_115_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_115_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_115_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_115_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_115_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_115_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_115_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_116_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_116_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_116_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_116_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_116_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_116_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_116_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_116_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_116_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_117_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_117_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_117_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_117_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_117_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_117_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_117_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_117_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_117_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_118_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_118_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_118_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_118_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_118_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_118_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_118_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_118_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_118_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_119_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_119_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_119_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_119_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_119_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_119_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_119_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_119_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_119_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_120_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_120_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_120_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_120_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_120_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_120_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_120_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_120_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_120_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_121_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_121_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_121_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_121_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_121_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_121_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_121_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_121_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_121_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_122_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_122_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_122_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_122_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_122_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_122_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_122_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_122_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_122_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_123_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_123_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_123_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_123_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_123_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_123_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_123_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_123_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_123_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_124_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_124_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_124_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_124_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_124_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_124_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_124_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_124_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_124_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_125_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_125_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_125_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_125_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_125_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_125_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_125_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_125_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_125_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_126_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_126_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_126_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_126_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_126_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_126_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_126_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_126_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_126_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_127_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_127_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_127_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_127_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_127_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_127_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_127_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_127_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_127_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_128_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_128_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_128_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_128_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_128_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_128_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_128_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_128_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_128_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_129_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_129_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_129_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_129_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_129_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_129_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_129_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_129_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_129_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_130_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_130_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_130_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_130_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_130_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_130_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_130_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_130_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_130_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_131_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_131_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_131_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_131_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_131_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_131_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_131_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_131_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_131_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_132_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_132_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_132_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_132_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_132_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_132_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_132_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_132_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_132_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_133_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_133_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_133_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_133_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_133_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_133_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_133_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_133_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_133_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_134_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_134_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_134_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_134_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_134_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_134_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_134_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_134_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_134_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_135_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_135_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_135_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_135_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_135_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_135_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_135_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_135_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_135_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_136_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_136_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_136_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_136_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_136_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_136_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_136_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_136_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_136_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_137_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_137_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_137_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_137_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_137_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_137_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_137_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_137_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_137_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_138_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_138_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_138_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_138_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_138_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_138_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_138_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_138_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_138_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_139_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_139_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_139_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_139_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_139_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_139_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_139_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_139_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_139_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_140_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_140_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_140_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_140_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_140_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_140_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_140_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_140_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_140_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_141_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_141_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_141_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_141_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_141_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_141_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_141_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_141_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_141_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_142_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_142_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_142_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_142_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_142_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_142_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_142_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_142_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_142_ppm_out_res)
  );
  PriorityMuxModule_5 ghv_write_datas_143_ppm ( // @[PriorityMuxGen.scala 136:25]
    .s2_new_bit_0_sel(ghv_write_datas_143_ppm_s2_new_bit_0_sel),
    .s2_new_bit_0_src(ghv_write_datas_143_ppm_s2_new_bit_0_src),
    .s1_new_bit_0_sel(ghv_write_datas_143_ppm_s1_new_bit_0_sel),
    .s1_new_bit_0_src(ghv_write_datas_143_ppm_s1_new_bit_0_src),
    .s3_new_bit_0_sel(ghv_write_datas_143_ppm_s3_new_bit_0_sel),
    .s3_new_bit_0_src(ghv_write_datas_143_ppm_s3_new_bit_0_src),
    .redirect_new_bit_0_src(ghv_write_datas_143_ppm_redirect_new_bit_0_src),
    .out_res(ghv_write_datas_143_ppm_out_res)
  );
  assign io_bpu_to_ftq_resp_valid = _io_bpu_to_ftq_resp_valid_T_3 | _io_bpu_to_ftq_resp_valid_T_4; // @[BPU.scala 383:28]
  assign io_bpu_to_ftq_resp_bits_s1_pc = predictors_io_out_s1_pc; // @[BPU.scala 385:28]
  assign io_bpu_to_ftq_resp_bits_s1_full_pred_br_taken_mask_0 = predictors_io_out_s1_full_pred_br_taken_mask_0; // @[BPU.scala 385:28]
  assign io_bpu_to_ftq_resp_bits_s1_full_pred_br_taken_mask_1 = predictors_io_out_s1_full_pred_br_taken_mask_1; // @[BPU.scala 385:28]
  assign io_bpu_to_ftq_resp_bits_s1_full_pred_slot_valids_0 = predictors_io_out_s1_full_pred_slot_valids_0; // @[BPU.scala 385:28]
  assign io_bpu_to_ftq_resp_bits_s1_full_pred_slot_valids_1 = predictors_io_out_s1_full_pred_slot_valids_1; // @[BPU.scala 385:28]
  assign io_bpu_to_ftq_resp_bits_s1_full_pred_targets_0 = predictors_io_out_s1_full_pred_targets_0; // @[BPU.scala 385:28]
  assign io_bpu_to_ftq_resp_bits_s1_full_pred_targets_1 = predictors_io_out_s1_full_pred_targets_1; // @[BPU.scala 385:28]
  assign io_bpu_to_ftq_resp_bits_s1_full_pred_offsets_0 = predictors_io_out_s1_full_pred_offsets_0; // @[BPU.scala 385:28]
  assign io_bpu_to_ftq_resp_bits_s1_full_pred_offsets_1 = predictors_io_out_s1_full_pred_offsets_1; // @[BPU.scala 385:28]
  assign io_bpu_to_ftq_resp_bits_s1_full_pred_fallThroughAddr = predictors_io_out_s1_full_pred_fallThroughAddr; // @[BPU.scala 385:28]
  assign io_bpu_to_ftq_resp_bits_s1_full_pred_fallThroughErr = predictors_io_out_s1_full_pred_fallThroughErr; // @[BPU.scala 385:28]
  assign io_bpu_to_ftq_resp_bits_s1_full_pred_is_br_sharing = predictors_io_out_s1_full_pred_is_br_sharing; // @[BPU.scala 385:28]
  assign io_bpu_to_ftq_resp_bits_s1_full_pred_hit = predictors_io_out_s1_full_pred_hit; // @[BPU.scala 385:28]
  assign io_bpu_to_ftq_resp_bits_s2_pc = predictors_io_out_s2_pc; // @[BPU.scala 385:28]
  assign io_bpu_to_ftq_resp_bits_s2_valid = s2_valid & _s3_valid_T; // @[BPU.scala 592:47]
  assign io_bpu_to_ftq_resp_bits_s2_hasRedirect = s2_valid & (s2_redirect_s1_last_pred_vec_0 |
    s2_redirect_s1_last_pred_vec_1 | s2_redirect_s1_last_pred_vec_2 | s2_redirect_s1_last_pred_vec_3); // @[BPU.scala 503:26]
  assign io_bpu_to_ftq_resp_bits_s2_ftq_idx_flag = s2_ftq_idx_flag; // @[BPU.scala 594:38]
  assign io_bpu_to_ftq_resp_bits_s2_ftq_idx_value = s2_ftq_idx_value; // @[BPU.scala 594:38]
  assign io_bpu_to_ftq_resp_bits_s2_full_pred_br_taken_mask_0 = predictors_io_out_s2_full_pred_br_taken_mask_0; // @[BPU.scala 385:28]
  assign io_bpu_to_ftq_resp_bits_s2_full_pred_br_taken_mask_1 = predictors_io_out_s2_full_pred_br_taken_mask_1; // @[BPU.scala 385:28]
  assign io_bpu_to_ftq_resp_bits_s2_full_pred_slot_valids_0 = predictors_io_out_s2_full_pred_slot_valids_0; // @[BPU.scala 385:28]
  assign io_bpu_to_ftq_resp_bits_s2_full_pred_slot_valids_1 = predictors_io_out_s2_full_pred_slot_valids_1; // @[BPU.scala 385:28]
  assign io_bpu_to_ftq_resp_bits_s2_full_pred_targets_0 = predictors_io_out_s2_full_pred_targets_0; // @[BPU.scala 385:28]
  assign io_bpu_to_ftq_resp_bits_s2_full_pred_targets_1 = predictors_io_out_s2_full_pred_targets_1; // @[BPU.scala 385:28]
  assign io_bpu_to_ftq_resp_bits_s2_full_pred_offsets_0 = predictors_io_out_s2_full_pred_offsets_0; // @[BPU.scala 385:28]
  assign io_bpu_to_ftq_resp_bits_s2_full_pred_offsets_1 = predictors_io_out_s2_full_pred_offsets_1; // @[BPU.scala 385:28]
  assign io_bpu_to_ftq_resp_bits_s2_full_pred_fallThroughAddr = predictors_io_out_s2_full_pred_fallThroughAddr; // @[BPU.scala 385:28]
  assign io_bpu_to_ftq_resp_bits_s2_full_pred_fallThroughErr = predictors_io_out_s2_full_pred_fallThroughErr; // @[BPU.scala 385:28]
  assign io_bpu_to_ftq_resp_bits_s2_full_pred_is_br_sharing = predictors_io_out_s2_full_pred_is_br_sharing; // @[BPU.scala 385:28]
  assign io_bpu_to_ftq_resp_bits_s2_full_pred_hit = predictors_io_out_s2_full_pred_hit; // @[BPU.scala 385:28]
  assign io_bpu_to_ftq_resp_bits_s3_pc = predictors_io_out_s3_pc; // @[BPU.scala 385:28]
  assign io_bpu_to_ftq_resp_bits_s3_valid = s3_valid & ~io_ftq_to_bpu_redirect_valid; // @[BPU.scala 595:47]
  assign io_bpu_to_ftq_resp_bits_s3_hasRedirect = s3_valid & _s3_redirect_T_1; // @[BPU.scala 568:26]
  assign io_bpu_to_ftq_resp_bits_s3_ftq_idx_flag = s3_ftq_idx_flag; // @[BPU.scala 597:38]
  assign io_bpu_to_ftq_resp_bits_s3_ftq_idx_value = s3_ftq_idx_value; // @[BPU.scala 597:38]
  assign io_bpu_to_ftq_resp_bits_s3_full_pred_br_taken_mask_0 = predictors_io_out_s3_full_pred_br_taken_mask_0; // @[BPU.scala 385:28]
  assign io_bpu_to_ftq_resp_bits_s3_full_pred_br_taken_mask_1 = predictors_io_out_s3_full_pred_br_taken_mask_1; // @[BPU.scala 385:28]
  assign io_bpu_to_ftq_resp_bits_s3_full_pred_slot_valids_0 = predictors_io_out_s3_full_pred_slot_valids_0; // @[BPU.scala 385:28]
  assign io_bpu_to_ftq_resp_bits_s3_full_pred_slot_valids_1 = predictors_io_out_s3_full_pred_slot_valids_1; // @[BPU.scala 385:28]
  assign io_bpu_to_ftq_resp_bits_s3_full_pred_targets_0 = predictors_io_out_s3_full_pred_targets_0; // @[BPU.scala 385:28]
  assign io_bpu_to_ftq_resp_bits_s3_full_pred_targets_1 = predictors_io_out_s3_full_pred_targets_1; // @[BPU.scala 385:28]
  assign io_bpu_to_ftq_resp_bits_s3_full_pred_offsets_0 = predictors_io_out_s3_full_pred_offsets_0; // @[BPU.scala 385:28]
  assign io_bpu_to_ftq_resp_bits_s3_full_pred_offsets_1 = predictors_io_out_s3_full_pred_offsets_1; // @[BPU.scala 385:28]
  assign io_bpu_to_ftq_resp_bits_s3_full_pred_fallThroughAddr = predictors_io_out_s3_full_pred_fallThroughAddr; // @[BPU.scala 385:28]
  assign io_bpu_to_ftq_resp_bits_s3_full_pred_fallThroughErr = predictors_io_out_s3_full_pred_fallThroughErr; // @[BPU.scala 385:28]
  assign io_bpu_to_ftq_resp_bits_s3_full_pred_is_br_sharing = predictors_io_out_s3_full_pred_is_br_sharing; // @[BPU.scala 385:28]
  assign io_bpu_to_ftq_resp_bits_s3_full_pred_hit = predictors_io_out_s3_full_pred_hit; // @[BPU.scala 385:28]
  assign io_bpu_to_ftq_resp_bits_last_stage_meta = predictors_io_out_last_stage_meta; // @[BPU.scala 385:28]
  assign io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_17_folded_hist = s3_folded_gh_hist_17_folded_hist
    ; // @[BPU.scala 386:60]
  assign io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_16_folded_hist = s3_folded_gh_hist_16_folded_hist
    ; // @[BPU.scala 386:60]
  assign io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_15_folded_hist = s3_folded_gh_hist_15_folded_hist
    ; // @[BPU.scala 386:60]
  assign io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_14_folded_hist = s3_folded_gh_hist_14_folded_hist
    ; // @[BPU.scala 386:60]
  assign io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_13_folded_hist = s3_folded_gh_hist_13_folded_hist
    ; // @[BPU.scala 386:60]
  assign io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_12_folded_hist = s3_folded_gh_hist_12_folded_hist
    ; // @[BPU.scala 386:60]
  assign io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_11_folded_hist = s3_folded_gh_hist_11_folded_hist
    ; // @[BPU.scala 386:60]
  assign io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_10_folded_hist = s3_folded_gh_hist_10_folded_hist
    ; // @[BPU.scala 386:60]
  assign io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_9_folded_hist = s3_folded_gh_hist_9_folded_hist; // @[BPU.scala 386:60]
  assign io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_8_folded_hist = s3_folded_gh_hist_8_folded_hist; // @[BPU.scala 386:60]
  assign io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_7_folded_hist = s3_folded_gh_hist_7_folded_hist; // @[BPU.scala 386:60]
  assign io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_6_folded_hist = s3_folded_gh_hist_6_folded_hist; // @[BPU.scala 386:60]
  assign io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_5_folded_hist = s3_folded_gh_hist_5_folded_hist; // @[BPU.scala 386:60]
  assign io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_4_folded_hist = s3_folded_gh_hist_4_folded_hist; // @[BPU.scala 386:60]
  assign io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_3_folded_hist = s3_folded_gh_hist_3_folded_hist; // @[BPU.scala 386:60]
  assign io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_2_folded_hist = s3_folded_gh_hist_2_folded_hist; // @[BPU.scala 386:60]
  assign io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_1_folded_hist = s3_folded_gh_hist_1_folded_hist; // @[BPU.scala 386:60]
  assign io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_0_folded_hist = s3_folded_gh_hist_0_folded_hist; // @[BPU.scala 386:60]
  assign io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_5_bits_0 = s3_ahead_fh_oldest_bits_afhob_5_bits_0; // @[BPU.scala 389:60]
  assign io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_5_bits_1 = s3_ahead_fh_oldest_bits_afhob_5_bits_1; // @[BPU.scala 389:60]
  assign io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_5_bits_2 = s3_ahead_fh_oldest_bits_afhob_5_bits_2; // @[BPU.scala 389:60]
  assign io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_5_bits_3 = s3_ahead_fh_oldest_bits_afhob_5_bits_3; // @[BPU.scala 389:60]
  assign io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_4_bits_0 = s3_ahead_fh_oldest_bits_afhob_4_bits_0; // @[BPU.scala 389:60]
  assign io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_4_bits_1 = s3_ahead_fh_oldest_bits_afhob_4_bits_1; // @[BPU.scala 389:60]
  assign io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_4_bits_2 = s3_ahead_fh_oldest_bits_afhob_4_bits_2; // @[BPU.scala 389:60]
  assign io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_4_bits_3 = s3_ahead_fh_oldest_bits_afhob_4_bits_3; // @[BPU.scala 389:60]
  assign io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_3_bits_0 = s3_ahead_fh_oldest_bits_afhob_3_bits_0; // @[BPU.scala 389:60]
  assign io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_3_bits_1 = s3_ahead_fh_oldest_bits_afhob_3_bits_1; // @[BPU.scala 389:60]
  assign io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_3_bits_2 = s3_ahead_fh_oldest_bits_afhob_3_bits_2; // @[BPU.scala 389:60]
  assign io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_3_bits_3 = s3_ahead_fh_oldest_bits_afhob_3_bits_3; // @[BPU.scala 389:60]
  assign io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_2_bits_0 = s3_ahead_fh_oldest_bits_afhob_2_bits_0; // @[BPU.scala 389:60]
  assign io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_2_bits_1 = s3_ahead_fh_oldest_bits_afhob_2_bits_1; // @[BPU.scala 389:60]
  assign io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_2_bits_2 = s3_ahead_fh_oldest_bits_afhob_2_bits_2; // @[BPU.scala 389:60]
  assign io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_2_bits_3 = s3_ahead_fh_oldest_bits_afhob_2_bits_3; // @[BPU.scala 389:60]
  assign io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_1_bits_0 = s3_ahead_fh_oldest_bits_afhob_1_bits_0; // @[BPU.scala 389:60]
  assign io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_1_bits_1 = s3_ahead_fh_oldest_bits_afhob_1_bits_1; // @[BPU.scala 389:60]
  assign io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_1_bits_2 = s3_ahead_fh_oldest_bits_afhob_1_bits_2; // @[BPU.scala 389:60]
  assign io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_1_bits_3 = s3_ahead_fh_oldest_bits_afhob_1_bits_3; // @[BPU.scala 389:60]
  assign io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_0_bits_0 = s3_ahead_fh_oldest_bits_afhob_0_bits_0; // @[BPU.scala 389:60]
  assign io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_0_bits_1 = s3_ahead_fh_oldest_bits_afhob_0_bits_1; // @[BPU.scala 389:60]
  assign io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_0_bits_2 = s3_ahead_fh_oldest_bits_afhob_0_bits_2; // @[BPU.scala 389:60]
  assign io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_0_bits_3 = s3_ahead_fh_oldest_bits_afhob_0_bits_3; // @[BPU.scala 389:60]
  assign io_bpu_to_ftq_resp_bits_last_stage_spec_info_lastBrNumOH = s3_last_br_num_oh; // @[BPU.scala 388:60]
  assign io_bpu_to_ftq_resp_bits_last_stage_spec_info_histPtr_flag = s3_ghist_ptr_flag; // @[BPU.scala 387:60]
  assign io_bpu_to_ftq_resp_bits_last_stage_spec_info_histPtr_value = s3_ghist_ptr_value; // @[BPU.scala 387:60]
  assign io_bpu_to_ftq_resp_bits_last_stage_spec_info_rasSp = predictors_io_out_last_stage_spec_info_rasSp; // @[BPU.scala 385:28]
  assign io_bpu_to_ftq_resp_bits_last_stage_spec_info_rasTop_retAddr =
    predictors_io_out_last_stage_spec_info_rasTop_retAddr; // @[BPU.scala 385:28]
  assign io_bpu_to_ftq_resp_bits_last_stage_spec_info_rasTop_ctr = predictors_io_out_last_stage_spec_info_rasTop_ctr; // @[BPU.scala 385:28]
  assign io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_valid = predictors_io_out_last_stage_ftb_entry_valid; // @[BPU.scala 385:28]
  assign io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_brSlots_0_offset =
    predictors_io_out_last_stage_ftb_entry_brSlots_0_offset; // @[BPU.scala 385:28]
  assign io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_brSlots_0_lower =
    predictors_io_out_last_stage_ftb_entry_brSlots_0_lower; // @[BPU.scala 385:28]
  assign io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_brSlots_0_tarStat =
    predictors_io_out_last_stage_ftb_entry_brSlots_0_tarStat; // @[BPU.scala 385:28]
  assign io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_brSlots_0_sharing =
    predictors_io_out_last_stage_ftb_entry_brSlots_0_sharing; // @[BPU.scala 385:28]
  assign io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_brSlots_0_valid =
    predictors_io_out_last_stage_ftb_entry_brSlots_0_valid; // @[BPU.scala 385:28]
  assign io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_tailSlot_offset =
    predictors_io_out_last_stage_ftb_entry_tailSlot_offset; // @[BPU.scala 385:28]
  assign io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_tailSlot_lower =
    predictors_io_out_last_stage_ftb_entry_tailSlot_lower; // @[BPU.scala 385:28]
  assign io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_tailSlot_tarStat =
    predictors_io_out_last_stage_ftb_entry_tailSlot_tarStat; // @[BPU.scala 385:28]
  assign io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_tailSlot_sharing =
    predictors_io_out_last_stage_ftb_entry_tailSlot_sharing; // @[BPU.scala 385:28]
  assign io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_tailSlot_valid =
    predictors_io_out_last_stage_ftb_entry_tailSlot_valid; // @[BPU.scala 385:28]
  assign io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_pftAddr = predictors_io_out_last_stage_ftb_entry_pftAddr; // @[BPU.scala 385:28]
  assign io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_carry = predictors_io_out_last_stage_ftb_entry_carry; // @[BPU.scala 385:28]
  assign io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_isCall = predictors_io_out_last_stage_ftb_entry_isCall; // @[BPU.scala 385:28]
  assign io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_isRet = predictors_io_out_last_stage_ftb_entry_isRet; // @[BPU.scala 385:28]
  assign io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_isJalr = predictors_io_out_last_stage_ftb_entry_isJalr; // @[BPU.scala 385:28]
  assign io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_last_may_be_rvi_call =
    predictors_io_out_last_stage_ftb_entry_last_may_be_rvi_call; // @[BPU.scala 385:28]
  assign io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_always_taken_0 =
    predictors_io_out_last_stage_ftb_entry_always_taken_0; // @[BPU.scala 385:28]
  assign io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_always_taken_1 =
    predictors_io_out_last_stage_ftb_entry_always_taken_1; // @[BPU.scala 385:28]
  assign io_perf_0_value = io_perf_0_value_REG_1; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_1_value = io_perf_1_value_REG_1; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_2_value = io_perf_2_value_REG_1; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_3_value = io_perf_3_value_REG_1; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_4_value = io_perf_4_value_REG_1; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_5_value = io_perf_5_value_REG_1; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_6_value = io_perf_6_value_REG_1; // @[PerfCounterUtils.scala 188:17]
  assign ctrl_delay_clock = clock;
  assign ctrl_delay_io_in_ubtb_enable = io_ctrl_ubtb_enable; // @[Hold.scala 98:17]
  assign ctrl_delay_io_in_btb_enable = io_ctrl_btb_enable; // @[Hold.scala 98:17]
  assign ctrl_delay_io_in_tage_enable = io_ctrl_tage_enable; // @[Hold.scala 98:17]
  assign ctrl_delay_io_in_sc_enable = io_ctrl_sc_enable; // @[Hold.scala 98:17]
  assign ctrl_delay_io_in_ras_enable = io_ctrl_ras_enable; // @[Hold.scala 98:17]
  assign predictors_clock = clock;
  assign predictors_reset = reset;
  assign predictors_io_reset_vector = io_reset_vector; // @[BPU.scala 249:30]
  assign predictors_io_in_bits_s0_pc = s0_pc_ppm_out_res; // @[BPU.scala 257:19 667:17]
  assign predictors_io_in_bits_folded_hist_hist_17_folded_hist = s0_folded_gh_ppm_out_res_hist_17_folded_hist; // @[BPU.scala 266:26 668:17]
  assign predictors_io_in_bits_folded_hist_hist_16_folded_hist = s0_folded_gh_ppm_out_res_hist_16_folded_hist; // @[BPU.scala 266:26 668:17]
  assign predictors_io_in_bits_folded_hist_hist_15_folded_hist = s0_folded_gh_ppm_out_res_hist_15_folded_hist; // @[BPU.scala 266:26 668:17]
  assign predictors_io_in_bits_folded_hist_hist_14_folded_hist = s0_folded_gh_ppm_out_res_hist_14_folded_hist; // @[BPU.scala 266:26 668:17]
  assign predictors_io_in_bits_folded_hist_hist_13_folded_hist = s0_folded_gh_ppm_out_res_hist_13_folded_hist; // @[BPU.scala 266:26 668:17]
  assign predictors_io_in_bits_folded_hist_hist_12_folded_hist = s0_folded_gh_ppm_out_res_hist_12_folded_hist; // @[BPU.scala 266:26 668:17]
  assign predictors_io_in_bits_folded_hist_hist_10_folded_hist = s0_folded_gh_ppm_out_res_hist_10_folded_hist; // @[BPU.scala 266:26 668:17]
  assign predictors_io_in_bits_folded_hist_hist_9_folded_hist = s0_folded_gh_ppm_out_res_hist_9_folded_hist; // @[BPU.scala 266:26 668:17]
  assign predictors_io_in_bits_folded_hist_hist_8_folded_hist = s0_folded_gh_ppm_out_res_hist_8_folded_hist; // @[BPU.scala 266:26 668:17]
  assign predictors_io_in_bits_folded_hist_hist_7_folded_hist = s0_folded_gh_ppm_out_res_hist_7_folded_hist; // @[BPU.scala 266:26 668:17]
  assign predictors_io_in_bits_folded_hist_hist_6_folded_hist = s0_folded_gh_ppm_out_res_hist_6_folded_hist; // @[BPU.scala 266:26 668:17]
  assign predictors_io_in_bits_folded_hist_hist_5_folded_hist = s0_folded_gh_ppm_out_res_hist_5_folded_hist; // @[BPU.scala 266:26 668:17]
  assign predictors_io_in_bits_folded_hist_hist_4_folded_hist = s0_folded_gh_ppm_out_res_hist_4_folded_hist; // @[BPU.scala 266:26 668:17]
  assign predictors_io_in_bits_folded_hist_hist_3_folded_hist = s0_folded_gh_ppm_out_res_hist_3_folded_hist; // @[BPU.scala 266:26 668:17]
  assign predictors_io_in_bits_folded_hist_hist_2_folded_hist = s0_folded_gh_ppm_out_res_hist_2_folded_hist; // @[BPU.scala 266:26 668:17]
  assign predictors_io_in_bits_folded_hist_hist_1_folded_hist = s0_folded_gh_ppm_out_res_hist_1_folded_hist; // @[BPU.scala 266:26 668:17]
  assign predictors_io_in_bits_folded_hist_hist_0_folded_hist = s0_folded_gh_ppm_out_res_hist_0_folded_hist; // @[BPU.scala 266:26 668:17]
  assign predictors_io_ctrl_ubtb_enable = ctrl_delay_io_out_ubtb_enable; // @[BPU.scala 248:22]
  assign predictors_io_ctrl_btb_enable = ctrl_delay_io_out_btb_enable; // @[BPU.scala 248:22]
  assign predictors_io_ctrl_tage_enable = ctrl_delay_io_out_tage_enable; // @[BPU.scala 248:22]
  assign predictors_io_ctrl_sc_enable = ctrl_delay_io_out_sc_enable; // @[BPU.scala 248:22]
  assign predictors_io_ctrl_ras_enable = ctrl_delay_io_out_ras_enable; // @[BPU.scala 248:22]
  assign predictors_io_s0_fire = s1_components_ready & s1_ready; // @[BPU.scala 344:34]
  assign predictors_io_s1_fire = s1_valid & s2_ready & io_bpu_to_ftq_resp_ready; // @[BPU.scala 349:58]
  assign predictors_io_s2_fire = s2_valid; // @[BPU.scala 251:48 362:11]
  assign predictors_io_s3_fire = s3_valid; // @[BPU.scala 251:48 371:11]
  assign predictors_io_s3_redirect = s3_valid & _s3_redirect_T_1; // @[BPU.scala 568:26]
  assign predictors_io_update_valid = predictors_io_update_REG_valid; // @[BPU.scala 601:24]
  assign predictors_io_update_bits_pc = predictors_io_update_REG_bits_pc; // @[BPU.scala 601:24]
  assign predictors_io_update_bits_spec_info_folded_hist_hist_17_folded_hist =
    predictors_io_update_REG_bits_spec_info_folded_hist_hist_17_folded_hist; // @[BPU.scala 601:24]
  assign predictors_io_update_bits_spec_info_folded_hist_hist_16_folded_hist =
    predictors_io_update_REG_bits_spec_info_folded_hist_hist_16_folded_hist; // @[BPU.scala 601:24]
  assign predictors_io_update_bits_spec_info_folded_hist_hist_15_folded_hist =
    predictors_io_update_REG_bits_spec_info_folded_hist_hist_15_folded_hist; // @[BPU.scala 601:24]
  assign predictors_io_update_bits_spec_info_folded_hist_hist_14_folded_hist =
    predictors_io_update_REG_bits_spec_info_folded_hist_hist_14_folded_hist; // @[BPU.scala 601:24]
  assign predictors_io_update_bits_spec_info_folded_hist_hist_13_folded_hist =
    predictors_io_update_REG_bits_spec_info_folded_hist_hist_13_folded_hist; // @[BPU.scala 601:24]
  assign predictors_io_update_bits_spec_info_folded_hist_hist_12_folded_hist =
    predictors_io_update_REG_bits_spec_info_folded_hist_hist_12_folded_hist; // @[BPU.scala 601:24]
  assign predictors_io_update_bits_spec_info_folded_hist_hist_10_folded_hist =
    predictors_io_update_REG_bits_spec_info_folded_hist_hist_10_folded_hist; // @[BPU.scala 601:24]
  assign predictors_io_update_bits_spec_info_folded_hist_hist_9_folded_hist =
    predictors_io_update_REG_bits_spec_info_folded_hist_hist_9_folded_hist; // @[BPU.scala 601:24]
  assign predictors_io_update_bits_spec_info_folded_hist_hist_8_folded_hist =
    predictors_io_update_REG_bits_spec_info_folded_hist_hist_8_folded_hist; // @[BPU.scala 601:24]
  assign predictors_io_update_bits_spec_info_folded_hist_hist_7_folded_hist =
    predictors_io_update_REG_bits_spec_info_folded_hist_hist_7_folded_hist; // @[BPU.scala 601:24]
  assign predictors_io_update_bits_spec_info_folded_hist_hist_6_folded_hist =
    predictors_io_update_REG_bits_spec_info_folded_hist_hist_6_folded_hist; // @[BPU.scala 601:24]
  assign predictors_io_update_bits_spec_info_folded_hist_hist_5_folded_hist =
    predictors_io_update_REG_bits_spec_info_folded_hist_hist_5_folded_hist; // @[BPU.scala 601:24]
  assign predictors_io_update_bits_spec_info_folded_hist_hist_4_folded_hist =
    predictors_io_update_REG_bits_spec_info_folded_hist_hist_4_folded_hist; // @[BPU.scala 601:24]
  assign predictors_io_update_bits_spec_info_folded_hist_hist_3_folded_hist =
    predictors_io_update_REG_bits_spec_info_folded_hist_hist_3_folded_hist; // @[BPU.scala 601:24]
  assign predictors_io_update_bits_spec_info_folded_hist_hist_2_folded_hist =
    predictors_io_update_REG_bits_spec_info_folded_hist_hist_2_folded_hist; // @[BPU.scala 601:24]
  assign predictors_io_update_bits_spec_info_folded_hist_hist_1_folded_hist =
    predictors_io_update_REG_bits_spec_info_folded_hist_hist_1_folded_hist; // @[BPU.scala 601:24]
  assign predictors_io_update_bits_spec_info_folded_hist_hist_0_folded_hist =
    predictors_io_update_REG_bits_spec_info_folded_hist_hist_0_folded_hist; // @[BPU.scala 601:24]
  assign predictors_io_update_bits_ftb_entry_valid = predictors_io_update_REG_bits_ftb_entry_valid; // @[BPU.scala 601:24]
  assign predictors_io_update_bits_ftb_entry_brSlots_0_offset = predictors_io_update_REG_bits_ftb_entry_brSlots_0_offset
    ; // @[BPU.scala 601:24]
  assign predictors_io_update_bits_ftb_entry_brSlots_0_lower = predictors_io_update_REG_bits_ftb_entry_brSlots_0_lower; // @[BPU.scala 601:24]
  assign predictors_io_update_bits_ftb_entry_brSlots_0_tarStat =
    predictors_io_update_REG_bits_ftb_entry_brSlots_0_tarStat; // @[BPU.scala 601:24]
  assign predictors_io_update_bits_ftb_entry_brSlots_0_sharing =
    predictors_io_update_REG_bits_ftb_entry_brSlots_0_sharing; // @[BPU.scala 601:24]
  assign predictors_io_update_bits_ftb_entry_brSlots_0_valid = predictors_io_update_REG_bits_ftb_entry_brSlots_0_valid; // @[BPU.scala 601:24]
  assign predictors_io_update_bits_ftb_entry_tailSlot_offset = predictors_io_update_REG_bits_ftb_entry_tailSlot_offset; // @[BPU.scala 601:24]
  assign predictors_io_update_bits_ftb_entry_tailSlot_lower = predictors_io_update_REG_bits_ftb_entry_tailSlot_lower; // @[BPU.scala 601:24]
  assign predictors_io_update_bits_ftb_entry_tailSlot_tarStat = predictors_io_update_REG_bits_ftb_entry_tailSlot_tarStat
    ; // @[BPU.scala 601:24]
  assign predictors_io_update_bits_ftb_entry_tailSlot_sharing = predictors_io_update_REG_bits_ftb_entry_tailSlot_sharing
    ; // @[BPU.scala 601:24]
  assign predictors_io_update_bits_ftb_entry_tailSlot_valid = predictors_io_update_REG_bits_ftb_entry_tailSlot_valid; // @[BPU.scala 601:24]
  assign predictors_io_update_bits_ftb_entry_pftAddr = predictors_io_update_REG_bits_ftb_entry_pftAddr; // @[BPU.scala 601:24]
  assign predictors_io_update_bits_ftb_entry_carry = predictors_io_update_REG_bits_ftb_entry_carry; // @[BPU.scala 601:24]
  assign predictors_io_update_bits_ftb_entry_isCall = predictors_io_update_REG_bits_ftb_entry_isCall; // @[BPU.scala 601:24]
  assign predictors_io_update_bits_ftb_entry_isRet = predictors_io_update_REG_bits_ftb_entry_isRet; // @[BPU.scala 601:24]
  assign predictors_io_update_bits_ftb_entry_isJalr = predictors_io_update_REG_bits_ftb_entry_isJalr; // @[BPU.scala 601:24]
  assign predictors_io_update_bits_ftb_entry_last_may_be_rvi_call =
    predictors_io_update_REG_bits_ftb_entry_last_may_be_rvi_call; // @[BPU.scala 601:24]
  assign predictors_io_update_bits_ftb_entry_always_taken_0 = predictors_io_update_REG_bits_ftb_entry_always_taken_0; // @[BPU.scala 601:24]
  assign predictors_io_update_bits_ftb_entry_always_taken_1 = predictors_io_update_REG_bits_ftb_entry_always_taken_1; // @[BPU.scala 601:24]
  assign predictors_io_update_bits_br_taken_mask_0 = predictors_io_update_REG_bits_br_taken_mask_0; // @[BPU.scala 601:24]
  assign predictors_io_update_bits_br_taken_mask_1 = predictors_io_update_REG_bits_br_taken_mask_1; // @[BPU.scala 601:24]
  assign predictors_io_update_bits_jmp_taken = predictors_io_update_REG_bits_jmp_taken; // @[BPU.scala 601:24]
  assign predictors_io_update_bits_mispred_mask_0 = predictors_io_update_REG_bits_mispred_mask_0; // @[BPU.scala 601:24]
  assign predictors_io_update_bits_mispred_mask_1 = predictors_io_update_REG_bits_mispred_mask_1; // @[BPU.scala 601:24]
  assign predictors_io_update_bits_mispred_mask_2 = predictors_io_update_REG_bits_mispred_mask_2; // @[BPU.scala 601:24]
  assign predictors_io_update_bits_old_entry = predictors_io_update_REG_bits_old_entry; // @[BPU.scala 601:24]
  assign predictors_io_update_bits_meta = predictors_io_update_REG_bits_meta; // @[BPU.scala 601:24]
  assign predictors_io_update_bits_full_target = predictors_io_update_REG_bits_full_target; // @[BPU.scala 601:24]
  assign predictors_io_redirect_valid = do_redirect_valid; // @[BPU.scala 603:26]
  assign predictors_io_redirect_bits_level = do_redirect_bits_level; // @[BPU.scala 603:26]
  assign predictors_io_redirect_bits_cfiUpdate_pc = do_redirect_bits_cfiUpdate_pc; // @[BPU.scala 603:26]
  assign predictors_io_redirect_bits_cfiUpdate_pd_isRVC = do_redirect_bits_cfiUpdate_pd_isRVC; // @[BPU.scala 603:26]
  assign predictors_io_redirect_bits_cfiUpdate_pd_isCall = do_redirect_bits_cfiUpdate_pd_isCall; // @[BPU.scala 603:26]
  assign predictors_io_redirect_bits_cfiUpdate_pd_isRet = do_redirect_bits_cfiUpdate_pd_isRet; // @[BPU.scala 603:26]
  assign predictors_io_redirect_bits_cfiUpdate_rasSp = do_redirect_bits_cfiUpdate_rasSp; // @[BPU.scala 603:26]
  assign predictors_io_redirect_bits_cfiUpdate_rasEntry_retAddr = do_redirect_bits_cfiUpdate_rasEntry_retAddr; // @[BPU.scala 603:26]
  assign predictors_io_redirect_bits_cfiUpdate_rasEntry_ctr = do_redirect_bits_cfiUpdate_rasEntry_ctr; // @[BPU.scala 603:26]
  assign reset_vector_delay_clock = clock;
  assign reset_vector_delay_io_in = io_reset_vector; // @[Hold.scala 98:17]
  assign s0_pc_ppm_s2_target_sel = s2_redirect & (~s3_redirect & ~do_redirect_valid); // @[PriorityMuxGen.scala 121:41]
  assign s0_pc_ppm_s2_target_src = _s2_redirect_s1_last_pred_vec_T_5 | _s2_redirect_s1_last_pred_vec_T_3; // @[Mux.scala 27:73]
  assign s0_pc_ppm_s1_target_sel = s1_valid & (~s2_redirect & ~s3_redirect & ~do_redirect_valid); // @[PriorityMuxGen.scala 121:41]
  assign s0_pc_ppm_s1_target_src = _T_59 | _T_57; // @[Mux.scala 27:73]
  assign s0_pc_ppm_s3_target_sel = s3_redirect & ~do_redirect_valid; // @[PriorityMuxGen.scala 121:41]
  assign s0_pc_ppm_s3_target_src = _s3_redirect_on_target_T_5 | _s3_redirect_on_target_T_3; // @[Mux.scala 27:73]
  assign s0_pc_ppm_redirect_target_sel = do_redirect_valid; // @[PriorityMuxGen.scala 121:41]
  assign s0_pc_ppm_redirect_target_src = do_redirect_bits_cfiUpdate_target; // @[PriorityMuxGen.scala 140:24]
  assign s0_pc_ppm_stallPC_src = s0_pc_reg; // @[PriorityMuxGen.scala 140:24]
  assign s0_folded_gh_ppm_s2_FGH_sel = s2_redirect & (~s3_redirect & ~do_redirect_valid); // @[PriorityMuxGen.scala 121:41]
  assign s0_folded_gh_ppm_s2_FGH_src_hist_17_folded_hist = _s2_predicted_fh_T_149 | _s2_predicted_fh_T_148; // @[Mux.scala 27:73]
  assign s0_folded_gh_ppm_s2_FGH_src_hist_16_folded_hist = _s2_predicted_fh_T_144 | _s2_predicted_fh_T_143; // @[Mux.scala 27:73]
  assign s0_folded_gh_ppm_s2_FGH_src_hist_15_folded_hist = _s2_predicted_fh_T_139 | _s2_predicted_fh_T_138; // @[Mux.scala 27:73]
  assign s0_folded_gh_ppm_s2_FGH_src_hist_14_folded_hist = _s2_predicted_fh_T_134 | _s2_predicted_fh_T_133; // @[Mux.scala 27:73]
  assign s0_folded_gh_ppm_s2_FGH_src_hist_13_folded_hist = _s2_predicted_fh_T_129 | _s2_predicted_fh_T_128; // @[Mux.scala 27:73]
  assign s0_folded_gh_ppm_s2_FGH_src_hist_12_folded_hist = _s2_predicted_fh_T_124 | _s2_predicted_fh_T_123; // @[Mux.scala 27:73]
  assign s0_folded_gh_ppm_s2_FGH_src_hist_11_folded_hist = _s2_predicted_fh_T_119 | _s2_predicted_fh_T_118; // @[Mux.scala 27:73]
  assign s0_folded_gh_ppm_s2_FGH_src_hist_10_folded_hist = _s2_predicted_fh_T_114 | _s2_predicted_fh_T_113; // @[Mux.scala 27:73]
  assign s0_folded_gh_ppm_s2_FGH_src_hist_9_folded_hist = _s2_predicted_fh_T_109 | _s2_predicted_fh_T_108; // @[Mux.scala 27:73]
  assign s0_folded_gh_ppm_s2_FGH_src_hist_8_folded_hist = _s2_predicted_fh_T_104 | _s2_predicted_fh_T_103; // @[Mux.scala 27:73]
  assign s0_folded_gh_ppm_s2_FGH_src_hist_7_folded_hist = _s2_predicted_fh_T_99 | _s2_predicted_fh_T_98; // @[Mux.scala 27:73]
  assign s0_folded_gh_ppm_s2_FGH_src_hist_6_folded_hist = _s2_predicted_fh_T_94 | _s2_predicted_fh_T_93; // @[Mux.scala 27:73]
  assign s0_folded_gh_ppm_s2_FGH_src_hist_5_folded_hist = _s2_predicted_fh_T_89 | _s2_predicted_fh_T_88; // @[Mux.scala 27:73]
  assign s0_folded_gh_ppm_s2_FGH_src_hist_4_folded_hist = _s2_predicted_fh_T_84 | _s2_predicted_fh_T_83; // @[Mux.scala 27:73]
  assign s0_folded_gh_ppm_s2_FGH_src_hist_3_folded_hist = _s2_predicted_fh_T_79 | _s2_predicted_fh_T_78; // @[Mux.scala 27:73]
  assign s0_folded_gh_ppm_s2_FGH_src_hist_2_folded_hist = _s2_predicted_fh_T_74 | _s2_predicted_fh_T_73; // @[Mux.scala 27:73]
  assign s0_folded_gh_ppm_s2_FGH_src_hist_1_folded_hist = _s2_predicted_fh_T_69 | _s2_predicted_fh_T_68; // @[Mux.scala 27:73]
  assign s0_folded_gh_ppm_s2_FGH_src_hist_0_folded_hist = _s2_predicted_fh_T_64 | _s2_predicted_fh_T_63; // @[Mux.scala 27:73]
  assign s0_folded_gh_ppm_s1_FGH_sel = s1_valid & (~s2_redirect & ~s3_redirect & ~do_redirect_valid); // @[PriorityMuxGen.scala 121:41]
  assign s0_folded_gh_ppm_s1_FGH_src_hist_17_folded_hist = _s1_predicted_fh_T_149 | _s1_predicted_fh_T_148; // @[Mux.scala 27:73]
  assign s0_folded_gh_ppm_s1_FGH_src_hist_16_folded_hist = _s1_predicted_fh_T_144 | _s1_predicted_fh_T_143; // @[Mux.scala 27:73]
  assign s0_folded_gh_ppm_s1_FGH_src_hist_15_folded_hist = _s1_predicted_fh_T_139 | _s1_predicted_fh_T_138; // @[Mux.scala 27:73]
  assign s0_folded_gh_ppm_s1_FGH_src_hist_14_folded_hist = _s1_predicted_fh_T_134 | _s1_predicted_fh_T_133; // @[Mux.scala 27:73]
  assign s0_folded_gh_ppm_s1_FGH_src_hist_13_folded_hist = _s1_predicted_fh_T_129 | _s1_predicted_fh_T_128; // @[Mux.scala 27:73]
  assign s0_folded_gh_ppm_s1_FGH_src_hist_12_folded_hist = _s1_predicted_fh_T_124 | _s1_predicted_fh_T_123; // @[Mux.scala 27:73]
  assign s0_folded_gh_ppm_s1_FGH_src_hist_11_folded_hist = _s1_predicted_fh_T_119 | _s1_predicted_fh_T_118; // @[Mux.scala 27:73]
  assign s0_folded_gh_ppm_s1_FGH_src_hist_10_folded_hist = _s1_predicted_fh_T_114 | _s1_predicted_fh_T_113; // @[Mux.scala 27:73]
  assign s0_folded_gh_ppm_s1_FGH_src_hist_9_folded_hist = _s1_predicted_fh_T_109 | _s1_predicted_fh_T_108; // @[Mux.scala 27:73]
  assign s0_folded_gh_ppm_s1_FGH_src_hist_8_folded_hist = _s1_predicted_fh_T_104 | _s1_predicted_fh_T_103; // @[Mux.scala 27:73]
  assign s0_folded_gh_ppm_s1_FGH_src_hist_7_folded_hist = _s1_predicted_fh_T_99 | _s1_predicted_fh_T_98; // @[Mux.scala 27:73]
  assign s0_folded_gh_ppm_s1_FGH_src_hist_6_folded_hist = _s1_predicted_fh_T_94 | _s1_predicted_fh_T_93; // @[Mux.scala 27:73]
  assign s0_folded_gh_ppm_s1_FGH_src_hist_5_folded_hist = _s1_predicted_fh_T_89 | _s1_predicted_fh_T_88; // @[Mux.scala 27:73]
  assign s0_folded_gh_ppm_s1_FGH_src_hist_4_folded_hist = _s1_predicted_fh_T_84 | _s1_predicted_fh_T_83; // @[Mux.scala 27:73]
  assign s0_folded_gh_ppm_s1_FGH_src_hist_3_folded_hist = _s1_predicted_fh_T_79 | _s1_predicted_fh_T_78; // @[Mux.scala 27:73]
  assign s0_folded_gh_ppm_s1_FGH_src_hist_2_folded_hist = _s1_predicted_fh_T_74 | _s1_predicted_fh_T_73; // @[Mux.scala 27:73]
  assign s0_folded_gh_ppm_s1_FGH_src_hist_1_folded_hist = _s1_predicted_fh_T_69 | _s1_predicted_fh_T_68; // @[Mux.scala 27:73]
  assign s0_folded_gh_ppm_s1_FGH_src_hist_0_folded_hist = _s1_predicted_fh_T_64 | _s1_predicted_fh_T_63; // @[Mux.scala 27:73]
  assign s0_folded_gh_ppm_s3_FGH_sel = s3_redirect & ~do_redirect_valid; // @[PriorityMuxGen.scala 121:41]
  assign s0_folded_gh_ppm_s3_FGH_src_hist_17_folded_hist = _s3_predicted_fh_T_149 | _s3_predicted_fh_T_148; // @[Mux.scala 27:73]
  assign s0_folded_gh_ppm_s3_FGH_src_hist_16_folded_hist = _s3_predicted_fh_T_144 | _s3_predicted_fh_T_143; // @[Mux.scala 27:73]
  assign s0_folded_gh_ppm_s3_FGH_src_hist_15_folded_hist = _s3_predicted_fh_T_139 | _s3_predicted_fh_T_138; // @[Mux.scala 27:73]
  assign s0_folded_gh_ppm_s3_FGH_src_hist_14_folded_hist = _s3_predicted_fh_T_134 | _s3_predicted_fh_T_133; // @[Mux.scala 27:73]
  assign s0_folded_gh_ppm_s3_FGH_src_hist_13_folded_hist = _s3_predicted_fh_T_129 | _s3_predicted_fh_T_128; // @[Mux.scala 27:73]
  assign s0_folded_gh_ppm_s3_FGH_src_hist_12_folded_hist = _s3_predicted_fh_T_124 | _s3_predicted_fh_T_123; // @[Mux.scala 27:73]
  assign s0_folded_gh_ppm_s3_FGH_src_hist_11_folded_hist = _s3_predicted_fh_T_119 | _s3_predicted_fh_T_118; // @[Mux.scala 27:73]
  assign s0_folded_gh_ppm_s3_FGH_src_hist_10_folded_hist = _s3_predicted_fh_T_114 | _s3_predicted_fh_T_113; // @[Mux.scala 27:73]
  assign s0_folded_gh_ppm_s3_FGH_src_hist_9_folded_hist = _s3_predicted_fh_T_109 | _s3_predicted_fh_T_108; // @[Mux.scala 27:73]
  assign s0_folded_gh_ppm_s3_FGH_src_hist_8_folded_hist = _s3_predicted_fh_T_104 | _s3_predicted_fh_T_103; // @[Mux.scala 27:73]
  assign s0_folded_gh_ppm_s3_FGH_src_hist_7_folded_hist = _s3_predicted_fh_T_99 | _s3_predicted_fh_T_98; // @[Mux.scala 27:73]
  assign s0_folded_gh_ppm_s3_FGH_src_hist_6_folded_hist = _s3_predicted_fh_T_94 | _s3_predicted_fh_T_93; // @[Mux.scala 27:73]
  assign s0_folded_gh_ppm_s3_FGH_src_hist_5_folded_hist = _s3_predicted_fh_T_89 | _s3_predicted_fh_T_88; // @[Mux.scala 27:73]
  assign s0_folded_gh_ppm_s3_FGH_src_hist_4_folded_hist = _s3_predicted_fh_T_84 | _s3_predicted_fh_T_83; // @[Mux.scala 27:73]
  assign s0_folded_gh_ppm_s3_FGH_src_hist_3_folded_hist = _s3_predicted_fh_T_79 | _s3_predicted_fh_T_78; // @[Mux.scala 27:73]
  assign s0_folded_gh_ppm_s3_FGH_src_hist_2_folded_hist = _s3_predicted_fh_T_74 | _s3_predicted_fh_T_73; // @[Mux.scala 27:73]
  assign s0_folded_gh_ppm_s3_FGH_src_hist_1_folded_hist = _s3_predicted_fh_T_69 | _s3_predicted_fh_T_68; // @[Mux.scala 27:73]
  assign s0_folded_gh_ppm_s3_FGH_src_hist_0_folded_hist = _s3_predicted_fh_T_64 | _s3_predicted_fh_T_63; // @[Mux.scala 27:73]
  assign s0_folded_gh_ppm_redirect_FGHT_sel = do_redirect_valid; // @[PriorityMuxGen.scala 121:41]
  assign s0_folded_gh_ppm_redirect_FGHT_src_hist_17_folded_hist = 2'h2 == do_redirect_bits_cfiUpdate_shift ?
    updated_fh_res_hist_17_new_folded_hist_2 : _GEN_11764; // @[PriorityMuxGen.scala 140:{24,24}]
  assign s0_folded_gh_ppm_redirect_FGHT_src_hist_16_folded_hist = 2'h2 == do_redirect_bits_cfiUpdate_shift ?
    updated_fh_res_hist_16_new_folded_hist_2 : _GEN_11761; // @[PriorityMuxGen.scala 140:{24,24}]
  assign s0_folded_gh_ppm_redirect_FGHT_src_hist_15_folded_hist = 2'h2 == do_redirect_bits_cfiUpdate_shift ?
    updated_fh_res_hist_15_new_folded_hist_2 : _GEN_11758; // @[PriorityMuxGen.scala 140:{24,24}]
  assign s0_folded_gh_ppm_redirect_FGHT_src_hist_14_folded_hist = 2'h2 == do_redirect_bits_cfiUpdate_shift ?
    updated_fh_res_hist_14_new_folded_hist_2 : _GEN_11755; // @[PriorityMuxGen.scala 140:{24,24}]
  assign s0_folded_gh_ppm_redirect_FGHT_src_hist_13_folded_hist = 2'h2 == do_redirect_bits_cfiUpdate_shift ?
    updated_fh_res_hist_13_new_folded_hist_2 : _GEN_11752; // @[PriorityMuxGen.scala 140:{24,24}]
  assign s0_folded_gh_ppm_redirect_FGHT_src_hist_12_folded_hist = 2'h2 == do_redirect_bits_cfiUpdate_shift ?
    updated_fh_res_hist_12_new_folded_hist_2 : _GEN_11749; // @[PriorityMuxGen.scala 140:{24,24}]
  assign s0_folded_gh_ppm_redirect_FGHT_src_hist_11_folded_hist = 2'h2 == do_redirect_bits_cfiUpdate_shift ?
    updated_fh_res_hist_11_new_folded_hist_2 : _GEN_11746; // @[PriorityMuxGen.scala 140:{24,24}]
  assign s0_folded_gh_ppm_redirect_FGHT_src_hist_10_folded_hist = 2'h2 == do_redirect_bits_cfiUpdate_shift ?
    updated_fh_res_hist_10_new_folded_hist_2 : _GEN_11743; // @[PriorityMuxGen.scala 140:{24,24}]
  assign s0_folded_gh_ppm_redirect_FGHT_src_hist_9_folded_hist = 2'h2 == do_redirect_bits_cfiUpdate_shift ?
    updated_fh_res_hist_9_new_folded_hist_2 : _GEN_11740; // @[PriorityMuxGen.scala 140:{24,24}]
  assign s0_folded_gh_ppm_redirect_FGHT_src_hist_8_folded_hist = 2'h2 == do_redirect_bits_cfiUpdate_shift ?
    updated_fh_res_hist_8_new_folded_hist_2 : _GEN_11737; // @[PriorityMuxGen.scala 140:{24,24}]
  assign s0_folded_gh_ppm_redirect_FGHT_src_hist_7_folded_hist = 2'h2 == do_redirect_bits_cfiUpdate_shift ?
    updated_fh_res_hist_7_new_folded_hist_2 : _GEN_11734; // @[PriorityMuxGen.scala 140:{24,24}]
  assign s0_folded_gh_ppm_redirect_FGHT_src_hist_6_folded_hist = 2'h2 == do_redirect_bits_cfiUpdate_shift ?
    updated_fh_res_hist_6_new_folded_hist_2 : _GEN_11731; // @[PriorityMuxGen.scala 140:{24,24}]
  assign s0_folded_gh_ppm_redirect_FGHT_src_hist_5_folded_hist = 2'h2 == do_redirect_bits_cfiUpdate_shift ?
    updated_fh_res_hist_5_new_folded_hist_2 : _GEN_11728; // @[PriorityMuxGen.scala 140:{24,24}]
  assign s0_folded_gh_ppm_redirect_FGHT_src_hist_4_folded_hist = 2'h2 == do_redirect_bits_cfiUpdate_shift ?
    updated_fh_res_hist_4_new_folded_hist_2 : _GEN_11725; // @[PriorityMuxGen.scala 140:{24,24}]
  assign s0_folded_gh_ppm_redirect_FGHT_src_hist_3_folded_hist = 2'h2 == do_redirect_bits_cfiUpdate_shift ?
    updated_fh_res_hist_3_new_folded_hist_2 : _GEN_11722; // @[PriorityMuxGen.scala 140:{24,24}]
  assign s0_folded_gh_ppm_redirect_FGHT_src_hist_2_folded_hist = 2'h2 == do_redirect_bits_cfiUpdate_shift ?
    updated_fh_res_hist_2_new_folded_hist_2 : _GEN_11719; // @[PriorityMuxGen.scala 140:{24,24}]
  assign s0_folded_gh_ppm_redirect_FGHT_src_hist_1_folded_hist = 2'h2 == do_redirect_bits_cfiUpdate_shift ?
    updated_fh_res_hist_1_new_folded_hist_2 : _GEN_11716; // @[PriorityMuxGen.scala 140:{24,24}]
  assign s0_folded_gh_ppm_redirect_FGHT_src_hist_0_folded_hist = 2'h2 == do_redirect_bits_cfiUpdate_shift ?
    updated_fh_res_hist_0_new_folded_hist_2 : _GEN_11713; // @[PriorityMuxGen.scala 140:{24,24}]
  assign s0_folded_gh_ppm_stallFGH_src_hist_17_folded_hist = s0_folded_gh_reg_hist_17_folded_hist; // @[PriorityMuxGen.scala 140:24]
  assign s0_folded_gh_ppm_stallFGH_src_hist_16_folded_hist = s0_folded_gh_reg_hist_16_folded_hist; // @[PriorityMuxGen.scala 140:24]
  assign s0_folded_gh_ppm_stallFGH_src_hist_15_folded_hist = s0_folded_gh_reg_hist_15_folded_hist; // @[PriorityMuxGen.scala 140:24]
  assign s0_folded_gh_ppm_stallFGH_src_hist_14_folded_hist = s0_folded_gh_reg_hist_14_folded_hist; // @[PriorityMuxGen.scala 140:24]
  assign s0_folded_gh_ppm_stallFGH_src_hist_13_folded_hist = s0_folded_gh_reg_hist_13_folded_hist; // @[PriorityMuxGen.scala 140:24]
  assign s0_folded_gh_ppm_stallFGH_src_hist_12_folded_hist = s0_folded_gh_reg_hist_12_folded_hist; // @[PriorityMuxGen.scala 140:24]
  assign s0_folded_gh_ppm_stallFGH_src_hist_11_folded_hist = s0_folded_gh_reg_hist_11_folded_hist; // @[PriorityMuxGen.scala 140:24]
  assign s0_folded_gh_ppm_stallFGH_src_hist_10_folded_hist = s0_folded_gh_reg_hist_10_folded_hist; // @[PriorityMuxGen.scala 140:24]
  assign s0_folded_gh_ppm_stallFGH_src_hist_9_folded_hist = s0_folded_gh_reg_hist_9_folded_hist; // @[PriorityMuxGen.scala 140:24]
  assign s0_folded_gh_ppm_stallFGH_src_hist_8_folded_hist = s0_folded_gh_reg_hist_8_folded_hist; // @[PriorityMuxGen.scala 140:24]
  assign s0_folded_gh_ppm_stallFGH_src_hist_7_folded_hist = s0_folded_gh_reg_hist_7_folded_hist; // @[PriorityMuxGen.scala 140:24]
  assign s0_folded_gh_ppm_stallFGH_src_hist_6_folded_hist = s0_folded_gh_reg_hist_6_folded_hist; // @[PriorityMuxGen.scala 140:24]
  assign s0_folded_gh_ppm_stallFGH_src_hist_5_folded_hist = s0_folded_gh_reg_hist_5_folded_hist; // @[PriorityMuxGen.scala 140:24]
  assign s0_folded_gh_ppm_stallFGH_src_hist_4_folded_hist = s0_folded_gh_reg_hist_4_folded_hist; // @[PriorityMuxGen.scala 140:24]
  assign s0_folded_gh_ppm_stallFGH_src_hist_3_folded_hist = s0_folded_gh_reg_hist_3_folded_hist; // @[PriorityMuxGen.scala 140:24]
  assign s0_folded_gh_ppm_stallFGH_src_hist_2_folded_hist = s0_folded_gh_reg_hist_2_folded_hist; // @[PriorityMuxGen.scala 140:24]
  assign s0_folded_gh_ppm_stallFGH_src_hist_1_folded_hist = s0_folded_gh_reg_hist_1_folded_hist; // @[PriorityMuxGen.scala 140:24]
  assign s0_folded_gh_ppm_stallFGH_src_hist_0_folded_hist = s0_folded_gh_reg_hist_0_folded_hist; // @[PriorityMuxGen.scala 140:24]
  assign s0_ghist_ptr_ppm_s2_GHPtr_sel = s2_redirect & (~s3_redirect & ~do_redirect_valid); // @[PriorityMuxGen.scala 121:41]
  assign s0_ghist_ptr_ppm_s2_GHPtr_src_flag = _s2_redirect_s1_last_pred_vec_T_12 &
    s2_possible_predicted_ghist_ptrs_0_flag | _s2_redirect_s1_last_pred_vec_T_40 &
    s2_possible_predicted_ghist_ptrs_1_flag | _s2_redirect_s1_last_pred_vec_T_68 &
    s2_possible_predicted_ghist_ptrs_2_flag; // @[Mux.scala 27:73]
  assign s0_ghist_ptr_ppm_s2_GHPtr_src_value = _s2_predicted_ghist_ptr_T_64 | _s2_predicted_ghist_ptr_T_63; // @[Mux.scala 27:73]
  assign s0_ghist_ptr_ppm_s1_GHPtr_sel = s1_valid & (~s2_redirect & ~s3_redirect & ~do_redirect_valid); // @[PriorityMuxGen.scala 121:41]
  assign s0_ghist_ptr_ppm_s1_GHPtr_src_flag = _s1_predicted_ghist_ptr_T_4 & s1_possible_predicted_ghist_ptrs_0_flag |
    _s1_predicted_ghist_ptr_T_32 & s1_possible_predicted_ghist_ptrs_1_flag | _s1_predicted_ghist_ptr_T_60 &
    s1_possible_predicted_ghist_ptrs_2_flag; // @[Mux.scala 27:73]
  assign s0_ghist_ptr_ppm_s1_GHPtr_src_value = _s1_predicted_ghist_ptr_T_64 | _s1_predicted_ghist_ptr_T_63; // @[Mux.scala 27:73]
  assign s0_ghist_ptr_ppm_s3_GHPtr_sel = s3_redirect & ~do_redirect_valid; // @[PriorityMuxGen.scala 121:41]
  assign s0_ghist_ptr_ppm_s3_GHPtr_src_flag = _s3_predicted_ghist_ptr_T_4 & s3_possible_predicted_ghist_ptrs_0_flag |
    _s3_predicted_ghist_ptr_T_32 & s3_possible_predicted_ghist_ptrs_1_flag | _s3_predicted_ghist_ptr_T_60 &
    s3_possible_predicted_ghist_ptrs_2_flag; // @[Mux.scala 27:73]
  assign s0_ghist_ptr_ppm_s3_GHPtr_src_value = _s3_predicted_ghist_ptr_T_64 | _s3_predicted_ghist_ptr_T_63; // @[Mux.scala 27:73]
  assign s0_ghist_ptr_ppm_redirect_GHPtr_sel = do_redirect_valid; // @[PriorityMuxGen.scala 121:41]
  assign s0_ghist_ptr_ppm_redirect_GHPtr_src_flag = ~updated_ptr_flipped_new_ptr_flag; // @[CircularQueuePtr.scala 56:21]
  assign s0_ghist_ptr_ppm_redirect_GHPtr_src_value = _updated_ptr_flipped_new_ptr_new_ptr_value_T_1[7:0]; // @[CircularQueuePtr.scala 37:23 45:21]
  assign s0_ghist_ptr_ppm_stallGHPtr_src_flag = s0_ghist_ptr_reg_flag; // @[PriorityMuxGen.scala 140:24]
  assign s0_ghist_ptr_ppm_stallGHPtr_src_value = s0_ghist_ptr_reg_value; // @[PriorityMuxGen.scala 140:24]
  assign s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_sel = s2_redirect & (~s3_redirect & ~do_redirect_valid); // @[PriorityMuxGen.scala 121:41]
  assign s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_src_afhob_5_bits_0 = 8'h8f == new_ptr_31_value ? ghv_143 : _GEN_5478; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_src_afhob_5_bits_1 = 8'h8f == new_ptr_27_value ? ghv_143 : _GEN_5622; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_src_afhob_5_bits_2 = 8'h8f == new_ptr_25_value ? ghv_143 : _GEN_5766; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_src_afhob_5_bits_3 = 8'h8f == new_ptr_20_value ? ghv_143 : _GEN_5910; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_src_afhob_4_bits_0 = 8'h8f == new_ptr_33_value ? ghv_143 : _GEN_3462; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_src_afhob_4_bits_1 = 8'h8f == new_ptr_26_value ? ghv_143 : _GEN_3606; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_src_afhob_4_bits_2 = 8'h8f == new_ptr_21_value ? ghv_143 : _GEN_5190; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_src_afhob_4_bits_3 = 8'h8f == new_ptr_38_value ? ghv_143 : _GEN_5334; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_src_afhob_3_bits_0 = 8'h8f == new_ptr_39_value ? ghv_143 : _GEN_4758; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_src_afhob_3_bits_1 = 8'h8f == new_ptr_23_value ? ghv_143 : _GEN_4902; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_src_afhob_3_bits_2 = 8'h8f == new_ptr_30_value ? ghv_143 : _GEN_5046; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_src_afhob_3_bits_3 = 8'h8f == new_ptr_32_value ? ghv_143 : _GEN_3750; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_src_afhob_2_bits_0 = 8'h8f == new_ptr_34_value ? ghv_143 : _GEN_4182; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_src_afhob_2_bits_1 = 8'h8f == new_ptr_37_value ? ghv_143 : _GEN_4326; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_src_afhob_2_bits_2 = 8'h8f == new_ptr_24_value ? ghv_143 : _GEN_4470; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_src_afhob_2_bits_3 = 8'h8f == new_ptr_28_value ? ghv_143 : _GEN_4614; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_src_afhob_1_bits_0 = 8'h8f == new_ptr_32_value ? ghv_143 : _GEN_3750; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_src_afhob_1_bits_1 = 8'h8f == new_ptr_35_value ? ghv_143 : _GEN_3894; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_src_afhob_1_bits_2 = 8'h8f == new_ptr_22_value ? ghv_143 : _GEN_4038; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_src_afhob_1_bits_3 = 8'h8f == new_ptr_29_value ? ghv_143 : _GEN_3174; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_src_afhob_0_bits_0 = 8'h8f == new_ptr_29_value ? ghv_143 : _GEN_3174; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_src_afhob_0_bits_1 = 8'h8f == new_ptr_36_value ? ghv_143 : _GEN_3318; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_src_afhob_0_bits_2 = 8'h8f == new_ptr_33_value ? ghv_143 : _GEN_3462; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_s2_AFHOB_src_afhob_0_bits_3 = 8'h8f == new_ptr_26_value ? ghv_143 : _GEN_3606; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_sel = s1_valid & (~s2_redirect & ~s3_redirect & ~do_redirect_valid); // @[PriorityMuxGen.scala 121:41]
  assign s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_src_afhob_5_bits_0 = 8'h8f == new_ptr_11_value ? ghv_143 : _GEN_2595; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_src_afhob_5_bits_1 = 8'h8f == new_ptr_7_value ? ghv_143 : _GEN_2739; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_src_afhob_5_bits_2 = 8'h8f == new_ptr_5_value ? ghv_143 : _GEN_2883; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_src_afhob_5_bits_3 = 8'h8f == new_ptr_value ? ghv_143 : _GEN_3027; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_src_afhob_4_bits_0 = 8'h8f == new_ptr_13_value ? ghv_143 : _GEN_579; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_src_afhob_4_bits_1 = 8'h8f == new_ptr_6_value ? ghv_143 : _GEN_723; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_src_afhob_4_bits_2 = 8'h8f == new_ptr_1_value ? ghv_143 : _GEN_2307; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_src_afhob_4_bits_3 = 8'h8f == new_ptr_18_value ? ghv_143 : _GEN_2451; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_src_afhob_3_bits_0 = 8'h8f == new_ptr_19_value ? ghv_143 : _GEN_1875; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_src_afhob_3_bits_1 = 8'h8f == new_ptr_3_value ? ghv_143 : _GEN_2019; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_src_afhob_3_bits_2 = 8'h8f == new_ptr_10_value ? ghv_143 : _GEN_2163; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_src_afhob_3_bits_3 = 8'h8f == new_ptr_12_value ? ghv_143 : _GEN_867; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_src_afhob_2_bits_0 = 8'h8f == new_ptr_14_value ? ghv_143 : _GEN_1299; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_src_afhob_2_bits_1 = 8'h8f == new_ptr_17_value ? ghv_143 : _GEN_1443; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_src_afhob_2_bits_2 = 8'h8f == new_ptr_4_value ? ghv_143 : _GEN_1587; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_src_afhob_2_bits_3 = 8'h8f == new_ptr_8_value ? ghv_143 : _GEN_1731; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_src_afhob_1_bits_0 = 8'h8f == new_ptr_12_value ? ghv_143 : _GEN_867; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_src_afhob_1_bits_1 = 8'h8f == new_ptr_15_value ? ghv_143 : _GEN_1011; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_src_afhob_1_bits_2 = 8'h8f == new_ptr_2_value ? ghv_143 : _GEN_1155; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_src_afhob_1_bits_3 = 8'h8f == new_ptr_9_value ? ghv_143 : _GEN_291; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_src_afhob_0_bits_0 = 8'h8f == new_ptr_9_value ? ghv_143 : _GEN_291; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_src_afhob_0_bits_1 = 8'h8f == new_ptr_16_value ? ghv_143 : _GEN_435; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_src_afhob_0_bits_2 = 8'h8f == new_ptr_13_value ? ghv_143 : _GEN_579; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_s1_AFHOB_src_afhob_0_bits_3 = 8'h8f == new_ptr_6_value ? ghv_143 : _GEN_723; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_sel = s3_redirect & ~do_redirect_valid; // @[PriorityMuxGen.scala 121:41]
  assign s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_src_afhob_5_bits_0 = 8'h8f == new_ptr_51_value ? ghv_143 : _GEN_8365; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_src_afhob_5_bits_1 = 8'h8f == new_ptr_47_value ? ghv_143 : _GEN_8509; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_src_afhob_5_bits_2 = 8'h8f == new_ptr_45_value ? ghv_143 : _GEN_8653; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_src_afhob_5_bits_3 = 8'h8f == new_ptr_40_value ? ghv_143 : _GEN_8797; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_src_afhob_4_bits_0 = 8'h8f == new_ptr_53_value ? ghv_143 : _GEN_6349; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_src_afhob_4_bits_1 = 8'h8f == new_ptr_46_value ? ghv_143 : _GEN_6493; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_src_afhob_4_bits_2 = 8'h8f == new_ptr_41_value ? ghv_143 : _GEN_8077; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_src_afhob_4_bits_3 = 8'h8f == new_ptr_58_value ? ghv_143 : _GEN_8221; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_src_afhob_3_bits_0 = 8'h8f == new_ptr_59_value ? ghv_143 : _GEN_7645; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_src_afhob_3_bits_1 = 8'h8f == new_ptr_43_value ? ghv_143 : _GEN_7789; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_src_afhob_3_bits_2 = 8'h8f == new_ptr_50_value ? ghv_143 : _GEN_7933; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_src_afhob_3_bits_3 = 8'h8f == new_ptr_52_value ? ghv_143 : _GEN_6637; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_src_afhob_2_bits_0 = 8'h8f == new_ptr_54_value ? ghv_143 : _GEN_7069; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_src_afhob_2_bits_1 = 8'h8f == new_ptr_57_value ? ghv_143 : _GEN_7213; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_src_afhob_2_bits_2 = 8'h8f == new_ptr_44_value ? ghv_143 : _GEN_7357; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_src_afhob_2_bits_3 = 8'h8f == new_ptr_48_value ? ghv_143 : _GEN_7501; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_src_afhob_1_bits_0 = 8'h8f == new_ptr_52_value ? ghv_143 : _GEN_6637; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_src_afhob_1_bits_1 = 8'h8f == new_ptr_55_value ? ghv_143 : _GEN_6781; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_src_afhob_1_bits_2 = 8'h8f == new_ptr_42_value ? ghv_143 : _GEN_6925; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_src_afhob_1_bits_3 = 8'h8f == new_ptr_49_value ? ghv_143 : _GEN_6061; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_src_afhob_0_bits_0 = 8'h8f == new_ptr_49_value ? ghv_143 : _GEN_6061; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_src_afhob_0_bits_1 = 8'h8f == new_ptr_56_value ? ghv_143 : _GEN_6205; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_src_afhob_0_bits_2 = 8'h8f == new_ptr_53_value ? ghv_143 : _GEN_6349; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_s3_AFHOB_src_afhob_0_bits_3 = 8'h8f == new_ptr_46_value ? ghv_143 : _GEN_6493; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_sel = do_redirect_valid; // @[PriorityMuxGen.scala 121:41]
  assign s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_src_afhob_5_bits_0 = 8'h8f == new_ptr_71_value ? ghv_143 :
    _GEN_11275; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_src_afhob_5_bits_1 = 8'h8f == new_ptr_67_value ? ghv_143 :
    _GEN_11419; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_src_afhob_5_bits_2 = 8'h8f == new_ptr_65_value ? ghv_143 :
    _GEN_11563; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_src_afhob_5_bits_3 = 8'h8f == new_ptr_60_value ? ghv_143 :
    _GEN_11707; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_src_afhob_4_bits_0 = 8'h8f == new_ptr_73_value ? ghv_143 : _GEN_9259
    ; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_src_afhob_4_bits_1 = 8'h8f == new_ptr_66_value ? ghv_143 : _GEN_9403
    ; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_src_afhob_4_bits_2 = 8'h8f == new_ptr_61_value ? ghv_143 :
    _GEN_10987; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_src_afhob_4_bits_3 = 8'h8f == new_ptr_78_value ? ghv_143 :
    _GEN_11131; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_src_afhob_3_bits_0 = 8'h8f == new_ptr_79_value ? ghv_143 :
    _GEN_10555; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_src_afhob_3_bits_1 = 8'h8f == new_ptr_63_value ? ghv_143 :
    _GEN_10699; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_src_afhob_3_bits_2 = 8'h8f == new_ptr_70_value ? ghv_143 :
    _GEN_10843; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_src_afhob_3_bits_3 = 8'h8f == new_ptr_72_value ? ghv_143 : _GEN_9547
    ; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_src_afhob_2_bits_0 = 8'h8f == new_ptr_74_value ? ghv_143 : _GEN_9979
    ; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_src_afhob_2_bits_1 = 8'h8f == new_ptr_77_value ? ghv_143 :
    _GEN_10123; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_src_afhob_2_bits_2 = 8'h8f == new_ptr_64_value ? ghv_143 :
    _GEN_10267; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_src_afhob_2_bits_3 = 8'h8f == new_ptr_68_value ? ghv_143 :
    _GEN_10411; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_src_afhob_1_bits_0 = 8'h8f == new_ptr_72_value ? ghv_143 : _GEN_9547
    ; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_src_afhob_1_bits_1 = 8'h8f == new_ptr_75_value ? ghv_143 : _GEN_9691
    ; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_src_afhob_1_bits_2 = 8'h8f == new_ptr_62_value ? ghv_143 : _GEN_9835
    ; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_src_afhob_1_bits_3 = 8'h8f == new_ptr_69_value ? ghv_143 : _GEN_8971
    ; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_src_afhob_0_bits_0 = 8'h8f == new_ptr_69_value ? ghv_143 : _GEN_8971
    ; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_src_afhob_0_bits_1 = 8'h8f == new_ptr_76_value ? ghv_143 : _GEN_9115
    ; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_src_afhob_0_bits_2 = 8'h8f == new_ptr_73_value ? ghv_143 : _GEN_9259
    ; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_redirect_AFHOB_src_afhob_0_bits_3 = 8'h8f == new_ptr_66_value ? ghv_143 : _GEN_9403
    ; // @[FrontendBundle.scala 329:{20,20}]
  assign s0_ahead_fh_oldest_bits_ppm_stallAFHOB_src_afhob_5_bits_0 = s0_ahead_fh_oldest_bits_reg_afhob_5_bits_0; // @[PriorityMuxGen.scala 140:24]
  assign s0_ahead_fh_oldest_bits_ppm_stallAFHOB_src_afhob_5_bits_1 = s0_ahead_fh_oldest_bits_reg_afhob_5_bits_1; // @[PriorityMuxGen.scala 140:24]
  assign s0_ahead_fh_oldest_bits_ppm_stallAFHOB_src_afhob_5_bits_2 = s0_ahead_fh_oldest_bits_reg_afhob_5_bits_2; // @[PriorityMuxGen.scala 140:24]
  assign s0_ahead_fh_oldest_bits_ppm_stallAFHOB_src_afhob_5_bits_3 = s0_ahead_fh_oldest_bits_reg_afhob_5_bits_3; // @[PriorityMuxGen.scala 140:24]
  assign s0_ahead_fh_oldest_bits_ppm_stallAFHOB_src_afhob_4_bits_0 = s0_ahead_fh_oldest_bits_reg_afhob_4_bits_0; // @[PriorityMuxGen.scala 140:24]
  assign s0_ahead_fh_oldest_bits_ppm_stallAFHOB_src_afhob_4_bits_1 = s0_ahead_fh_oldest_bits_reg_afhob_4_bits_1; // @[PriorityMuxGen.scala 140:24]
  assign s0_ahead_fh_oldest_bits_ppm_stallAFHOB_src_afhob_4_bits_2 = s0_ahead_fh_oldest_bits_reg_afhob_4_bits_2; // @[PriorityMuxGen.scala 140:24]
  assign s0_ahead_fh_oldest_bits_ppm_stallAFHOB_src_afhob_4_bits_3 = s0_ahead_fh_oldest_bits_reg_afhob_4_bits_3; // @[PriorityMuxGen.scala 140:24]
  assign s0_ahead_fh_oldest_bits_ppm_stallAFHOB_src_afhob_3_bits_0 = s0_ahead_fh_oldest_bits_reg_afhob_3_bits_0; // @[PriorityMuxGen.scala 140:24]
  assign s0_ahead_fh_oldest_bits_ppm_stallAFHOB_src_afhob_3_bits_1 = s0_ahead_fh_oldest_bits_reg_afhob_3_bits_1; // @[PriorityMuxGen.scala 140:24]
  assign s0_ahead_fh_oldest_bits_ppm_stallAFHOB_src_afhob_3_bits_2 = s0_ahead_fh_oldest_bits_reg_afhob_3_bits_2; // @[PriorityMuxGen.scala 140:24]
  assign s0_ahead_fh_oldest_bits_ppm_stallAFHOB_src_afhob_3_bits_3 = s0_ahead_fh_oldest_bits_reg_afhob_3_bits_3; // @[PriorityMuxGen.scala 140:24]
  assign s0_ahead_fh_oldest_bits_ppm_stallAFHOB_src_afhob_2_bits_0 = s0_ahead_fh_oldest_bits_reg_afhob_2_bits_0; // @[PriorityMuxGen.scala 140:24]
  assign s0_ahead_fh_oldest_bits_ppm_stallAFHOB_src_afhob_2_bits_1 = s0_ahead_fh_oldest_bits_reg_afhob_2_bits_1; // @[PriorityMuxGen.scala 140:24]
  assign s0_ahead_fh_oldest_bits_ppm_stallAFHOB_src_afhob_2_bits_2 = s0_ahead_fh_oldest_bits_reg_afhob_2_bits_2; // @[PriorityMuxGen.scala 140:24]
  assign s0_ahead_fh_oldest_bits_ppm_stallAFHOB_src_afhob_2_bits_3 = s0_ahead_fh_oldest_bits_reg_afhob_2_bits_3; // @[PriorityMuxGen.scala 140:24]
  assign s0_ahead_fh_oldest_bits_ppm_stallAFHOB_src_afhob_1_bits_0 = s0_ahead_fh_oldest_bits_reg_afhob_1_bits_0; // @[PriorityMuxGen.scala 140:24]
  assign s0_ahead_fh_oldest_bits_ppm_stallAFHOB_src_afhob_1_bits_1 = s0_ahead_fh_oldest_bits_reg_afhob_1_bits_1; // @[PriorityMuxGen.scala 140:24]
  assign s0_ahead_fh_oldest_bits_ppm_stallAFHOB_src_afhob_1_bits_2 = s0_ahead_fh_oldest_bits_reg_afhob_1_bits_2; // @[PriorityMuxGen.scala 140:24]
  assign s0_ahead_fh_oldest_bits_ppm_stallAFHOB_src_afhob_1_bits_3 = s0_ahead_fh_oldest_bits_reg_afhob_1_bits_3; // @[PriorityMuxGen.scala 140:24]
  assign s0_ahead_fh_oldest_bits_ppm_stallAFHOB_src_afhob_0_bits_0 = s0_ahead_fh_oldest_bits_reg_afhob_0_bits_0; // @[PriorityMuxGen.scala 140:24]
  assign s0_ahead_fh_oldest_bits_ppm_stallAFHOB_src_afhob_0_bits_1 = s0_ahead_fh_oldest_bits_reg_afhob_0_bits_1; // @[PriorityMuxGen.scala 140:24]
  assign s0_ahead_fh_oldest_bits_ppm_stallAFHOB_src_afhob_0_bits_2 = s0_ahead_fh_oldest_bits_reg_afhob_0_bits_2; // @[PriorityMuxGen.scala 140:24]
  assign s0_ahead_fh_oldest_bits_ppm_stallAFHOB_src_afhob_0_bits_3 = s0_ahead_fh_oldest_bits_reg_afhob_0_bits_3; // @[PriorityMuxGen.scala 140:24]
  assign s0_last_br_num_oh_ppm_s2_BrNumOH_sel = s2_redirect & (~s3_redirect & ~do_redirect_valid); // @[PriorityMuxGen.scala 121:41]
  assign s0_last_br_num_oh_ppm_s2_BrNumOH_src = {s2_redirect_s1_last_pred_vec_hi,_s2_redirect_s1_last_pred_vec_T_12}; // @[BPU.scala 508:60]
  assign s0_last_br_num_oh_ppm_s1_BrNumOH_sel = s1_valid & (~s2_redirect & ~s3_redirect & ~do_redirect_valid); // @[PriorityMuxGen.scala 121:41]
  assign s0_last_br_num_oh_ppm_s1_BrNumOH_src = {hi,_s1_predicted_ghist_ptr_T_4}; // @[BPU.scala 435:57]
  assign s0_last_br_num_oh_ppm_s3_BrNumOH_sel = s3_redirect & ~do_redirect_valid; // @[PriorityMuxGen.scala 121:41]
  assign s0_last_br_num_oh_ppm_s3_BrNumOH_src = {hi_2,_s3_predicted_ghist_ptr_T_4}; // @[BPU.scala 579:60]
  assign s0_last_br_num_oh_ppm_redirect_BrNumOH_sel = do_redirect_valid; // @[PriorityMuxGen.scala 121:41]
  assign s0_last_br_num_oh_ppm_redirect_BrNumOH_src = _thisBrNumOH_T[2:0]; // @[OneHot.scala 64:27]
  assign s0_last_br_num_oh_ppm_stallBrNumOH_src = s0_last_br_num_oh_reg; // @[PriorityMuxGen.scala 140:24]
  assign ghv_write_datas_0_ppm_s2_new_bit_0_sel = _T_385 & (~_T_666 & ~_T_812); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_0_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_26 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_53 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_0_ppm_s1_new_bit_0_sel = _T_123 & (~_T_385 & ~_T_666 & ~_T_812); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_0_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_26 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_53 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_0_ppm_s3_new_bit_0_sel = _T_666 & ~_T_812; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_0_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_26 & _s3_redirect_on_br_taken_T_5 | _s3_ghv_wens_T_53
     & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_0_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_1 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_3 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_1_ppm_s2_new_bit_0_sel = _T_386 & (~_T_667 & ~_T_813); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_1_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_80 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_107 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_1_ppm_s1_new_bit_0_sel = _T_124 & (~_T_386 & ~_T_667 & ~_T_813); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_1_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_80 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_107 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_1_ppm_s3_new_bit_0_sel = _T_667 & ~_T_813; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_1_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_80 & _s3_redirect_on_br_taken_T_5 | _s3_ghv_wens_T_107
     & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_1_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_5 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_7 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_2_ppm_s2_new_bit_0_sel = _T_387 & (~_T_668 & ~_T_814); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_2_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_134 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_161 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_2_ppm_s1_new_bit_0_sel = _T_125 & (~_T_387 & ~_T_668 & ~_T_814); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_2_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_134 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_161 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_2_ppm_s3_new_bit_0_sel = _T_668 & ~_T_814; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_2_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_134 & _s3_redirect_on_br_taken_T_5 | _s3_ghv_wens_T_161
     & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_2_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_9 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_11 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_3_ppm_s2_new_bit_0_sel = _T_388 & (~_T_669 & ~_T_815); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_3_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_188 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_215 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_3_ppm_s1_new_bit_0_sel = _T_126 & (~_T_388 & ~_T_669 & ~_T_815); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_3_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_188 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_215 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_3_ppm_s3_new_bit_0_sel = _T_669 & ~_T_815; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_3_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_188 & _s3_redirect_on_br_taken_T_5 | _s3_ghv_wens_T_215
     & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_3_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_13 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_15 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_4_ppm_s2_new_bit_0_sel = _T_389 & (~_T_670 & ~_T_816); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_4_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_242 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_269 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_4_ppm_s1_new_bit_0_sel = _T_127 & (~_T_389 & ~_T_670 & ~_T_816); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_4_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_242 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_269 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_4_ppm_s3_new_bit_0_sel = _T_670 & ~_T_816; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_4_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_242 & _s3_redirect_on_br_taken_T_5 | _s3_ghv_wens_T_269
     & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_4_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_17 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_19 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_5_ppm_s2_new_bit_0_sel = _T_390 & (~_T_671 & ~_T_817); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_5_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_296 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_323 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_5_ppm_s1_new_bit_0_sel = _T_128 & (~_T_390 & ~_T_671 & ~_T_817); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_5_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_296 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_323 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_5_ppm_s3_new_bit_0_sel = _T_671 & ~_T_817; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_5_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_296 & _s3_redirect_on_br_taken_T_5 | _s3_ghv_wens_T_323
     & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_5_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_21 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_23 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_6_ppm_s2_new_bit_0_sel = _T_391 & (~_T_672 & ~_T_818); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_6_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_350 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_377 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_6_ppm_s1_new_bit_0_sel = _T_129 & (~_T_391 & ~_T_672 & ~_T_818); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_6_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_350 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_377 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_6_ppm_s3_new_bit_0_sel = _T_672 & ~_T_818; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_6_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_350 & _s3_redirect_on_br_taken_T_5 | _s3_ghv_wens_T_377
     & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_6_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_25 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_27 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_7_ppm_s2_new_bit_0_sel = _T_392 & (~_T_673 & ~_T_819); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_7_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_404 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_431 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_7_ppm_s1_new_bit_0_sel = _T_130 & (~_T_392 & ~_T_673 & ~_T_819); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_7_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_404 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_431 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_7_ppm_s3_new_bit_0_sel = _T_673 & ~_T_819; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_7_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_404 & _s3_redirect_on_br_taken_T_5 | _s3_ghv_wens_T_431
     & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_7_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_29 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_31 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_8_ppm_s2_new_bit_0_sel = _T_393 & (~_T_674 & ~_T_820); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_8_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_458 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_485 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_8_ppm_s1_new_bit_0_sel = _T_131 & (~_T_393 & ~_T_674 & ~_T_820); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_8_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_458 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_485 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_8_ppm_s3_new_bit_0_sel = _T_674 & ~_T_820; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_8_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_458 & _s3_redirect_on_br_taken_T_5 | _s3_ghv_wens_T_485
     & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_8_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_33 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_35 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_9_ppm_s2_new_bit_0_sel = _T_394 & (~_T_675 & ~_T_821); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_9_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_512 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_539 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_9_ppm_s1_new_bit_0_sel = _T_132 & (~_T_394 & ~_T_675 & ~_T_821); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_9_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_512 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_539 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_9_ppm_s3_new_bit_0_sel = _T_675 & ~_T_821; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_9_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_512 & _s3_redirect_on_br_taken_T_5 | _s3_ghv_wens_T_539
     & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_9_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_37 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_39 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_10_ppm_s2_new_bit_0_sel = _T_395 & (~_T_676 & ~_T_822); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_10_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_566 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_593 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_10_ppm_s1_new_bit_0_sel = _T_133 & (~_T_395 & ~_T_676 & ~_T_822); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_10_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_566 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_593 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_10_ppm_s3_new_bit_0_sel = _T_676 & ~_T_822; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_10_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_566 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_593 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_10_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_41 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_43 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_11_ppm_s2_new_bit_0_sel = _T_396 & (~_T_677 & ~_T_823); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_11_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_620 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_647 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_11_ppm_s1_new_bit_0_sel = _T_134 & (~_T_396 & ~_T_677 & ~_T_823); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_11_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_620 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_647 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_11_ppm_s3_new_bit_0_sel = _T_677 & ~_T_823; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_11_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_620 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_647 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_11_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_45 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_47 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_12_ppm_s2_new_bit_0_sel = _T_397 & (~_T_678 & ~_T_824); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_12_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_674 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_701 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_12_ppm_s1_new_bit_0_sel = _T_135 & (~_T_397 & ~_T_678 & ~_T_824); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_12_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_674 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_701 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_12_ppm_s3_new_bit_0_sel = _T_678 & ~_T_824; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_12_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_674 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_701 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_12_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_49 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_51 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_13_ppm_s2_new_bit_0_sel = _T_398 & (~_T_679 & ~_T_825); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_13_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_728 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_755 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_13_ppm_s1_new_bit_0_sel = _T_136 & (~_T_398 & ~_T_679 & ~_T_825); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_13_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_728 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_755 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_13_ppm_s3_new_bit_0_sel = _T_679 & ~_T_825; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_13_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_728 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_755 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_13_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_53 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_55 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_14_ppm_s2_new_bit_0_sel = _T_399 & (~_T_680 & ~_T_826); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_14_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_782 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_809 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_14_ppm_s1_new_bit_0_sel = _T_137 & (~_T_399 & ~_T_680 & ~_T_826); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_14_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_782 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_809 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_14_ppm_s3_new_bit_0_sel = _T_680 & ~_T_826; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_14_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_782 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_809 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_14_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_57 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_59 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_15_ppm_s2_new_bit_0_sel = _T_400 & (~_T_681 & ~_T_827); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_15_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_836 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_863 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_15_ppm_s1_new_bit_0_sel = _T_138 & (~_T_400 & ~_T_681 & ~_T_827); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_15_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_836 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_863 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_15_ppm_s3_new_bit_0_sel = _T_681 & ~_T_827; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_15_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_836 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_863 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_15_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_61 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_63 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_16_ppm_s2_new_bit_0_sel = _T_401 & (~_T_682 & ~_T_828); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_16_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_890 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_917 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_16_ppm_s1_new_bit_0_sel = _T_139 & (~_T_401 & ~_T_682 & ~_T_828); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_16_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_890 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_917 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_16_ppm_s3_new_bit_0_sel = _T_682 & ~_T_828; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_16_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_890 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_917 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_16_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_65 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_67 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_17_ppm_s2_new_bit_0_sel = _T_402 & (~_T_683 & ~_T_829); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_17_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_944 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_971 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_17_ppm_s1_new_bit_0_sel = _T_140 & (~_T_402 & ~_T_683 & ~_T_829); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_17_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_944 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_971 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_17_ppm_s3_new_bit_0_sel = _T_683 & ~_T_829; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_17_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_944 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_971 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_17_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_69 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_71 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_18_ppm_s2_new_bit_0_sel = _T_403 & (~_T_684 & ~_T_830); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_18_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_998 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_1025 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_18_ppm_s1_new_bit_0_sel = _T_141 & (~_T_403 & ~_T_684 & ~_T_830); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_18_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_998 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_1025 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_18_ppm_s3_new_bit_0_sel = _T_684 & ~_T_830; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_18_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_998 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_1025 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_18_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_73 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_75 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_19_ppm_s2_new_bit_0_sel = _T_404 & (~_T_685 & ~_T_831); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_19_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_1052 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_1079 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_19_ppm_s1_new_bit_0_sel = _T_142 & (~_T_404 & ~_T_685 & ~_T_831); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_19_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_1052 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_1079 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_19_ppm_s3_new_bit_0_sel = _T_685 & ~_T_831; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_19_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_1052 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_1079 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_19_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_77 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_79 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_20_ppm_s2_new_bit_0_sel = _T_405 & (~_T_686 & ~_T_832); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_20_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_1106 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_1133 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_20_ppm_s1_new_bit_0_sel = _T_143 & (~_T_405 & ~_T_686 & ~_T_832); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_20_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_1106 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_1133 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_20_ppm_s3_new_bit_0_sel = _T_686 & ~_T_832; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_20_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_1106 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_1133 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_20_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_81 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_83 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_21_ppm_s2_new_bit_0_sel = _T_406 & (~_T_687 & ~_T_833); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_21_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_1160 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_1187 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_21_ppm_s1_new_bit_0_sel = _T_144 & (~_T_406 & ~_T_687 & ~_T_833); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_21_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_1160 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_1187 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_21_ppm_s3_new_bit_0_sel = _T_687 & ~_T_833; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_21_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_1160 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_1187 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_21_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_85 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_87 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_22_ppm_s2_new_bit_0_sel = _T_407 & (~_T_688 & ~_T_834); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_22_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_1214 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_1241 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_22_ppm_s1_new_bit_0_sel = _T_145 & (~_T_407 & ~_T_688 & ~_T_834); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_22_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_1214 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_1241 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_22_ppm_s3_new_bit_0_sel = _T_688 & ~_T_834; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_22_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_1214 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_1241 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_22_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_89 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_91 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_23_ppm_s2_new_bit_0_sel = _T_408 & (~_T_689 & ~_T_835); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_23_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_1268 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_1295 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_23_ppm_s1_new_bit_0_sel = _T_146 & (~_T_408 & ~_T_689 & ~_T_835); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_23_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_1268 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_1295 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_23_ppm_s3_new_bit_0_sel = _T_689 & ~_T_835; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_23_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_1268 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_1295 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_23_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_93 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_95 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_24_ppm_s2_new_bit_0_sel = _T_409 & (~_T_690 & ~_T_836); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_24_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_1322 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_1349 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_24_ppm_s1_new_bit_0_sel = _T_147 & (~_T_409 & ~_T_690 & ~_T_836); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_24_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_1322 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_1349 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_24_ppm_s3_new_bit_0_sel = _T_690 & ~_T_836; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_24_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_1322 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_1349 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_24_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_97 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_99 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_25_ppm_s2_new_bit_0_sel = _T_410 & (~_T_691 & ~_T_837); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_25_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_1376 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_1403 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_25_ppm_s1_new_bit_0_sel = _T_148 & (~_T_410 & ~_T_691 & ~_T_837); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_25_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_1376 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_1403 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_25_ppm_s3_new_bit_0_sel = _T_691 & ~_T_837; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_25_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_1376 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_1403 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_25_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_101 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_103 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_26_ppm_s2_new_bit_0_sel = _T_411 & (~_T_692 & ~_T_838); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_26_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_1430 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_1457 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_26_ppm_s1_new_bit_0_sel = _T_149 & (~_T_411 & ~_T_692 & ~_T_838); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_26_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_1430 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_1457 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_26_ppm_s3_new_bit_0_sel = _T_692 & ~_T_838; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_26_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_1430 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_1457 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_26_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_105 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_107 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_27_ppm_s2_new_bit_0_sel = _T_412 & (~_T_693 & ~_T_839); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_27_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_1484 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_1511 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_27_ppm_s1_new_bit_0_sel = _T_150 & (~_T_412 & ~_T_693 & ~_T_839); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_27_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_1484 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_1511 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_27_ppm_s3_new_bit_0_sel = _T_693 & ~_T_839; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_27_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_1484 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_1511 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_27_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_109 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_111 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_28_ppm_s2_new_bit_0_sel = _T_413 & (~_T_694 & ~_T_840); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_28_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_1538 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_1565 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_28_ppm_s1_new_bit_0_sel = _T_151 & (~_T_413 & ~_T_694 & ~_T_840); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_28_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_1538 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_1565 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_28_ppm_s3_new_bit_0_sel = _T_694 & ~_T_840; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_28_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_1538 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_1565 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_28_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_113 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_115 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_29_ppm_s2_new_bit_0_sel = _T_414 & (~_T_695 & ~_T_841); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_29_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_1592 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_1619 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_29_ppm_s1_new_bit_0_sel = _T_152 & (~_T_414 & ~_T_695 & ~_T_841); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_29_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_1592 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_1619 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_29_ppm_s3_new_bit_0_sel = _T_695 & ~_T_841; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_29_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_1592 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_1619 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_29_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_117 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_119 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_30_ppm_s2_new_bit_0_sel = _T_415 & (~_T_696 & ~_T_842); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_30_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_1646 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_1673 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_30_ppm_s1_new_bit_0_sel = _T_153 & (~_T_415 & ~_T_696 & ~_T_842); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_30_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_1646 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_1673 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_30_ppm_s3_new_bit_0_sel = _T_696 & ~_T_842; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_30_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_1646 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_1673 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_30_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_121 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_123 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_31_ppm_s2_new_bit_0_sel = _T_416 & (~_T_697 & ~_T_843); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_31_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_1700 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_1727 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_31_ppm_s1_new_bit_0_sel = _T_154 & (~_T_416 & ~_T_697 & ~_T_843); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_31_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_1700 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_1727 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_31_ppm_s3_new_bit_0_sel = _T_697 & ~_T_843; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_31_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_1700 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_1727 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_31_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_125 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_127 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_32_ppm_s2_new_bit_0_sel = _T_417 & (~_T_698 & ~_T_844); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_32_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_1754 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_1781 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_32_ppm_s1_new_bit_0_sel = _T_155 & (~_T_417 & ~_T_698 & ~_T_844); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_32_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_1754 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_1781 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_32_ppm_s3_new_bit_0_sel = _T_698 & ~_T_844; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_32_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_1754 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_1781 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_32_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_129 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_131 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_33_ppm_s2_new_bit_0_sel = _T_418 & (~_T_699 & ~_T_845); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_33_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_1808 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_1835 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_33_ppm_s1_new_bit_0_sel = _T_156 & (~_T_418 & ~_T_699 & ~_T_845); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_33_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_1808 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_1835 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_33_ppm_s3_new_bit_0_sel = _T_699 & ~_T_845; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_33_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_1808 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_1835 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_33_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_133 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_135 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_34_ppm_s2_new_bit_0_sel = _T_419 & (~_T_700 & ~_T_846); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_34_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_1862 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_1889 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_34_ppm_s1_new_bit_0_sel = _T_157 & (~_T_419 & ~_T_700 & ~_T_846); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_34_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_1862 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_1889 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_34_ppm_s3_new_bit_0_sel = _T_700 & ~_T_846; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_34_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_1862 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_1889 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_34_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_137 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_139 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_35_ppm_s2_new_bit_0_sel = _T_420 & (~_T_701 & ~_T_847); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_35_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_1916 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_1943 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_35_ppm_s1_new_bit_0_sel = _T_158 & (~_T_420 & ~_T_701 & ~_T_847); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_35_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_1916 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_1943 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_35_ppm_s3_new_bit_0_sel = _T_701 & ~_T_847; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_35_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_1916 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_1943 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_35_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_141 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_143 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_36_ppm_s2_new_bit_0_sel = _T_421 & (~_T_702 & ~_T_848); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_36_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_1970 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_1997 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_36_ppm_s1_new_bit_0_sel = _T_159 & (~_T_421 & ~_T_702 & ~_T_848); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_36_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_1970 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_1997 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_36_ppm_s3_new_bit_0_sel = _T_702 & ~_T_848; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_36_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_1970 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_1997 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_36_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_145 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_147 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_37_ppm_s2_new_bit_0_sel = _T_422 & (~_T_703 & ~_T_849); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_37_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_2024 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_2051 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_37_ppm_s1_new_bit_0_sel = _T_160 & (~_T_422 & ~_T_703 & ~_T_849); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_37_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_2024 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_2051 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_37_ppm_s3_new_bit_0_sel = _T_703 & ~_T_849; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_37_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_2024 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_2051 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_37_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_149 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_151 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_38_ppm_s2_new_bit_0_sel = _T_423 & (~_T_704 & ~_T_850); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_38_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_2078 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_2105 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_38_ppm_s1_new_bit_0_sel = _T_161 & (~_T_423 & ~_T_704 & ~_T_850); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_38_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_2078 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_2105 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_38_ppm_s3_new_bit_0_sel = _T_704 & ~_T_850; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_38_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_2078 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_2105 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_38_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_153 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_155 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_39_ppm_s2_new_bit_0_sel = _T_424 & (~_T_705 & ~_T_851); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_39_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_2132 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_2159 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_39_ppm_s1_new_bit_0_sel = _T_162 & (~_T_424 & ~_T_705 & ~_T_851); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_39_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_2132 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_2159 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_39_ppm_s3_new_bit_0_sel = _T_705 & ~_T_851; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_39_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_2132 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_2159 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_39_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_157 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_159 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_40_ppm_s2_new_bit_0_sel = _T_425 & (~_T_706 & ~_T_852); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_40_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_2186 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_2213 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_40_ppm_s1_new_bit_0_sel = _T_163 & (~_T_425 & ~_T_706 & ~_T_852); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_40_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_2186 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_2213 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_40_ppm_s3_new_bit_0_sel = _T_706 & ~_T_852; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_40_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_2186 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_2213 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_40_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_161 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_163 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_41_ppm_s2_new_bit_0_sel = _T_426 & (~_T_707 & ~_T_853); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_41_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_2240 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_2267 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_41_ppm_s1_new_bit_0_sel = _T_164 & (~_T_426 & ~_T_707 & ~_T_853); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_41_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_2240 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_2267 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_41_ppm_s3_new_bit_0_sel = _T_707 & ~_T_853; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_41_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_2240 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_2267 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_41_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_165 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_167 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_42_ppm_s2_new_bit_0_sel = _T_427 & (~_T_708 & ~_T_854); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_42_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_2294 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_2321 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_42_ppm_s1_new_bit_0_sel = _T_165 & (~_T_427 & ~_T_708 & ~_T_854); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_42_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_2294 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_2321 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_42_ppm_s3_new_bit_0_sel = _T_708 & ~_T_854; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_42_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_2294 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_2321 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_42_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_169 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_171 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_43_ppm_s2_new_bit_0_sel = _T_428 & (~_T_709 & ~_T_855); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_43_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_2348 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_2375 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_43_ppm_s1_new_bit_0_sel = _T_166 & (~_T_428 & ~_T_709 & ~_T_855); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_43_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_2348 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_2375 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_43_ppm_s3_new_bit_0_sel = _T_709 & ~_T_855; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_43_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_2348 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_2375 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_43_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_173 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_175 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_44_ppm_s2_new_bit_0_sel = _T_429 & (~_T_710 & ~_T_856); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_44_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_2402 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_2429 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_44_ppm_s1_new_bit_0_sel = _T_167 & (~_T_429 & ~_T_710 & ~_T_856); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_44_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_2402 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_2429 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_44_ppm_s3_new_bit_0_sel = _T_710 & ~_T_856; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_44_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_2402 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_2429 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_44_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_177 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_179 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_45_ppm_s2_new_bit_0_sel = _T_430 & (~_T_711 & ~_T_857); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_45_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_2456 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_2483 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_45_ppm_s1_new_bit_0_sel = _T_168 & (~_T_430 & ~_T_711 & ~_T_857); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_45_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_2456 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_2483 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_45_ppm_s3_new_bit_0_sel = _T_711 & ~_T_857; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_45_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_2456 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_2483 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_45_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_181 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_183 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_46_ppm_s2_new_bit_0_sel = _T_431 & (~_T_712 & ~_T_858); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_46_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_2510 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_2537 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_46_ppm_s1_new_bit_0_sel = _T_169 & (~_T_431 & ~_T_712 & ~_T_858); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_46_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_2510 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_2537 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_46_ppm_s3_new_bit_0_sel = _T_712 & ~_T_858; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_46_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_2510 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_2537 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_46_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_185 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_187 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_47_ppm_s2_new_bit_0_sel = _T_432 & (~_T_713 & ~_T_859); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_47_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_2564 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_2591 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_47_ppm_s1_new_bit_0_sel = _T_170 & (~_T_432 & ~_T_713 & ~_T_859); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_47_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_2564 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_2591 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_47_ppm_s3_new_bit_0_sel = _T_713 & ~_T_859; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_47_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_2564 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_2591 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_47_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_189 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_191 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_48_ppm_s2_new_bit_0_sel = _T_433 & (~_T_714 & ~_T_860); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_48_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_2618 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_2645 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_48_ppm_s1_new_bit_0_sel = _T_171 & (~_T_433 & ~_T_714 & ~_T_860); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_48_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_2618 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_2645 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_48_ppm_s3_new_bit_0_sel = _T_714 & ~_T_860; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_48_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_2618 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_2645 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_48_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_193 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_195 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_49_ppm_s2_new_bit_0_sel = _T_434 & (~_T_715 & ~_T_861); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_49_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_2672 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_2699 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_49_ppm_s1_new_bit_0_sel = _T_172 & (~_T_434 & ~_T_715 & ~_T_861); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_49_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_2672 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_2699 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_49_ppm_s3_new_bit_0_sel = _T_715 & ~_T_861; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_49_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_2672 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_2699 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_49_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_197 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_199 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_50_ppm_s2_new_bit_0_sel = _T_435 & (~_T_716 & ~_T_862); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_50_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_2726 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_2753 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_50_ppm_s1_new_bit_0_sel = _T_173 & (~_T_435 & ~_T_716 & ~_T_862); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_50_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_2726 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_2753 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_50_ppm_s3_new_bit_0_sel = _T_716 & ~_T_862; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_50_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_2726 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_2753 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_50_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_201 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_203 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_51_ppm_s2_new_bit_0_sel = _T_436 & (~_T_717 & ~_T_863); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_51_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_2780 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_2807 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_51_ppm_s1_new_bit_0_sel = _T_174 & (~_T_436 & ~_T_717 & ~_T_863); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_51_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_2780 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_2807 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_51_ppm_s3_new_bit_0_sel = _T_717 & ~_T_863; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_51_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_2780 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_2807 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_51_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_205 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_207 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_52_ppm_s2_new_bit_0_sel = _T_437 & (~_T_718 & ~_T_864); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_52_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_2834 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_2861 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_52_ppm_s1_new_bit_0_sel = _T_175 & (~_T_437 & ~_T_718 & ~_T_864); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_52_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_2834 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_2861 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_52_ppm_s3_new_bit_0_sel = _T_718 & ~_T_864; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_52_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_2834 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_2861 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_52_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_209 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_211 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_53_ppm_s2_new_bit_0_sel = _T_438 & (~_T_719 & ~_T_865); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_53_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_2888 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_2915 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_53_ppm_s1_new_bit_0_sel = _T_176 & (~_T_438 & ~_T_719 & ~_T_865); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_53_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_2888 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_2915 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_53_ppm_s3_new_bit_0_sel = _T_719 & ~_T_865; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_53_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_2888 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_2915 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_53_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_213 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_215 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_54_ppm_s2_new_bit_0_sel = _T_439 & (~_T_720 & ~_T_866); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_54_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_2942 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_2969 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_54_ppm_s1_new_bit_0_sel = _T_177 & (~_T_439 & ~_T_720 & ~_T_866); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_54_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_2942 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_2969 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_54_ppm_s3_new_bit_0_sel = _T_720 & ~_T_866; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_54_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_2942 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_2969 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_54_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_217 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_219 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_55_ppm_s2_new_bit_0_sel = _T_440 & (~_T_721 & ~_T_867); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_55_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_2996 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_3023 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_55_ppm_s1_new_bit_0_sel = _T_178 & (~_T_440 & ~_T_721 & ~_T_867); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_55_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_2996 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_3023 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_55_ppm_s3_new_bit_0_sel = _T_721 & ~_T_867; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_55_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_2996 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_3023 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_55_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_221 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_223 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_56_ppm_s2_new_bit_0_sel = _T_441 & (~_T_722 & ~_T_868); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_56_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_3050 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_3077 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_56_ppm_s1_new_bit_0_sel = _T_179 & (~_T_441 & ~_T_722 & ~_T_868); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_56_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_3050 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_3077 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_56_ppm_s3_new_bit_0_sel = _T_722 & ~_T_868; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_56_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_3050 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_3077 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_56_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_225 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_227 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_57_ppm_s2_new_bit_0_sel = _T_442 & (~_T_723 & ~_T_869); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_57_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_3104 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_3131 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_57_ppm_s1_new_bit_0_sel = _T_180 & (~_T_442 & ~_T_723 & ~_T_869); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_57_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_3104 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_3131 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_57_ppm_s3_new_bit_0_sel = _T_723 & ~_T_869; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_57_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_3104 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_3131 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_57_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_229 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_231 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_58_ppm_s2_new_bit_0_sel = _T_443 & (~_T_724 & ~_T_870); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_58_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_3158 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_3185 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_58_ppm_s1_new_bit_0_sel = _T_181 & (~_T_443 & ~_T_724 & ~_T_870); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_58_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_3158 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_3185 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_58_ppm_s3_new_bit_0_sel = _T_724 & ~_T_870; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_58_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_3158 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_3185 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_58_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_233 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_235 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_59_ppm_s2_new_bit_0_sel = _T_444 & (~_T_725 & ~_T_871); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_59_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_3212 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_3239 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_59_ppm_s1_new_bit_0_sel = _T_182 & (~_T_444 & ~_T_725 & ~_T_871); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_59_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_3212 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_3239 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_59_ppm_s3_new_bit_0_sel = _T_725 & ~_T_871; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_59_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_3212 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_3239 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_59_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_237 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_239 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_60_ppm_s2_new_bit_0_sel = _T_445 & (~_T_726 & ~_T_872); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_60_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_3266 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_3293 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_60_ppm_s1_new_bit_0_sel = _T_183 & (~_T_445 & ~_T_726 & ~_T_872); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_60_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_3266 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_3293 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_60_ppm_s3_new_bit_0_sel = _T_726 & ~_T_872; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_60_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_3266 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_3293 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_60_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_241 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_243 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_61_ppm_s2_new_bit_0_sel = _T_446 & (~_T_727 & ~_T_873); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_61_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_3320 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_3347 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_61_ppm_s1_new_bit_0_sel = _T_184 & (~_T_446 & ~_T_727 & ~_T_873); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_61_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_3320 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_3347 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_61_ppm_s3_new_bit_0_sel = _T_727 & ~_T_873; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_61_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_3320 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_3347 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_61_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_245 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_247 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_62_ppm_s2_new_bit_0_sel = _T_447 & (~_T_728 & ~_T_874); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_62_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_3374 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_3401 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_62_ppm_s1_new_bit_0_sel = _T_185 & (~_T_447 & ~_T_728 & ~_T_874); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_62_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_3374 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_3401 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_62_ppm_s3_new_bit_0_sel = _T_728 & ~_T_874; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_62_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_3374 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_3401 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_62_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_249 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_251 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_63_ppm_s2_new_bit_0_sel = _T_448 & (~_T_729 & ~_T_875); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_63_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_3428 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_3455 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_63_ppm_s1_new_bit_0_sel = _T_186 & (~_T_448 & ~_T_729 & ~_T_875); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_63_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_3428 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_3455 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_63_ppm_s3_new_bit_0_sel = _T_729 & ~_T_875; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_63_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_3428 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_3455 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_63_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_253 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_255 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_64_ppm_s2_new_bit_0_sel = _T_449 & (~_T_730 & ~_T_876); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_64_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_3482 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_3509 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_64_ppm_s1_new_bit_0_sel = _T_187 & (~_T_449 & ~_T_730 & ~_T_876); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_64_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_3482 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_3509 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_64_ppm_s3_new_bit_0_sel = _T_730 & ~_T_876; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_64_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_3482 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_3509 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_64_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_257 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_259 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_65_ppm_s2_new_bit_0_sel = _T_450 & (~_T_731 & ~_T_877); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_65_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_3536 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_3563 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_65_ppm_s1_new_bit_0_sel = _T_188 & (~_T_450 & ~_T_731 & ~_T_877); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_65_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_3536 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_3563 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_65_ppm_s3_new_bit_0_sel = _T_731 & ~_T_877; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_65_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_3536 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_3563 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_65_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_261 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_263 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_66_ppm_s2_new_bit_0_sel = _T_451 & (~_T_732 & ~_T_878); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_66_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_3590 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_3617 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_66_ppm_s1_new_bit_0_sel = _T_189 & (~_T_451 & ~_T_732 & ~_T_878); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_66_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_3590 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_3617 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_66_ppm_s3_new_bit_0_sel = _T_732 & ~_T_878; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_66_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_3590 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_3617 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_66_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_265 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_267 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_67_ppm_s2_new_bit_0_sel = _T_452 & (~_T_733 & ~_T_879); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_67_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_3644 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_3671 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_67_ppm_s1_new_bit_0_sel = _T_190 & (~_T_452 & ~_T_733 & ~_T_879); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_67_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_3644 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_3671 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_67_ppm_s3_new_bit_0_sel = _T_733 & ~_T_879; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_67_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_3644 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_3671 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_67_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_269 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_271 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_68_ppm_s2_new_bit_0_sel = _T_453 & (~_T_734 & ~_T_880); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_68_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_3698 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_3725 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_68_ppm_s1_new_bit_0_sel = _T_191 & (~_T_453 & ~_T_734 & ~_T_880); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_68_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_3698 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_3725 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_68_ppm_s3_new_bit_0_sel = _T_734 & ~_T_880; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_68_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_3698 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_3725 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_68_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_273 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_275 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_69_ppm_s2_new_bit_0_sel = _T_454 & (~_T_735 & ~_T_881); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_69_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_3752 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_3779 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_69_ppm_s1_new_bit_0_sel = _T_192 & (~_T_454 & ~_T_735 & ~_T_881); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_69_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_3752 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_3779 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_69_ppm_s3_new_bit_0_sel = _T_735 & ~_T_881; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_69_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_3752 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_3779 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_69_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_277 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_279 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_70_ppm_s2_new_bit_0_sel = _T_455 & (~_T_736 & ~_T_882); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_70_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_3806 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_3833 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_70_ppm_s1_new_bit_0_sel = _T_193 & (~_T_455 & ~_T_736 & ~_T_882); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_70_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_3806 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_3833 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_70_ppm_s3_new_bit_0_sel = _T_736 & ~_T_882; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_70_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_3806 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_3833 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_70_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_281 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_283 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_71_ppm_s2_new_bit_0_sel = _T_456 & (~_T_737 & ~_T_883); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_71_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_3860 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_3887 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_71_ppm_s1_new_bit_0_sel = _T_194 & (~_T_456 & ~_T_737 & ~_T_883); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_71_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_3860 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_3887 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_71_ppm_s3_new_bit_0_sel = _T_737 & ~_T_883; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_71_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_3860 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_3887 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_71_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_285 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_287 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_72_ppm_s2_new_bit_0_sel = _T_457 & (~_T_738 & ~_T_884); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_72_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_3914 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_3941 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_72_ppm_s1_new_bit_0_sel = _T_195 & (~_T_457 & ~_T_738 & ~_T_884); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_72_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_3914 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_3941 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_72_ppm_s3_new_bit_0_sel = _T_738 & ~_T_884; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_72_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_3914 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_3941 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_72_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_289 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_291 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_73_ppm_s2_new_bit_0_sel = _T_458 & (~_T_739 & ~_T_885); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_73_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_3968 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_3995 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_73_ppm_s1_new_bit_0_sel = _T_196 & (~_T_458 & ~_T_739 & ~_T_885); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_73_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_3968 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_3995 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_73_ppm_s3_new_bit_0_sel = _T_739 & ~_T_885; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_73_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_3968 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_3995 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_73_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_293 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_295 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_74_ppm_s2_new_bit_0_sel = _T_459 & (~_T_740 & ~_T_886); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_74_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_4022 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_4049 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_74_ppm_s1_new_bit_0_sel = _T_197 & (~_T_459 & ~_T_740 & ~_T_886); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_74_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_4022 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_4049 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_74_ppm_s3_new_bit_0_sel = _T_740 & ~_T_886; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_74_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_4022 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_4049 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_74_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_297 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_299 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_75_ppm_s2_new_bit_0_sel = _T_460 & (~_T_741 & ~_T_887); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_75_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_4076 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_4103 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_75_ppm_s1_new_bit_0_sel = _T_198 & (~_T_460 & ~_T_741 & ~_T_887); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_75_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_4076 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_4103 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_75_ppm_s3_new_bit_0_sel = _T_741 & ~_T_887; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_75_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_4076 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_4103 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_75_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_301 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_303 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_76_ppm_s2_new_bit_0_sel = _T_461 & (~_T_742 & ~_T_888); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_76_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_4130 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_4157 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_76_ppm_s1_new_bit_0_sel = _T_199 & (~_T_461 & ~_T_742 & ~_T_888); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_76_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_4130 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_4157 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_76_ppm_s3_new_bit_0_sel = _T_742 & ~_T_888; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_76_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_4130 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_4157 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_76_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_305 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_307 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_77_ppm_s2_new_bit_0_sel = _T_462 & (~_T_743 & ~_T_889); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_77_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_4184 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_4211 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_77_ppm_s1_new_bit_0_sel = _T_200 & (~_T_462 & ~_T_743 & ~_T_889); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_77_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_4184 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_4211 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_77_ppm_s3_new_bit_0_sel = _T_743 & ~_T_889; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_77_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_4184 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_4211 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_77_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_309 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_311 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_78_ppm_s2_new_bit_0_sel = _T_463 & (~_T_744 & ~_T_890); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_78_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_4238 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_4265 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_78_ppm_s1_new_bit_0_sel = _T_201 & (~_T_463 & ~_T_744 & ~_T_890); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_78_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_4238 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_4265 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_78_ppm_s3_new_bit_0_sel = _T_744 & ~_T_890; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_78_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_4238 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_4265 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_78_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_313 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_315 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_79_ppm_s2_new_bit_0_sel = _T_464 & (~_T_745 & ~_T_891); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_79_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_4292 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_4319 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_79_ppm_s1_new_bit_0_sel = _T_202 & (~_T_464 & ~_T_745 & ~_T_891); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_79_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_4292 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_4319 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_79_ppm_s3_new_bit_0_sel = _T_745 & ~_T_891; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_79_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_4292 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_4319 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_79_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_317 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_319 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_80_ppm_s2_new_bit_0_sel = _T_465 & (~_T_746 & ~_T_892); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_80_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_4346 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_4373 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_80_ppm_s1_new_bit_0_sel = _T_203 & (~_T_465 & ~_T_746 & ~_T_892); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_80_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_4346 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_4373 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_80_ppm_s3_new_bit_0_sel = _T_746 & ~_T_892; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_80_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_4346 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_4373 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_80_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_321 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_323 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_81_ppm_s2_new_bit_0_sel = _T_466 & (~_T_747 & ~_T_893); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_81_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_4400 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_4427 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_81_ppm_s1_new_bit_0_sel = _T_204 & (~_T_466 & ~_T_747 & ~_T_893); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_81_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_4400 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_4427 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_81_ppm_s3_new_bit_0_sel = _T_747 & ~_T_893; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_81_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_4400 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_4427 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_81_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_325 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_327 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_82_ppm_s2_new_bit_0_sel = _T_467 & (~_T_748 & ~_T_894); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_82_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_4454 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_4481 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_82_ppm_s1_new_bit_0_sel = _T_205 & (~_T_467 & ~_T_748 & ~_T_894); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_82_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_4454 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_4481 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_82_ppm_s3_new_bit_0_sel = _T_748 & ~_T_894; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_82_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_4454 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_4481 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_82_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_329 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_331 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_83_ppm_s2_new_bit_0_sel = _T_468 & (~_T_749 & ~_T_895); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_83_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_4508 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_4535 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_83_ppm_s1_new_bit_0_sel = _T_206 & (~_T_468 & ~_T_749 & ~_T_895); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_83_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_4508 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_4535 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_83_ppm_s3_new_bit_0_sel = _T_749 & ~_T_895; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_83_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_4508 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_4535 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_83_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_333 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_335 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_84_ppm_s2_new_bit_0_sel = _T_469 & (~_T_750 & ~_T_896); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_84_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_4562 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_4589 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_84_ppm_s1_new_bit_0_sel = _T_207 & (~_T_469 & ~_T_750 & ~_T_896); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_84_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_4562 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_4589 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_84_ppm_s3_new_bit_0_sel = _T_750 & ~_T_896; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_84_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_4562 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_4589 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_84_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_337 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_339 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_85_ppm_s2_new_bit_0_sel = _T_470 & (~_T_751 & ~_T_897); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_85_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_4616 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_4643 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_85_ppm_s1_new_bit_0_sel = _T_208 & (~_T_470 & ~_T_751 & ~_T_897); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_85_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_4616 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_4643 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_85_ppm_s3_new_bit_0_sel = _T_751 & ~_T_897; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_85_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_4616 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_4643 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_85_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_341 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_343 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_86_ppm_s2_new_bit_0_sel = _T_471 & (~_T_752 & ~_T_898); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_86_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_4670 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_4697 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_86_ppm_s1_new_bit_0_sel = _T_209 & (~_T_471 & ~_T_752 & ~_T_898); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_86_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_4670 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_4697 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_86_ppm_s3_new_bit_0_sel = _T_752 & ~_T_898; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_86_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_4670 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_4697 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_86_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_345 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_347 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_87_ppm_s2_new_bit_0_sel = _T_472 & (~_T_753 & ~_T_899); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_87_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_4724 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_4751 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_87_ppm_s1_new_bit_0_sel = _T_210 & (~_T_472 & ~_T_753 & ~_T_899); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_87_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_4724 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_4751 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_87_ppm_s3_new_bit_0_sel = _T_753 & ~_T_899; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_87_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_4724 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_4751 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_87_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_349 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_351 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_88_ppm_s2_new_bit_0_sel = _T_473 & (~_T_754 & ~_T_900); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_88_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_4778 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_4805 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_88_ppm_s1_new_bit_0_sel = _T_211 & (~_T_473 & ~_T_754 & ~_T_900); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_88_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_4778 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_4805 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_88_ppm_s3_new_bit_0_sel = _T_754 & ~_T_900; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_88_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_4778 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_4805 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_88_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_353 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_355 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_89_ppm_s2_new_bit_0_sel = _T_474 & (~_T_755 & ~_T_901); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_89_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_4832 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_4859 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_89_ppm_s1_new_bit_0_sel = _T_212 & (~_T_474 & ~_T_755 & ~_T_901); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_89_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_4832 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_4859 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_89_ppm_s3_new_bit_0_sel = _T_755 & ~_T_901; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_89_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_4832 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_4859 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_89_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_357 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_359 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_90_ppm_s2_new_bit_0_sel = _T_475 & (~_T_756 & ~_T_902); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_90_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_4886 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_4913 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_90_ppm_s1_new_bit_0_sel = _T_213 & (~_T_475 & ~_T_756 & ~_T_902); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_90_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_4886 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_4913 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_90_ppm_s3_new_bit_0_sel = _T_756 & ~_T_902; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_90_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_4886 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_4913 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_90_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_361 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_363 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_91_ppm_s2_new_bit_0_sel = _T_476 & (~_T_757 & ~_T_903); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_91_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_4940 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_4967 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_91_ppm_s1_new_bit_0_sel = _T_214 & (~_T_476 & ~_T_757 & ~_T_903); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_91_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_4940 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_4967 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_91_ppm_s3_new_bit_0_sel = _T_757 & ~_T_903; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_91_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_4940 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_4967 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_91_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_365 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_367 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_92_ppm_s2_new_bit_0_sel = _T_477 & (~_T_758 & ~_T_904); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_92_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_4994 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_5021 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_92_ppm_s1_new_bit_0_sel = _T_215 & (~_T_477 & ~_T_758 & ~_T_904); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_92_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_4994 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_5021 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_92_ppm_s3_new_bit_0_sel = _T_758 & ~_T_904; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_92_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_4994 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_5021 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_92_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_369 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_371 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_93_ppm_s2_new_bit_0_sel = _T_478 & (~_T_759 & ~_T_905); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_93_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_5048 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_5075 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_93_ppm_s1_new_bit_0_sel = _T_216 & (~_T_478 & ~_T_759 & ~_T_905); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_93_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_5048 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_5075 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_93_ppm_s3_new_bit_0_sel = _T_759 & ~_T_905; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_93_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_5048 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_5075 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_93_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_373 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_375 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_94_ppm_s2_new_bit_0_sel = _T_479 & (~_T_760 & ~_T_906); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_94_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_5102 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_5129 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_94_ppm_s1_new_bit_0_sel = _T_217 & (~_T_479 & ~_T_760 & ~_T_906); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_94_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_5102 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_5129 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_94_ppm_s3_new_bit_0_sel = _T_760 & ~_T_906; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_94_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_5102 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_5129 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_94_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_377 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_379 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_95_ppm_s2_new_bit_0_sel = _T_480 & (~_T_761 & ~_T_907); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_95_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_5156 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_5183 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_95_ppm_s1_new_bit_0_sel = _T_218 & (~_T_480 & ~_T_761 & ~_T_907); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_95_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_5156 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_5183 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_95_ppm_s3_new_bit_0_sel = _T_761 & ~_T_907; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_95_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_5156 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_5183 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_95_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_381 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_383 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_96_ppm_s2_new_bit_0_sel = _T_481 & (~_T_762 & ~_T_908); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_96_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_5210 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_5237 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_96_ppm_s1_new_bit_0_sel = _T_219 & (~_T_481 & ~_T_762 & ~_T_908); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_96_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_5210 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_5237 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_96_ppm_s3_new_bit_0_sel = _T_762 & ~_T_908; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_96_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_5210 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_5237 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_96_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_385 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_387 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_97_ppm_s2_new_bit_0_sel = _T_482 & (~_T_763 & ~_T_909); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_97_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_5264 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_5291 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_97_ppm_s1_new_bit_0_sel = _T_220 & (~_T_482 & ~_T_763 & ~_T_909); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_97_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_5264 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_5291 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_97_ppm_s3_new_bit_0_sel = _T_763 & ~_T_909; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_97_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_5264 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_5291 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_97_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_389 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_391 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_98_ppm_s2_new_bit_0_sel = _T_483 & (~_T_764 & ~_T_910); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_98_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_5318 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_5345 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_98_ppm_s1_new_bit_0_sel = _T_221 & (~_T_483 & ~_T_764 & ~_T_910); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_98_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_5318 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_5345 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_98_ppm_s3_new_bit_0_sel = _T_764 & ~_T_910; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_98_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_5318 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_5345 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_98_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_393 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_395 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_99_ppm_s2_new_bit_0_sel = _T_484 & (~_T_765 & ~_T_911); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_99_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_5372 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_5399 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_99_ppm_s1_new_bit_0_sel = _T_222 & (~_T_484 & ~_T_765 & ~_T_911); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_99_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_5372 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_5399 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_99_ppm_s3_new_bit_0_sel = _T_765 & ~_T_911; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_99_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_5372 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_5399 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_99_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_397 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_399 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_100_ppm_s2_new_bit_0_sel = _T_485 & (~_T_766 & ~_T_912); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_100_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_5426 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_5453 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_100_ppm_s1_new_bit_0_sel = _T_223 & (~_T_485 & ~_T_766 & ~_T_912); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_100_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_5426 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_5453 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_100_ppm_s3_new_bit_0_sel = _T_766 & ~_T_912; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_100_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_5426 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_5453 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_100_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_401 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_403 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_101_ppm_s2_new_bit_0_sel = _T_486 & (~_T_767 & ~_T_913); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_101_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_5480 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_5507 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_101_ppm_s1_new_bit_0_sel = _T_224 & (~_T_486 & ~_T_767 & ~_T_913); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_101_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_5480 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_5507 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_101_ppm_s3_new_bit_0_sel = _T_767 & ~_T_913; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_101_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_5480 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_5507 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_101_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_405 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_407 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_102_ppm_s2_new_bit_0_sel = _T_487 & (~_T_768 & ~_T_914); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_102_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_5534 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_5561 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_102_ppm_s1_new_bit_0_sel = _T_225 & (~_T_487 & ~_T_768 & ~_T_914); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_102_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_5534 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_5561 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_102_ppm_s3_new_bit_0_sel = _T_768 & ~_T_914; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_102_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_5534 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_5561 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_102_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_409 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_411 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_103_ppm_s2_new_bit_0_sel = _T_488 & (~_T_769 & ~_T_915); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_103_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_5588 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_5615 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_103_ppm_s1_new_bit_0_sel = _T_226 & (~_T_488 & ~_T_769 & ~_T_915); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_103_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_5588 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_5615 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_103_ppm_s3_new_bit_0_sel = _T_769 & ~_T_915; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_103_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_5588 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_5615 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_103_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_413 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_415 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_104_ppm_s2_new_bit_0_sel = _T_489 & (~_T_770 & ~_T_916); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_104_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_5642 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_5669 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_104_ppm_s1_new_bit_0_sel = _T_227 & (~_T_489 & ~_T_770 & ~_T_916); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_104_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_5642 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_5669 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_104_ppm_s3_new_bit_0_sel = _T_770 & ~_T_916; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_104_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_5642 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_5669 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_104_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_417 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_419 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_105_ppm_s2_new_bit_0_sel = _T_490 & (~_T_771 & ~_T_917); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_105_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_5696 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_5723 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_105_ppm_s1_new_bit_0_sel = _T_228 & (~_T_490 & ~_T_771 & ~_T_917); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_105_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_5696 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_5723 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_105_ppm_s3_new_bit_0_sel = _T_771 & ~_T_917; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_105_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_5696 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_5723 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_105_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_421 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_423 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_106_ppm_s2_new_bit_0_sel = _T_491 & (~_T_772 & ~_T_918); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_106_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_5750 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_5777 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_106_ppm_s1_new_bit_0_sel = _T_229 & (~_T_491 & ~_T_772 & ~_T_918); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_106_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_5750 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_5777 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_106_ppm_s3_new_bit_0_sel = _T_772 & ~_T_918; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_106_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_5750 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_5777 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_106_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_425 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_427 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_107_ppm_s2_new_bit_0_sel = _T_492 & (~_T_773 & ~_T_919); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_107_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_5804 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_5831 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_107_ppm_s1_new_bit_0_sel = _T_230 & (~_T_492 & ~_T_773 & ~_T_919); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_107_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_5804 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_5831 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_107_ppm_s3_new_bit_0_sel = _T_773 & ~_T_919; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_107_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_5804 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_5831 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_107_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_429 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_431 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_108_ppm_s2_new_bit_0_sel = _T_493 & (~_T_774 & ~_T_920); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_108_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_5858 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_5885 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_108_ppm_s1_new_bit_0_sel = _T_231 & (~_T_493 & ~_T_774 & ~_T_920); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_108_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_5858 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_5885 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_108_ppm_s3_new_bit_0_sel = _T_774 & ~_T_920; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_108_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_5858 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_5885 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_108_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_433 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_435 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_109_ppm_s2_new_bit_0_sel = _T_494 & (~_T_775 & ~_T_921); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_109_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_5912 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_5939 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_109_ppm_s1_new_bit_0_sel = _T_232 & (~_T_494 & ~_T_775 & ~_T_921); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_109_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_5912 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_5939 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_109_ppm_s3_new_bit_0_sel = _T_775 & ~_T_921; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_109_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_5912 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_5939 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_109_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_437 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_439 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_110_ppm_s2_new_bit_0_sel = _T_495 & (~_T_776 & ~_T_922); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_110_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_5966 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_5993 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_110_ppm_s1_new_bit_0_sel = _T_233 & (~_T_495 & ~_T_776 & ~_T_922); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_110_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_5966 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_5993 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_110_ppm_s3_new_bit_0_sel = _T_776 & ~_T_922; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_110_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_5966 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_5993 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_110_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_441 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_443 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_111_ppm_s2_new_bit_0_sel = _T_496 & (~_T_777 & ~_T_923); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_111_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_6020 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_6047 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_111_ppm_s1_new_bit_0_sel = _T_234 & (~_T_496 & ~_T_777 & ~_T_923); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_111_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_6020 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_6047 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_111_ppm_s3_new_bit_0_sel = _T_777 & ~_T_923; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_111_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_6020 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_6047 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_111_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_445 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_447 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_112_ppm_s2_new_bit_0_sel = _T_497 & (~_T_778 & ~_T_924); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_112_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_6074 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_6101 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_112_ppm_s1_new_bit_0_sel = _T_235 & (~_T_497 & ~_T_778 & ~_T_924); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_112_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_6074 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_6101 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_112_ppm_s3_new_bit_0_sel = _T_778 & ~_T_924; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_112_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_6074 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_6101 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_112_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_449 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_451 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_113_ppm_s2_new_bit_0_sel = _T_498 & (~_T_779 & ~_T_925); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_113_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_6128 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_6155 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_113_ppm_s1_new_bit_0_sel = _T_236 & (~_T_498 & ~_T_779 & ~_T_925); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_113_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_6128 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_6155 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_113_ppm_s3_new_bit_0_sel = _T_779 & ~_T_925; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_113_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_6128 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_6155 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_113_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_453 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_455 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_114_ppm_s2_new_bit_0_sel = _T_499 & (~_T_780 & ~_T_926); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_114_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_6182 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_6209 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_114_ppm_s1_new_bit_0_sel = _T_237 & (~_T_499 & ~_T_780 & ~_T_926); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_114_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_6182 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_6209 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_114_ppm_s3_new_bit_0_sel = _T_780 & ~_T_926; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_114_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_6182 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_6209 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_114_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_457 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_459 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_115_ppm_s2_new_bit_0_sel = _T_500 & (~_T_781 & ~_T_927); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_115_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_6236 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_6263 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_115_ppm_s1_new_bit_0_sel = _T_238 & (~_T_500 & ~_T_781 & ~_T_927); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_115_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_6236 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_6263 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_115_ppm_s3_new_bit_0_sel = _T_781 & ~_T_927; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_115_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_6236 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_6263 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_115_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_461 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_463 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_116_ppm_s2_new_bit_0_sel = _T_501 & (~_T_782 & ~_T_928); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_116_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_6290 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_6317 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_116_ppm_s1_new_bit_0_sel = _T_239 & (~_T_501 & ~_T_782 & ~_T_928); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_116_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_6290 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_6317 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_116_ppm_s3_new_bit_0_sel = _T_782 & ~_T_928; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_116_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_6290 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_6317 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_116_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_465 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_467 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_117_ppm_s2_new_bit_0_sel = _T_502 & (~_T_783 & ~_T_929); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_117_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_6344 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_6371 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_117_ppm_s1_new_bit_0_sel = _T_240 & (~_T_502 & ~_T_783 & ~_T_929); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_117_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_6344 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_6371 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_117_ppm_s3_new_bit_0_sel = _T_783 & ~_T_929; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_117_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_6344 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_6371 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_117_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_469 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_471 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_118_ppm_s2_new_bit_0_sel = _T_503 & (~_T_784 & ~_T_930); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_118_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_6398 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_6425 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_118_ppm_s1_new_bit_0_sel = _T_241 & (~_T_503 & ~_T_784 & ~_T_930); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_118_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_6398 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_6425 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_118_ppm_s3_new_bit_0_sel = _T_784 & ~_T_930; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_118_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_6398 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_6425 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_118_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_473 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_475 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_119_ppm_s2_new_bit_0_sel = _T_504 & (~_T_785 & ~_T_931); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_119_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_6452 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_6479 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_119_ppm_s1_new_bit_0_sel = _T_242 & (~_T_504 & ~_T_785 & ~_T_931); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_119_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_6452 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_6479 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_119_ppm_s3_new_bit_0_sel = _T_785 & ~_T_931; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_119_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_6452 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_6479 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_119_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_477 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_479 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_120_ppm_s2_new_bit_0_sel = _T_505 & (~_T_786 & ~_T_932); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_120_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_6506 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_6533 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_120_ppm_s1_new_bit_0_sel = _T_243 & (~_T_505 & ~_T_786 & ~_T_932); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_120_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_6506 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_6533 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_120_ppm_s3_new_bit_0_sel = _T_786 & ~_T_932; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_120_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_6506 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_6533 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_120_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_481 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_483 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_121_ppm_s2_new_bit_0_sel = _T_506 & (~_T_787 & ~_T_933); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_121_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_6560 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_6587 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_121_ppm_s1_new_bit_0_sel = _T_244 & (~_T_506 & ~_T_787 & ~_T_933); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_121_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_6560 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_6587 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_121_ppm_s3_new_bit_0_sel = _T_787 & ~_T_933; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_121_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_6560 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_6587 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_121_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_485 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_487 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_122_ppm_s2_new_bit_0_sel = _T_507 & (~_T_788 & ~_T_934); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_122_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_6614 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_6641 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_122_ppm_s1_new_bit_0_sel = _T_245 & (~_T_507 & ~_T_788 & ~_T_934); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_122_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_6614 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_6641 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_122_ppm_s3_new_bit_0_sel = _T_788 & ~_T_934; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_122_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_6614 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_6641 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_122_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_489 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_491 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_123_ppm_s2_new_bit_0_sel = _T_508 & (~_T_789 & ~_T_935); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_123_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_6668 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_6695 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_123_ppm_s1_new_bit_0_sel = _T_246 & (~_T_508 & ~_T_789 & ~_T_935); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_123_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_6668 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_6695 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_123_ppm_s3_new_bit_0_sel = _T_789 & ~_T_935; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_123_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_6668 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_6695 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_123_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_493 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_495 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_124_ppm_s2_new_bit_0_sel = _T_509 & (~_T_790 & ~_T_936); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_124_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_6722 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_6749 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_124_ppm_s1_new_bit_0_sel = _T_247 & (~_T_509 & ~_T_790 & ~_T_936); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_124_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_6722 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_6749 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_124_ppm_s3_new_bit_0_sel = _T_790 & ~_T_936; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_124_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_6722 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_6749 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_124_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_497 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_499 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_125_ppm_s2_new_bit_0_sel = _T_510 & (~_T_791 & ~_T_937); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_125_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_6776 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_6803 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_125_ppm_s1_new_bit_0_sel = _T_248 & (~_T_510 & ~_T_791 & ~_T_937); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_125_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_6776 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_6803 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_125_ppm_s3_new_bit_0_sel = _T_791 & ~_T_937; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_125_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_6776 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_6803 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_125_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_501 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_503 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_126_ppm_s2_new_bit_0_sel = _T_511 & (~_T_792 & ~_T_938); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_126_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_6830 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_6857 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_126_ppm_s1_new_bit_0_sel = _T_249 & (~_T_511 & ~_T_792 & ~_T_938); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_126_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_6830 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_6857 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_126_ppm_s3_new_bit_0_sel = _T_792 & ~_T_938; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_126_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_6830 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_6857 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_126_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_505 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_507 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_127_ppm_s2_new_bit_0_sel = _T_512 & (~_T_793 & ~_T_939); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_127_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_6884 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_6911 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_127_ppm_s1_new_bit_0_sel = _T_250 & (~_T_512 & ~_T_793 & ~_T_939); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_127_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_6884 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_6911 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_127_ppm_s3_new_bit_0_sel = _T_793 & ~_T_939; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_127_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_6884 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_6911 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_127_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_509 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_511 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_128_ppm_s2_new_bit_0_sel = _T_513 & (~_T_794 & ~_T_940); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_128_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_6938 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_6965 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_128_ppm_s1_new_bit_0_sel = _T_251 & (~_T_513 & ~_T_794 & ~_T_940); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_128_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_6938 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_6965 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_128_ppm_s3_new_bit_0_sel = _T_794 & ~_T_940; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_128_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_6938 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_6965 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_128_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_513 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_515 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_129_ppm_s2_new_bit_0_sel = _T_514 & (~_T_795 & ~_T_941); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_129_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_6992 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_7019 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_129_ppm_s1_new_bit_0_sel = _T_252 & (~_T_514 & ~_T_795 & ~_T_941); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_129_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_6992 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_7019 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_129_ppm_s3_new_bit_0_sel = _T_795 & ~_T_941; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_129_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_6992 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_7019 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_129_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_517 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_519 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_130_ppm_s2_new_bit_0_sel = _T_515 & (~_T_796 & ~_T_942); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_130_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_7046 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_7073 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_130_ppm_s1_new_bit_0_sel = _T_253 & (~_T_515 & ~_T_796 & ~_T_942); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_130_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_7046 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_7073 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_130_ppm_s3_new_bit_0_sel = _T_796 & ~_T_942; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_130_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_7046 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_7073 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_130_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_521 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_523 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_131_ppm_s2_new_bit_0_sel = _T_516 & (~_T_797 & ~_T_943); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_131_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_7100 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_7127 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_131_ppm_s1_new_bit_0_sel = _T_254 & (~_T_516 & ~_T_797 & ~_T_943); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_131_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_7100 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_7127 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_131_ppm_s3_new_bit_0_sel = _T_797 & ~_T_943; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_131_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_7100 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_7127 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_131_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_525 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_527 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_132_ppm_s2_new_bit_0_sel = _T_517 & (~_T_798 & ~_T_944); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_132_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_7154 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_7181 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_132_ppm_s1_new_bit_0_sel = _T_255 & (~_T_517 & ~_T_798 & ~_T_944); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_132_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_7154 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_7181 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_132_ppm_s3_new_bit_0_sel = _T_798 & ~_T_944; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_132_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_7154 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_7181 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_132_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_529 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_531 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_133_ppm_s2_new_bit_0_sel = _T_518 & (~_T_799 & ~_T_945); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_133_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_7208 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_7235 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_133_ppm_s1_new_bit_0_sel = _T_256 & (~_T_518 & ~_T_799 & ~_T_945); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_133_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_7208 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_7235 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_133_ppm_s3_new_bit_0_sel = _T_799 & ~_T_945; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_133_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_7208 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_7235 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_133_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_533 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_535 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_134_ppm_s2_new_bit_0_sel = _T_519 & (~_T_800 & ~_T_946); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_134_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_7262 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_7289 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_134_ppm_s1_new_bit_0_sel = _T_257 & (~_T_519 & ~_T_800 & ~_T_946); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_134_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_7262 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_7289 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_134_ppm_s3_new_bit_0_sel = _T_800 & ~_T_946; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_134_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_7262 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_7289 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_134_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_537 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_539 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_135_ppm_s2_new_bit_0_sel = _T_520 & (~_T_801 & ~_T_947); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_135_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_7316 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_7343 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_135_ppm_s1_new_bit_0_sel = _T_258 & (~_T_520 & ~_T_801 & ~_T_947); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_135_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_7316 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_7343 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_135_ppm_s3_new_bit_0_sel = _T_801 & ~_T_947; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_135_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_7316 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_7343 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_135_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_541 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_543 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_136_ppm_s2_new_bit_0_sel = _T_521 & (~_T_802 & ~_T_948); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_136_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_7370 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_7397 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_136_ppm_s1_new_bit_0_sel = _T_259 & (~_T_521 & ~_T_802 & ~_T_948); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_136_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_7370 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_7397 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_136_ppm_s3_new_bit_0_sel = _T_802 & ~_T_948; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_136_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_7370 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_7397 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_136_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_545 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_547 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_137_ppm_s2_new_bit_0_sel = _T_522 & (~_T_803 & ~_T_949); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_137_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_7424 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_7451 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_137_ppm_s1_new_bit_0_sel = _T_260 & (~_T_522 & ~_T_803 & ~_T_949); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_137_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_7424 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_7451 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_137_ppm_s3_new_bit_0_sel = _T_803 & ~_T_949; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_137_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_7424 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_7451 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_137_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_549 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_551 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_138_ppm_s2_new_bit_0_sel = _T_523 & (~_T_804 & ~_T_950); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_138_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_7478 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_7505 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_138_ppm_s1_new_bit_0_sel = _T_261 & (~_T_523 & ~_T_804 & ~_T_950); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_138_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_7478 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_7505 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_138_ppm_s3_new_bit_0_sel = _T_804 & ~_T_950; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_138_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_7478 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_7505 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_138_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_553 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_555 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_139_ppm_s2_new_bit_0_sel = _T_524 & (~_T_805 & ~_T_951); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_139_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_7532 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_7559 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_139_ppm_s1_new_bit_0_sel = _T_262 & (~_T_524 & ~_T_805 & ~_T_951); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_139_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_7532 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_7559 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_139_ppm_s3_new_bit_0_sel = _T_805 & ~_T_951; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_139_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_7532 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_7559 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_139_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_557 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_559 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_140_ppm_s2_new_bit_0_sel = _T_525 & (~_T_806 & ~_T_952); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_140_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_7586 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_7613 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_140_ppm_s1_new_bit_0_sel = _T_263 & (~_T_525 & ~_T_806 & ~_T_952); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_140_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_7586 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_7613 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_140_ppm_s3_new_bit_0_sel = _T_806 & ~_T_952; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_140_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_7586 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_7613 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_140_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_561 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_563 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_141_ppm_s2_new_bit_0_sel = _T_526 & (~_T_807 & ~_T_953); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_141_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_7640 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_7667 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_141_ppm_s1_new_bit_0_sel = _T_264 & (~_T_526 & ~_T_807 & ~_T_953); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_141_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_7640 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_7667 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_141_ppm_s3_new_bit_0_sel = _T_807 & ~_T_953; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_141_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_7640 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_7667 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_141_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_565 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_567 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_142_ppm_s2_new_bit_0_sel = _T_527 & (~_T_808 & ~_T_954); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_142_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_7694 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_7721 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_142_ppm_s1_new_bit_0_sel = _T_265 & (~_T_527 & ~_T_808 & ~_T_954); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_142_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_7694 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_7721 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_142_ppm_s3_new_bit_0_sel = _T_808 & ~_T_954; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_142_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_7694 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_7721 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_142_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_569 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_571 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  assign ghv_write_datas_143_ppm_s2_new_bit_0_sel = _T_528 & (~_T_809 & ~_T_955); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_143_ppm_s2_new_bit_0_src = _s2_ghv_wens_T_7748 & s2_redirect_s1_last_pred_vec_selVecOH_0 |
    _s2_ghv_wens_T_7775 & _s2_redirect_s1_last_pred_vec_T_63; // @[Mux.scala 27:73]
  assign ghv_write_datas_143_ppm_s1_new_bit_0_sel = _T_266 & (~_T_528 & ~_T_809 & ~_T_955); // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_143_ppm_s1_new_bit_0_src = _s1_ghv_wens_T_7748 & _s1_possible_predicted_fhs_T_135 |
    _s1_ghv_wens_T_7775 & _s1_possible_predicted_fhs_T_203; // @[Mux.scala 27:73]
  assign ghv_write_datas_143_ppm_s3_new_bit_0_sel = _T_809 & ~_T_955; // @[PriorityMuxGen.scala 121:41]
  assign ghv_write_datas_143_ppm_s3_new_bit_0_src = _s3_ghv_wens_T_7748 & _s3_redirect_on_br_taken_T_5 |
    _s3_ghv_wens_T_7775 & _s3_redirect_on_br_taken_T_9; // @[Mux.scala 27:73]
  assign ghv_write_datas_143_ppm_redirect_new_bit_0_src = _redirect_ghv_wens_T_573 & real_br_taken_mask_0 |
    _redirect_ghv_wens_T_575 & real_br_taken_mask_1; // @[Mux.scala 27:73]
  always @(posedge clock) begin
    if (REG_1) begin // @[BPU.scala 259:58]
      s0_pc_reg <= {{3'd0}, reset_vector_delay_io_out}; // @[BPU.scala 260:15]
    end else begin
      s0_pc_reg <= s0_pc; // @[BPU.scala 258:26]
    end
    REG <= reset; // @[BPU.scala 259:31]
    REG_1 <= REG & ~reset; // @[BPU.scala 259:39]
    if (s1_fire) begin // @[Reg.scala 17:18]
      s2_ftq_idx_flag <= io_ftq_to_bpu_enq_ptr_flag; // @[Reg.scala 17:22]
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      s2_ftq_idx_value <= io_ftq_to_bpu_enq_ptr_value; // @[Reg.scala 17:22]
    end
    if (s2_valid) begin // @[Reg.scala 17:18]
      s3_ftq_idx_flag <= s2_ftq_idx_flag; // @[Reg.scala 17:22]
    end
    if (s2_valid) begin // @[Reg.scala 17:18]
      s3_ftq_idx_value <= s2_ftq_idx_value; // @[Reg.scala 17:22]
    end
    predictors_io_update_REG_valid <= io_ftq_to_bpu_update_valid; // @[BPU.scala 601:34]
    predictors_io_update_REG_bits_pc <= io_ftq_to_bpu_update_bits_pc; // @[BPU.scala 601:34]
    predictors_io_update_REG_bits_spec_info_folded_hist_hist_17_folded_hist <=
      io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_17_folded_hist; // @[BPU.scala 601:34]
    predictors_io_update_REG_bits_spec_info_folded_hist_hist_16_folded_hist <=
      io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_16_folded_hist; // @[BPU.scala 601:34]
    predictors_io_update_REG_bits_spec_info_folded_hist_hist_15_folded_hist <=
      io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_15_folded_hist; // @[BPU.scala 601:34]
    predictors_io_update_REG_bits_spec_info_folded_hist_hist_14_folded_hist <=
      io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_14_folded_hist; // @[BPU.scala 601:34]
    predictors_io_update_REG_bits_spec_info_folded_hist_hist_13_folded_hist <=
      io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_13_folded_hist; // @[BPU.scala 601:34]
    predictors_io_update_REG_bits_spec_info_folded_hist_hist_12_folded_hist <=
      io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_12_folded_hist; // @[BPU.scala 601:34]
    predictors_io_update_REG_bits_spec_info_folded_hist_hist_10_folded_hist <=
      io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_10_folded_hist; // @[BPU.scala 601:34]
    predictors_io_update_REG_bits_spec_info_folded_hist_hist_9_folded_hist <=
      io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_9_folded_hist; // @[BPU.scala 601:34]
    predictors_io_update_REG_bits_spec_info_folded_hist_hist_8_folded_hist <=
      io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_8_folded_hist; // @[BPU.scala 601:34]
    predictors_io_update_REG_bits_spec_info_folded_hist_hist_7_folded_hist <=
      io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_7_folded_hist; // @[BPU.scala 601:34]
    predictors_io_update_REG_bits_spec_info_folded_hist_hist_6_folded_hist <=
      io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_6_folded_hist; // @[BPU.scala 601:34]
    predictors_io_update_REG_bits_spec_info_folded_hist_hist_5_folded_hist <=
      io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_5_folded_hist; // @[BPU.scala 601:34]
    predictors_io_update_REG_bits_spec_info_folded_hist_hist_4_folded_hist <=
      io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_4_folded_hist; // @[BPU.scala 601:34]
    predictors_io_update_REG_bits_spec_info_folded_hist_hist_3_folded_hist <=
      io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_3_folded_hist; // @[BPU.scala 601:34]
    predictors_io_update_REG_bits_spec_info_folded_hist_hist_2_folded_hist <=
      io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_2_folded_hist; // @[BPU.scala 601:34]
    predictors_io_update_REG_bits_spec_info_folded_hist_hist_1_folded_hist <=
      io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_1_folded_hist; // @[BPU.scala 601:34]
    predictors_io_update_REG_bits_spec_info_folded_hist_hist_0_folded_hist <=
      io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_0_folded_hist; // @[BPU.scala 601:34]
    predictors_io_update_REG_bits_ftb_entry_valid <= io_ftq_to_bpu_update_bits_ftb_entry_valid; // @[BPU.scala 601:34]
    predictors_io_update_REG_bits_ftb_entry_brSlots_0_offset <= io_ftq_to_bpu_update_bits_ftb_entry_brSlots_0_offset; // @[BPU.scala 601:34]
    predictors_io_update_REG_bits_ftb_entry_brSlots_0_lower <= io_ftq_to_bpu_update_bits_ftb_entry_brSlots_0_lower; // @[BPU.scala 601:34]
    predictors_io_update_REG_bits_ftb_entry_brSlots_0_tarStat <= io_ftq_to_bpu_update_bits_ftb_entry_brSlots_0_tarStat; // @[BPU.scala 601:34]
    predictors_io_update_REG_bits_ftb_entry_brSlots_0_sharing <= io_ftq_to_bpu_update_bits_ftb_entry_brSlots_0_sharing; // @[BPU.scala 601:34]
    predictors_io_update_REG_bits_ftb_entry_brSlots_0_valid <= io_ftq_to_bpu_update_bits_ftb_entry_brSlots_0_valid; // @[BPU.scala 601:34]
    predictors_io_update_REG_bits_ftb_entry_tailSlot_offset <= io_ftq_to_bpu_update_bits_ftb_entry_tailSlot_offset; // @[BPU.scala 601:34]
    predictors_io_update_REG_bits_ftb_entry_tailSlot_lower <= io_ftq_to_bpu_update_bits_ftb_entry_tailSlot_lower; // @[BPU.scala 601:34]
    predictors_io_update_REG_bits_ftb_entry_tailSlot_tarStat <= io_ftq_to_bpu_update_bits_ftb_entry_tailSlot_tarStat; // @[BPU.scala 601:34]
    predictors_io_update_REG_bits_ftb_entry_tailSlot_sharing <= io_ftq_to_bpu_update_bits_ftb_entry_tailSlot_sharing; // @[BPU.scala 601:34]
    predictors_io_update_REG_bits_ftb_entry_tailSlot_valid <= io_ftq_to_bpu_update_bits_ftb_entry_tailSlot_valid; // @[BPU.scala 601:34]
    predictors_io_update_REG_bits_ftb_entry_pftAddr <= io_ftq_to_bpu_update_bits_ftb_entry_pftAddr; // @[BPU.scala 601:34]
    predictors_io_update_REG_bits_ftb_entry_carry <= io_ftq_to_bpu_update_bits_ftb_entry_carry; // @[BPU.scala 601:34]
    predictors_io_update_REG_bits_ftb_entry_isCall <= io_ftq_to_bpu_update_bits_ftb_entry_isCall; // @[BPU.scala 601:34]
    predictors_io_update_REG_bits_ftb_entry_isRet <= io_ftq_to_bpu_update_bits_ftb_entry_isRet; // @[BPU.scala 601:34]
    predictors_io_update_REG_bits_ftb_entry_isJalr <= io_ftq_to_bpu_update_bits_ftb_entry_isJalr; // @[BPU.scala 601:34]
    predictors_io_update_REG_bits_ftb_entry_last_may_be_rvi_call <=
      io_ftq_to_bpu_update_bits_ftb_entry_last_may_be_rvi_call; // @[BPU.scala 601:34]
    predictors_io_update_REG_bits_ftb_entry_always_taken_0 <= io_ftq_to_bpu_update_bits_ftb_entry_always_taken_0; // @[BPU.scala 601:34]
    predictors_io_update_REG_bits_ftb_entry_always_taken_1 <= io_ftq_to_bpu_update_bits_ftb_entry_always_taken_1; // @[BPU.scala 601:34]
    predictors_io_update_REG_bits_br_taken_mask_0 <= io_ftq_to_bpu_update_bits_br_taken_mask_0; // @[BPU.scala 601:34]
    predictors_io_update_REG_bits_br_taken_mask_1 <= io_ftq_to_bpu_update_bits_br_taken_mask_1; // @[BPU.scala 601:34]
    predictors_io_update_REG_bits_jmp_taken <= io_ftq_to_bpu_update_bits_jmp_taken; // @[BPU.scala 601:34]
    predictors_io_update_REG_bits_mispred_mask_0 <= io_ftq_to_bpu_update_bits_mispred_mask_0; // @[BPU.scala 601:34]
    predictors_io_update_REG_bits_mispred_mask_1 <= io_ftq_to_bpu_update_bits_mispred_mask_1; // @[BPU.scala 601:34]
    predictors_io_update_REG_bits_mispred_mask_2 <= io_ftq_to_bpu_update_bits_mispred_mask_2; // @[BPU.scala 601:34]
    predictors_io_update_REG_bits_old_entry <= io_ftq_to_bpu_update_bits_old_entry; // @[BPU.scala 601:34]
    predictors_io_update_REG_bits_meta <= io_ftq_to_bpu_update_bits_meta; // @[BPU.scala 601:34]
    predictors_io_update_REG_bits_full_target <= io_ftq_to_bpu_update_bits_full_target; // @[BPU.scala 601:34]
    io_perf_0_value_REG <= predictors_io_perf_0_value; // @[PerfCounterUtils.scala 188:35]
    io_perf_0_value_REG_1 <= io_perf_0_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_1_value_REG <= predictors_io_perf_1_value; // @[PerfCounterUtils.scala 188:35]
    io_perf_1_value_REG_1 <= io_perf_1_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_2_value_REG <= predictors_io_perf_2_value; // @[PerfCounterUtils.scala 188:35]
    io_perf_2_value_REG_1 <= io_perf_2_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_3_value_REG <= predictors_io_perf_3_value; // @[PerfCounterUtils.scala 188:35]
    io_perf_3_value_REG_1 <= io_perf_3_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_4_value_REG <= predictors_io_perf_4_value; // @[PerfCounterUtils.scala 188:35]
    io_perf_4_value_REG_1 <= io_perf_4_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_5_value_REG <= predictors_io_perf_5_value; // @[PerfCounterUtils.scala 188:35]
    io_perf_5_value_REG_1 <= io_perf_5_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_6_value_REG <= predictors_io_perf_6_value; // @[PerfCounterUtils.scala 188:35]
    io_perf_6_value_REG_1 <= io_perf_6_value_REG; // @[PerfCounterUtils.scala 188:27]
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 355:29]
      s1_valid <= 1'h0; // @[BPU.scala 355:40]
    end else if (io_ftq_to_bpu_redirect_valid) begin
      s1_valid <= 1'h0;
    end else begin
      s1_valid <= _GEN_141;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 364:24]
      s2_valid <= 1'h0; // @[BPU.scala 364:35]
    end else if (s2_flush) begin // @[BPU.scala 365:24]
      s2_valid <= 1'h0; // @[BPU.scala 365:35]
    end else if (s1_fire) begin // @[BPU.scala 366:24]
      s2_valid <= ~s1_flush; // @[BPU.scala 366:35]
    end else if (s2_valid) begin // @[BPU.scala 252:45]
      s2_valid <= 1'h0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 373:24]
      s3_valid <= 1'h0; // @[BPU.scala 373:35]
    end else if (io_ftq_to_bpu_redirect_valid) begin // @[BPU.scala 374:24]
      s3_valid <= 1'h0; // @[BPU.scala 374:35]
    end else if (s2_valid) begin // @[BPU.scala 375:24]
      s3_valid <= ~s2_flush; // @[BPU.scala 375:35]
    end else if (s3_valid) begin // @[BPU.scala 252:45]
      s3_valid <= 1'h0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 266:26 668:17]
      s0_folded_gh_reg_hist_17_folded_hist <= 8'h0;
    end else begin
      s0_folded_gh_reg_hist_17_folded_hist <= s0_folded_gh_ppm_out_res_hist_17_folded_hist;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 266:26 668:17]
      s0_folded_gh_reg_hist_16_folded_hist <= 8'h0;
    end else begin
      s0_folded_gh_reg_hist_16_folded_hist <= s0_folded_gh_ppm_out_res_hist_16_folded_hist;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 266:26 668:17]
      s0_folded_gh_reg_hist_15_folded_hist <= 11'h0;
    end else begin
      s0_folded_gh_reg_hist_15_folded_hist <= s0_folded_gh_ppm_out_res_hist_15_folded_hist;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 266:26 668:17]
      s0_folded_gh_reg_hist_14_folded_hist <= 7'h0;
    end else begin
      s0_folded_gh_reg_hist_14_folded_hist <= s0_folded_gh_ppm_out_res_hist_14_folded_hist;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 266:26 668:17]
      s0_folded_gh_reg_hist_13_folded_hist <= 7'h0;
    end else begin
      s0_folded_gh_reg_hist_13_folded_hist <= s0_folded_gh_ppm_out_res_hist_13_folded_hist;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 266:26 668:17]
      s0_folded_gh_reg_hist_12_folded_hist <= 7'h0;
    end else begin
      s0_folded_gh_reg_hist_12_folded_hist <= s0_folded_gh_ppm_out_res_hist_12_folded_hist;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 266:26 668:17]
      s0_folded_gh_reg_hist_11_folded_hist <= 8'h0;
    end else begin
      s0_folded_gh_reg_hist_11_folded_hist <= s0_folded_gh_ppm_out_res_hist_11_folded_hist;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 266:26 668:17]
      s0_folded_gh_reg_hist_10_folded_hist <= 9'h0;
    end else begin
      s0_folded_gh_reg_hist_10_folded_hist <= s0_folded_gh_ppm_out_res_hist_10_folded_hist;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 266:26 668:17]
      s0_folded_gh_reg_hist_9_folded_hist <= 7'h0;
    end else begin
      s0_folded_gh_reg_hist_9_folded_hist <= s0_folded_gh_ppm_out_res_hist_9_folded_hist;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 266:26 668:17]
      s0_folded_gh_reg_hist_8_folded_hist <= 8'h0;
    end else begin
      s0_folded_gh_reg_hist_8_folded_hist <= s0_folded_gh_ppm_out_res_hist_8_folded_hist;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 266:26 668:17]
      s0_folded_gh_reg_hist_7_folded_hist <= 9'h0;
    end else begin
      s0_folded_gh_reg_hist_7_folded_hist <= s0_folded_gh_ppm_out_res_hist_7_folded_hist;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 266:26 668:17]
      s0_folded_gh_reg_hist_6_folded_hist <= 9'h0;
    end else begin
      s0_folded_gh_reg_hist_6_folded_hist <= s0_folded_gh_ppm_out_res_hist_6_folded_hist;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 266:26 668:17]
      s0_folded_gh_reg_hist_5_folded_hist <= 11'h0;
    end else begin
      s0_folded_gh_reg_hist_5_folded_hist <= s0_folded_gh_ppm_out_res_hist_5_folded_hist;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 266:26 668:17]
      s0_folded_gh_reg_hist_4_folded_hist <= 4'h0;
    end else begin
      s0_folded_gh_reg_hist_4_folded_hist <= s0_folded_gh_ppm_out_res_hist_4_folded_hist;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 266:26 668:17]
      s0_folded_gh_reg_hist_3_folded_hist <= 11'h0;
    end else begin
      s0_folded_gh_reg_hist_3_folded_hist <= s0_folded_gh_ppm_out_res_hist_3_folded_hist;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 266:26 668:17]
      s0_folded_gh_reg_hist_2_folded_hist <= 8'h0;
    end else begin
      s0_folded_gh_reg_hist_2_folded_hist <= s0_folded_gh_ppm_out_res_hist_2_folded_hist;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 266:26 668:17]
      s0_folded_gh_reg_hist_1_folded_hist <= 8'h0;
    end else begin
      s0_folded_gh_reg_hist_1_folded_hist <= s0_folded_gh_ppm_out_res_hist_1_folded_hist;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 266:26 668:17]
      s0_folded_gh_reg_hist_0_folded_hist <= 8'h0;
    end else begin
      s0_folded_gh_reg_hist_0_folded_hist <= s0_folded_gh_ppm_out_res_hist_0_folded_hist;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s1_folded_gh_hist_17_folded_hist <= 8'h0; // @[Reg.scala 29:22]
    end else if (s0_fire) begin // @[Reg.scala 28:20]
      s1_folded_gh_hist_17_folded_hist <= s0_folded_gh_hist_17_folded_hist;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s1_folded_gh_hist_16_folded_hist <= 8'h0; // @[Reg.scala 29:22]
    end else if (s0_fire) begin // @[Reg.scala 28:20]
      s1_folded_gh_hist_16_folded_hist <= s0_folded_gh_hist_16_folded_hist;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s1_folded_gh_hist_15_folded_hist <= 11'h0; // @[Reg.scala 29:22]
    end else if (s0_fire) begin // @[Reg.scala 28:20]
      s1_folded_gh_hist_15_folded_hist <= s0_folded_gh_hist_15_folded_hist;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s1_folded_gh_hist_14_folded_hist <= 7'h0; // @[Reg.scala 29:22]
    end else if (s0_fire) begin // @[Reg.scala 28:20]
      s1_folded_gh_hist_14_folded_hist <= s0_folded_gh_hist_14_folded_hist;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s1_folded_gh_hist_13_folded_hist <= 7'h0; // @[Reg.scala 29:22]
    end else if (s0_fire) begin // @[Reg.scala 28:20]
      s1_folded_gh_hist_13_folded_hist <= s0_folded_gh_hist_13_folded_hist;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s1_folded_gh_hist_12_folded_hist <= 7'h0; // @[Reg.scala 29:22]
    end else if (s0_fire) begin // @[Reg.scala 28:20]
      s1_folded_gh_hist_12_folded_hist <= s0_folded_gh_hist_12_folded_hist;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s1_folded_gh_hist_11_folded_hist <= 8'h0; // @[Reg.scala 29:22]
    end else if (s0_fire) begin // @[Reg.scala 28:20]
      s1_folded_gh_hist_11_folded_hist <= s0_folded_gh_hist_11_folded_hist;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s1_folded_gh_hist_10_folded_hist <= 9'h0; // @[Reg.scala 29:22]
    end else if (s0_fire) begin // @[Reg.scala 28:20]
      s1_folded_gh_hist_10_folded_hist <= s0_folded_gh_hist_10_folded_hist;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s1_folded_gh_hist_9_folded_hist <= 7'h0; // @[Reg.scala 29:22]
    end else if (s0_fire) begin // @[Reg.scala 28:20]
      s1_folded_gh_hist_9_folded_hist <= s0_folded_gh_hist_9_folded_hist;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s1_folded_gh_hist_8_folded_hist <= 8'h0; // @[Reg.scala 29:22]
    end else if (s0_fire) begin // @[Reg.scala 28:20]
      s1_folded_gh_hist_8_folded_hist <= s0_folded_gh_hist_8_folded_hist;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s1_folded_gh_hist_7_folded_hist <= 9'h0; // @[Reg.scala 29:22]
    end else if (s0_fire) begin // @[Reg.scala 28:20]
      s1_folded_gh_hist_7_folded_hist <= s0_folded_gh_hist_7_folded_hist;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s1_folded_gh_hist_6_folded_hist <= 9'h0; // @[Reg.scala 29:22]
    end else if (s0_fire) begin // @[Reg.scala 28:20]
      s1_folded_gh_hist_6_folded_hist <= s0_folded_gh_hist_6_folded_hist;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s1_folded_gh_hist_5_folded_hist <= 11'h0; // @[Reg.scala 29:22]
    end else if (s0_fire) begin // @[Reg.scala 28:20]
      s1_folded_gh_hist_5_folded_hist <= s0_folded_gh_hist_5_folded_hist;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s1_folded_gh_hist_4_folded_hist <= 4'h0; // @[Reg.scala 29:22]
    end else if (s0_fire) begin // @[Reg.scala 28:20]
      s1_folded_gh_hist_4_folded_hist <= s0_folded_gh_hist_4_folded_hist;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s1_folded_gh_hist_3_folded_hist <= 11'h0; // @[Reg.scala 29:22]
    end else if (s0_fire) begin // @[Reg.scala 28:20]
      s1_folded_gh_hist_3_folded_hist <= s0_folded_gh_hist_3_folded_hist;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s1_folded_gh_hist_2_folded_hist <= 8'h0; // @[Reg.scala 29:22]
    end else if (s0_fire) begin // @[Reg.scala 28:20]
      s1_folded_gh_hist_2_folded_hist <= s0_folded_gh_hist_2_folded_hist;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s1_folded_gh_hist_1_folded_hist <= 8'h0; // @[Reg.scala 29:22]
    end else if (s0_fire) begin // @[Reg.scala 28:20]
      s1_folded_gh_hist_1_folded_hist <= s0_folded_gh_hist_1_folded_hist;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s1_folded_gh_hist_0_folded_hist <= 8'h0; // @[Reg.scala 29:22]
    end else if (s0_fire) begin // @[Reg.scala 28:20]
      s1_folded_gh_hist_0_folded_hist <= s0_folded_gh_hist_0_folded_hist;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s2_folded_gh_hist_17_folded_hist <= 8'h0; // @[Reg.scala 29:22]
    end else if (s1_fire) begin // @[Reg.scala 28:20]
      s2_folded_gh_hist_17_folded_hist <= s1_folded_gh_hist_17_folded_hist;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s2_folded_gh_hist_16_folded_hist <= 8'h0; // @[Reg.scala 29:22]
    end else if (s1_fire) begin // @[Reg.scala 28:20]
      s2_folded_gh_hist_16_folded_hist <= s1_folded_gh_hist_16_folded_hist;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s2_folded_gh_hist_15_folded_hist <= 11'h0; // @[Reg.scala 29:22]
    end else if (s1_fire) begin // @[Reg.scala 28:20]
      s2_folded_gh_hist_15_folded_hist <= s1_folded_gh_hist_15_folded_hist;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s2_folded_gh_hist_14_folded_hist <= 7'h0; // @[Reg.scala 29:22]
    end else if (s1_fire) begin // @[Reg.scala 28:20]
      s2_folded_gh_hist_14_folded_hist <= s1_folded_gh_hist_14_folded_hist;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s2_folded_gh_hist_13_folded_hist <= 7'h0; // @[Reg.scala 29:22]
    end else if (s1_fire) begin // @[Reg.scala 28:20]
      s2_folded_gh_hist_13_folded_hist <= s1_folded_gh_hist_13_folded_hist;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s2_folded_gh_hist_12_folded_hist <= 7'h0; // @[Reg.scala 29:22]
    end else if (s1_fire) begin // @[Reg.scala 28:20]
      s2_folded_gh_hist_12_folded_hist <= s1_folded_gh_hist_12_folded_hist;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s2_folded_gh_hist_11_folded_hist <= 8'h0; // @[Reg.scala 29:22]
    end else if (s1_fire) begin // @[Reg.scala 28:20]
      s2_folded_gh_hist_11_folded_hist <= s1_folded_gh_hist_11_folded_hist;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s2_folded_gh_hist_10_folded_hist <= 9'h0; // @[Reg.scala 29:22]
    end else if (s1_fire) begin // @[Reg.scala 28:20]
      s2_folded_gh_hist_10_folded_hist <= s1_folded_gh_hist_10_folded_hist;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s2_folded_gh_hist_9_folded_hist <= 7'h0; // @[Reg.scala 29:22]
    end else if (s1_fire) begin // @[Reg.scala 28:20]
      s2_folded_gh_hist_9_folded_hist <= s1_folded_gh_hist_9_folded_hist;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s2_folded_gh_hist_8_folded_hist <= 8'h0; // @[Reg.scala 29:22]
    end else if (s1_fire) begin // @[Reg.scala 28:20]
      s2_folded_gh_hist_8_folded_hist <= s1_folded_gh_hist_8_folded_hist;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s2_folded_gh_hist_7_folded_hist <= 9'h0; // @[Reg.scala 29:22]
    end else if (s1_fire) begin // @[Reg.scala 28:20]
      s2_folded_gh_hist_7_folded_hist <= s1_folded_gh_hist_7_folded_hist;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s2_folded_gh_hist_6_folded_hist <= 9'h0; // @[Reg.scala 29:22]
    end else if (s1_fire) begin // @[Reg.scala 28:20]
      s2_folded_gh_hist_6_folded_hist <= s1_folded_gh_hist_6_folded_hist;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s2_folded_gh_hist_5_folded_hist <= 11'h0; // @[Reg.scala 29:22]
    end else if (s1_fire) begin // @[Reg.scala 28:20]
      s2_folded_gh_hist_5_folded_hist <= s1_folded_gh_hist_5_folded_hist;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s2_folded_gh_hist_4_folded_hist <= 4'h0; // @[Reg.scala 29:22]
    end else if (s1_fire) begin // @[Reg.scala 28:20]
      s2_folded_gh_hist_4_folded_hist <= s1_folded_gh_hist_4_folded_hist;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s2_folded_gh_hist_3_folded_hist <= 11'h0; // @[Reg.scala 29:22]
    end else if (s1_fire) begin // @[Reg.scala 28:20]
      s2_folded_gh_hist_3_folded_hist <= s1_folded_gh_hist_3_folded_hist;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s2_folded_gh_hist_2_folded_hist <= 8'h0; // @[Reg.scala 29:22]
    end else if (s1_fire) begin // @[Reg.scala 28:20]
      s2_folded_gh_hist_2_folded_hist <= s1_folded_gh_hist_2_folded_hist;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s2_folded_gh_hist_1_folded_hist <= 8'h0; // @[Reg.scala 29:22]
    end else if (s1_fire) begin // @[Reg.scala 28:20]
      s2_folded_gh_hist_1_folded_hist <= s1_folded_gh_hist_1_folded_hist;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s2_folded_gh_hist_0_folded_hist <= 8'h0; // @[Reg.scala 29:22]
    end else if (s1_fire) begin // @[Reg.scala 28:20]
      s2_folded_gh_hist_0_folded_hist <= s1_folded_gh_hist_0_folded_hist;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s3_folded_gh_hist_17_folded_hist <= 8'h0; // @[Reg.scala 29:22]
    end else if (s2_valid) begin // @[Reg.scala 28:20]
      s3_folded_gh_hist_17_folded_hist <= s2_folded_gh_hist_17_folded_hist;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s3_folded_gh_hist_16_folded_hist <= 8'h0; // @[Reg.scala 29:22]
    end else if (s2_valid) begin // @[Reg.scala 28:20]
      s3_folded_gh_hist_16_folded_hist <= s2_folded_gh_hist_16_folded_hist;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s3_folded_gh_hist_15_folded_hist <= 11'h0; // @[Reg.scala 29:22]
    end else if (s2_valid) begin // @[Reg.scala 28:20]
      s3_folded_gh_hist_15_folded_hist <= s2_folded_gh_hist_15_folded_hist;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s3_folded_gh_hist_14_folded_hist <= 7'h0; // @[Reg.scala 29:22]
    end else if (s2_valid) begin // @[Reg.scala 28:20]
      s3_folded_gh_hist_14_folded_hist <= s2_folded_gh_hist_14_folded_hist;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s3_folded_gh_hist_13_folded_hist <= 7'h0; // @[Reg.scala 29:22]
    end else if (s2_valid) begin // @[Reg.scala 28:20]
      s3_folded_gh_hist_13_folded_hist <= s2_folded_gh_hist_13_folded_hist;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s3_folded_gh_hist_12_folded_hist <= 7'h0; // @[Reg.scala 29:22]
    end else if (s2_valid) begin // @[Reg.scala 28:20]
      s3_folded_gh_hist_12_folded_hist <= s2_folded_gh_hist_12_folded_hist;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s3_folded_gh_hist_11_folded_hist <= 8'h0; // @[Reg.scala 29:22]
    end else if (s2_valid) begin // @[Reg.scala 28:20]
      s3_folded_gh_hist_11_folded_hist <= s2_folded_gh_hist_11_folded_hist;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s3_folded_gh_hist_10_folded_hist <= 9'h0; // @[Reg.scala 29:22]
    end else if (s2_valid) begin // @[Reg.scala 28:20]
      s3_folded_gh_hist_10_folded_hist <= s2_folded_gh_hist_10_folded_hist;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s3_folded_gh_hist_9_folded_hist <= 7'h0; // @[Reg.scala 29:22]
    end else if (s2_valid) begin // @[Reg.scala 28:20]
      s3_folded_gh_hist_9_folded_hist <= s2_folded_gh_hist_9_folded_hist;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s3_folded_gh_hist_8_folded_hist <= 8'h0; // @[Reg.scala 29:22]
    end else if (s2_valid) begin // @[Reg.scala 28:20]
      s3_folded_gh_hist_8_folded_hist <= s2_folded_gh_hist_8_folded_hist;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s3_folded_gh_hist_7_folded_hist <= 9'h0; // @[Reg.scala 29:22]
    end else if (s2_valid) begin // @[Reg.scala 28:20]
      s3_folded_gh_hist_7_folded_hist <= s2_folded_gh_hist_7_folded_hist;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s3_folded_gh_hist_6_folded_hist <= 9'h0; // @[Reg.scala 29:22]
    end else if (s2_valid) begin // @[Reg.scala 28:20]
      s3_folded_gh_hist_6_folded_hist <= s2_folded_gh_hist_6_folded_hist;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s3_folded_gh_hist_5_folded_hist <= 11'h0; // @[Reg.scala 29:22]
    end else if (s2_valid) begin // @[Reg.scala 28:20]
      s3_folded_gh_hist_5_folded_hist <= s2_folded_gh_hist_5_folded_hist;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s3_folded_gh_hist_4_folded_hist <= 4'h0; // @[Reg.scala 29:22]
    end else if (s2_valid) begin // @[Reg.scala 28:20]
      s3_folded_gh_hist_4_folded_hist <= s2_folded_gh_hist_4_folded_hist;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s3_folded_gh_hist_3_folded_hist <= 11'h0; // @[Reg.scala 29:22]
    end else if (s2_valid) begin // @[Reg.scala 28:20]
      s3_folded_gh_hist_3_folded_hist <= s2_folded_gh_hist_3_folded_hist;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s3_folded_gh_hist_2_folded_hist <= 8'h0; // @[Reg.scala 29:22]
    end else if (s2_valid) begin // @[Reg.scala 28:20]
      s3_folded_gh_hist_2_folded_hist <= s2_folded_gh_hist_2_folded_hist;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s3_folded_gh_hist_1_folded_hist <= 8'h0; // @[Reg.scala 29:22]
    end else if (s2_valid) begin // @[Reg.scala 28:20]
      s3_folded_gh_hist_1_folded_hist <= s2_folded_gh_hist_1_folded_hist;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s3_folded_gh_hist_0_folded_hist <= 8'h0; // @[Reg.scala 29:22]
    end else if (s2_valid) begin // @[Reg.scala 28:20]
      s3_folded_gh_hist_0_folded_hist <= s2_folded_gh_hist_0_folded_hist;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 272:31 671:21]
      s0_last_br_num_oh_reg <= 3'h0;
    end else begin
      s0_last_br_num_oh_reg <= s0_last_br_num_oh_ppm_out_res;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s1_last_br_num_oh <= 3'h0; // @[Reg.scala 29:22]
    end else if (s0_fire) begin // @[Reg.scala 28:20]
      s1_last_br_num_oh <= s0_last_br_num_oh;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s2_last_br_num_oh <= 3'h0; // @[Reg.scala 29:22]
    end else if (s1_fire) begin // @[Reg.scala 28:20]
      s2_last_br_num_oh <= s1_last_br_num_oh;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s3_last_br_num_oh <= 3'h0; // @[Reg.scala 29:22]
    end else if (s2_valid) begin // @[Reg.scala 28:20]
      s3_last_br_num_oh <= s2_last_br_num_oh;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 278:37 670:27]
      s0_ahead_fh_oldest_bits_reg_afhob_5_bits_0 <= 1'h0;
    end else begin
      s0_ahead_fh_oldest_bits_reg_afhob_5_bits_0 <= s0_ahead_fh_oldest_bits_ppm_out_res_afhob_5_bits_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 278:37 670:27]
      s0_ahead_fh_oldest_bits_reg_afhob_5_bits_1 <= 1'h0;
    end else begin
      s0_ahead_fh_oldest_bits_reg_afhob_5_bits_1 <= s0_ahead_fh_oldest_bits_ppm_out_res_afhob_5_bits_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 278:37 670:27]
      s0_ahead_fh_oldest_bits_reg_afhob_5_bits_2 <= 1'h0;
    end else begin
      s0_ahead_fh_oldest_bits_reg_afhob_5_bits_2 <= s0_ahead_fh_oldest_bits_ppm_out_res_afhob_5_bits_2;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 278:37 670:27]
      s0_ahead_fh_oldest_bits_reg_afhob_5_bits_3 <= 1'h0;
    end else begin
      s0_ahead_fh_oldest_bits_reg_afhob_5_bits_3 <= s0_ahead_fh_oldest_bits_ppm_out_res_afhob_5_bits_3;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 278:37 670:27]
      s0_ahead_fh_oldest_bits_reg_afhob_4_bits_0 <= 1'h0;
    end else begin
      s0_ahead_fh_oldest_bits_reg_afhob_4_bits_0 <= s0_ahead_fh_oldest_bits_ppm_out_res_afhob_4_bits_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 278:37 670:27]
      s0_ahead_fh_oldest_bits_reg_afhob_4_bits_1 <= 1'h0;
    end else begin
      s0_ahead_fh_oldest_bits_reg_afhob_4_bits_1 <= s0_ahead_fh_oldest_bits_ppm_out_res_afhob_4_bits_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 278:37 670:27]
      s0_ahead_fh_oldest_bits_reg_afhob_4_bits_2 <= 1'h0;
    end else begin
      s0_ahead_fh_oldest_bits_reg_afhob_4_bits_2 <= s0_ahead_fh_oldest_bits_ppm_out_res_afhob_4_bits_2;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 278:37 670:27]
      s0_ahead_fh_oldest_bits_reg_afhob_4_bits_3 <= 1'h0;
    end else begin
      s0_ahead_fh_oldest_bits_reg_afhob_4_bits_3 <= s0_ahead_fh_oldest_bits_ppm_out_res_afhob_4_bits_3;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 278:37 670:27]
      s0_ahead_fh_oldest_bits_reg_afhob_3_bits_0 <= 1'h0;
    end else begin
      s0_ahead_fh_oldest_bits_reg_afhob_3_bits_0 <= s0_ahead_fh_oldest_bits_ppm_out_res_afhob_3_bits_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 278:37 670:27]
      s0_ahead_fh_oldest_bits_reg_afhob_3_bits_1 <= 1'h0;
    end else begin
      s0_ahead_fh_oldest_bits_reg_afhob_3_bits_1 <= s0_ahead_fh_oldest_bits_ppm_out_res_afhob_3_bits_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 278:37 670:27]
      s0_ahead_fh_oldest_bits_reg_afhob_3_bits_2 <= 1'h0;
    end else begin
      s0_ahead_fh_oldest_bits_reg_afhob_3_bits_2 <= s0_ahead_fh_oldest_bits_ppm_out_res_afhob_3_bits_2;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 278:37 670:27]
      s0_ahead_fh_oldest_bits_reg_afhob_3_bits_3 <= 1'h0;
    end else begin
      s0_ahead_fh_oldest_bits_reg_afhob_3_bits_3 <= s0_ahead_fh_oldest_bits_ppm_out_res_afhob_3_bits_3;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 278:37 670:27]
      s0_ahead_fh_oldest_bits_reg_afhob_2_bits_0 <= 1'h0;
    end else begin
      s0_ahead_fh_oldest_bits_reg_afhob_2_bits_0 <= s0_ahead_fh_oldest_bits_ppm_out_res_afhob_2_bits_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 278:37 670:27]
      s0_ahead_fh_oldest_bits_reg_afhob_2_bits_1 <= 1'h0;
    end else begin
      s0_ahead_fh_oldest_bits_reg_afhob_2_bits_1 <= s0_ahead_fh_oldest_bits_ppm_out_res_afhob_2_bits_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 278:37 670:27]
      s0_ahead_fh_oldest_bits_reg_afhob_2_bits_2 <= 1'h0;
    end else begin
      s0_ahead_fh_oldest_bits_reg_afhob_2_bits_2 <= s0_ahead_fh_oldest_bits_ppm_out_res_afhob_2_bits_2;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 278:37 670:27]
      s0_ahead_fh_oldest_bits_reg_afhob_2_bits_3 <= 1'h0;
    end else begin
      s0_ahead_fh_oldest_bits_reg_afhob_2_bits_3 <= s0_ahead_fh_oldest_bits_ppm_out_res_afhob_2_bits_3;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 278:37 670:27]
      s0_ahead_fh_oldest_bits_reg_afhob_1_bits_0 <= 1'h0;
    end else begin
      s0_ahead_fh_oldest_bits_reg_afhob_1_bits_0 <= s0_ahead_fh_oldest_bits_ppm_out_res_afhob_1_bits_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 278:37 670:27]
      s0_ahead_fh_oldest_bits_reg_afhob_1_bits_1 <= 1'h0;
    end else begin
      s0_ahead_fh_oldest_bits_reg_afhob_1_bits_1 <= s0_ahead_fh_oldest_bits_ppm_out_res_afhob_1_bits_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 278:37 670:27]
      s0_ahead_fh_oldest_bits_reg_afhob_1_bits_2 <= 1'h0;
    end else begin
      s0_ahead_fh_oldest_bits_reg_afhob_1_bits_2 <= s0_ahead_fh_oldest_bits_ppm_out_res_afhob_1_bits_2;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 278:37 670:27]
      s0_ahead_fh_oldest_bits_reg_afhob_1_bits_3 <= 1'h0;
    end else begin
      s0_ahead_fh_oldest_bits_reg_afhob_1_bits_3 <= s0_ahead_fh_oldest_bits_ppm_out_res_afhob_1_bits_3;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 278:37 670:27]
      s0_ahead_fh_oldest_bits_reg_afhob_0_bits_0 <= 1'h0;
    end else begin
      s0_ahead_fh_oldest_bits_reg_afhob_0_bits_0 <= s0_ahead_fh_oldest_bits_ppm_out_res_afhob_0_bits_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 278:37 670:27]
      s0_ahead_fh_oldest_bits_reg_afhob_0_bits_1 <= 1'h0;
    end else begin
      s0_ahead_fh_oldest_bits_reg_afhob_0_bits_1 <= s0_ahead_fh_oldest_bits_ppm_out_res_afhob_0_bits_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 278:37 670:27]
      s0_ahead_fh_oldest_bits_reg_afhob_0_bits_2 <= 1'h0;
    end else begin
      s0_ahead_fh_oldest_bits_reg_afhob_0_bits_2 <= s0_ahead_fh_oldest_bits_ppm_out_res_afhob_0_bits_2;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 278:37 670:27]
      s0_ahead_fh_oldest_bits_reg_afhob_0_bits_3 <= 1'h0;
    end else begin
      s0_ahead_fh_oldest_bits_reg_afhob_0_bits_3 <= s0_ahead_fh_oldest_bits_ppm_out_res_afhob_0_bits_3;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s1_ahead_fh_oldest_bits_afhob_5_bits_0 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s0_fire) begin // @[Reg.scala 28:20]
      s1_ahead_fh_oldest_bits_afhob_5_bits_0 <= s0_ahead_fh_oldest_bits_afhob_5_bits_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s1_ahead_fh_oldest_bits_afhob_5_bits_1 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s0_fire) begin // @[Reg.scala 28:20]
      s1_ahead_fh_oldest_bits_afhob_5_bits_1 <= s0_ahead_fh_oldest_bits_afhob_5_bits_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s1_ahead_fh_oldest_bits_afhob_5_bits_2 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s0_fire) begin // @[Reg.scala 28:20]
      s1_ahead_fh_oldest_bits_afhob_5_bits_2 <= s0_ahead_fh_oldest_bits_afhob_5_bits_2;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s1_ahead_fh_oldest_bits_afhob_5_bits_3 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s0_fire) begin // @[Reg.scala 28:20]
      s1_ahead_fh_oldest_bits_afhob_5_bits_3 <= s0_ahead_fh_oldest_bits_afhob_5_bits_3;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s1_ahead_fh_oldest_bits_afhob_4_bits_0 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s0_fire) begin // @[Reg.scala 28:20]
      s1_ahead_fh_oldest_bits_afhob_4_bits_0 <= s0_ahead_fh_oldest_bits_afhob_4_bits_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s1_ahead_fh_oldest_bits_afhob_4_bits_1 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s0_fire) begin // @[Reg.scala 28:20]
      s1_ahead_fh_oldest_bits_afhob_4_bits_1 <= s0_ahead_fh_oldest_bits_afhob_4_bits_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s1_ahead_fh_oldest_bits_afhob_4_bits_2 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s0_fire) begin // @[Reg.scala 28:20]
      s1_ahead_fh_oldest_bits_afhob_4_bits_2 <= s0_ahead_fh_oldest_bits_afhob_4_bits_2;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s1_ahead_fh_oldest_bits_afhob_4_bits_3 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s0_fire) begin // @[Reg.scala 28:20]
      s1_ahead_fh_oldest_bits_afhob_4_bits_3 <= s0_ahead_fh_oldest_bits_afhob_4_bits_3;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s1_ahead_fh_oldest_bits_afhob_3_bits_0 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s0_fire) begin // @[Reg.scala 28:20]
      s1_ahead_fh_oldest_bits_afhob_3_bits_0 <= s0_ahead_fh_oldest_bits_afhob_3_bits_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s1_ahead_fh_oldest_bits_afhob_3_bits_1 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s0_fire) begin // @[Reg.scala 28:20]
      s1_ahead_fh_oldest_bits_afhob_3_bits_1 <= s0_ahead_fh_oldest_bits_afhob_3_bits_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s1_ahead_fh_oldest_bits_afhob_3_bits_2 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s0_fire) begin // @[Reg.scala 28:20]
      s1_ahead_fh_oldest_bits_afhob_3_bits_2 <= s0_ahead_fh_oldest_bits_afhob_3_bits_2;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s1_ahead_fh_oldest_bits_afhob_3_bits_3 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s0_fire) begin // @[Reg.scala 28:20]
      s1_ahead_fh_oldest_bits_afhob_3_bits_3 <= s0_ahead_fh_oldest_bits_afhob_3_bits_3;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s1_ahead_fh_oldest_bits_afhob_2_bits_0 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s0_fire) begin // @[Reg.scala 28:20]
      s1_ahead_fh_oldest_bits_afhob_2_bits_0 <= s0_ahead_fh_oldest_bits_afhob_2_bits_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s1_ahead_fh_oldest_bits_afhob_2_bits_1 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s0_fire) begin // @[Reg.scala 28:20]
      s1_ahead_fh_oldest_bits_afhob_2_bits_1 <= s0_ahead_fh_oldest_bits_afhob_2_bits_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s1_ahead_fh_oldest_bits_afhob_2_bits_2 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s0_fire) begin // @[Reg.scala 28:20]
      s1_ahead_fh_oldest_bits_afhob_2_bits_2 <= s0_ahead_fh_oldest_bits_afhob_2_bits_2;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s1_ahead_fh_oldest_bits_afhob_2_bits_3 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s0_fire) begin // @[Reg.scala 28:20]
      s1_ahead_fh_oldest_bits_afhob_2_bits_3 <= s0_ahead_fh_oldest_bits_afhob_2_bits_3;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s1_ahead_fh_oldest_bits_afhob_1_bits_0 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s0_fire) begin // @[Reg.scala 28:20]
      s1_ahead_fh_oldest_bits_afhob_1_bits_0 <= s0_ahead_fh_oldest_bits_afhob_1_bits_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s1_ahead_fh_oldest_bits_afhob_1_bits_1 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s0_fire) begin // @[Reg.scala 28:20]
      s1_ahead_fh_oldest_bits_afhob_1_bits_1 <= s0_ahead_fh_oldest_bits_afhob_1_bits_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s1_ahead_fh_oldest_bits_afhob_1_bits_2 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s0_fire) begin // @[Reg.scala 28:20]
      s1_ahead_fh_oldest_bits_afhob_1_bits_2 <= s0_ahead_fh_oldest_bits_afhob_1_bits_2;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s1_ahead_fh_oldest_bits_afhob_1_bits_3 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s0_fire) begin // @[Reg.scala 28:20]
      s1_ahead_fh_oldest_bits_afhob_1_bits_3 <= s0_ahead_fh_oldest_bits_afhob_1_bits_3;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s1_ahead_fh_oldest_bits_afhob_0_bits_0 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s0_fire) begin // @[Reg.scala 28:20]
      s1_ahead_fh_oldest_bits_afhob_0_bits_0 <= s0_ahead_fh_oldest_bits_afhob_0_bits_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s1_ahead_fh_oldest_bits_afhob_0_bits_1 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s0_fire) begin // @[Reg.scala 28:20]
      s1_ahead_fh_oldest_bits_afhob_0_bits_1 <= s0_ahead_fh_oldest_bits_afhob_0_bits_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s1_ahead_fh_oldest_bits_afhob_0_bits_2 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s0_fire) begin // @[Reg.scala 28:20]
      s1_ahead_fh_oldest_bits_afhob_0_bits_2 <= s0_ahead_fh_oldest_bits_afhob_0_bits_2;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s1_ahead_fh_oldest_bits_afhob_0_bits_3 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s0_fire) begin // @[Reg.scala 28:20]
      s1_ahead_fh_oldest_bits_afhob_0_bits_3 <= s0_ahead_fh_oldest_bits_afhob_0_bits_3;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s2_ahead_fh_oldest_bits_afhob_5_bits_0 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s1_fire) begin // @[Reg.scala 28:20]
      s2_ahead_fh_oldest_bits_afhob_5_bits_0 <= s1_ahead_fh_oldest_bits_afhob_5_bits_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s2_ahead_fh_oldest_bits_afhob_5_bits_1 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s1_fire) begin // @[Reg.scala 28:20]
      s2_ahead_fh_oldest_bits_afhob_5_bits_1 <= s1_ahead_fh_oldest_bits_afhob_5_bits_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s2_ahead_fh_oldest_bits_afhob_5_bits_2 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s1_fire) begin // @[Reg.scala 28:20]
      s2_ahead_fh_oldest_bits_afhob_5_bits_2 <= s1_ahead_fh_oldest_bits_afhob_5_bits_2;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s2_ahead_fh_oldest_bits_afhob_5_bits_3 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s1_fire) begin // @[Reg.scala 28:20]
      s2_ahead_fh_oldest_bits_afhob_5_bits_3 <= s1_ahead_fh_oldest_bits_afhob_5_bits_3;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s2_ahead_fh_oldest_bits_afhob_4_bits_0 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s1_fire) begin // @[Reg.scala 28:20]
      s2_ahead_fh_oldest_bits_afhob_4_bits_0 <= s1_ahead_fh_oldest_bits_afhob_4_bits_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s2_ahead_fh_oldest_bits_afhob_4_bits_1 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s1_fire) begin // @[Reg.scala 28:20]
      s2_ahead_fh_oldest_bits_afhob_4_bits_1 <= s1_ahead_fh_oldest_bits_afhob_4_bits_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s2_ahead_fh_oldest_bits_afhob_4_bits_2 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s1_fire) begin // @[Reg.scala 28:20]
      s2_ahead_fh_oldest_bits_afhob_4_bits_2 <= s1_ahead_fh_oldest_bits_afhob_4_bits_2;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s2_ahead_fh_oldest_bits_afhob_4_bits_3 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s1_fire) begin // @[Reg.scala 28:20]
      s2_ahead_fh_oldest_bits_afhob_4_bits_3 <= s1_ahead_fh_oldest_bits_afhob_4_bits_3;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s2_ahead_fh_oldest_bits_afhob_3_bits_0 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s1_fire) begin // @[Reg.scala 28:20]
      s2_ahead_fh_oldest_bits_afhob_3_bits_0 <= s1_ahead_fh_oldest_bits_afhob_3_bits_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s2_ahead_fh_oldest_bits_afhob_3_bits_1 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s1_fire) begin // @[Reg.scala 28:20]
      s2_ahead_fh_oldest_bits_afhob_3_bits_1 <= s1_ahead_fh_oldest_bits_afhob_3_bits_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s2_ahead_fh_oldest_bits_afhob_3_bits_2 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s1_fire) begin // @[Reg.scala 28:20]
      s2_ahead_fh_oldest_bits_afhob_3_bits_2 <= s1_ahead_fh_oldest_bits_afhob_3_bits_2;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s2_ahead_fh_oldest_bits_afhob_3_bits_3 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s1_fire) begin // @[Reg.scala 28:20]
      s2_ahead_fh_oldest_bits_afhob_3_bits_3 <= s1_ahead_fh_oldest_bits_afhob_3_bits_3;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s2_ahead_fh_oldest_bits_afhob_2_bits_0 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s1_fire) begin // @[Reg.scala 28:20]
      s2_ahead_fh_oldest_bits_afhob_2_bits_0 <= s1_ahead_fh_oldest_bits_afhob_2_bits_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s2_ahead_fh_oldest_bits_afhob_2_bits_1 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s1_fire) begin // @[Reg.scala 28:20]
      s2_ahead_fh_oldest_bits_afhob_2_bits_1 <= s1_ahead_fh_oldest_bits_afhob_2_bits_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s2_ahead_fh_oldest_bits_afhob_2_bits_2 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s1_fire) begin // @[Reg.scala 28:20]
      s2_ahead_fh_oldest_bits_afhob_2_bits_2 <= s1_ahead_fh_oldest_bits_afhob_2_bits_2;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s2_ahead_fh_oldest_bits_afhob_2_bits_3 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s1_fire) begin // @[Reg.scala 28:20]
      s2_ahead_fh_oldest_bits_afhob_2_bits_3 <= s1_ahead_fh_oldest_bits_afhob_2_bits_3;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s2_ahead_fh_oldest_bits_afhob_1_bits_0 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s1_fire) begin // @[Reg.scala 28:20]
      s2_ahead_fh_oldest_bits_afhob_1_bits_0 <= s1_ahead_fh_oldest_bits_afhob_1_bits_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s2_ahead_fh_oldest_bits_afhob_1_bits_1 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s1_fire) begin // @[Reg.scala 28:20]
      s2_ahead_fh_oldest_bits_afhob_1_bits_1 <= s1_ahead_fh_oldest_bits_afhob_1_bits_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s2_ahead_fh_oldest_bits_afhob_1_bits_2 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s1_fire) begin // @[Reg.scala 28:20]
      s2_ahead_fh_oldest_bits_afhob_1_bits_2 <= s1_ahead_fh_oldest_bits_afhob_1_bits_2;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s2_ahead_fh_oldest_bits_afhob_1_bits_3 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s1_fire) begin // @[Reg.scala 28:20]
      s2_ahead_fh_oldest_bits_afhob_1_bits_3 <= s1_ahead_fh_oldest_bits_afhob_1_bits_3;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s2_ahead_fh_oldest_bits_afhob_0_bits_0 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s1_fire) begin // @[Reg.scala 28:20]
      s2_ahead_fh_oldest_bits_afhob_0_bits_0 <= s1_ahead_fh_oldest_bits_afhob_0_bits_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s2_ahead_fh_oldest_bits_afhob_0_bits_1 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s1_fire) begin // @[Reg.scala 28:20]
      s2_ahead_fh_oldest_bits_afhob_0_bits_1 <= s1_ahead_fh_oldest_bits_afhob_0_bits_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s2_ahead_fh_oldest_bits_afhob_0_bits_2 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s1_fire) begin // @[Reg.scala 28:20]
      s2_ahead_fh_oldest_bits_afhob_0_bits_2 <= s1_ahead_fh_oldest_bits_afhob_0_bits_2;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s2_ahead_fh_oldest_bits_afhob_0_bits_3 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s1_fire) begin // @[Reg.scala 28:20]
      s2_ahead_fh_oldest_bits_afhob_0_bits_3 <= s1_ahead_fh_oldest_bits_afhob_0_bits_3;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s3_ahead_fh_oldest_bits_afhob_5_bits_0 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s2_valid) begin // @[Reg.scala 28:20]
      s3_ahead_fh_oldest_bits_afhob_5_bits_0 <= s2_ahead_fh_oldest_bits_afhob_5_bits_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s3_ahead_fh_oldest_bits_afhob_5_bits_1 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s2_valid) begin // @[Reg.scala 28:20]
      s3_ahead_fh_oldest_bits_afhob_5_bits_1 <= s2_ahead_fh_oldest_bits_afhob_5_bits_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s3_ahead_fh_oldest_bits_afhob_5_bits_2 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s2_valid) begin // @[Reg.scala 28:20]
      s3_ahead_fh_oldest_bits_afhob_5_bits_2 <= s2_ahead_fh_oldest_bits_afhob_5_bits_2;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s3_ahead_fh_oldest_bits_afhob_5_bits_3 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s2_valid) begin // @[Reg.scala 28:20]
      s3_ahead_fh_oldest_bits_afhob_5_bits_3 <= s2_ahead_fh_oldest_bits_afhob_5_bits_3;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s3_ahead_fh_oldest_bits_afhob_4_bits_0 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s2_valid) begin // @[Reg.scala 28:20]
      s3_ahead_fh_oldest_bits_afhob_4_bits_0 <= s2_ahead_fh_oldest_bits_afhob_4_bits_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s3_ahead_fh_oldest_bits_afhob_4_bits_1 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s2_valid) begin // @[Reg.scala 28:20]
      s3_ahead_fh_oldest_bits_afhob_4_bits_1 <= s2_ahead_fh_oldest_bits_afhob_4_bits_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s3_ahead_fh_oldest_bits_afhob_4_bits_2 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s2_valid) begin // @[Reg.scala 28:20]
      s3_ahead_fh_oldest_bits_afhob_4_bits_2 <= s2_ahead_fh_oldest_bits_afhob_4_bits_2;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s3_ahead_fh_oldest_bits_afhob_4_bits_3 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s2_valid) begin // @[Reg.scala 28:20]
      s3_ahead_fh_oldest_bits_afhob_4_bits_3 <= s2_ahead_fh_oldest_bits_afhob_4_bits_3;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s3_ahead_fh_oldest_bits_afhob_3_bits_0 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s2_valid) begin // @[Reg.scala 28:20]
      s3_ahead_fh_oldest_bits_afhob_3_bits_0 <= s2_ahead_fh_oldest_bits_afhob_3_bits_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s3_ahead_fh_oldest_bits_afhob_3_bits_1 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s2_valid) begin // @[Reg.scala 28:20]
      s3_ahead_fh_oldest_bits_afhob_3_bits_1 <= s2_ahead_fh_oldest_bits_afhob_3_bits_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s3_ahead_fh_oldest_bits_afhob_3_bits_2 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s2_valid) begin // @[Reg.scala 28:20]
      s3_ahead_fh_oldest_bits_afhob_3_bits_2 <= s2_ahead_fh_oldest_bits_afhob_3_bits_2;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s3_ahead_fh_oldest_bits_afhob_3_bits_3 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s2_valid) begin // @[Reg.scala 28:20]
      s3_ahead_fh_oldest_bits_afhob_3_bits_3 <= s2_ahead_fh_oldest_bits_afhob_3_bits_3;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s3_ahead_fh_oldest_bits_afhob_2_bits_0 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s2_valid) begin // @[Reg.scala 28:20]
      s3_ahead_fh_oldest_bits_afhob_2_bits_0 <= s2_ahead_fh_oldest_bits_afhob_2_bits_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s3_ahead_fh_oldest_bits_afhob_2_bits_1 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s2_valid) begin // @[Reg.scala 28:20]
      s3_ahead_fh_oldest_bits_afhob_2_bits_1 <= s2_ahead_fh_oldest_bits_afhob_2_bits_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s3_ahead_fh_oldest_bits_afhob_2_bits_2 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s2_valid) begin // @[Reg.scala 28:20]
      s3_ahead_fh_oldest_bits_afhob_2_bits_2 <= s2_ahead_fh_oldest_bits_afhob_2_bits_2;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s3_ahead_fh_oldest_bits_afhob_2_bits_3 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s2_valid) begin // @[Reg.scala 28:20]
      s3_ahead_fh_oldest_bits_afhob_2_bits_3 <= s2_ahead_fh_oldest_bits_afhob_2_bits_3;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s3_ahead_fh_oldest_bits_afhob_1_bits_0 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s2_valid) begin // @[Reg.scala 28:20]
      s3_ahead_fh_oldest_bits_afhob_1_bits_0 <= s2_ahead_fh_oldest_bits_afhob_1_bits_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s3_ahead_fh_oldest_bits_afhob_1_bits_1 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s2_valid) begin // @[Reg.scala 28:20]
      s3_ahead_fh_oldest_bits_afhob_1_bits_1 <= s2_ahead_fh_oldest_bits_afhob_1_bits_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s3_ahead_fh_oldest_bits_afhob_1_bits_2 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s2_valid) begin // @[Reg.scala 28:20]
      s3_ahead_fh_oldest_bits_afhob_1_bits_2 <= s2_ahead_fh_oldest_bits_afhob_1_bits_2;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s3_ahead_fh_oldest_bits_afhob_1_bits_3 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s2_valid) begin // @[Reg.scala 28:20]
      s3_ahead_fh_oldest_bits_afhob_1_bits_3 <= s2_ahead_fh_oldest_bits_afhob_1_bits_3;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s3_ahead_fh_oldest_bits_afhob_0_bits_0 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s2_valid) begin // @[Reg.scala 28:20]
      s3_ahead_fh_oldest_bits_afhob_0_bits_0 <= s2_ahead_fh_oldest_bits_afhob_0_bits_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s3_ahead_fh_oldest_bits_afhob_0_bits_1 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s2_valid) begin // @[Reg.scala 28:20]
      s3_ahead_fh_oldest_bits_afhob_0_bits_1 <= s2_ahead_fh_oldest_bits_afhob_0_bits_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s3_ahead_fh_oldest_bits_afhob_0_bits_2 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s2_valid) begin // @[Reg.scala 28:20]
      s3_ahead_fh_oldest_bits_afhob_0_bits_2 <= s2_ahead_fh_oldest_bits_afhob_0_bits_2;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s3_ahead_fh_oldest_bits_afhob_0_bits_3 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s2_valid) begin // @[Reg.scala 28:20]
      s3_ahead_fh_oldest_bits_afhob_0_bits_3 <= s2_ahead_fh_oldest_bits_afhob_0_bits_3;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_0 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_0) begin // @[BPU.scala 293:20]
      ghv_0 <= ghv_write_datas_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_1 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_1) begin // @[BPU.scala 293:20]
      ghv_1 <= ghv_write_datas_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_2 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_2) begin // @[BPU.scala 293:20]
      ghv_2 <= ghv_write_datas_2;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_3 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_3) begin // @[BPU.scala 293:20]
      ghv_3 <= ghv_write_datas_3;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_4 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_4) begin // @[BPU.scala 293:20]
      ghv_4 <= ghv_write_datas_4;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_5 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_5) begin // @[BPU.scala 293:20]
      ghv_5 <= ghv_write_datas_5;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_6 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_6) begin // @[BPU.scala 293:20]
      ghv_6 <= ghv_write_datas_6;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_7 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_7) begin // @[BPU.scala 293:20]
      ghv_7 <= ghv_write_datas_7;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_8 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_8) begin // @[BPU.scala 293:20]
      ghv_8 <= ghv_write_datas_8;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_9 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_9) begin // @[BPU.scala 293:20]
      ghv_9 <= ghv_write_datas_9;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_10 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_10) begin // @[BPU.scala 293:20]
      ghv_10 <= ghv_write_datas_10;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_11 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_11) begin // @[BPU.scala 293:20]
      ghv_11 <= ghv_write_datas_11;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_12 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_12) begin // @[BPU.scala 293:20]
      ghv_12 <= ghv_write_datas_12;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_13 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_13) begin // @[BPU.scala 293:20]
      ghv_13 <= ghv_write_datas_13;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_14 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_14) begin // @[BPU.scala 293:20]
      ghv_14 <= ghv_write_datas_14;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_15 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_15) begin // @[BPU.scala 293:20]
      ghv_15 <= ghv_write_datas_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_16 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_16) begin // @[BPU.scala 293:20]
      ghv_16 <= ghv_write_datas_16;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_17 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_17) begin // @[BPU.scala 293:20]
      ghv_17 <= ghv_write_datas_17;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_18 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_18) begin // @[BPU.scala 293:20]
      ghv_18 <= ghv_write_datas_18;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_19 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_19) begin // @[BPU.scala 293:20]
      ghv_19 <= ghv_write_datas_19;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_20 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_20) begin // @[BPU.scala 293:20]
      ghv_20 <= ghv_write_datas_20;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_21 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_21) begin // @[BPU.scala 293:20]
      ghv_21 <= ghv_write_datas_21;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_22 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_22) begin // @[BPU.scala 293:20]
      ghv_22 <= ghv_write_datas_22;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_23 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_23) begin // @[BPU.scala 293:20]
      ghv_23 <= ghv_write_datas_23;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_24 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_24) begin // @[BPU.scala 293:20]
      ghv_24 <= ghv_write_datas_24;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_25 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_25) begin // @[BPU.scala 293:20]
      ghv_25 <= ghv_write_datas_25;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_26 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_26) begin // @[BPU.scala 293:20]
      ghv_26 <= ghv_write_datas_26;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_27 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_27) begin // @[BPU.scala 293:20]
      ghv_27 <= ghv_write_datas_27;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_28 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_28) begin // @[BPU.scala 293:20]
      ghv_28 <= ghv_write_datas_28;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_29 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_29) begin // @[BPU.scala 293:20]
      ghv_29 <= ghv_write_datas_29;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_30 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_30) begin // @[BPU.scala 293:20]
      ghv_30 <= ghv_write_datas_30;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_31 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_31) begin // @[BPU.scala 293:20]
      ghv_31 <= ghv_write_datas_31;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_32 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_32) begin // @[BPU.scala 293:20]
      ghv_32 <= ghv_write_datas_32;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_33 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_33) begin // @[BPU.scala 293:20]
      ghv_33 <= ghv_write_datas_33;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_34 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_34) begin // @[BPU.scala 293:20]
      ghv_34 <= ghv_write_datas_34;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_35 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_35) begin // @[BPU.scala 293:20]
      ghv_35 <= ghv_write_datas_35;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_36 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_36) begin // @[BPU.scala 293:20]
      ghv_36 <= ghv_write_datas_36;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_37 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_37) begin // @[BPU.scala 293:20]
      ghv_37 <= ghv_write_datas_37;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_38 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_38) begin // @[BPU.scala 293:20]
      ghv_38 <= ghv_write_datas_38;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_39 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_39) begin // @[BPU.scala 293:20]
      ghv_39 <= ghv_write_datas_39;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_40 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_40) begin // @[BPU.scala 293:20]
      ghv_40 <= ghv_write_datas_40;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_41 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_41) begin // @[BPU.scala 293:20]
      ghv_41 <= ghv_write_datas_41;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_42 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_42) begin // @[BPU.scala 293:20]
      ghv_42 <= ghv_write_datas_42;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_43 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_43) begin // @[BPU.scala 293:20]
      ghv_43 <= ghv_write_datas_43;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_44 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_44) begin // @[BPU.scala 293:20]
      ghv_44 <= ghv_write_datas_44;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_45 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_45) begin // @[BPU.scala 293:20]
      ghv_45 <= ghv_write_datas_45;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_46 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_46) begin // @[BPU.scala 293:20]
      ghv_46 <= ghv_write_datas_46;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_47 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_47) begin // @[BPU.scala 293:20]
      ghv_47 <= ghv_write_datas_47;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_48 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_48) begin // @[BPU.scala 293:20]
      ghv_48 <= ghv_write_datas_48;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_49 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_49) begin // @[BPU.scala 293:20]
      ghv_49 <= ghv_write_datas_49;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_50 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_50) begin // @[BPU.scala 293:20]
      ghv_50 <= ghv_write_datas_50;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_51 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_51) begin // @[BPU.scala 293:20]
      ghv_51 <= ghv_write_datas_51;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_52 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_52) begin // @[BPU.scala 293:20]
      ghv_52 <= ghv_write_datas_52;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_53 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_53) begin // @[BPU.scala 293:20]
      ghv_53 <= ghv_write_datas_53;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_54 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_54) begin // @[BPU.scala 293:20]
      ghv_54 <= ghv_write_datas_54;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_55 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_55) begin // @[BPU.scala 293:20]
      ghv_55 <= ghv_write_datas_55;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_56 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_56) begin // @[BPU.scala 293:20]
      ghv_56 <= ghv_write_datas_56;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_57 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_57) begin // @[BPU.scala 293:20]
      ghv_57 <= ghv_write_datas_57;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_58 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_58) begin // @[BPU.scala 293:20]
      ghv_58 <= ghv_write_datas_58;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_59 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_59) begin // @[BPU.scala 293:20]
      ghv_59 <= ghv_write_datas_59;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_60 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_60) begin // @[BPU.scala 293:20]
      ghv_60 <= ghv_write_datas_60;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_61 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_61) begin // @[BPU.scala 293:20]
      ghv_61 <= ghv_write_datas_61;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_62 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_62) begin // @[BPU.scala 293:20]
      ghv_62 <= ghv_write_datas_62;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_63 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_63) begin // @[BPU.scala 293:20]
      ghv_63 <= ghv_write_datas_63;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_64 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_64) begin // @[BPU.scala 293:20]
      ghv_64 <= ghv_write_datas_64;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_65 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_65) begin // @[BPU.scala 293:20]
      ghv_65 <= ghv_write_datas_65;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_66 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_66) begin // @[BPU.scala 293:20]
      ghv_66 <= ghv_write_datas_66;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_67 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_67) begin // @[BPU.scala 293:20]
      ghv_67 <= ghv_write_datas_67;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_68 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_68) begin // @[BPU.scala 293:20]
      ghv_68 <= ghv_write_datas_68;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_69 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_69) begin // @[BPU.scala 293:20]
      ghv_69 <= ghv_write_datas_69;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_70 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_70) begin // @[BPU.scala 293:20]
      ghv_70 <= ghv_write_datas_70;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_71 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_71) begin // @[BPU.scala 293:20]
      ghv_71 <= ghv_write_datas_71;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_72 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_72) begin // @[BPU.scala 293:20]
      ghv_72 <= ghv_write_datas_72;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_73 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_73) begin // @[BPU.scala 293:20]
      ghv_73 <= ghv_write_datas_73;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_74 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_74) begin // @[BPU.scala 293:20]
      ghv_74 <= ghv_write_datas_74;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_75 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_75) begin // @[BPU.scala 293:20]
      ghv_75 <= ghv_write_datas_75;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_76 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_76) begin // @[BPU.scala 293:20]
      ghv_76 <= ghv_write_datas_76;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_77 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_77) begin // @[BPU.scala 293:20]
      ghv_77 <= ghv_write_datas_77;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_78 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_78) begin // @[BPU.scala 293:20]
      ghv_78 <= ghv_write_datas_78;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_79 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_79) begin // @[BPU.scala 293:20]
      ghv_79 <= ghv_write_datas_79;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_80 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_80) begin // @[BPU.scala 293:20]
      ghv_80 <= ghv_write_datas_80;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_81 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_81) begin // @[BPU.scala 293:20]
      ghv_81 <= ghv_write_datas_81;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_82 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_82) begin // @[BPU.scala 293:20]
      ghv_82 <= ghv_write_datas_82;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_83 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_83) begin // @[BPU.scala 293:20]
      ghv_83 <= ghv_write_datas_83;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_84 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_84) begin // @[BPU.scala 293:20]
      ghv_84 <= ghv_write_datas_84;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_85 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_85) begin // @[BPU.scala 293:20]
      ghv_85 <= ghv_write_datas_85;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_86 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_86) begin // @[BPU.scala 293:20]
      ghv_86 <= ghv_write_datas_86;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_87 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_87) begin // @[BPU.scala 293:20]
      ghv_87 <= ghv_write_datas_87;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_88 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_88) begin // @[BPU.scala 293:20]
      ghv_88 <= ghv_write_datas_88;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_89 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_89) begin // @[BPU.scala 293:20]
      ghv_89 <= ghv_write_datas_89;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_90 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_90) begin // @[BPU.scala 293:20]
      ghv_90 <= ghv_write_datas_90;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_91 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_91) begin // @[BPU.scala 293:20]
      ghv_91 <= ghv_write_datas_91;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_92 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_92) begin // @[BPU.scala 293:20]
      ghv_92 <= ghv_write_datas_92;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_93 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_93) begin // @[BPU.scala 293:20]
      ghv_93 <= ghv_write_datas_93;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_94 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_94) begin // @[BPU.scala 293:20]
      ghv_94 <= ghv_write_datas_94;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_95 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_95) begin // @[BPU.scala 293:20]
      ghv_95 <= ghv_write_datas_95;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_96 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_96) begin // @[BPU.scala 293:20]
      ghv_96 <= ghv_write_datas_96;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_97 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_97) begin // @[BPU.scala 293:20]
      ghv_97 <= ghv_write_datas_97;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_98 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_98) begin // @[BPU.scala 293:20]
      ghv_98 <= ghv_write_datas_98;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_99 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_99) begin // @[BPU.scala 293:20]
      ghv_99 <= ghv_write_datas_99;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_100 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_100) begin // @[BPU.scala 293:20]
      ghv_100 <= ghv_write_datas_100;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_101 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_101) begin // @[BPU.scala 293:20]
      ghv_101 <= ghv_write_datas_101;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_102 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_102) begin // @[BPU.scala 293:20]
      ghv_102 <= ghv_write_datas_102;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_103 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_103) begin // @[BPU.scala 293:20]
      ghv_103 <= ghv_write_datas_103;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_104 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_104) begin // @[BPU.scala 293:20]
      ghv_104 <= ghv_write_datas_104;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_105 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_105) begin // @[BPU.scala 293:20]
      ghv_105 <= ghv_write_datas_105;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_106 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_106) begin // @[BPU.scala 293:20]
      ghv_106 <= ghv_write_datas_106;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_107 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_107) begin // @[BPU.scala 293:20]
      ghv_107 <= ghv_write_datas_107;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_108 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_108) begin // @[BPU.scala 293:20]
      ghv_108 <= ghv_write_datas_108;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_109 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_109) begin // @[BPU.scala 293:20]
      ghv_109 <= ghv_write_datas_109;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_110 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_110) begin // @[BPU.scala 293:20]
      ghv_110 <= ghv_write_datas_110;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_111 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_111) begin // @[BPU.scala 293:20]
      ghv_111 <= ghv_write_datas_111;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_112 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_112) begin // @[BPU.scala 293:20]
      ghv_112 <= ghv_write_datas_112;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_113 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_113) begin // @[BPU.scala 293:20]
      ghv_113 <= ghv_write_datas_113;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_114 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_114) begin // @[BPU.scala 293:20]
      ghv_114 <= ghv_write_datas_114;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_115 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_115) begin // @[BPU.scala 293:20]
      ghv_115 <= ghv_write_datas_115;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_116 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_116) begin // @[BPU.scala 293:20]
      ghv_116 <= ghv_write_datas_116;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_117 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_117) begin // @[BPU.scala 293:20]
      ghv_117 <= ghv_write_datas_117;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_118 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_118) begin // @[BPU.scala 293:20]
      ghv_118 <= ghv_write_datas_118;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_119 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_119) begin // @[BPU.scala 293:20]
      ghv_119 <= ghv_write_datas_119;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_120 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_120) begin // @[BPU.scala 293:20]
      ghv_120 <= ghv_write_datas_120;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_121 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_121) begin // @[BPU.scala 293:20]
      ghv_121 <= ghv_write_datas_121;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_122 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_122) begin // @[BPU.scala 293:20]
      ghv_122 <= ghv_write_datas_122;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_123 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_123) begin // @[BPU.scala 293:20]
      ghv_123 <= ghv_write_datas_123;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_124 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_124) begin // @[BPU.scala 293:20]
      ghv_124 <= ghv_write_datas_124;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_125 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_125) begin // @[BPU.scala 293:20]
      ghv_125 <= ghv_write_datas_125;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_126 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_126) begin // @[BPU.scala 293:20]
      ghv_126 <= ghv_write_datas_126;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_127 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_127) begin // @[BPU.scala 293:20]
      ghv_127 <= ghv_write_datas_127;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_128 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_128) begin // @[BPU.scala 293:20]
      ghv_128 <= ghv_write_datas_128;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_129 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_129) begin // @[BPU.scala 293:20]
      ghv_129 <= ghv_write_datas_129;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_130 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_130) begin // @[BPU.scala 293:20]
      ghv_130 <= ghv_write_datas_130;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_131 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_131) begin // @[BPU.scala 293:20]
      ghv_131 <= ghv_write_datas_131;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_132 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_132) begin // @[BPU.scala 293:20]
      ghv_132 <= ghv_write_datas_132;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_133 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_133) begin // @[BPU.scala 293:20]
      ghv_133 <= ghv_write_datas_133;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_134 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_134) begin // @[BPU.scala 293:20]
      ghv_134 <= ghv_write_datas_134;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_135 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_135) begin // @[BPU.scala 293:20]
      ghv_135 <= ghv_write_datas_135;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_136 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_136) begin // @[BPU.scala 293:20]
      ghv_136 <= ghv_write_datas_136;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_137 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_137) begin // @[BPU.scala 293:20]
      ghv_137 <= ghv_write_datas_137;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_138 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_138) begin // @[BPU.scala 293:20]
      ghv_138 <= ghv_write_datas_138;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_139 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_139) begin // @[BPU.scala 293:20]
      ghv_139 <= ghv_write_datas_139;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_140 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_140) begin // @[BPU.scala 293:20]
      ghv_140 <= ghv_write_datas_140;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_141 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_141) begin // @[BPU.scala 293:20]
      ghv_141 <= ghv_write_datas_141;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_142 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_142) begin // @[BPU.scala 293:20]
      ghv_142 <= ghv_write_datas_142;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 675:24]
      ghv_143 <= 1'h0; // @[BPU.scala 676:14]
    end else if (ghv_wens_143) begin // @[BPU.scala 293:20]
      ghv_143 <= ghv_write_datas_143;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 303:26 669:17]
      s0_ghist_ptr_reg_flag <= 1'h0;
    end else begin
      s0_ghist_ptr_reg_flag <= s0_ghist_ptr_ppm_out_res_flag;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 303:26 669:17]
      s0_ghist_ptr_reg_value <= 8'h0;
    end else begin
      s0_ghist_ptr_reg_value <= s0_ghist_ptr_ppm_out_res_value;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s1_ghist_ptr_flag <= 1'h0; // @[Reg.scala 29:22]
    end else if (s0_fire) begin // @[Reg.scala 28:20]
      s1_ghist_ptr_flag <= s0_ghist_ptr_flag;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s1_ghist_ptr_value <= 8'h0; // @[Reg.scala 29:22]
    end else if (s0_fire) begin // @[Reg.scala 28:20]
      s1_ghist_ptr_value <= s0_ghist_ptr_value;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s2_ghist_ptr_flag <= 1'h0; // @[Reg.scala 29:22]
    end else if (s1_fire) begin // @[Reg.scala 28:20]
      s2_ghist_ptr_flag <= s1_ghist_ptr_flag;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s2_ghist_ptr_value <= 8'h0; // @[Reg.scala 29:22]
    end else if (s1_fire) begin // @[Reg.scala 28:20]
      s2_ghist_ptr_value <= s1_ghist_ptr_value;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s3_ghist_ptr_flag <= 1'h0; // @[Reg.scala 29:22]
    end else if (s2_valid) begin // @[Reg.scala 28:20]
      s3_ghist_ptr_flag <= s2_ghist_ptr_flag;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      s3_ghist_ptr_value <= 8'h0; // @[Reg.scala 29:22]
    end else if (s2_valid) begin // @[Reg.scala 28:20]
      s3_ghist_ptr_value <= s2_ghist_ptr_value;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 332:28]
      do_redirect_valid <= 1'h0; // @[BPU.scala 332:28]
    end else begin
      do_redirect_valid <= io_ftq_to_bpu_redirect_valid; // @[BPU.scala 332:28]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 332:28]
      do_redirect_bits_level <= 1'h0; // @[BPU.scala 332:28]
    end else begin
      do_redirect_bits_level <= io_ftq_to_bpu_redirect_bits_level; // @[BPU.scala 332:28]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 332:28]
      do_redirect_bits_cfiUpdate_pc <= 39'h0; // @[BPU.scala 332:28]
    end else begin
      do_redirect_bits_cfiUpdate_pc <= io_ftq_to_bpu_redirect_bits_cfiUpdate_pc; // @[BPU.scala 332:28]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 332:28]
      do_redirect_bits_cfiUpdate_pd_isRVC <= 1'h0; // @[BPU.scala 332:28]
    end else begin
      do_redirect_bits_cfiUpdate_pd_isRVC <= io_ftq_to_bpu_redirect_bits_cfiUpdate_pd_isRVC; // @[BPU.scala 332:28]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 332:28]
      do_redirect_bits_cfiUpdate_pd_isCall <= 1'h0; // @[BPU.scala 332:28]
    end else begin
      do_redirect_bits_cfiUpdate_pd_isCall <= io_ftq_to_bpu_redirect_bits_cfiUpdate_pd_isCall; // @[BPU.scala 332:28]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 332:28]
      do_redirect_bits_cfiUpdate_pd_isRet <= 1'h0; // @[BPU.scala 332:28]
    end else begin
      do_redirect_bits_cfiUpdate_pd_isRet <= io_ftq_to_bpu_redirect_bits_cfiUpdate_pd_isRet; // @[BPU.scala 332:28]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 332:28]
      do_redirect_bits_cfiUpdate_rasSp <= 5'h0; // @[BPU.scala 332:28]
    end else begin
      do_redirect_bits_cfiUpdate_rasSp <= io_ftq_to_bpu_redirect_bits_cfiUpdate_rasSp; // @[BPU.scala 332:28]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 332:28]
      do_redirect_bits_cfiUpdate_rasEntry_retAddr <= 39'h0; // @[BPU.scala 332:28]
    end else begin
      do_redirect_bits_cfiUpdate_rasEntry_retAddr <= io_ftq_to_bpu_redirect_bits_cfiUpdate_rasEntry_retAddr; // @[BPU.scala 332:28]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 332:28]
      do_redirect_bits_cfiUpdate_rasEntry_ctr <= 8'h0; // @[BPU.scala 332:28]
    end else begin
      do_redirect_bits_cfiUpdate_rasEntry_ctr <= io_ftq_to_bpu_redirect_bits_cfiUpdate_rasEntry_ctr; // @[BPU.scala 332:28]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 332:28]
      do_redirect_bits_cfiUpdate_folded_hist_hist_17_folded_hist <= 8'h0; // @[BPU.scala 332:28]
    end else begin
      do_redirect_bits_cfiUpdate_folded_hist_hist_17_folded_hist <=
        io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_17_folded_hist; // @[BPU.scala 332:28]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 332:28]
      do_redirect_bits_cfiUpdate_folded_hist_hist_16_folded_hist <= 8'h0; // @[BPU.scala 332:28]
    end else begin
      do_redirect_bits_cfiUpdate_folded_hist_hist_16_folded_hist <=
        io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_16_folded_hist; // @[BPU.scala 332:28]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 332:28]
      do_redirect_bits_cfiUpdate_folded_hist_hist_15_folded_hist <= 11'h0; // @[BPU.scala 332:28]
    end else begin
      do_redirect_bits_cfiUpdate_folded_hist_hist_15_folded_hist <=
        io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_15_folded_hist; // @[BPU.scala 332:28]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 332:28]
      do_redirect_bits_cfiUpdate_folded_hist_hist_14_folded_hist <= 7'h0; // @[BPU.scala 332:28]
    end else begin
      do_redirect_bits_cfiUpdate_folded_hist_hist_14_folded_hist <=
        io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_14_folded_hist; // @[BPU.scala 332:28]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 332:28]
      do_redirect_bits_cfiUpdate_folded_hist_hist_13_folded_hist <= 7'h0; // @[BPU.scala 332:28]
    end else begin
      do_redirect_bits_cfiUpdate_folded_hist_hist_13_folded_hist <=
        io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_13_folded_hist; // @[BPU.scala 332:28]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 332:28]
      do_redirect_bits_cfiUpdate_folded_hist_hist_12_folded_hist <= 7'h0; // @[BPU.scala 332:28]
    end else begin
      do_redirect_bits_cfiUpdate_folded_hist_hist_12_folded_hist <=
        io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_12_folded_hist; // @[BPU.scala 332:28]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 332:28]
      do_redirect_bits_cfiUpdate_folded_hist_hist_11_folded_hist <= 8'h0; // @[BPU.scala 332:28]
    end else begin
      do_redirect_bits_cfiUpdate_folded_hist_hist_11_folded_hist <=
        io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_11_folded_hist; // @[BPU.scala 332:28]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 332:28]
      do_redirect_bits_cfiUpdate_folded_hist_hist_10_folded_hist <= 9'h0; // @[BPU.scala 332:28]
    end else begin
      do_redirect_bits_cfiUpdate_folded_hist_hist_10_folded_hist <=
        io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_10_folded_hist; // @[BPU.scala 332:28]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 332:28]
      do_redirect_bits_cfiUpdate_folded_hist_hist_9_folded_hist <= 7'h0; // @[BPU.scala 332:28]
    end else begin
      do_redirect_bits_cfiUpdate_folded_hist_hist_9_folded_hist <=
        io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_9_folded_hist; // @[BPU.scala 332:28]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 332:28]
      do_redirect_bits_cfiUpdate_folded_hist_hist_8_folded_hist <= 8'h0; // @[BPU.scala 332:28]
    end else begin
      do_redirect_bits_cfiUpdate_folded_hist_hist_8_folded_hist <=
        io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_8_folded_hist; // @[BPU.scala 332:28]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 332:28]
      do_redirect_bits_cfiUpdate_folded_hist_hist_7_folded_hist <= 9'h0; // @[BPU.scala 332:28]
    end else begin
      do_redirect_bits_cfiUpdate_folded_hist_hist_7_folded_hist <=
        io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_7_folded_hist; // @[BPU.scala 332:28]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 332:28]
      do_redirect_bits_cfiUpdate_folded_hist_hist_6_folded_hist <= 9'h0; // @[BPU.scala 332:28]
    end else begin
      do_redirect_bits_cfiUpdate_folded_hist_hist_6_folded_hist <=
        io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_6_folded_hist; // @[BPU.scala 332:28]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 332:28]
      do_redirect_bits_cfiUpdate_folded_hist_hist_5_folded_hist <= 11'h0; // @[BPU.scala 332:28]
    end else begin
      do_redirect_bits_cfiUpdate_folded_hist_hist_5_folded_hist <=
        io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_5_folded_hist; // @[BPU.scala 332:28]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 332:28]
      do_redirect_bits_cfiUpdate_folded_hist_hist_4_folded_hist <= 4'h0; // @[BPU.scala 332:28]
    end else begin
      do_redirect_bits_cfiUpdate_folded_hist_hist_4_folded_hist <=
        io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_4_folded_hist; // @[BPU.scala 332:28]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 332:28]
      do_redirect_bits_cfiUpdate_folded_hist_hist_3_folded_hist <= 11'h0; // @[BPU.scala 332:28]
    end else begin
      do_redirect_bits_cfiUpdate_folded_hist_hist_3_folded_hist <=
        io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_3_folded_hist; // @[BPU.scala 332:28]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 332:28]
      do_redirect_bits_cfiUpdate_folded_hist_hist_2_folded_hist <= 8'h0; // @[BPU.scala 332:28]
    end else begin
      do_redirect_bits_cfiUpdate_folded_hist_hist_2_folded_hist <=
        io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_2_folded_hist; // @[BPU.scala 332:28]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 332:28]
      do_redirect_bits_cfiUpdate_folded_hist_hist_1_folded_hist <= 8'h0; // @[BPU.scala 332:28]
    end else begin
      do_redirect_bits_cfiUpdate_folded_hist_hist_1_folded_hist <=
        io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_1_folded_hist; // @[BPU.scala 332:28]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 332:28]
      do_redirect_bits_cfiUpdate_folded_hist_hist_0_folded_hist <= 8'h0; // @[BPU.scala 332:28]
    end else begin
      do_redirect_bits_cfiUpdate_folded_hist_hist_0_folded_hist <=
        io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_0_folded_hist; // @[BPU.scala 332:28]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 332:28]
      do_redirect_bits_cfiUpdate_afhob_afhob_5_bits_0 <= 1'h0; // @[BPU.scala 332:28]
    end else begin
      do_redirect_bits_cfiUpdate_afhob_afhob_5_bits_0 <= io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_5_bits_0; // @[BPU.scala 332:28]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 332:28]
      do_redirect_bits_cfiUpdate_afhob_afhob_5_bits_1 <= 1'h0; // @[BPU.scala 332:28]
    end else begin
      do_redirect_bits_cfiUpdate_afhob_afhob_5_bits_1 <= io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_5_bits_1; // @[BPU.scala 332:28]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 332:28]
      do_redirect_bits_cfiUpdate_afhob_afhob_5_bits_2 <= 1'h0; // @[BPU.scala 332:28]
    end else begin
      do_redirect_bits_cfiUpdate_afhob_afhob_5_bits_2 <= io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_5_bits_2; // @[BPU.scala 332:28]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 332:28]
      do_redirect_bits_cfiUpdate_afhob_afhob_5_bits_3 <= 1'h0; // @[BPU.scala 332:28]
    end else begin
      do_redirect_bits_cfiUpdate_afhob_afhob_5_bits_3 <= io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_5_bits_3; // @[BPU.scala 332:28]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 332:28]
      do_redirect_bits_cfiUpdate_afhob_afhob_4_bits_0 <= 1'h0; // @[BPU.scala 332:28]
    end else begin
      do_redirect_bits_cfiUpdate_afhob_afhob_4_bits_0 <= io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_4_bits_0; // @[BPU.scala 332:28]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 332:28]
      do_redirect_bits_cfiUpdate_afhob_afhob_4_bits_1 <= 1'h0; // @[BPU.scala 332:28]
    end else begin
      do_redirect_bits_cfiUpdate_afhob_afhob_4_bits_1 <= io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_4_bits_1; // @[BPU.scala 332:28]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 332:28]
      do_redirect_bits_cfiUpdate_afhob_afhob_4_bits_2 <= 1'h0; // @[BPU.scala 332:28]
    end else begin
      do_redirect_bits_cfiUpdate_afhob_afhob_4_bits_2 <= io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_4_bits_2; // @[BPU.scala 332:28]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 332:28]
      do_redirect_bits_cfiUpdate_afhob_afhob_3_bits_0 <= 1'h0; // @[BPU.scala 332:28]
    end else begin
      do_redirect_bits_cfiUpdate_afhob_afhob_3_bits_0 <= io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_3_bits_0; // @[BPU.scala 332:28]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 332:28]
      do_redirect_bits_cfiUpdate_afhob_afhob_3_bits_1 <= 1'h0; // @[BPU.scala 332:28]
    end else begin
      do_redirect_bits_cfiUpdate_afhob_afhob_3_bits_1 <= io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_3_bits_1; // @[BPU.scala 332:28]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 332:28]
      do_redirect_bits_cfiUpdate_afhob_afhob_3_bits_2 <= 1'h0; // @[BPU.scala 332:28]
    end else begin
      do_redirect_bits_cfiUpdate_afhob_afhob_3_bits_2 <= io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_3_bits_2; // @[BPU.scala 332:28]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 332:28]
      do_redirect_bits_cfiUpdate_afhob_afhob_3_bits_3 <= 1'h0; // @[BPU.scala 332:28]
    end else begin
      do_redirect_bits_cfiUpdate_afhob_afhob_3_bits_3 <= io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_3_bits_3; // @[BPU.scala 332:28]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 332:28]
      do_redirect_bits_cfiUpdate_afhob_afhob_2_bits_0 <= 1'h0; // @[BPU.scala 332:28]
    end else begin
      do_redirect_bits_cfiUpdate_afhob_afhob_2_bits_0 <= io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_2_bits_0; // @[BPU.scala 332:28]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 332:28]
      do_redirect_bits_cfiUpdate_afhob_afhob_2_bits_1 <= 1'h0; // @[BPU.scala 332:28]
    end else begin
      do_redirect_bits_cfiUpdate_afhob_afhob_2_bits_1 <= io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_2_bits_1; // @[BPU.scala 332:28]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 332:28]
      do_redirect_bits_cfiUpdate_afhob_afhob_2_bits_2 <= 1'h0; // @[BPU.scala 332:28]
    end else begin
      do_redirect_bits_cfiUpdate_afhob_afhob_2_bits_2 <= io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_2_bits_2; // @[BPU.scala 332:28]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 332:28]
      do_redirect_bits_cfiUpdate_afhob_afhob_2_bits_3 <= 1'h0; // @[BPU.scala 332:28]
    end else begin
      do_redirect_bits_cfiUpdate_afhob_afhob_2_bits_3 <= io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_2_bits_3; // @[BPU.scala 332:28]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 332:28]
      do_redirect_bits_cfiUpdate_afhob_afhob_1_bits_0 <= 1'h0; // @[BPU.scala 332:28]
    end else begin
      do_redirect_bits_cfiUpdate_afhob_afhob_1_bits_0 <= io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_1_bits_0; // @[BPU.scala 332:28]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 332:28]
      do_redirect_bits_cfiUpdate_afhob_afhob_1_bits_1 <= 1'h0; // @[BPU.scala 332:28]
    end else begin
      do_redirect_bits_cfiUpdate_afhob_afhob_1_bits_1 <= io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_1_bits_1; // @[BPU.scala 332:28]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 332:28]
      do_redirect_bits_cfiUpdate_afhob_afhob_1_bits_2 <= 1'h0; // @[BPU.scala 332:28]
    end else begin
      do_redirect_bits_cfiUpdate_afhob_afhob_1_bits_2 <= io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_1_bits_2; // @[BPU.scala 332:28]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 332:28]
      do_redirect_bits_cfiUpdate_afhob_afhob_1_bits_3 <= 1'h0; // @[BPU.scala 332:28]
    end else begin
      do_redirect_bits_cfiUpdate_afhob_afhob_1_bits_3 <= io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_1_bits_3; // @[BPU.scala 332:28]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 332:28]
      do_redirect_bits_cfiUpdate_afhob_afhob_0_bits_0 <= 1'h0; // @[BPU.scala 332:28]
    end else begin
      do_redirect_bits_cfiUpdate_afhob_afhob_0_bits_0 <= io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_0_bits_0; // @[BPU.scala 332:28]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 332:28]
      do_redirect_bits_cfiUpdate_afhob_afhob_0_bits_1 <= 1'h0; // @[BPU.scala 332:28]
    end else begin
      do_redirect_bits_cfiUpdate_afhob_afhob_0_bits_1 <= io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_0_bits_1; // @[BPU.scala 332:28]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 332:28]
      do_redirect_bits_cfiUpdate_afhob_afhob_0_bits_2 <= 1'h0; // @[BPU.scala 332:28]
    end else begin
      do_redirect_bits_cfiUpdate_afhob_afhob_0_bits_2 <= io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_0_bits_2; // @[BPU.scala 332:28]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 332:28]
      do_redirect_bits_cfiUpdate_afhob_afhob_0_bits_3 <= 1'h0; // @[BPU.scala 332:28]
    end else begin
      do_redirect_bits_cfiUpdate_afhob_afhob_0_bits_3 <= io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_0_bits_3; // @[BPU.scala 332:28]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 332:28]
      do_redirect_bits_cfiUpdate_lastBrNumOH <= 3'h0; // @[BPU.scala 332:28]
    end else begin
      do_redirect_bits_cfiUpdate_lastBrNumOH <= io_ftq_to_bpu_redirect_bits_cfiUpdate_lastBrNumOH; // @[BPU.scala 332:28]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 332:28]
      do_redirect_bits_cfiUpdate_histPtr_flag <= 1'h0; // @[BPU.scala 332:28]
    end else begin
      do_redirect_bits_cfiUpdate_histPtr_flag <= io_ftq_to_bpu_redirect_bits_cfiUpdate_histPtr_flag; // @[BPU.scala 332:28]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 332:28]
      do_redirect_bits_cfiUpdate_histPtr_value <= 8'h0; // @[BPU.scala 332:28]
    end else begin
      do_redirect_bits_cfiUpdate_histPtr_value <= io_ftq_to_bpu_redirect_bits_cfiUpdate_histPtr_value; // @[BPU.scala 332:28]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 332:28]
      do_redirect_bits_cfiUpdate_target <= 39'h0; // @[BPU.scala 332:28]
    end else begin
      do_redirect_bits_cfiUpdate_target <= io_ftq_to_bpu_redirect_bits_cfiUpdate_target; // @[BPU.scala 332:28]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 332:28]
      do_redirect_bits_cfiUpdate_taken <= 1'h0; // @[BPU.scala 332:28]
    end else begin
      do_redirect_bits_cfiUpdate_taken <= io_ftq_to_bpu_redirect_bits_cfiUpdate_taken; // @[BPU.scala 332:28]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 332:28]
      do_redirect_bits_cfiUpdate_shift <= 2'h0; // @[BPU.scala 332:28]
    end else begin
      do_redirect_bits_cfiUpdate_shift <= io_ftq_to_bpu_redirect_bits_cfiUpdate_shift; // @[BPU.scala 332:28]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BPU.scala 332:28]
      do_redirect_bits_cfiUpdate_addIntoHist <= 1'h0; // @[BPU.scala 332:28]
    end else begin
      do_redirect_bits_cfiUpdate_addIntoHist <= io_ftq_to_bpu_redirect_bits_cfiUpdate_addIntoHist; // @[BPU.scala 332:28]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      previous_s2_pred_full_pred_br_taken_mask_1 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s2_valid) begin // @[Reg.scala 28:20]
      previous_s2_pred_full_pred_br_taken_mask_1 <= predictors_io_out_s2_full_pred_br_taken_mask_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      previous_s2_pred_full_pred_slot_valids_1 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s2_valid) begin // @[Reg.scala 28:20]
      previous_s2_pred_full_pred_slot_valids_1 <= predictors_io_out_s2_full_pred_slot_valids_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      previous_s2_pred_full_pred_is_br_sharing <= 1'h0; // @[Reg.scala 29:22]
    end else if (s2_valid) begin // @[Reg.scala 28:20]
      previous_s2_pred_full_pred_is_br_sharing <= predictors_io_out_s2_full_pred_is_br_sharing;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      previous_s2_pred_full_pred_hit <= 1'h0; // @[Reg.scala 29:22]
    end else if (s2_valid) begin // @[Reg.scala 28:20]
      previous_s2_pred_full_pred_hit <= predictors_io_out_s2_full_pred_hit;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      previous_s2_pred_full_pred_slot_valids_0 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s2_valid) begin // @[Reg.scala 28:20]
      previous_s2_pred_full_pred_slot_valids_0 <= predictors_io_out_s2_full_pred_slot_valids_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      previous_s2_pred_full_pred_br_taken_mask_0 <= 1'h0; // @[Reg.scala 29:22]
    end else if (s2_valid) begin // @[Reg.scala 28:20]
      previous_s2_pred_full_pred_br_taken_mask_0 <= predictors_io_out_s2_full_pred_br_taken_mask_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      previous_s2_pred_full_pred_targets_0 <= 39'h0; // @[Reg.scala 29:22]
    end else if (s2_valid) begin // @[Reg.scala 28:20]
      previous_s2_pred_full_pred_targets_0 <= predictors_io_out_s2_full_pred_targets_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      previous_s2_pred_full_pred_targets_1 <= 39'h0; // @[Reg.scala 29:22]
    end else if (s2_valid) begin // @[Reg.scala 28:20]
      previous_s2_pred_full_pred_targets_1 <= predictors_io_out_s2_full_pred_targets_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      previous_s2_pred_full_pred_fallThroughAddr <= 39'h0; // @[Reg.scala 29:22]
    end else if (s2_valid) begin // @[Reg.scala 28:20]
      previous_s2_pred_full_pred_fallThroughAddr <= predictors_io_out_s2_full_pred_fallThroughAddr;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      previous_s2_pred_pc <= 39'h0; // @[Reg.scala 29:22]
    end else if (s2_valid) begin // @[Reg.scala 28:20]
      previous_s2_pred_pc <= predictors_io_out_s2_pc;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      previous_s1_pred_info_target <= 39'h0; // @[Reg.scala 29:22]
    end else if (s1_fire) begin // @[Reg.scala 28:20]
      previous_s1_pred_info_target <= _T_60;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      previous_s1_pred_info_lastBrPosOH <= 3'h0; // @[Reg.scala 29:22]
    end else if (s1_fire) begin // @[Reg.scala 28:20]
      previous_s1_pred_info_lastBrPosOH <= _T_122;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      previous_s1_pred_info_taken <= 1'h0; // @[Reg.scala 29:22]
    end else if (s1_fire) begin // @[Reg.scala 28:20]
      previous_s1_pred_info_taken <= cfiIndex_valid;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      previous_s1_pred_info_cfiIndex <= 3'h0; // @[Reg.scala 29:22]
    end else if (s1_fire) begin // @[Reg.scala 28:20]
      previous_s1_pred_info_cfiIndex <= cfiIndex_bits;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  s1_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  s2_valid = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  s3_valid = _RAND_2[0:0];
  _RAND_3 = {2{`RANDOM}};
  s0_pc_reg = _RAND_3[38:0];
  _RAND_4 = {1{`RANDOM}};
  REG = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  REG_1 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  s0_folded_gh_reg_hist_17_folded_hist = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  s0_folded_gh_reg_hist_16_folded_hist = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  s0_folded_gh_reg_hist_15_folded_hist = _RAND_8[10:0];
  _RAND_9 = {1{`RANDOM}};
  s0_folded_gh_reg_hist_14_folded_hist = _RAND_9[6:0];
  _RAND_10 = {1{`RANDOM}};
  s0_folded_gh_reg_hist_13_folded_hist = _RAND_10[6:0];
  _RAND_11 = {1{`RANDOM}};
  s0_folded_gh_reg_hist_12_folded_hist = _RAND_11[6:0];
  _RAND_12 = {1{`RANDOM}};
  s0_folded_gh_reg_hist_11_folded_hist = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  s0_folded_gh_reg_hist_10_folded_hist = _RAND_13[8:0];
  _RAND_14 = {1{`RANDOM}};
  s0_folded_gh_reg_hist_9_folded_hist = _RAND_14[6:0];
  _RAND_15 = {1{`RANDOM}};
  s0_folded_gh_reg_hist_8_folded_hist = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  s0_folded_gh_reg_hist_7_folded_hist = _RAND_16[8:0];
  _RAND_17 = {1{`RANDOM}};
  s0_folded_gh_reg_hist_6_folded_hist = _RAND_17[8:0];
  _RAND_18 = {1{`RANDOM}};
  s0_folded_gh_reg_hist_5_folded_hist = _RAND_18[10:0];
  _RAND_19 = {1{`RANDOM}};
  s0_folded_gh_reg_hist_4_folded_hist = _RAND_19[3:0];
  _RAND_20 = {1{`RANDOM}};
  s0_folded_gh_reg_hist_3_folded_hist = _RAND_20[10:0];
  _RAND_21 = {1{`RANDOM}};
  s0_folded_gh_reg_hist_2_folded_hist = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  s0_folded_gh_reg_hist_1_folded_hist = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  s0_folded_gh_reg_hist_0_folded_hist = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  s1_folded_gh_hist_17_folded_hist = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  s1_folded_gh_hist_16_folded_hist = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  s1_folded_gh_hist_15_folded_hist = _RAND_26[10:0];
  _RAND_27 = {1{`RANDOM}};
  s1_folded_gh_hist_14_folded_hist = _RAND_27[6:0];
  _RAND_28 = {1{`RANDOM}};
  s1_folded_gh_hist_13_folded_hist = _RAND_28[6:0];
  _RAND_29 = {1{`RANDOM}};
  s1_folded_gh_hist_12_folded_hist = _RAND_29[6:0];
  _RAND_30 = {1{`RANDOM}};
  s1_folded_gh_hist_11_folded_hist = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  s1_folded_gh_hist_10_folded_hist = _RAND_31[8:0];
  _RAND_32 = {1{`RANDOM}};
  s1_folded_gh_hist_9_folded_hist = _RAND_32[6:0];
  _RAND_33 = {1{`RANDOM}};
  s1_folded_gh_hist_8_folded_hist = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  s1_folded_gh_hist_7_folded_hist = _RAND_34[8:0];
  _RAND_35 = {1{`RANDOM}};
  s1_folded_gh_hist_6_folded_hist = _RAND_35[8:0];
  _RAND_36 = {1{`RANDOM}};
  s1_folded_gh_hist_5_folded_hist = _RAND_36[10:0];
  _RAND_37 = {1{`RANDOM}};
  s1_folded_gh_hist_4_folded_hist = _RAND_37[3:0];
  _RAND_38 = {1{`RANDOM}};
  s1_folded_gh_hist_3_folded_hist = _RAND_38[10:0];
  _RAND_39 = {1{`RANDOM}};
  s1_folded_gh_hist_2_folded_hist = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  s1_folded_gh_hist_1_folded_hist = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  s1_folded_gh_hist_0_folded_hist = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  s2_folded_gh_hist_17_folded_hist = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  s2_folded_gh_hist_16_folded_hist = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  s2_folded_gh_hist_15_folded_hist = _RAND_44[10:0];
  _RAND_45 = {1{`RANDOM}};
  s2_folded_gh_hist_14_folded_hist = _RAND_45[6:0];
  _RAND_46 = {1{`RANDOM}};
  s2_folded_gh_hist_13_folded_hist = _RAND_46[6:0];
  _RAND_47 = {1{`RANDOM}};
  s2_folded_gh_hist_12_folded_hist = _RAND_47[6:0];
  _RAND_48 = {1{`RANDOM}};
  s2_folded_gh_hist_11_folded_hist = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  s2_folded_gh_hist_10_folded_hist = _RAND_49[8:0];
  _RAND_50 = {1{`RANDOM}};
  s2_folded_gh_hist_9_folded_hist = _RAND_50[6:0];
  _RAND_51 = {1{`RANDOM}};
  s2_folded_gh_hist_8_folded_hist = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  s2_folded_gh_hist_7_folded_hist = _RAND_52[8:0];
  _RAND_53 = {1{`RANDOM}};
  s2_folded_gh_hist_6_folded_hist = _RAND_53[8:0];
  _RAND_54 = {1{`RANDOM}};
  s2_folded_gh_hist_5_folded_hist = _RAND_54[10:0];
  _RAND_55 = {1{`RANDOM}};
  s2_folded_gh_hist_4_folded_hist = _RAND_55[3:0];
  _RAND_56 = {1{`RANDOM}};
  s2_folded_gh_hist_3_folded_hist = _RAND_56[10:0];
  _RAND_57 = {1{`RANDOM}};
  s2_folded_gh_hist_2_folded_hist = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  s2_folded_gh_hist_1_folded_hist = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  s2_folded_gh_hist_0_folded_hist = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  s3_folded_gh_hist_17_folded_hist = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  s3_folded_gh_hist_16_folded_hist = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  s3_folded_gh_hist_15_folded_hist = _RAND_62[10:0];
  _RAND_63 = {1{`RANDOM}};
  s3_folded_gh_hist_14_folded_hist = _RAND_63[6:0];
  _RAND_64 = {1{`RANDOM}};
  s3_folded_gh_hist_13_folded_hist = _RAND_64[6:0];
  _RAND_65 = {1{`RANDOM}};
  s3_folded_gh_hist_12_folded_hist = _RAND_65[6:0];
  _RAND_66 = {1{`RANDOM}};
  s3_folded_gh_hist_11_folded_hist = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  s3_folded_gh_hist_10_folded_hist = _RAND_67[8:0];
  _RAND_68 = {1{`RANDOM}};
  s3_folded_gh_hist_9_folded_hist = _RAND_68[6:0];
  _RAND_69 = {1{`RANDOM}};
  s3_folded_gh_hist_8_folded_hist = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  s3_folded_gh_hist_7_folded_hist = _RAND_70[8:0];
  _RAND_71 = {1{`RANDOM}};
  s3_folded_gh_hist_6_folded_hist = _RAND_71[8:0];
  _RAND_72 = {1{`RANDOM}};
  s3_folded_gh_hist_5_folded_hist = _RAND_72[10:0];
  _RAND_73 = {1{`RANDOM}};
  s3_folded_gh_hist_4_folded_hist = _RAND_73[3:0];
  _RAND_74 = {1{`RANDOM}};
  s3_folded_gh_hist_3_folded_hist = _RAND_74[10:0];
  _RAND_75 = {1{`RANDOM}};
  s3_folded_gh_hist_2_folded_hist = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  s3_folded_gh_hist_1_folded_hist = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  s3_folded_gh_hist_0_folded_hist = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  s0_last_br_num_oh_reg = _RAND_78[2:0];
  _RAND_79 = {1{`RANDOM}};
  s1_last_br_num_oh = _RAND_79[2:0];
  _RAND_80 = {1{`RANDOM}};
  s2_last_br_num_oh = _RAND_80[2:0];
  _RAND_81 = {1{`RANDOM}};
  s3_last_br_num_oh = _RAND_81[2:0];
  _RAND_82 = {1{`RANDOM}};
  s0_ahead_fh_oldest_bits_reg_afhob_5_bits_0 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  s0_ahead_fh_oldest_bits_reg_afhob_5_bits_1 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  s0_ahead_fh_oldest_bits_reg_afhob_5_bits_2 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  s0_ahead_fh_oldest_bits_reg_afhob_5_bits_3 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  s0_ahead_fh_oldest_bits_reg_afhob_4_bits_0 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  s0_ahead_fh_oldest_bits_reg_afhob_4_bits_1 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  s0_ahead_fh_oldest_bits_reg_afhob_4_bits_2 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  s0_ahead_fh_oldest_bits_reg_afhob_4_bits_3 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  s0_ahead_fh_oldest_bits_reg_afhob_3_bits_0 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  s0_ahead_fh_oldest_bits_reg_afhob_3_bits_1 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  s0_ahead_fh_oldest_bits_reg_afhob_3_bits_2 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  s0_ahead_fh_oldest_bits_reg_afhob_3_bits_3 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  s0_ahead_fh_oldest_bits_reg_afhob_2_bits_0 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  s0_ahead_fh_oldest_bits_reg_afhob_2_bits_1 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  s0_ahead_fh_oldest_bits_reg_afhob_2_bits_2 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  s0_ahead_fh_oldest_bits_reg_afhob_2_bits_3 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  s0_ahead_fh_oldest_bits_reg_afhob_1_bits_0 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  s0_ahead_fh_oldest_bits_reg_afhob_1_bits_1 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  s0_ahead_fh_oldest_bits_reg_afhob_1_bits_2 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  s0_ahead_fh_oldest_bits_reg_afhob_1_bits_3 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  s0_ahead_fh_oldest_bits_reg_afhob_0_bits_0 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  s0_ahead_fh_oldest_bits_reg_afhob_0_bits_1 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  s0_ahead_fh_oldest_bits_reg_afhob_0_bits_2 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  s0_ahead_fh_oldest_bits_reg_afhob_0_bits_3 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  s1_ahead_fh_oldest_bits_afhob_5_bits_0 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  s1_ahead_fh_oldest_bits_afhob_5_bits_1 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  s1_ahead_fh_oldest_bits_afhob_5_bits_2 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  s1_ahead_fh_oldest_bits_afhob_5_bits_3 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  s1_ahead_fh_oldest_bits_afhob_4_bits_0 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  s1_ahead_fh_oldest_bits_afhob_4_bits_1 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  s1_ahead_fh_oldest_bits_afhob_4_bits_2 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  s1_ahead_fh_oldest_bits_afhob_4_bits_3 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  s1_ahead_fh_oldest_bits_afhob_3_bits_0 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  s1_ahead_fh_oldest_bits_afhob_3_bits_1 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  s1_ahead_fh_oldest_bits_afhob_3_bits_2 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  s1_ahead_fh_oldest_bits_afhob_3_bits_3 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  s1_ahead_fh_oldest_bits_afhob_2_bits_0 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  s1_ahead_fh_oldest_bits_afhob_2_bits_1 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  s1_ahead_fh_oldest_bits_afhob_2_bits_2 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  s1_ahead_fh_oldest_bits_afhob_2_bits_3 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  s1_ahead_fh_oldest_bits_afhob_1_bits_0 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  s1_ahead_fh_oldest_bits_afhob_1_bits_1 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  s1_ahead_fh_oldest_bits_afhob_1_bits_2 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  s1_ahead_fh_oldest_bits_afhob_1_bits_3 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  s1_ahead_fh_oldest_bits_afhob_0_bits_0 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  s1_ahead_fh_oldest_bits_afhob_0_bits_1 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  s1_ahead_fh_oldest_bits_afhob_0_bits_2 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  s1_ahead_fh_oldest_bits_afhob_0_bits_3 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  s2_ahead_fh_oldest_bits_afhob_5_bits_0 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  s2_ahead_fh_oldest_bits_afhob_5_bits_1 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  s2_ahead_fh_oldest_bits_afhob_5_bits_2 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  s2_ahead_fh_oldest_bits_afhob_5_bits_3 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  s2_ahead_fh_oldest_bits_afhob_4_bits_0 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  s2_ahead_fh_oldest_bits_afhob_4_bits_1 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  s2_ahead_fh_oldest_bits_afhob_4_bits_2 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  s2_ahead_fh_oldest_bits_afhob_4_bits_3 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  s2_ahead_fh_oldest_bits_afhob_3_bits_0 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  s2_ahead_fh_oldest_bits_afhob_3_bits_1 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  s2_ahead_fh_oldest_bits_afhob_3_bits_2 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  s2_ahead_fh_oldest_bits_afhob_3_bits_3 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  s2_ahead_fh_oldest_bits_afhob_2_bits_0 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  s2_ahead_fh_oldest_bits_afhob_2_bits_1 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  s2_ahead_fh_oldest_bits_afhob_2_bits_2 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  s2_ahead_fh_oldest_bits_afhob_2_bits_3 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  s2_ahead_fh_oldest_bits_afhob_1_bits_0 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  s2_ahead_fh_oldest_bits_afhob_1_bits_1 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  s2_ahead_fh_oldest_bits_afhob_1_bits_2 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  s2_ahead_fh_oldest_bits_afhob_1_bits_3 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  s2_ahead_fh_oldest_bits_afhob_0_bits_0 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  s2_ahead_fh_oldest_bits_afhob_0_bits_1 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  s2_ahead_fh_oldest_bits_afhob_0_bits_2 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  s2_ahead_fh_oldest_bits_afhob_0_bits_3 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  s3_ahead_fh_oldest_bits_afhob_5_bits_0 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  s3_ahead_fh_oldest_bits_afhob_5_bits_1 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  s3_ahead_fh_oldest_bits_afhob_5_bits_2 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  s3_ahead_fh_oldest_bits_afhob_5_bits_3 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  s3_ahead_fh_oldest_bits_afhob_4_bits_0 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  s3_ahead_fh_oldest_bits_afhob_4_bits_1 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  s3_ahead_fh_oldest_bits_afhob_4_bits_2 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  s3_ahead_fh_oldest_bits_afhob_4_bits_3 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  s3_ahead_fh_oldest_bits_afhob_3_bits_0 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  s3_ahead_fh_oldest_bits_afhob_3_bits_1 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  s3_ahead_fh_oldest_bits_afhob_3_bits_2 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  s3_ahead_fh_oldest_bits_afhob_3_bits_3 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  s3_ahead_fh_oldest_bits_afhob_2_bits_0 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  s3_ahead_fh_oldest_bits_afhob_2_bits_1 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  s3_ahead_fh_oldest_bits_afhob_2_bits_2 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  s3_ahead_fh_oldest_bits_afhob_2_bits_3 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  s3_ahead_fh_oldest_bits_afhob_1_bits_0 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  s3_ahead_fh_oldest_bits_afhob_1_bits_1 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  s3_ahead_fh_oldest_bits_afhob_1_bits_2 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  s3_ahead_fh_oldest_bits_afhob_1_bits_3 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  s3_ahead_fh_oldest_bits_afhob_0_bits_0 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  s3_ahead_fh_oldest_bits_afhob_0_bits_1 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  s3_ahead_fh_oldest_bits_afhob_0_bits_2 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  s3_ahead_fh_oldest_bits_afhob_0_bits_3 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  ghv_0 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  ghv_1 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  ghv_2 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  ghv_3 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  ghv_4 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  ghv_5 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  ghv_6 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  ghv_7 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  ghv_8 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  ghv_9 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  ghv_10 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  ghv_11 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  ghv_12 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  ghv_13 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  ghv_14 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  ghv_15 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  ghv_16 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  ghv_17 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  ghv_18 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  ghv_19 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  ghv_20 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  ghv_21 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  ghv_22 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  ghv_23 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  ghv_24 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  ghv_25 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  ghv_26 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  ghv_27 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  ghv_28 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  ghv_29 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  ghv_30 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  ghv_31 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  ghv_32 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  ghv_33 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  ghv_34 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  ghv_35 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  ghv_36 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  ghv_37 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  ghv_38 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  ghv_39 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  ghv_40 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  ghv_41 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  ghv_42 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  ghv_43 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  ghv_44 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  ghv_45 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  ghv_46 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  ghv_47 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  ghv_48 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  ghv_49 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  ghv_50 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  ghv_51 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  ghv_52 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  ghv_53 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  ghv_54 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  ghv_55 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  ghv_56 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  ghv_57 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  ghv_58 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  ghv_59 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  ghv_60 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  ghv_61 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  ghv_62 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  ghv_63 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  ghv_64 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  ghv_65 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  ghv_66 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  ghv_67 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  ghv_68 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  ghv_69 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  ghv_70 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  ghv_71 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  ghv_72 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  ghv_73 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  ghv_74 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  ghv_75 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  ghv_76 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  ghv_77 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  ghv_78 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  ghv_79 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  ghv_80 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  ghv_81 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  ghv_82 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  ghv_83 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  ghv_84 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  ghv_85 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  ghv_86 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  ghv_87 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  ghv_88 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  ghv_89 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  ghv_90 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  ghv_91 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  ghv_92 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  ghv_93 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  ghv_94 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  ghv_95 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  ghv_96 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  ghv_97 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  ghv_98 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  ghv_99 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  ghv_100 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  ghv_101 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  ghv_102 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  ghv_103 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  ghv_104 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  ghv_105 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  ghv_106 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  ghv_107 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  ghv_108 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  ghv_109 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  ghv_110 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  ghv_111 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  ghv_112 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  ghv_113 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  ghv_114 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  ghv_115 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  ghv_116 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  ghv_117 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  ghv_118 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  ghv_119 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  ghv_120 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  ghv_121 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  ghv_122 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  ghv_123 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  ghv_124 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  ghv_125 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  ghv_126 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  ghv_127 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  ghv_128 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  ghv_129 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  ghv_130 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  ghv_131 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  ghv_132 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  ghv_133 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  ghv_134 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  ghv_135 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  ghv_136 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  ghv_137 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  ghv_138 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  ghv_139 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  ghv_140 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  ghv_141 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  ghv_142 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  ghv_143 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  s0_ghist_ptr_reg_flag = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  s0_ghist_ptr_reg_value = _RAND_323[7:0];
  _RAND_324 = {1{`RANDOM}};
  s1_ghist_ptr_flag = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  s1_ghist_ptr_value = _RAND_325[7:0];
  _RAND_326 = {1{`RANDOM}};
  s2_ghist_ptr_flag = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  s2_ghist_ptr_value = _RAND_327[7:0];
  _RAND_328 = {1{`RANDOM}};
  s3_ghist_ptr_flag = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  s3_ghist_ptr_value = _RAND_329[7:0];
  _RAND_330 = {1{`RANDOM}};
  do_redirect_valid = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  do_redirect_bits_level = _RAND_331[0:0];
  _RAND_332 = {2{`RANDOM}};
  do_redirect_bits_cfiUpdate_pc = _RAND_332[38:0];
  _RAND_333 = {1{`RANDOM}};
  do_redirect_bits_cfiUpdate_pd_isRVC = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  do_redirect_bits_cfiUpdate_pd_isCall = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  do_redirect_bits_cfiUpdate_pd_isRet = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  do_redirect_bits_cfiUpdate_rasSp = _RAND_336[4:0];
  _RAND_337 = {2{`RANDOM}};
  do_redirect_bits_cfiUpdate_rasEntry_retAddr = _RAND_337[38:0];
  _RAND_338 = {1{`RANDOM}};
  do_redirect_bits_cfiUpdate_rasEntry_ctr = _RAND_338[7:0];
  _RAND_339 = {1{`RANDOM}};
  do_redirect_bits_cfiUpdate_folded_hist_hist_17_folded_hist = _RAND_339[7:0];
  _RAND_340 = {1{`RANDOM}};
  do_redirect_bits_cfiUpdate_folded_hist_hist_16_folded_hist = _RAND_340[7:0];
  _RAND_341 = {1{`RANDOM}};
  do_redirect_bits_cfiUpdate_folded_hist_hist_15_folded_hist = _RAND_341[10:0];
  _RAND_342 = {1{`RANDOM}};
  do_redirect_bits_cfiUpdate_folded_hist_hist_14_folded_hist = _RAND_342[6:0];
  _RAND_343 = {1{`RANDOM}};
  do_redirect_bits_cfiUpdate_folded_hist_hist_13_folded_hist = _RAND_343[6:0];
  _RAND_344 = {1{`RANDOM}};
  do_redirect_bits_cfiUpdate_folded_hist_hist_12_folded_hist = _RAND_344[6:0];
  _RAND_345 = {1{`RANDOM}};
  do_redirect_bits_cfiUpdate_folded_hist_hist_11_folded_hist = _RAND_345[7:0];
  _RAND_346 = {1{`RANDOM}};
  do_redirect_bits_cfiUpdate_folded_hist_hist_10_folded_hist = _RAND_346[8:0];
  _RAND_347 = {1{`RANDOM}};
  do_redirect_bits_cfiUpdate_folded_hist_hist_9_folded_hist = _RAND_347[6:0];
  _RAND_348 = {1{`RANDOM}};
  do_redirect_bits_cfiUpdate_folded_hist_hist_8_folded_hist = _RAND_348[7:0];
  _RAND_349 = {1{`RANDOM}};
  do_redirect_bits_cfiUpdate_folded_hist_hist_7_folded_hist = _RAND_349[8:0];
  _RAND_350 = {1{`RANDOM}};
  do_redirect_bits_cfiUpdate_folded_hist_hist_6_folded_hist = _RAND_350[8:0];
  _RAND_351 = {1{`RANDOM}};
  do_redirect_bits_cfiUpdate_folded_hist_hist_5_folded_hist = _RAND_351[10:0];
  _RAND_352 = {1{`RANDOM}};
  do_redirect_bits_cfiUpdate_folded_hist_hist_4_folded_hist = _RAND_352[3:0];
  _RAND_353 = {1{`RANDOM}};
  do_redirect_bits_cfiUpdate_folded_hist_hist_3_folded_hist = _RAND_353[10:0];
  _RAND_354 = {1{`RANDOM}};
  do_redirect_bits_cfiUpdate_folded_hist_hist_2_folded_hist = _RAND_354[7:0];
  _RAND_355 = {1{`RANDOM}};
  do_redirect_bits_cfiUpdate_folded_hist_hist_1_folded_hist = _RAND_355[7:0];
  _RAND_356 = {1{`RANDOM}};
  do_redirect_bits_cfiUpdate_folded_hist_hist_0_folded_hist = _RAND_356[7:0];
  _RAND_357 = {1{`RANDOM}};
  do_redirect_bits_cfiUpdate_afhob_afhob_5_bits_0 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  do_redirect_bits_cfiUpdate_afhob_afhob_5_bits_1 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  do_redirect_bits_cfiUpdate_afhob_afhob_5_bits_2 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  do_redirect_bits_cfiUpdate_afhob_afhob_5_bits_3 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  do_redirect_bits_cfiUpdate_afhob_afhob_4_bits_0 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  do_redirect_bits_cfiUpdate_afhob_afhob_4_bits_1 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  do_redirect_bits_cfiUpdate_afhob_afhob_4_bits_2 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  do_redirect_bits_cfiUpdate_afhob_afhob_3_bits_0 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  do_redirect_bits_cfiUpdate_afhob_afhob_3_bits_1 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  do_redirect_bits_cfiUpdate_afhob_afhob_3_bits_2 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  do_redirect_bits_cfiUpdate_afhob_afhob_3_bits_3 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  do_redirect_bits_cfiUpdate_afhob_afhob_2_bits_0 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  do_redirect_bits_cfiUpdate_afhob_afhob_2_bits_1 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  do_redirect_bits_cfiUpdate_afhob_afhob_2_bits_2 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  do_redirect_bits_cfiUpdate_afhob_afhob_2_bits_3 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  do_redirect_bits_cfiUpdate_afhob_afhob_1_bits_0 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  do_redirect_bits_cfiUpdate_afhob_afhob_1_bits_1 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  do_redirect_bits_cfiUpdate_afhob_afhob_1_bits_2 = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  do_redirect_bits_cfiUpdate_afhob_afhob_1_bits_3 = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  do_redirect_bits_cfiUpdate_afhob_afhob_0_bits_0 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  do_redirect_bits_cfiUpdate_afhob_afhob_0_bits_1 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  do_redirect_bits_cfiUpdate_afhob_afhob_0_bits_2 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  do_redirect_bits_cfiUpdate_afhob_afhob_0_bits_3 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  do_redirect_bits_cfiUpdate_lastBrNumOH = _RAND_380[2:0];
  _RAND_381 = {1{`RANDOM}};
  do_redirect_bits_cfiUpdate_histPtr_flag = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  do_redirect_bits_cfiUpdate_histPtr_value = _RAND_382[7:0];
  _RAND_383 = {2{`RANDOM}};
  do_redirect_bits_cfiUpdate_target = _RAND_383[38:0];
  _RAND_384 = {1{`RANDOM}};
  do_redirect_bits_cfiUpdate_taken = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  do_redirect_bits_cfiUpdate_shift = _RAND_385[1:0];
  _RAND_386 = {1{`RANDOM}};
  do_redirect_bits_cfiUpdate_addIntoHist = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  previous_s2_pred_full_pred_br_taken_mask_1 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  previous_s2_pred_full_pred_slot_valids_1 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  previous_s2_pred_full_pred_is_br_sharing = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  previous_s2_pred_full_pred_hit = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  previous_s2_pred_full_pred_slot_valids_0 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  previous_s2_pred_full_pred_br_taken_mask_0 = _RAND_392[0:0];
  _RAND_393 = {2{`RANDOM}};
  previous_s2_pred_full_pred_targets_0 = _RAND_393[38:0];
  _RAND_394 = {2{`RANDOM}};
  previous_s2_pred_full_pred_targets_1 = _RAND_394[38:0];
  _RAND_395 = {2{`RANDOM}};
  previous_s2_pred_full_pred_fallThroughAddr = _RAND_395[38:0];
  _RAND_396 = {2{`RANDOM}};
  previous_s2_pred_pc = _RAND_396[38:0];
  _RAND_397 = {2{`RANDOM}};
  previous_s1_pred_info_target = _RAND_397[38:0];
  _RAND_398 = {1{`RANDOM}};
  previous_s1_pred_info_lastBrPosOH = _RAND_398[2:0];
  _RAND_399 = {1{`RANDOM}};
  previous_s1_pred_info_taken = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  previous_s1_pred_info_cfiIndex = _RAND_400[2:0];
  _RAND_401 = {1{`RANDOM}};
  s2_ftq_idx_flag = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  s2_ftq_idx_value = _RAND_402[2:0];
  _RAND_403 = {1{`RANDOM}};
  s3_ftq_idx_flag = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  s3_ftq_idx_value = _RAND_404[2:0];
  _RAND_405 = {1{`RANDOM}};
  predictors_io_update_REG_valid = _RAND_405[0:0];
  _RAND_406 = {2{`RANDOM}};
  predictors_io_update_REG_bits_pc = _RAND_406[38:0];
  _RAND_407 = {1{`RANDOM}};
  predictors_io_update_REG_bits_spec_info_folded_hist_hist_17_folded_hist = _RAND_407[7:0];
  _RAND_408 = {1{`RANDOM}};
  predictors_io_update_REG_bits_spec_info_folded_hist_hist_16_folded_hist = _RAND_408[7:0];
  _RAND_409 = {1{`RANDOM}};
  predictors_io_update_REG_bits_spec_info_folded_hist_hist_15_folded_hist = _RAND_409[10:0];
  _RAND_410 = {1{`RANDOM}};
  predictors_io_update_REG_bits_spec_info_folded_hist_hist_14_folded_hist = _RAND_410[6:0];
  _RAND_411 = {1{`RANDOM}};
  predictors_io_update_REG_bits_spec_info_folded_hist_hist_13_folded_hist = _RAND_411[6:0];
  _RAND_412 = {1{`RANDOM}};
  predictors_io_update_REG_bits_spec_info_folded_hist_hist_12_folded_hist = _RAND_412[6:0];
  _RAND_413 = {1{`RANDOM}};
  predictors_io_update_REG_bits_spec_info_folded_hist_hist_10_folded_hist = _RAND_413[8:0];
  _RAND_414 = {1{`RANDOM}};
  predictors_io_update_REG_bits_spec_info_folded_hist_hist_9_folded_hist = _RAND_414[6:0];
  _RAND_415 = {1{`RANDOM}};
  predictors_io_update_REG_bits_spec_info_folded_hist_hist_8_folded_hist = _RAND_415[7:0];
  _RAND_416 = {1{`RANDOM}};
  predictors_io_update_REG_bits_spec_info_folded_hist_hist_7_folded_hist = _RAND_416[8:0];
  _RAND_417 = {1{`RANDOM}};
  predictors_io_update_REG_bits_spec_info_folded_hist_hist_6_folded_hist = _RAND_417[8:0];
  _RAND_418 = {1{`RANDOM}};
  predictors_io_update_REG_bits_spec_info_folded_hist_hist_5_folded_hist = _RAND_418[10:0];
  _RAND_419 = {1{`RANDOM}};
  predictors_io_update_REG_bits_spec_info_folded_hist_hist_4_folded_hist = _RAND_419[3:0];
  _RAND_420 = {1{`RANDOM}};
  predictors_io_update_REG_bits_spec_info_folded_hist_hist_3_folded_hist = _RAND_420[10:0];
  _RAND_421 = {1{`RANDOM}};
  predictors_io_update_REG_bits_spec_info_folded_hist_hist_2_folded_hist = _RAND_421[7:0];
  _RAND_422 = {1{`RANDOM}};
  predictors_io_update_REG_bits_spec_info_folded_hist_hist_1_folded_hist = _RAND_422[7:0];
  _RAND_423 = {1{`RANDOM}};
  predictors_io_update_REG_bits_spec_info_folded_hist_hist_0_folded_hist = _RAND_423[7:0];
  _RAND_424 = {1{`RANDOM}};
  predictors_io_update_REG_bits_ftb_entry_valid = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  predictors_io_update_REG_bits_ftb_entry_brSlots_0_offset = _RAND_425[2:0];
  _RAND_426 = {1{`RANDOM}};
  predictors_io_update_REG_bits_ftb_entry_brSlots_0_lower = _RAND_426[11:0];
  _RAND_427 = {1{`RANDOM}};
  predictors_io_update_REG_bits_ftb_entry_brSlots_0_tarStat = _RAND_427[1:0];
  _RAND_428 = {1{`RANDOM}};
  predictors_io_update_REG_bits_ftb_entry_brSlots_0_sharing = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  predictors_io_update_REG_bits_ftb_entry_brSlots_0_valid = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  predictors_io_update_REG_bits_ftb_entry_tailSlot_offset = _RAND_430[2:0];
  _RAND_431 = {1{`RANDOM}};
  predictors_io_update_REG_bits_ftb_entry_tailSlot_lower = _RAND_431[19:0];
  _RAND_432 = {1{`RANDOM}};
  predictors_io_update_REG_bits_ftb_entry_tailSlot_tarStat = _RAND_432[1:0];
  _RAND_433 = {1{`RANDOM}};
  predictors_io_update_REG_bits_ftb_entry_tailSlot_sharing = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  predictors_io_update_REG_bits_ftb_entry_tailSlot_valid = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  predictors_io_update_REG_bits_ftb_entry_pftAddr = _RAND_435[2:0];
  _RAND_436 = {1{`RANDOM}};
  predictors_io_update_REG_bits_ftb_entry_carry = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  predictors_io_update_REG_bits_ftb_entry_isCall = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  predictors_io_update_REG_bits_ftb_entry_isRet = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  predictors_io_update_REG_bits_ftb_entry_isJalr = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  predictors_io_update_REG_bits_ftb_entry_last_may_be_rvi_call = _RAND_440[0:0];
  _RAND_441 = {1{`RANDOM}};
  predictors_io_update_REG_bits_ftb_entry_always_taken_0 = _RAND_441[0:0];
  _RAND_442 = {1{`RANDOM}};
  predictors_io_update_REG_bits_ftb_entry_always_taken_1 = _RAND_442[0:0];
  _RAND_443 = {1{`RANDOM}};
  predictors_io_update_REG_bits_br_taken_mask_0 = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  predictors_io_update_REG_bits_br_taken_mask_1 = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  predictors_io_update_REG_bits_jmp_taken = _RAND_445[0:0];
  _RAND_446 = {1{`RANDOM}};
  predictors_io_update_REG_bits_mispred_mask_0 = _RAND_446[0:0];
  _RAND_447 = {1{`RANDOM}};
  predictors_io_update_REG_bits_mispred_mask_1 = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  predictors_io_update_REG_bits_mispred_mask_2 = _RAND_448[0:0];
  _RAND_449 = {1{`RANDOM}};
  predictors_io_update_REG_bits_old_entry = _RAND_449[0:0];
  _RAND_450 = {8{`RANDOM}};
  predictors_io_update_REG_bits_meta = _RAND_450[255:0];
  _RAND_451 = {2{`RANDOM}};
  predictors_io_update_REG_bits_full_target = _RAND_451[38:0];
  _RAND_452 = {1{`RANDOM}};
  io_perf_0_value_REG = _RAND_452[5:0];
  _RAND_453 = {1{`RANDOM}};
  io_perf_0_value_REG_1 = _RAND_453[5:0];
  _RAND_454 = {1{`RANDOM}};
  io_perf_1_value_REG = _RAND_454[5:0];
  _RAND_455 = {1{`RANDOM}};
  io_perf_1_value_REG_1 = _RAND_455[5:0];
  _RAND_456 = {1{`RANDOM}};
  io_perf_2_value_REG = _RAND_456[5:0];
  _RAND_457 = {1{`RANDOM}};
  io_perf_2_value_REG_1 = _RAND_457[5:0];
  _RAND_458 = {1{`RANDOM}};
  io_perf_3_value_REG = _RAND_458[5:0];
  _RAND_459 = {1{`RANDOM}};
  io_perf_3_value_REG_1 = _RAND_459[5:0];
  _RAND_460 = {1{`RANDOM}};
  io_perf_4_value_REG = _RAND_460[5:0];
  _RAND_461 = {1{`RANDOM}};
  io_perf_4_value_REG_1 = _RAND_461[5:0];
  _RAND_462 = {1{`RANDOM}};
  io_perf_5_value_REG = _RAND_462[5:0];
  _RAND_463 = {1{`RANDOM}};
  io_perf_5_value_REG_1 = _RAND_463[5:0];
  _RAND_464 = {1{`RANDOM}};
  io_perf_6_value_REG = _RAND_464[5:0];
  _RAND_465 = {1{`RANDOM}};
  io_perf_6_value_REG_1 = _RAND_465[5:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    s1_valid = 1'h0;
  end
  if (reset) begin
    s2_valid = 1'h0;
  end
  if (reset) begin
    s3_valid = 1'h0;
  end
  if (reset) begin
    s0_folded_gh_reg_hist_17_folded_hist = 8'h0;
  end
  if (reset) begin
    s0_folded_gh_reg_hist_16_folded_hist = 8'h0;
  end
  if (reset) begin
    s0_folded_gh_reg_hist_15_folded_hist = 11'h0;
  end
  if (reset) begin
    s0_folded_gh_reg_hist_14_folded_hist = 7'h0;
  end
  if (reset) begin
    s0_folded_gh_reg_hist_13_folded_hist = 7'h0;
  end
  if (reset) begin
    s0_folded_gh_reg_hist_12_folded_hist = 7'h0;
  end
  if (reset) begin
    s0_folded_gh_reg_hist_11_folded_hist = 8'h0;
  end
  if (reset) begin
    s0_folded_gh_reg_hist_10_folded_hist = 9'h0;
  end
  if (reset) begin
    s0_folded_gh_reg_hist_9_folded_hist = 7'h0;
  end
  if (reset) begin
    s0_folded_gh_reg_hist_8_folded_hist = 8'h0;
  end
  if (reset) begin
    s0_folded_gh_reg_hist_7_folded_hist = 9'h0;
  end
  if (reset) begin
    s0_folded_gh_reg_hist_6_folded_hist = 9'h0;
  end
  if (reset) begin
    s0_folded_gh_reg_hist_5_folded_hist = 11'h0;
  end
  if (reset) begin
    s0_folded_gh_reg_hist_4_folded_hist = 4'h0;
  end
  if (reset) begin
    s0_folded_gh_reg_hist_3_folded_hist = 11'h0;
  end
  if (reset) begin
    s0_folded_gh_reg_hist_2_folded_hist = 8'h0;
  end
  if (reset) begin
    s0_folded_gh_reg_hist_1_folded_hist = 8'h0;
  end
  if (reset) begin
    s0_folded_gh_reg_hist_0_folded_hist = 8'h0;
  end
  if (reset) begin
    s1_folded_gh_hist_17_folded_hist = 8'h0;
  end
  if (reset) begin
    s1_folded_gh_hist_16_folded_hist = 8'h0;
  end
  if (reset) begin
    s1_folded_gh_hist_15_folded_hist = 11'h0;
  end
  if (reset) begin
    s1_folded_gh_hist_14_folded_hist = 7'h0;
  end
  if (reset) begin
    s1_folded_gh_hist_13_folded_hist = 7'h0;
  end
  if (reset) begin
    s1_folded_gh_hist_12_folded_hist = 7'h0;
  end
  if (reset) begin
    s1_folded_gh_hist_11_folded_hist = 8'h0;
  end
  if (reset) begin
    s1_folded_gh_hist_10_folded_hist = 9'h0;
  end
  if (reset) begin
    s1_folded_gh_hist_9_folded_hist = 7'h0;
  end
  if (reset) begin
    s1_folded_gh_hist_8_folded_hist = 8'h0;
  end
  if (reset) begin
    s1_folded_gh_hist_7_folded_hist = 9'h0;
  end
  if (reset) begin
    s1_folded_gh_hist_6_folded_hist = 9'h0;
  end
  if (reset) begin
    s1_folded_gh_hist_5_folded_hist = 11'h0;
  end
  if (reset) begin
    s1_folded_gh_hist_4_folded_hist = 4'h0;
  end
  if (reset) begin
    s1_folded_gh_hist_3_folded_hist = 11'h0;
  end
  if (reset) begin
    s1_folded_gh_hist_2_folded_hist = 8'h0;
  end
  if (reset) begin
    s1_folded_gh_hist_1_folded_hist = 8'h0;
  end
  if (reset) begin
    s1_folded_gh_hist_0_folded_hist = 8'h0;
  end
  if (reset) begin
    s2_folded_gh_hist_17_folded_hist = 8'h0;
  end
  if (reset) begin
    s2_folded_gh_hist_16_folded_hist = 8'h0;
  end
  if (reset) begin
    s2_folded_gh_hist_15_folded_hist = 11'h0;
  end
  if (reset) begin
    s2_folded_gh_hist_14_folded_hist = 7'h0;
  end
  if (reset) begin
    s2_folded_gh_hist_13_folded_hist = 7'h0;
  end
  if (reset) begin
    s2_folded_gh_hist_12_folded_hist = 7'h0;
  end
  if (reset) begin
    s2_folded_gh_hist_11_folded_hist = 8'h0;
  end
  if (reset) begin
    s2_folded_gh_hist_10_folded_hist = 9'h0;
  end
  if (reset) begin
    s2_folded_gh_hist_9_folded_hist = 7'h0;
  end
  if (reset) begin
    s2_folded_gh_hist_8_folded_hist = 8'h0;
  end
  if (reset) begin
    s2_folded_gh_hist_7_folded_hist = 9'h0;
  end
  if (reset) begin
    s2_folded_gh_hist_6_folded_hist = 9'h0;
  end
  if (reset) begin
    s2_folded_gh_hist_5_folded_hist = 11'h0;
  end
  if (reset) begin
    s2_folded_gh_hist_4_folded_hist = 4'h0;
  end
  if (reset) begin
    s2_folded_gh_hist_3_folded_hist = 11'h0;
  end
  if (reset) begin
    s2_folded_gh_hist_2_folded_hist = 8'h0;
  end
  if (reset) begin
    s2_folded_gh_hist_1_folded_hist = 8'h0;
  end
  if (reset) begin
    s2_folded_gh_hist_0_folded_hist = 8'h0;
  end
  if (reset) begin
    s3_folded_gh_hist_17_folded_hist = 8'h0;
  end
  if (reset) begin
    s3_folded_gh_hist_16_folded_hist = 8'h0;
  end
  if (reset) begin
    s3_folded_gh_hist_15_folded_hist = 11'h0;
  end
  if (reset) begin
    s3_folded_gh_hist_14_folded_hist = 7'h0;
  end
  if (reset) begin
    s3_folded_gh_hist_13_folded_hist = 7'h0;
  end
  if (reset) begin
    s3_folded_gh_hist_12_folded_hist = 7'h0;
  end
  if (reset) begin
    s3_folded_gh_hist_11_folded_hist = 8'h0;
  end
  if (reset) begin
    s3_folded_gh_hist_10_folded_hist = 9'h0;
  end
  if (reset) begin
    s3_folded_gh_hist_9_folded_hist = 7'h0;
  end
  if (reset) begin
    s3_folded_gh_hist_8_folded_hist = 8'h0;
  end
  if (reset) begin
    s3_folded_gh_hist_7_folded_hist = 9'h0;
  end
  if (reset) begin
    s3_folded_gh_hist_6_folded_hist = 9'h0;
  end
  if (reset) begin
    s3_folded_gh_hist_5_folded_hist = 11'h0;
  end
  if (reset) begin
    s3_folded_gh_hist_4_folded_hist = 4'h0;
  end
  if (reset) begin
    s3_folded_gh_hist_3_folded_hist = 11'h0;
  end
  if (reset) begin
    s3_folded_gh_hist_2_folded_hist = 8'h0;
  end
  if (reset) begin
    s3_folded_gh_hist_1_folded_hist = 8'h0;
  end
  if (reset) begin
    s3_folded_gh_hist_0_folded_hist = 8'h0;
  end
  if (reset) begin
    s0_last_br_num_oh_reg = 3'h0;
  end
  if (reset) begin
    s1_last_br_num_oh = 3'h0;
  end
  if (reset) begin
    s2_last_br_num_oh = 3'h0;
  end
  if (reset) begin
    s3_last_br_num_oh = 3'h0;
  end
  if (reset) begin
    s0_ahead_fh_oldest_bits_reg_afhob_5_bits_0 = 1'h0;
  end
  if (reset) begin
    s0_ahead_fh_oldest_bits_reg_afhob_5_bits_1 = 1'h0;
  end
  if (reset) begin
    s0_ahead_fh_oldest_bits_reg_afhob_5_bits_2 = 1'h0;
  end
  if (reset) begin
    s0_ahead_fh_oldest_bits_reg_afhob_5_bits_3 = 1'h0;
  end
  if (reset) begin
    s0_ahead_fh_oldest_bits_reg_afhob_4_bits_0 = 1'h0;
  end
  if (reset) begin
    s0_ahead_fh_oldest_bits_reg_afhob_4_bits_1 = 1'h0;
  end
  if (reset) begin
    s0_ahead_fh_oldest_bits_reg_afhob_4_bits_2 = 1'h0;
  end
  if (reset) begin
    s0_ahead_fh_oldest_bits_reg_afhob_4_bits_3 = 1'h0;
  end
  if (reset) begin
    s0_ahead_fh_oldest_bits_reg_afhob_3_bits_0 = 1'h0;
  end
  if (reset) begin
    s0_ahead_fh_oldest_bits_reg_afhob_3_bits_1 = 1'h0;
  end
  if (reset) begin
    s0_ahead_fh_oldest_bits_reg_afhob_3_bits_2 = 1'h0;
  end
  if (reset) begin
    s0_ahead_fh_oldest_bits_reg_afhob_3_bits_3 = 1'h0;
  end
  if (reset) begin
    s0_ahead_fh_oldest_bits_reg_afhob_2_bits_0 = 1'h0;
  end
  if (reset) begin
    s0_ahead_fh_oldest_bits_reg_afhob_2_bits_1 = 1'h0;
  end
  if (reset) begin
    s0_ahead_fh_oldest_bits_reg_afhob_2_bits_2 = 1'h0;
  end
  if (reset) begin
    s0_ahead_fh_oldest_bits_reg_afhob_2_bits_3 = 1'h0;
  end
  if (reset) begin
    s0_ahead_fh_oldest_bits_reg_afhob_1_bits_0 = 1'h0;
  end
  if (reset) begin
    s0_ahead_fh_oldest_bits_reg_afhob_1_bits_1 = 1'h0;
  end
  if (reset) begin
    s0_ahead_fh_oldest_bits_reg_afhob_1_bits_2 = 1'h0;
  end
  if (reset) begin
    s0_ahead_fh_oldest_bits_reg_afhob_1_bits_3 = 1'h0;
  end
  if (reset) begin
    s0_ahead_fh_oldest_bits_reg_afhob_0_bits_0 = 1'h0;
  end
  if (reset) begin
    s0_ahead_fh_oldest_bits_reg_afhob_0_bits_1 = 1'h0;
  end
  if (reset) begin
    s0_ahead_fh_oldest_bits_reg_afhob_0_bits_2 = 1'h0;
  end
  if (reset) begin
    s0_ahead_fh_oldest_bits_reg_afhob_0_bits_3 = 1'h0;
  end
  if (reset) begin
    s1_ahead_fh_oldest_bits_afhob_5_bits_0 = 1'h0;
  end
  if (reset) begin
    s1_ahead_fh_oldest_bits_afhob_5_bits_1 = 1'h0;
  end
  if (reset) begin
    s1_ahead_fh_oldest_bits_afhob_5_bits_2 = 1'h0;
  end
  if (reset) begin
    s1_ahead_fh_oldest_bits_afhob_5_bits_3 = 1'h0;
  end
  if (reset) begin
    s1_ahead_fh_oldest_bits_afhob_4_bits_0 = 1'h0;
  end
  if (reset) begin
    s1_ahead_fh_oldest_bits_afhob_4_bits_1 = 1'h0;
  end
  if (reset) begin
    s1_ahead_fh_oldest_bits_afhob_4_bits_2 = 1'h0;
  end
  if (reset) begin
    s1_ahead_fh_oldest_bits_afhob_4_bits_3 = 1'h0;
  end
  if (reset) begin
    s1_ahead_fh_oldest_bits_afhob_3_bits_0 = 1'h0;
  end
  if (reset) begin
    s1_ahead_fh_oldest_bits_afhob_3_bits_1 = 1'h0;
  end
  if (reset) begin
    s1_ahead_fh_oldest_bits_afhob_3_bits_2 = 1'h0;
  end
  if (reset) begin
    s1_ahead_fh_oldest_bits_afhob_3_bits_3 = 1'h0;
  end
  if (reset) begin
    s1_ahead_fh_oldest_bits_afhob_2_bits_0 = 1'h0;
  end
  if (reset) begin
    s1_ahead_fh_oldest_bits_afhob_2_bits_1 = 1'h0;
  end
  if (reset) begin
    s1_ahead_fh_oldest_bits_afhob_2_bits_2 = 1'h0;
  end
  if (reset) begin
    s1_ahead_fh_oldest_bits_afhob_2_bits_3 = 1'h0;
  end
  if (reset) begin
    s1_ahead_fh_oldest_bits_afhob_1_bits_0 = 1'h0;
  end
  if (reset) begin
    s1_ahead_fh_oldest_bits_afhob_1_bits_1 = 1'h0;
  end
  if (reset) begin
    s1_ahead_fh_oldest_bits_afhob_1_bits_2 = 1'h0;
  end
  if (reset) begin
    s1_ahead_fh_oldest_bits_afhob_1_bits_3 = 1'h0;
  end
  if (reset) begin
    s1_ahead_fh_oldest_bits_afhob_0_bits_0 = 1'h0;
  end
  if (reset) begin
    s1_ahead_fh_oldest_bits_afhob_0_bits_1 = 1'h0;
  end
  if (reset) begin
    s1_ahead_fh_oldest_bits_afhob_0_bits_2 = 1'h0;
  end
  if (reset) begin
    s1_ahead_fh_oldest_bits_afhob_0_bits_3 = 1'h0;
  end
  if (reset) begin
    s2_ahead_fh_oldest_bits_afhob_5_bits_0 = 1'h0;
  end
  if (reset) begin
    s2_ahead_fh_oldest_bits_afhob_5_bits_1 = 1'h0;
  end
  if (reset) begin
    s2_ahead_fh_oldest_bits_afhob_5_bits_2 = 1'h0;
  end
  if (reset) begin
    s2_ahead_fh_oldest_bits_afhob_5_bits_3 = 1'h0;
  end
  if (reset) begin
    s2_ahead_fh_oldest_bits_afhob_4_bits_0 = 1'h0;
  end
  if (reset) begin
    s2_ahead_fh_oldest_bits_afhob_4_bits_1 = 1'h0;
  end
  if (reset) begin
    s2_ahead_fh_oldest_bits_afhob_4_bits_2 = 1'h0;
  end
  if (reset) begin
    s2_ahead_fh_oldest_bits_afhob_4_bits_3 = 1'h0;
  end
  if (reset) begin
    s2_ahead_fh_oldest_bits_afhob_3_bits_0 = 1'h0;
  end
  if (reset) begin
    s2_ahead_fh_oldest_bits_afhob_3_bits_1 = 1'h0;
  end
  if (reset) begin
    s2_ahead_fh_oldest_bits_afhob_3_bits_2 = 1'h0;
  end
  if (reset) begin
    s2_ahead_fh_oldest_bits_afhob_3_bits_3 = 1'h0;
  end
  if (reset) begin
    s2_ahead_fh_oldest_bits_afhob_2_bits_0 = 1'h0;
  end
  if (reset) begin
    s2_ahead_fh_oldest_bits_afhob_2_bits_1 = 1'h0;
  end
  if (reset) begin
    s2_ahead_fh_oldest_bits_afhob_2_bits_2 = 1'h0;
  end
  if (reset) begin
    s2_ahead_fh_oldest_bits_afhob_2_bits_3 = 1'h0;
  end
  if (reset) begin
    s2_ahead_fh_oldest_bits_afhob_1_bits_0 = 1'h0;
  end
  if (reset) begin
    s2_ahead_fh_oldest_bits_afhob_1_bits_1 = 1'h0;
  end
  if (reset) begin
    s2_ahead_fh_oldest_bits_afhob_1_bits_2 = 1'h0;
  end
  if (reset) begin
    s2_ahead_fh_oldest_bits_afhob_1_bits_3 = 1'h0;
  end
  if (reset) begin
    s2_ahead_fh_oldest_bits_afhob_0_bits_0 = 1'h0;
  end
  if (reset) begin
    s2_ahead_fh_oldest_bits_afhob_0_bits_1 = 1'h0;
  end
  if (reset) begin
    s2_ahead_fh_oldest_bits_afhob_0_bits_2 = 1'h0;
  end
  if (reset) begin
    s2_ahead_fh_oldest_bits_afhob_0_bits_3 = 1'h0;
  end
  if (reset) begin
    s3_ahead_fh_oldest_bits_afhob_5_bits_0 = 1'h0;
  end
  if (reset) begin
    s3_ahead_fh_oldest_bits_afhob_5_bits_1 = 1'h0;
  end
  if (reset) begin
    s3_ahead_fh_oldest_bits_afhob_5_bits_2 = 1'h0;
  end
  if (reset) begin
    s3_ahead_fh_oldest_bits_afhob_5_bits_3 = 1'h0;
  end
  if (reset) begin
    s3_ahead_fh_oldest_bits_afhob_4_bits_0 = 1'h0;
  end
  if (reset) begin
    s3_ahead_fh_oldest_bits_afhob_4_bits_1 = 1'h0;
  end
  if (reset) begin
    s3_ahead_fh_oldest_bits_afhob_4_bits_2 = 1'h0;
  end
  if (reset) begin
    s3_ahead_fh_oldest_bits_afhob_4_bits_3 = 1'h0;
  end
  if (reset) begin
    s3_ahead_fh_oldest_bits_afhob_3_bits_0 = 1'h0;
  end
  if (reset) begin
    s3_ahead_fh_oldest_bits_afhob_3_bits_1 = 1'h0;
  end
  if (reset) begin
    s3_ahead_fh_oldest_bits_afhob_3_bits_2 = 1'h0;
  end
  if (reset) begin
    s3_ahead_fh_oldest_bits_afhob_3_bits_3 = 1'h0;
  end
  if (reset) begin
    s3_ahead_fh_oldest_bits_afhob_2_bits_0 = 1'h0;
  end
  if (reset) begin
    s3_ahead_fh_oldest_bits_afhob_2_bits_1 = 1'h0;
  end
  if (reset) begin
    s3_ahead_fh_oldest_bits_afhob_2_bits_2 = 1'h0;
  end
  if (reset) begin
    s3_ahead_fh_oldest_bits_afhob_2_bits_3 = 1'h0;
  end
  if (reset) begin
    s3_ahead_fh_oldest_bits_afhob_1_bits_0 = 1'h0;
  end
  if (reset) begin
    s3_ahead_fh_oldest_bits_afhob_1_bits_1 = 1'h0;
  end
  if (reset) begin
    s3_ahead_fh_oldest_bits_afhob_1_bits_2 = 1'h0;
  end
  if (reset) begin
    s3_ahead_fh_oldest_bits_afhob_1_bits_3 = 1'h0;
  end
  if (reset) begin
    s3_ahead_fh_oldest_bits_afhob_0_bits_0 = 1'h0;
  end
  if (reset) begin
    s3_ahead_fh_oldest_bits_afhob_0_bits_1 = 1'h0;
  end
  if (reset) begin
    s3_ahead_fh_oldest_bits_afhob_0_bits_2 = 1'h0;
  end
  if (reset) begin
    s3_ahead_fh_oldest_bits_afhob_0_bits_3 = 1'h0;
  end
  if (reset) begin
    ghv_0 = 1'h0;
  end
  if (reset) begin
    ghv_1 = 1'h0;
  end
  if (reset) begin
    ghv_2 = 1'h0;
  end
  if (reset) begin
    ghv_3 = 1'h0;
  end
  if (reset) begin
    ghv_4 = 1'h0;
  end
  if (reset) begin
    ghv_5 = 1'h0;
  end
  if (reset) begin
    ghv_6 = 1'h0;
  end
  if (reset) begin
    ghv_7 = 1'h0;
  end
  if (reset) begin
    ghv_8 = 1'h0;
  end
  if (reset) begin
    ghv_9 = 1'h0;
  end
  if (reset) begin
    ghv_10 = 1'h0;
  end
  if (reset) begin
    ghv_11 = 1'h0;
  end
  if (reset) begin
    ghv_12 = 1'h0;
  end
  if (reset) begin
    ghv_13 = 1'h0;
  end
  if (reset) begin
    ghv_14 = 1'h0;
  end
  if (reset) begin
    ghv_15 = 1'h0;
  end
  if (reset) begin
    ghv_16 = 1'h0;
  end
  if (reset) begin
    ghv_17 = 1'h0;
  end
  if (reset) begin
    ghv_18 = 1'h0;
  end
  if (reset) begin
    ghv_19 = 1'h0;
  end
  if (reset) begin
    ghv_20 = 1'h0;
  end
  if (reset) begin
    ghv_21 = 1'h0;
  end
  if (reset) begin
    ghv_22 = 1'h0;
  end
  if (reset) begin
    ghv_23 = 1'h0;
  end
  if (reset) begin
    ghv_24 = 1'h0;
  end
  if (reset) begin
    ghv_25 = 1'h0;
  end
  if (reset) begin
    ghv_26 = 1'h0;
  end
  if (reset) begin
    ghv_27 = 1'h0;
  end
  if (reset) begin
    ghv_28 = 1'h0;
  end
  if (reset) begin
    ghv_29 = 1'h0;
  end
  if (reset) begin
    ghv_30 = 1'h0;
  end
  if (reset) begin
    ghv_31 = 1'h0;
  end
  if (reset) begin
    ghv_32 = 1'h0;
  end
  if (reset) begin
    ghv_33 = 1'h0;
  end
  if (reset) begin
    ghv_34 = 1'h0;
  end
  if (reset) begin
    ghv_35 = 1'h0;
  end
  if (reset) begin
    ghv_36 = 1'h0;
  end
  if (reset) begin
    ghv_37 = 1'h0;
  end
  if (reset) begin
    ghv_38 = 1'h0;
  end
  if (reset) begin
    ghv_39 = 1'h0;
  end
  if (reset) begin
    ghv_40 = 1'h0;
  end
  if (reset) begin
    ghv_41 = 1'h0;
  end
  if (reset) begin
    ghv_42 = 1'h0;
  end
  if (reset) begin
    ghv_43 = 1'h0;
  end
  if (reset) begin
    ghv_44 = 1'h0;
  end
  if (reset) begin
    ghv_45 = 1'h0;
  end
  if (reset) begin
    ghv_46 = 1'h0;
  end
  if (reset) begin
    ghv_47 = 1'h0;
  end
  if (reset) begin
    ghv_48 = 1'h0;
  end
  if (reset) begin
    ghv_49 = 1'h0;
  end
  if (reset) begin
    ghv_50 = 1'h0;
  end
  if (reset) begin
    ghv_51 = 1'h0;
  end
  if (reset) begin
    ghv_52 = 1'h0;
  end
  if (reset) begin
    ghv_53 = 1'h0;
  end
  if (reset) begin
    ghv_54 = 1'h0;
  end
  if (reset) begin
    ghv_55 = 1'h0;
  end
  if (reset) begin
    ghv_56 = 1'h0;
  end
  if (reset) begin
    ghv_57 = 1'h0;
  end
  if (reset) begin
    ghv_58 = 1'h0;
  end
  if (reset) begin
    ghv_59 = 1'h0;
  end
  if (reset) begin
    ghv_60 = 1'h0;
  end
  if (reset) begin
    ghv_61 = 1'h0;
  end
  if (reset) begin
    ghv_62 = 1'h0;
  end
  if (reset) begin
    ghv_63 = 1'h0;
  end
  if (reset) begin
    ghv_64 = 1'h0;
  end
  if (reset) begin
    ghv_65 = 1'h0;
  end
  if (reset) begin
    ghv_66 = 1'h0;
  end
  if (reset) begin
    ghv_67 = 1'h0;
  end
  if (reset) begin
    ghv_68 = 1'h0;
  end
  if (reset) begin
    ghv_69 = 1'h0;
  end
  if (reset) begin
    ghv_70 = 1'h0;
  end
  if (reset) begin
    ghv_71 = 1'h0;
  end
  if (reset) begin
    ghv_72 = 1'h0;
  end
  if (reset) begin
    ghv_73 = 1'h0;
  end
  if (reset) begin
    ghv_74 = 1'h0;
  end
  if (reset) begin
    ghv_75 = 1'h0;
  end
  if (reset) begin
    ghv_76 = 1'h0;
  end
  if (reset) begin
    ghv_77 = 1'h0;
  end
  if (reset) begin
    ghv_78 = 1'h0;
  end
  if (reset) begin
    ghv_79 = 1'h0;
  end
  if (reset) begin
    ghv_80 = 1'h0;
  end
  if (reset) begin
    ghv_81 = 1'h0;
  end
  if (reset) begin
    ghv_82 = 1'h0;
  end
  if (reset) begin
    ghv_83 = 1'h0;
  end
  if (reset) begin
    ghv_84 = 1'h0;
  end
  if (reset) begin
    ghv_85 = 1'h0;
  end
  if (reset) begin
    ghv_86 = 1'h0;
  end
  if (reset) begin
    ghv_87 = 1'h0;
  end
  if (reset) begin
    ghv_88 = 1'h0;
  end
  if (reset) begin
    ghv_89 = 1'h0;
  end
  if (reset) begin
    ghv_90 = 1'h0;
  end
  if (reset) begin
    ghv_91 = 1'h0;
  end
  if (reset) begin
    ghv_92 = 1'h0;
  end
  if (reset) begin
    ghv_93 = 1'h0;
  end
  if (reset) begin
    ghv_94 = 1'h0;
  end
  if (reset) begin
    ghv_95 = 1'h0;
  end
  if (reset) begin
    ghv_96 = 1'h0;
  end
  if (reset) begin
    ghv_97 = 1'h0;
  end
  if (reset) begin
    ghv_98 = 1'h0;
  end
  if (reset) begin
    ghv_99 = 1'h0;
  end
  if (reset) begin
    ghv_100 = 1'h0;
  end
  if (reset) begin
    ghv_101 = 1'h0;
  end
  if (reset) begin
    ghv_102 = 1'h0;
  end
  if (reset) begin
    ghv_103 = 1'h0;
  end
  if (reset) begin
    ghv_104 = 1'h0;
  end
  if (reset) begin
    ghv_105 = 1'h0;
  end
  if (reset) begin
    ghv_106 = 1'h0;
  end
  if (reset) begin
    ghv_107 = 1'h0;
  end
  if (reset) begin
    ghv_108 = 1'h0;
  end
  if (reset) begin
    ghv_109 = 1'h0;
  end
  if (reset) begin
    ghv_110 = 1'h0;
  end
  if (reset) begin
    ghv_111 = 1'h0;
  end
  if (reset) begin
    ghv_112 = 1'h0;
  end
  if (reset) begin
    ghv_113 = 1'h0;
  end
  if (reset) begin
    ghv_114 = 1'h0;
  end
  if (reset) begin
    ghv_115 = 1'h0;
  end
  if (reset) begin
    ghv_116 = 1'h0;
  end
  if (reset) begin
    ghv_117 = 1'h0;
  end
  if (reset) begin
    ghv_118 = 1'h0;
  end
  if (reset) begin
    ghv_119 = 1'h0;
  end
  if (reset) begin
    ghv_120 = 1'h0;
  end
  if (reset) begin
    ghv_121 = 1'h0;
  end
  if (reset) begin
    ghv_122 = 1'h0;
  end
  if (reset) begin
    ghv_123 = 1'h0;
  end
  if (reset) begin
    ghv_124 = 1'h0;
  end
  if (reset) begin
    ghv_125 = 1'h0;
  end
  if (reset) begin
    ghv_126 = 1'h0;
  end
  if (reset) begin
    ghv_127 = 1'h0;
  end
  if (reset) begin
    ghv_128 = 1'h0;
  end
  if (reset) begin
    ghv_129 = 1'h0;
  end
  if (reset) begin
    ghv_130 = 1'h0;
  end
  if (reset) begin
    ghv_131 = 1'h0;
  end
  if (reset) begin
    ghv_132 = 1'h0;
  end
  if (reset) begin
    ghv_133 = 1'h0;
  end
  if (reset) begin
    ghv_134 = 1'h0;
  end
  if (reset) begin
    ghv_135 = 1'h0;
  end
  if (reset) begin
    ghv_136 = 1'h0;
  end
  if (reset) begin
    ghv_137 = 1'h0;
  end
  if (reset) begin
    ghv_138 = 1'h0;
  end
  if (reset) begin
    ghv_139 = 1'h0;
  end
  if (reset) begin
    ghv_140 = 1'h0;
  end
  if (reset) begin
    ghv_141 = 1'h0;
  end
  if (reset) begin
    ghv_142 = 1'h0;
  end
  if (reset) begin
    ghv_143 = 1'h0;
  end
  if (reset) begin
    s0_ghist_ptr_reg_flag = 1'h0;
  end
  if (reset) begin
    s0_ghist_ptr_reg_value = 8'h0;
  end
  if (reset) begin
    s1_ghist_ptr_flag = 1'h0;
  end
  if (reset) begin
    s1_ghist_ptr_value = 8'h0;
  end
  if (reset) begin
    s2_ghist_ptr_flag = 1'h0;
  end
  if (reset) begin
    s2_ghist_ptr_value = 8'h0;
  end
  if (reset) begin
    s3_ghist_ptr_flag = 1'h0;
  end
  if (reset) begin
    s3_ghist_ptr_value = 8'h0;
  end
  if (reset) begin
    do_redirect_valid = 1'h0;
  end
  if (reset) begin
    do_redirect_bits_level = 1'h0;
  end
  if (reset) begin
    do_redirect_bits_cfiUpdate_pc = 39'h0;
  end
  if (reset) begin
    do_redirect_bits_cfiUpdate_pd_isRVC = 1'h0;
  end
  if (reset) begin
    do_redirect_bits_cfiUpdate_pd_isCall = 1'h0;
  end
  if (reset) begin
    do_redirect_bits_cfiUpdate_pd_isRet = 1'h0;
  end
  if (reset) begin
    do_redirect_bits_cfiUpdate_rasSp = 5'h0;
  end
  if (reset) begin
    do_redirect_bits_cfiUpdate_rasEntry_retAddr = 39'h0;
  end
  if (reset) begin
    do_redirect_bits_cfiUpdate_rasEntry_ctr = 8'h0;
  end
  if (reset) begin
    do_redirect_bits_cfiUpdate_folded_hist_hist_17_folded_hist = 8'h0;
  end
  if (reset) begin
    do_redirect_bits_cfiUpdate_folded_hist_hist_16_folded_hist = 8'h0;
  end
  if (reset) begin
    do_redirect_bits_cfiUpdate_folded_hist_hist_15_folded_hist = 11'h0;
  end
  if (reset) begin
    do_redirect_bits_cfiUpdate_folded_hist_hist_14_folded_hist = 7'h0;
  end
  if (reset) begin
    do_redirect_bits_cfiUpdate_folded_hist_hist_13_folded_hist = 7'h0;
  end
  if (reset) begin
    do_redirect_bits_cfiUpdate_folded_hist_hist_12_folded_hist = 7'h0;
  end
  if (reset) begin
    do_redirect_bits_cfiUpdate_folded_hist_hist_11_folded_hist = 8'h0;
  end
  if (reset) begin
    do_redirect_bits_cfiUpdate_folded_hist_hist_10_folded_hist = 9'h0;
  end
  if (reset) begin
    do_redirect_bits_cfiUpdate_folded_hist_hist_9_folded_hist = 7'h0;
  end
  if (reset) begin
    do_redirect_bits_cfiUpdate_folded_hist_hist_8_folded_hist = 8'h0;
  end
  if (reset) begin
    do_redirect_bits_cfiUpdate_folded_hist_hist_7_folded_hist = 9'h0;
  end
  if (reset) begin
    do_redirect_bits_cfiUpdate_folded_hist_hist_6_folded_hist = 9'h0;
  end
  if (reset) begin
    do_redirect_bits_cfiUpdate_folded_hist_hist_5_folded_hist = 11'h0;
  end
  if (reset) begin
    do_redirect_bits_cfiUpdate_folded_hist_hist_4_folded_hist = 4'h0;
  end
  if (reset) begin
    do_redirect_bits_cfiUpdate_folded_hist_hist_3_folded_hist = 11'h0;
  end
  if (reset) begin
    do_redirect_bits_cfiUpdate_folded_hist_hist_2_folded_hist = 8'h0;
  end
  if (reset) begin
    do_redirect_bits_cfiUpdate_folded_hist_hist_1_folded_hist = 8'h0;
  end
  if (reset) begin
    do_redirect_bits_cfiUpdate_folded_hist_hist_0_folded_hist = 8'h0;
  end
  if (reset) begin
    do_redirect_bits_cfiUpdate_afhob_afhob_5_bits_0 = 1'h0;
  end
  if (reset) begin
    do_redirect_bits_cfiUpdate_afhob_afhob_5_bits_1 = 1'h0;
  end
  if (reset) begin
    do_redirect_bits_cfiUpdate_afhob_afhob_5_bits_2 = 1'h0;
  end
  if (reset) begin
    do_redirect_bits_cfiUpdate_afhob_afhob_5_bits_3 = 1'h0;
  end
  if (reset) begin
    do_redirect_bits_cfiUpdate_afhob_afhob_4_bits_0 = 1'h0;
  end
  if (reset) begin
    do_redirect_bits_cfiUpdate_afhob_afhob_4_bits_1 = 1'h0;
  end
  if (reset) begin
    do_redirect_bits_cfiUpdate_afhob_afhob_4_bits_2 = 1'h0;
  end
  if (reset) begin
    do_redirect_bits_cfiUpdate_afhob_afhob_3_bits_0 = 1'h0;
  end
  if (reset) begin
    do_redirect_bits_cfiUpdate_afhob_afhob_3_bits_1 = 1'h0;
  end
  if (reset) begin
    do_redirect_bits_cfiUpdate_afhob_afhob_3_bits_2 = 1'h0;
  end
  if (reset) begin
    do_redirect_bits_cfiUpdate_afhob_afhob_3_bits_3 = 1'h0;
  end
  if (reset) begin
    do_redirect_bits_cfiUpdate_afhob_afhob_2_bits_0 = 1'h0;
  end
  if (reset) begin
    do_redirect_bits_cfiUpdate_afhob_afhob_2_bits_1 = 1'h0;
  end
  if (reset) begin
    do_redirect_bits_cfiUpdate_afhob_afhob_2_bits_2 = 1'h0;
  end
  if (reset) begin
    do_redirect_bits_cfiUpdate_afhob_afhob_2_bits_3 = 1'h0;
  end
  if (reset) begin
    do_redirect_bits_cfiUpdate_afhob_afhob_1_bits_0 = 1'h0;
  end
  if (reset) begin
    do_redirect_bits_cfiUpdate_afhob_afhob_1_bits_1 = 1'h0;
  end
  if (reset) begin
    do_redirect_bits_cfiUpdate_afhob_afhob_1_bits_2 = 1'h0;
  end
  if (reset) begin
    do_redirect_bits_cfiUpdate_afhob_afhob_1_bits_3 = 1'h0;
  end
  if (reset) begin
    do_redirect_bits_cfiUpdate_afhob_afhob_0_bits_0 = 1'h0;
  end
  if (reset) begin
    do_redirect_bits_cfiUpdate_afhob_afhob_0_bits_1 = 1'h0;
  end
  if (reset) begin
    do_redirect_bits_cfiUpdate_afhob_afhob_0_bits_2 = 1'h0;
  end
  if (reset) begin
    do_redirect_bits_cfiUpdate_afhob_afhob_0_bits_3 = 1'h0;
  end
  if (reset) begin
    do_redirect_bits_cfiUpdate_lastBrNumOH = 3'h0;
  end
  if (reset) begin
    do_redirect_bits_cfiUpdate_histPtr_flag = 1'h0;
  end
  if (reset) begin
    do_redirect_bits_cfiUpdate_histPtr_value = 8'h0;
  end
  if (reset) begin
    do_redirect_bits_cfiUpdate_target = 39'h0;
  end
  if (reset) begin
    do_redirect_bits_cfiUpdate_taken = 1'h0;
  end
  if (reset) begin
    do_redirect_bits_cfiUpdate_shift = 2'h0;
  end
  if (reset) begin
    do_redirect_bits_cfiUpdate_addIntoHist = 1'h0;
  end
  if (reset) begin
    previous_s2_pred_full_pred_br_taken_mask_1 = 1'h0;
  end
  if (reset) begin
    previous_s2_pred_full_pred_slot_valids_1 = 1'h0;
  end
  if (reset) begin
    previous_s2_pred_full_pred_is_br_sharing = 1'h0;
  end
  if (reset) begin
    previous_s2_pred_full_pred_hit = 1'h0;
  end
  if (reset) begin
    previous_s2_pred_full_pred_slot_valids_0 = 1'h0;
  end
  if (reset) begin
    previous_s2_pred_full_pred_br_taken_mask_0 = 1'h0;
  end
  if (reset) begin
    previous_s2_pred_full_pred_targets_0 = 39'h0;
  end
  if (reset) begin
    previous_s2_pred_full_pred_targets_1 = 39'h0;
  end
  if (reset) begin
    previous_s2_pred_full_pred_fallThroughAddr = 39'h0;
  end
  if (reset) begin
    previous_s2_pred_pc = 39'h0;
  end
  if (reset) begin
    previous_s1_pred_info_target = 39'h0;
  end
  if (reset) begin
    previous_s1_pred_info_lastBrPosOH = 3'h0;
  end
  if (reset) begin
    previous_s1_pred_info_taken = 1'h0;
  end
  if (reset) begin
    previous_s1_pred_info_cfiIndex = 3'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule

