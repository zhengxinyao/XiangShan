module PMPChecker(
  input  [1:0]  io_check_env_mode,
  input         io_check_env_pmp_0_cfg_l,
  input  [1:0]  io_check_env_pmp_0_cfg_a,
  input         io_check_env_pmp_0_cfg_x,
  input         io_check_env_pmp_0_cfg_w,
  input         io_check_env_pmp_0_cfg_r,
  input  [33:0] io_check_env_pmp_0_addr,
  input  [35:0] io_check_env_pmp_0_mask,
  input         io_check_env_pmp_1_cfg_l,
  input  [1:0]  io_check_env_pmp_1_cfg_a,
  input         io_check_env_pmp_1_cfg_x,
  input         io_check_env_pmp_1_cfg_w,
  input         io_check_env_pmp_1_cfg_r,
  input  [33:0] io_check_env_pmp_1_addr,
  input  [35:0] io_check_env_pmp_1_mask,
  input         io_check_env_pmp_2_cfg_l,
  input  [1:0]  io_check_env_pmp_2_cfg_a,
  input         io_check_env_pmp_2_cfg_x,
  input         io_check_env_pmp_2_cfg_w,
  input         io_check_env_pmp_2_cfg_r,
  input  [33:0] io_check_env_pmp_2_addr,
  input  [35:0] io_check_env_pmp_2_mask,
  input         io_check_env_pmp_3_cfg_l,
  input  [1:0]  io_check_env_pmp_3_cfg_a,
  input         io_check_env_pmp_3_cfg_x,
  input         io_check_env_pmp_3_cfg_w,
  input         io_check_env_pmp_3_cfg_r,
  input  [33:0] io_check_env_pmp_3_addr,
  input  [35:0] io_check_env_pmp_3_mask,
  input         io_check_env_pmp_4_cfg_l,
  input  [1:0]  io_check_env_pmp_4_cfg_a,
  input         io_check_env_pmp_4_cfg_x,
  input         io_check_env_pmp_4_cfg_w,
  input         io_check_env_pmp_4_cfg_r,
  input  [33:0] io_check_env_pmp_4_addr,
  input  [35:0] io_check_env_pmp_4_mask,
  input         io_check_env_pmp_5_cfg_l,
  input  [1:0]  io_check_env_pmp_5_cfg_a,
  input         io_check_env_pmp_5_cfg_x,
  input         io_check_env_pmp_5_cfg_w,
  input         io_check_env_pmp_5_cfg_r,
  input  [33:0] io_check_env_pmp_5_addr,
  input  [35:0] io_check_env_pmp_5_mask,
  input         io_check_env_pmp_6_cfg_l,
  input  [1:0]  io_check_env_pmp_6_cfg_a,
  input         io_check_env_pmp_6_cfg_x,
  input         io_check_env_pmp_6_cfg_w,
  input         io_check_env_pmp_6_cfg_r,
  input  [33:0] io_check_env_pmp_6_addr,
  input  [35:0] io_check_env_pmp_6_mask,
  input         io_check_env_pmp_7_cfg_l,
  input  [1:0]  io_check_env_pmp_7_cfg_a,
  input         io_check_env_pmp_7_cfg_x,
  input         io_check_env_pmp_7_cfg_w,
  input         io_check_env_pmp_7_cfg_r,
  input  [33:0] io_check_env_pmp_7_addr,
  input  [35:0] io_check_env_pmp_7_mask,
  input         io_check_env_pmp_8_cfg_l,
  input  [1:0]  io_check_env_pmp_8_cfg_a,
  input         io_check_env_pmp_8_cfg_x,
  input         io_check_env_pmp_8_cfg_w,
  input         io_check_env_pmp_8_cfg_r,
  input  [33:0] io_check_env_pmp_8_addr,
  input  [35:0] io_check_env_pmp_8_mask,
  input         io_check_env_pmp_9_cfg_l,
  input  [1:0]  io_check_env_pmp_9_cfg_a,
  input         io_check_env_pmp_9_cfg_x,
  input         io_check_env_pmp_9_cfg_w,
  input         io_check_env_pmp_9_cfg_r,
  input  [33:0] io_check_env_pmp_9_addr,
  input  [35:0] io_check_env_pmp_9_mask,
  input         io_check_env_pmp_10_cfg_l,
  input  [1:0]  io_check_env_pmp_10_cfg_a,
  input         io_check_env_pmp_10_cfg_x,
  input         io_check_env_pmp_10_cfg_w,
  input         io_check_env_pmp_10_cfg_r,
  input  [33:0] io_check_env_pmp_10_addr,
  input  [35:0] io_check_env_pmp_10_mask,
  input         io_check_env_pmp_11_cfg_l,
  input  [1:0]  io_check_env_pmp_11_cfg_a,
  input         io_check_env_pmp_11_cfg_x,
  input         io_check_env_pmp_11_cfg_w,
  input         io_check_env_pmp_11_cfg_r,
  input  [33:0] io_check_env_pmp_11_addr,
  input  [35:0] io_check_env_pmp_11_mask,
  input         io_check_env_pmp_12_cfg_l,
  input  [1:0]  io_check_env_pmp_12_cfg_a,
  input         io_check_env_pmp_12_cfg_x,
  input         io_check_env_pmp_12_cfg_w,
  input         io_check_env_pmp_12_cfg_r,
  input  [33:0] io_check_env_pmp_12_addr,
  input  [35:0] io_check_env_pmp_12_mask,
  input         io_check_env_pmp_13_cfg_l,
  input  [1:0]  io_check_env_pmp_13_cfg_a,
  input         io_check_env_pmp_13_cfg_x,
  input         io_check_env_pmp_13_cfg_w,
  input         io_check_env_pmp_13_cfg_r,
  input  [33:0] io_check_env_pmp_13_addr,
  input  [35:0] io_check_env_pmp_13_mask,
  input         io_check_env_pmp_14_cfg_l,
  input  [1:0]  io_check_env_pmp_14_cfg_a,
  input         io_check_env_pmp_14_cfg_x,
  input         io_check_env_pmp_14_cfg_w,
  input         io_check_env_pmp_14_cfg_r,
  input  [33:0] io_check_env_pmp_14_addr,
  input  [35:0] io_check_env_pmp_14_mask,
  input         io_check_env_pmp_15_cfg_l,
  input  [1:0]  io_check_env_pmp_15_cfg_a,
  input         io_check_env_pmp_15_cfg_x,
  input         io_check_env_pmp_15_cfg_w,
  input         io_check_env_pmp_15_cfg_r,
  input  [33:0] io_check_env_pmp_15_addr,
  input  [35:0] io_check_env_pmp_15_mask,
  input         io_check_env_pma_0_cfg_c,
  input         io_check_env_pma_0_cfg_atomic,
  input  [1:0]  io_check_env_pma_0_cfg_a,
  input         io_check_env_pma_0_cfg_x,
  input         io_check_env_pma_0_cfg_w,
  input         io_check_env_pma_0_cfg_r,
  input  [33:0] io_check_env_pma_0_addr,
  input  [35:0] io_check_env_pma_0_mask,
  input         io_check_env_pma_1_cfg_c,
  input         io_check_env_pma_1_cfg_atomic,
  input  [1:0]  io_check_env_pma_1_cfg_a,
  input         io_check_env_pma_1_cfg_x,
  input         io_check_env_pma_1_cfg_w,
  input         io_check_env_pma_1_cfg_r,
  input  [33:0] io_check_env_pma_1_addr,
  input  [35:0] io_check_env_pma_1_mask,
  input         io_check_env_pma_2_cfg_c,
  input         io_check_env_pma_2_cfg_atomic,
  input  [1:0]  io_check_env_pma_2_cfg_a,
  input         io_check_env_pma_2_cfg_x,
  input         io_check_env_pma_2_cfg_w,
  input         io_check_env_pma_2_cfg_r,
  input  [33:0] io_check_env_pma_2_addr,
  input  [35:0] io_check_env_pma_2_mask,
  input         io_check_env_pma_3_cfg_c,
  input         io_check_env_pma_3_cfg_atomic,
  input  [1:0]  io_check_env_pma_3_cfg_a,
  input         io_check_env_pma_3_cfg_x,
  input         io_check_env_pma_3_cfg_w,
  input         io_check_env_pma_3_cfg_r,
  input  [33:0] io_check_env_pma_3_addr,
  input  [35:0] io_check_env_pma_3_mask,
  input         io_check_env_pma_4_cfg_c,
  input         io_check_env_pma_4_cfg_atomic,
  input  [1:0]  io_check_env_pma_4_cfg_a,
  input         io_check_env_pma_4_cfg_x,
  input         io_check_env_pma_4_cfg_w,
  input         io_check_env_pma_4_cfg_r,
  input  [33:0] io_check_env_pma_4_addr,
  input  [35:0] io_check_env_pma_4_mask,
  input         io_check_env_pma_5_cfg_c,
  input         io_check_env_pma_5_cfg_atomic,
  input  [1:0]  io_check_env_pma_5_cfg_a,
  input         io_check_env_pma_5_cfg_x,
  input         io_check_env_pma_5_cfg_w,
  input         io_check_env_pma_5_cfg_r,
  input  [33:0] io_check_env_pma_5_addr,
  input  [35:0] io_check_env_pma_5_mask,
  input         io_check_env_pma_6_cfg_c,
  input         io_check_env_pma_6_cfg_atomic,
  input  [1:0]  io_check_env_pma_6_cfg_a,
  input         io_check_env_pma_6_cfg_x,
  input         io_check_env_pma_6_cfg_w,
  input         io_check_env_pma_6_cfg_r,
  input  [33:0] io_check_env_pma_6_addr,
  input  [35:0] io_check_env_pma_6_mask,
  input         io_check_env_pma_7_cfg_c,
  input         io_check_env_pma_7_cfg_atomic,
  input  [1:0]  io_check_env_pma_7_cfg_a,
  input         io_check_env_pma_7_cfg_x,
  input         io_check_env_pma_7_cfg_w,
  input         io_check_env_pma_7_cfg_r,
  input  [33:0] io_check_env_pma_7_addr,
  input  [35:0] io_check_env_pma_7_mask,
  input         io_check_env_pma_8_cfg_c,
  input         io_check_env_pma_8_cfg_atomic,
  input  [1:0]  io_check_env_pma_8_cfg_a,
  input         io_check_env_pma_8_cfg_x,
  input         io_check_env_pma_8_cfg_w,
  input         io_check_env_pma_8_cfg_r,
  input  [33:0] io_check_env_pma_8_addr,
  input  [35:0] io_check_env_pma_8_mask,
  input         io_check_env_pma_9_cfg_c,
  input         io_check_env_pma_9_cfg_atomic,
  input  [1:0]  io_check_env_pma_9_cfg_a,
  input         io_check_env_pma_9_cfg_x,
  input         io_check_env_pma_9_cfg_w,
  input         io_check_env_pma_9_cfg_r,
  input  [33:0] io_check_env_pma_9_addr,
  input  [35:0] io_check_env_pma_9_mask,
  input         io_check_env_pma_10_cfg_c,
  input         io_check_env_pma_10_cfg_atomic,
  input  [1:0]  io_check_env_pma_10_cfg_a,
  input         io_check_env_pma_10_cfg_x,
  input         io_check_env_pma_10_cfg_w,
  input         io_check_env_pma_10_cfg_r,
  input  [33:0] io_check_env_pma_10_addr,
  input  [35:0] io_check_env_pma_10_mask,
  input         io_check_env_pma_11_cfg_c,
  input         io_check_env_pma_11_cfg_atomic,
  input  [1:0]  io_check_env_pma_11_cfg_a,
  input         io_check_env_pma_11_cfg_x,
  input         io_check_env_pma_11_cfg_w,
  input         io_check_env_pma_11_cfg_r,
  input  [33:0] io_check_env_pma_11_addr,
  input  [35:0] io_check_env_pma_11_mask,
  input         io_check_env_pma_12_cfg_c,
  input         io_check_env_pma_12_cfg_atomic,
  input  [1:0]  io_check_env_pma_12_cfg_a,
  input         io_check_env_pma_12_cfg_x,
  input         io_check_env_pma_12_cfg_w,
  input         io_check_env_pma_12_cfg_r,
  input  [33:0] io_check_env_pma_12_addr,
  input  [35:0] io_check_env_pma_12_mask,
  input         io_check_env_pma_13_cfg_c,
  input         io_check_env_pma_13_cfg_atomic,
  input  [1:0]  io_check_env_pma_13_cfg_a,
  input         io_check_env_pma_13_cfg_x,
  input         io_check_env_pma_13_cfg_w,
  input         io_check_env_pma_13_cfg_r,
  input  [33:0] io_check_env_pma_13_addr,
  input  [35:0] io_check_env_pma_13_mask,
  input         io_check_env_pma_14_cfg_c,
  input         io_check_env_pma_14_cfg_atomic,
  input  [1:0]  io_check_env_pma_14_cfg_a,
  input         io_check_env_pma_14_cfg_x,
  input         io_check_env_pma_14_cfg_w,
  input         io_check_env_pma_14_cfg_r,
  input  [33:0] io_check_env_pma_14_addr,
  input  [35:0] io_check_env_pma_14_mask,
  input         io_check_env_pma_15_cfg_c,
  input         io_check_env_pma_15_cfg_atomic,
  input  [1:0]  io_check_env_pma_15_cfg_a,
  input         io_check_env_pma_15_cfg_x,
  input         io_check_env_pma_15_cfg_w,
  input         io_check_env_pma_15_cfg_r,
  input  [33:0] io_check_env_pma_15_addr,
  input  [35:0] io_check_env_pma_15_mask,
  input  [35:0] io_req_bits_addr,
  input  [2:0]  io_req_bits_cmd,
  output        io_resp_ld,
  output        io_resp_st,
  output        io_resp_instr,
  output        io_resp_mmio,
  output        io_resp_atomic
);
  wire  res_pmp_passThrough = io_check_env_mode > 2'h1; // @[PMP.scala 423:65]
  wire [35:0] _res_pmp_is_match_T_1 = {io_check_env_pmp_0_addr, 2'h0}; // @[PMP.scala 190:35]
  wire [35:0] _res_pmp_is_match_T_3 = _res_pmp_is_match_T_1 & 36'hffffff000; // @[PMP.scala 190:50]
  wire [35:0] _res_pmp_is_match_T_4 = ~io_check_env_pmp_0_mask; // @[PMP.scala 232:10]
  wire [35:0] _res_pmp_is_match_T_5 = io_req_bits_addr & _res_pmp_is_match_T_4; // @[PMP.scala 232:8]
  wire [35:0] _res_pmp_is_match_T_7 = _res_pmp_is_match_T_3 & _res_pmp_is_match_T_4; // @[PMP.scala 232:21]
  wire  _res_pmp_is_match_T_8 = _res_pmp_is_match_T_5 == _res_pmp_is_match_T_7; // @[PMP.scala 232:14]
  wire  _res_pmp_is_match_T_9 = io_check_env_pmp_0_cfg_a == 2'h1; // @[PMP.scala 53:15]
  wire  _res_pmp_is_match_T_18 = io_req_bits_addr < _res_pmp_is_match_T_3; // @[PMP.scala 210:14]
  wire  _res_pmp_is_match_T_20 = _res_pmp_is_match_T_9 & _res_pmp_is_match_T_18; // @[PMP.scala 200:10]
  wire  res_pmp_is_match = io_check_env_pmp_0_cfg_a[1] ? _res_pmp_is_match_T_8 : _res_pmp_is_match_T_20; // @[PMP.scala 199:8]
  wire  res_pmp_ignore = res_pmp_passThrough & ~io_check_env_pmp_0_cfg_l; // @[PMP.scala 434:32]
  wire  res_pmp_cur_cfg_r = io_check_env_pmp_0_cfg_r | res_pmp_ignore; // @[PMP.scala 438:42]
  wire  res_pmp_cur_cfg_w = io_check_env_pmp_0_cfg_w | res_pmp_ignore; // @[PMP.scala 439:42]
  wire  res_pmp_cur_cfg_x = io_check_env_pmp_0_cfg_x | res_pmp_ignore; // @[PMP.scala 440:42]
  wire [35:0] _res_pmp_is_match_T_22 = {io_check_env_pmp_1_addr, 2'h0}; // @[PMP.scala 190:35]
  wire [35:0] _res_pmp_is_match_T_24 = _res_pmp_is_match_T_22 & 36'hffffff000; // @[PMP.scala 190:50]
  wire [35:0] _res_pmp_is_match_T_25 = ~io_check_env_pmp_1_mask; // @[PMP.scala 232:10]
  wire [35:0] _res_pmp_is_match_T_26 = io_req_bits_addr & _res_pmp_is_match_T_25; // @[PMP.scala 232:8]
  wire [35:0] _res_pmp_is_match_T_28 = _res_pmp_is_match_T_24 & _res_pmp_is_match_T_25; // @[PMP.scala 232:21]
  wire  _res_pmp_is_match_T_29 = _res_pmp_is_match_T_26 == _res_pmp_is_match_T_28; // @[PMP.scala 232:14]
  wire  _res_pmp_is_match_T_30 = io_check_env_pmp_1_cfg_a == 2'h1; // @[PMP.scala 53:15]
  wire  _res_pmp_is_match_T_35 = ~_res_pmp_is_match_T_18; // @[PMP.scala 220:5]
  wire  _res_pmp_is_match_T_39 = io_req_bits_addr < _res_pmp_is_match_T_24; // @[PMP.scala 210:14]
  wire  _res_pmp_is_match_T_40 = _res_pmp_is_match_T_35 & _res_pmp_is_match_T_39; // @[PMP.scala 228:56]
  wire  _res_pmp_is_match_T_41 = _res_pmp_is_match_T_30 & _res_pmp_is_match_T_40; // @[PMP.scala 200:10]
  wire  res_pmp_is_match_1 = io_check_env_pmp_1_cfg_a[1] ? _res_pmp_is_match_T_29 : _res_pmp_is_match_T_41; // @[PMP.scala 199:8]
  wire  res_pmp_ignore_1 = res_pmp_passThrough & ~io_check_env_pmp_1_cfg_l; // @[PMP.scala 434:32]
  wire  res_pmp_cur_1_cfg_r = io_check_env_pmp_1_cfg_r | res_pmp_ignore_1; // @[PMP.scala 438:42]
  wire  res_pmp_cur_1_cfg_w = io_check_env_pmp_1_cfg_w | res_pmp_ignore_1; // @[PMP.scala 439:42]
  wire  res_pmp_cur_1_cfg_x = io_check_env_pmp_1_cfg_x | res_pmp_ignore_1; // @[PMP.scala 440:42]
  wire [35:0] _res_pmp_is_match_T_43 = {io_check_env_pmp_2_addr, 2'h0}; // @[PMP.scala 190:35]
  wire [35:0] _res_pmp_is_match_T_45 = _res_pmp_is_match_T_43 & 36'hffffff000; // @[PMP.scala 190:50]
  wire [35:0] _res_pmp_is_match_T_46 = ~io_check_env_pmp_2_mask; // @[PMP.scala 232:10]
  wire [35:0] _res_pmp_is_match_T_47 = io_req_bits_addr & _res_pmp_is_match_T_46; // @[PMP.scala 232:8]
  wire [35:0] _res_pmp_is_match_T_49 = _res_pmp_is_match_T_45 & _res_pmp_is_match_T_46; // @[PMP.scala 232:21]
  wire  _res_pmp_is_match_T_50 = _res_pmp_is_match_T_47 == _res_pmp_is_match_T_49; // @[PMP.scala 232:14]
  wire  _res_pmp_is_match_T_51 = io_check_env_pmp_2_cfg_a == 2'h1; // @[PMP.scala 53:15]
  wire  _res_pmp_is_match_T_56 = ~_res_pmp_is_match_T_39; // @[PMP.scala 220:5]
  wire  _res_pmp_is_match_T_60 = io_req_bits_addr < _res_pmp_is_match_T_45; // @[PMP.scala 210:14]
  wire  _res_pmp_is_match_T_61 = _res_pmp_is_match_T_56 & _res_pmp_is_match_T_60; // @[PMP.scala 228:56]
  wire  _res_pmp_is_match_T_62 = _res_pmp_is_match_T_51 & _res_pmp_is_match_T_61; // @[PMP.scala 200:10]
  wire  res_pmp_is_match_2 = io_check_env_pmp_2_cfg_a[1] ? _res_pmp_is_match_T_50 : _res_pmp_is_match_T_62; // @[PMP.scala 199:8]
  wire  res_pmp_ignore_2 = res_pmp_passThrough & ~io_check_env_pmp_2_cfg_l; // @[PMP.scala 434:32]
  wire  res_pmp_cur_2_cfg_r = io_check_env_pmp_2_cfg_r | res_pmp_ignore_2; // @[PMP.scala 438:42]
  wire  res_pmp_cur_2_cfg_w = io_check_env_pmp_2_cfg_w | res_pmp_ignore_2; // @[PMP.scala 439:42]
  wire  res_pmp_cur_2_cfg_x = io_check_env_pmp_2_cfg_x | res_pmp_ignore_2; // @[PMP.scala 440:42]
  wire [35:0] _res_pmp_is_match_T_64 = {io_check_env_pmp_3_addr, 2'h0}; // @[PMP.scala 190:35]
  wire [35:0] _res_pmp_is_match_T_66 = _res_pmp_is_match_T_64 & 36'hffffff000; // @[PMP.scala 190:50]
  wire [35:0] _res_pmp_is_match_T_67 = ~io_check_env_pmp_3_mask; // @[PMP.scala 232:10]
  wire [35:0] _res_pmp_is_match_T_68 = io_req_bits_addr & _res_pmp_is_match_T_67; // @[PMP.scala 232:8]
  wire [35:0] _res_pmp_is_match_T_70 = _res_pmp_is_match_T_66 & _res_pmp_is_match_T_67; // @[PMP.scala 232:21]
  wire  _res_pmp_is_match_T_71 = _res_pmp_is_match_T_68 == _res_pmp_is_match_T_70; // @[PMP.scala 232:14]
  wire  _res_pmp_is_match_T_72 = io_check_env_pmp_3_cfg_a == 2'h1; // @[PMP.scala 53:15]
  wire  _res_pmp_is_match_T_77 = ~_res_pmp_is_match_T_60; // @[PMP.scala 220:5]
  wire  _res_pmp_is_match_T_81 = io_req_bits_addr < _res_pmp_is_match_T_66; // @[PMP.scala 210:14]
  wire  _res_pmp_is_match_T_82 = _res_pmp_is_match_T_77 & _res_pmp_is_match_T_81; // @[PMP.scala 228:56]
  wire  _res_pmp_is_match_T_83 = _res_pmp_is_match_T_72 & _res_pmp_is_match_T_82; // @[PMP.scala 200:10]
  wire  res_pmp_is_match_3 = io_check_env_pmp_3_cfg_a[1] ? _res_pmp_is_match_T_71 : _res_pmp_is_match_T_83; // @[PMP.scala 199:8]
  wire  res_pmp_ignore_3 = res_pmp_passThrough & ~io_check_env_pmp_3_cfg_l; // @[PMP.scala 434:32]
  wire  res_pmp_cur_3_cfg_r = io_check_env_pmp_3_cfg_r | res_pmp_ignore_3; // @[PMP.scala 438:42]
  wire  res_pmp_cur_3_cfg_w = io_check_env_pmp_3_cfg_w | res_pmp_ignore_3; // @[PMP.scala 439:42]
  wire  res_pmp_cur_3_cfg_x = io_check_env_pmp_3_cfg_x | res_pmp_ignore_3; // @[PMP.scala 440:42]
  wire [35:0] _res_pmp_is_match_T_85 = {io_check_env_pmp_4_addr, 2'h0}; // @[PMP.scala 190:35]
  wire [35:0] _res_pmp_is_match_T_87 = _res_pmp_is_match_T_85 & 36'hffffff000; // @[PMP.scala 190:50]
  wire [35:0] _res_pmp_is_match_T_88 = ~io_check_env_pmp_4_mask; // @[PMP.scala 232:10]
  wire [35:0] _res_pmp_is_match_T_89 = io_req_bits_addr & _res_pmp_is_match_T_88; // @[PMP.scala 232:8]
  wire [35:0] _res_pmp_is_match_T_91 = _res_pmp_is_match_T_87 & _res_pmp_is_match_T_88; // @[PMP.scala 232:21]
  wire  _res_pmp_is_match_T_92 = _res_pmp_is_match_T_89 == _res_pmp_is_match_T_91; // @[PMP.scala 232:14]
  wire  _res_pmp_is_match_T_93 = io_check_env_pmp_4_cfg_a == 2'h1; // @[PMP.scala 53:15]
  wire  _res_pmp_is_match_T_98 = ~_res_pmp_is_match_T_81; // @[PMP.scala 220:5]
  wire  _res_pmp_is_match_T_102 = io_req_bits_addr < _res_pmp_is_match_T_87; // @[PMP.scala 210:14]
  wire  _res_pmp_is_match_T_103 = _res_pmp_is_match_T_98 & _res_pmp_is_match_T_102; // @[PMP.scala 228:56]
  wire  _res_pmp_is_match_T_104 = _res_pmp_is_match_T_93 & _res_pmp_is_match_T_103; // @[PMP.scala 200:10]
  wire  res_pmp_is_match_4 = io_check_env_pmp_4_cfg_a[1] ? _res_pmp_is_match_T_92 : _res_pmp_is_match_T_104; // @[PMP.scala 199:8]
  wire  res_pmp_ignore_4 = res_pmp_passThrough & ~io_check_env_pmp_4_cfg_l; // @[PMP.scala 434:32]
  wire  res_pmp_cur_4_cfg_r = io_check_env_pmp_4_cfg_r | res_pmp_ignore_4; // @[PMP.scala 438:42]
  wire  res_pmp_cur_4_cfg_w = io_check_env_pmp_4_cfg_w | res_pmp_ignore_4; // @[PMP.scala 439:42]
  wire  res_pmp_cur_4_cfg_x = io_check_env_pmp_4_cfg_x | res_pmp_ignore_4; // @[PMP.scala 440:42]
  wire [35:0] _res_pmp_is_match_T_106 = {io_check_env_pmp_5_addr, 2'h0}; // @[PMP.scala 190:35]
  wire [35:0] _res_pmp_is_match_T_108 = _res_pmp_is_match_T_106 & 36'hffffff000; // @[PMP.scala 190:50]
  wire [35:0] _res_pmp_is_match_T_109 = ~io_check_env_pmp_5_mask; // @[PMP.scala 232:10]
  wire [35:0] _res_pmp_is_match_T_110 = io_req_bits_addr & _res_pmp_is_match_T_109; // @[PMP.scala 232:8]
  wire [35:0] _res_pmp_is_match_T_112 = _res_pmp_is_match_T_108 & _res_pmp_is_match_T_109; // @[PMP.scala 232:21]
  wire  _res_pmp_is_match_T_113 = _res_pmp_is_match_T_110 == _res_pmp_is_match_T_112; // @[PMP.scala 232:14]
  wire  _res_pmp_is_match_T_114 = io_check_env_pmp_5_cfg_a == 2'h1; // @[PMP.scala 53:15]
  wire  _res_pmp_is_match_T_119 = ~_res_pmp_is_match_T_102; // @[PMP.scala 220:5]
  wire  _res_pmp_is_match_T_123 = io_req_bits_addr < _res_pmp_is_match_T_108; // @[PMP.scala 210:14]
  wire  _res_pmp_is_match_T_124 = _res_pmp_is_match_T_119 & _res_pmp_is_match_T_123; // @[PMP.scala 228:56]
  wire  _res_pmp_is_match_T_125 = _res_pmp_is_match_T_114 & _res_pmp_is_match_T_124; // @[PMP.scala 200:10]
  wire  res_pmp_is_match_5 = io_check_env_pmp_5_cfg_a[1] ? _res_pmp_is_match_T_113 : _res_pmp_is_match_T_125; // @[PMP.scala 199:8]
  wire  res_pmp_ignore_5 = res_pmp_passThrough & ~io_check_env_pmp_5_cfg_l; // @[PMP.scala 434:32]
  wire  res_pmp_cur_5_cfg_r = io_check_env_pmp_5_cfg_r | res_pmp_ignore_5; // @[PMP.scala 438:42]
  wire  res_pmp_cur_5_cfg_w = io_check_env_pmp_5_cfg_w | res_pmp_ignore_5; // @[PMP.scala 439:42]
  wire  res_pmp_cur_5_cfg_x = io_check_env_pmp_5_cfg_x | res_pmp_ignore_5; // @[PMP.scala 440:42]
  wire [35:0] _res_pmp_is_match_T_127 = {io_check_env_pmp_6_addr, 2'h0}; // @[PMP.scala 190:35]
  wire [35:0] _res_pmp_is_match_T_129 = _res_pmp_is_match_T_127 & 36'hffffff000; // @[PMP.scala 190:50]
  wire [35:0] _res_pmp_is_match_T_130 = ~io_check_env_pmp_6_mask; // @[PMP.scala 232:10]
  wire [35:0] _res_pmp_is_match_T_131 = io_req_bits_addr & _res_pmp_is_match_T_130; // @[PMP.scala 232:8]
  wire [35:0] _res_pmp_is_match_T_133 = _res_pmp_is_match_T_129 & _res_pmp_is_match_T_130; // @[PMP.scala 232:21]
  wire  _res_pmp_is_match_T_134 = _res_pmp_is_match_T_131 == _res_pmp_is_match_T_133; // @[PMP.scala 232:14]
  wire  _res_pmp_is_match_T_135 = io_check_env_pmp_6_cfg_a == 2'h1; // @[PMP.scala 53:15]
  wire  _res_pmp_is_match_T_140 = ~_res_pmp_is_match_T_123; // @[PMP.scala 220:5]
  wire  _res_pmp_is_match_T_144 = io_req_bits_addr < _res_pmp_is_match_T_129; // @[PMP.scala 210:14]
  wire  _res_pmp_is_match_T_145 = _res_pmp_is_match_T_140 & _res_pmp_is_match_T_144; // @[PMP.scala 228:56]
  wire  _res_pmp_is_match_T_146 = _res_pmp_is_match_T_135 & _res_pmp_is_match_T_145; // @[PMP.scala 200:10]
  wire  res_pmp_is_match_6 = io_check_env_pmp_6_cfg_a[1] ? _res_pmp_is_match_T_134 : _res_pmp_is_match_T_146; // @[PMP.scala 199:8]
  wire  res_pmp_ignore_6 = res_pmp_passThrough & ~io_check_env_pmp_6_cfg_l; // @[PMP.scala 434:32]
  wire  res_pmp_cur_6_cfg_r = io_check_env_pmp_6_cfg_r | res_pmp_ignore_6; // @[PMP.scala 438:42]
  wire  res_pmp_cur_6_cfg_w = io_check_env_pmp_6_cfg_w | res_pmp_ignore_6; // @[PMP.scala 439:42]
  wire  res_pmp_cur_6_cfg_x = io_check_env_pmp_6_cfg_x | res_pmp_ignore_6; // @[PMP.scala 440:42]
  wire [35:0] _res_pmp_is_match_T_148 = {io_check_env_pmp_7_addr, 2'h0}; // @[PMP.scala 190:35]
  wire [35:0] _res_pmp_is_match_T_150 = _res_pmp_is_match_T_148 & 36'hffffff000; // @[PMP.scala 190:50]
  wire [35:0] _res_pmp_is_match_T_151 = ~io_check_env_pmp_7_mask; // @[PMP.scala 232:10]
  wire [35:0] _res_pmp_is_match_T_152 = io_req_bits_addr & _res_pmp_is_match_T_151; // @[PMP.scala 232:8]
  wire [35:0] _res_pmp_is_match_T_154 = _res_pmp_is_match_T_150 & _res_pmp_is_match_T_151; // @[PMP.scala 232:21]
  wire  _res_pmp_is_match_T_155 = _res_pmp_is_match_T_152 == _res_pmp_is_match_T_154; // @[PMP.scala 232:14]
  wire  _res_pmp_is_match_T_156 = io_check_env_pmp_7_cfg_a == 2'h1; // @[PMP.scala 53:15]
  wire  _res_pmp_is_match_T_161 = ~_res_pmp_is_match_T_144; // @[PMP.scala 220:5]
  wire  _res_pmp_is_match_T_165 = io_req_bits_addr < _res_pmp_is_match_T_150; // @[PMP.scala 210:14]
  wire  _res_pmp_is_match_T_166 = _res_pmp_is_match_T_161 & _res_pmp_is_match_T_165; // @[PMP.scala 228:56]
  wire  _res_pmp_is_match_T_167 = _res_pmp_is_match_T_156 & _res_pmp_is_match_T_166; // @[PMP.scala 200:10]
  wire  res_pmp_is_match_7 = io_check_env_pmp_7_cfg_a[1] ? _res_pmp_is_match_T_155 : _res_pmp_is_match_T_167; // @[PMP.scala 199:8]
  wire  res_pmp_ignore_7 = res_pmp_passThrough & ~io_check_env_pmp_7_cfg_l; // @[PMP.scala 434:32]
  wire  res_pmp_cur_7_cfg_r = io_check_env_pmp_7_cfg_r | res_pmp_ignore_7; // @[PMP.scala 438:42]
  wire  res_pmp_cur_7_cfg_w = io_check_env_pmp_7_cfg_w | res_pmp_ignore_7; // @[PMP.scala 439:42]
  wire  res_pmp_cur_7_cfg_x = io_check_env_pmp_7_cfg_x | res_pmp_ignore_7; // @[PMP.scala 440:42]
  wire [35:0] _res_pmp_is_match_T_169 = {io_check_env_pmp_8_addr, 2'h0}; // @[PMP.scala 190:35]
  wire [35:0] _res_pmp_is_match_T_171 = _res_pmp_is_match_T_169 & 36'hffffff000; // @[PMP.scala 190:50]
  wire [35:0] _res_pmp_is_match_T_172 = ~io_check_env_pmp_8_mask; // @[PMP.scala 232:10]
  wire [35:0] _res_pmp_is_match_T_173 = io_req_bits_addr & _res_pmp_is_match_T_172; // @[PMP.scala 232:8]
  wire [35:0] _res_pmp_is_match_T_175 = _res_pmp_is_match_T_171 & _res_pmp_is_match_T_172; // @[PMP.scala 232:21]
  wire  _res_pmp_is_match_T_176 = _res_pmp_is_match_T_173 == _res_pmp_is_match_T_175; // @[PMP.scala 232:14]
  wire  _res_pmp_is_match_T_177 = io_check_env_pmp_8_cfg_a == 2'h1; // @[PMP.scala 53:15]
  wire  _res_pmp_is_match_T_182 = ~_res_pmp_is_match_T_165; // @[PMP.scala 220:5]
  wire  _res_pmp_is_match_T_186 = io_req_bits_addr < _res_pmp_is_match_T_171; // @[PMP.scala 210:14]
  wire  _res_pmp_is_match_T_187 = _res_pmp_is_match_T_182 & _res_pmp_is_match_T_186; // @[PMP.scala 228:56]
  wire  _res_pmp_is_match_T_188 = _res_pmp_is_match_T_177 & _res_pmp_is_match_T_187; // @[PMP.scala 200:10]
  wire  res_pmp_is_match_8 = io_check_env_pmp_8_cfg_a[1] ? _res_pmp_is_match_T_176 : _res_pmp_is_match_T_188; // @[PMP.scala 199:8]
  wire  res_pmp_ignore_8 = res_pmp_passThrough & ~io_check_env_pmp_8_cfg_l; // @[PMP.scala 434:32]
  wire  res_pmp_cur_8_cfg_r = io_check_env_pmp_8_cfg_r | res_pmp_ignore_8; // @[PMP.scala 438:42]
  wire  res_pmp_cur_8_cfg_w = io_check_env_pmp_8_cfg_w | res_pmp_ignore_8; // @[PMP.scala 439:42]
  wire  res_pmp_cur_8_cfg_x = io_check_env_pmp_8_cfg_x | res_pmp_ignore_8; // @[PMP.scala 440:42]
  wire [35:0] _res_pmp_is_match_T_190 = {io_check_env_pmp_9_addr, 2'h0}; // @[PMP.scala 190:35]
  wire [35:0] _res_pmp_is_match_T_192 = _res_pmp_is_match_T_190 & 36'hffffff000; // @[PMP.scala 190:50]
  wire [35:0] _res_pmp_is_match_T_193 = ~io_check_env_pmp_9_mask; // @[PMP.scala 232:10]
  wire [35:0] _res_pmp_is_match_T_194 = io_req_bits_addr & _res_pmp_is_match_T_193; // @[PMP.scala 232:8]
  wire [35:0] _res_pmp_is_match_T_196 = _res_pmp_is_match_T_192 & _res_pmp_is_match_T_193; // @[PMP.scala 232:21]
  wire  _res_pmp_is_match_T_197 = _res_pmp_is_match_T_194 == _res_pmp_is_match_T_196; // @[PMP.scala 232:14]
  wire  _res_pmp_is_match_T_198 = io_check_env_pmp_9_cfg_a == 2'h1; // @[PMP.scala 53:15]
  wire  _res_pmp_is_match_T_203 = ~_res_pmp_is_match_T_186; // @[PMP.scala 220:5]
  wire  _res_pmp_is_match_T_207 = io_req_bits_addr < _res_pmp_is_match_T_192; // @[PMP.scala 210:14]
  wire  _res_pmp_is_match_T_208 = _res_pmp_is_match_T_203 & _res_pmp_is_match_T_207; // @[PMP.scala 228:56]
  wire  _res_pmp_is_match_T_209 = _res_pmp_is_match_T_198 & _res_pmp_is_match_T_208; // @[PMP.scala 200:10]
  wire  res_pmp_is_match_9 = io_check_env_pmp_9_cfg_a[1] ? _res_pmp_is_match_T_197 : _res_pmp_is_match_T_209; // @[PMP.scala 199:8]
  wire  res_pmp_ignore_9 = res_pmp_passThrough & ~io_check_env_pmp_9_cfg_l; // @[PMP.scala 434:32]
  wire  res_pmp_cur_9_cfg_r = io_check_env_pmp_9_cfg_r | res_pmp_ignore_9; // @[PMP.scala 438:42]
  wire  res_pmp_cur_9_cfg_w = io_check_env_pmp_9_cfg_w | res_pmp_ignore_9; // @[PMP.scala 439:42]
  wire  res_pmp_cur_9_cfg_x = io_check_env_pmp_9_cfg_x | res_pmp_ignore_9; // @[PMP.scala 440:42]
  wire [35:0] _res_pmp_is_match_T_211 = {io_check_env_pmp_10_addr, 2'h0}; // @[PMP.scala 190:35]
  wire [35:0] _res_pmp_is_match_T_213 = _res_pmp_is_match_T_211 & 36'hffffff000; // @[PMP.scala 190:50]
  wire [35:0] _res_pmp_is_match_T_214 = ~io_check_env_pmp_10_mask; // @[PMP.scala 232:10]
  wire [35:0] _res_pmp_is_match_T_215 = io_req_bits_addr & _res_pmp_is_match_T_214; // @[PMP.scala 232:8]
  wire [35:0] _res_pmp_is_match_T_217 = _res_pmp_is_match_T_213 & _res_pmp_is_match_T_214; // @[PMP.scala 232:21]
  wire  _res_pmp_is_match_T_218 = _res_pmp_is_match_T_215 == _res_pmp_is_match_T_217; // @[PMP.scala 232:14]
  wire  _res_pmp_is_match_T_219 = io_check_env_pmp_10_cfg_a == 2'h1; // @[PMP.scala 53:15]
  wire  _res_pmp_is_match_T_224 = ~_res_pmp_is_match_T_207; // @[PMP.scala 220:5]
  wire  _res_pmp_is_match_T_228 = io_req_bits_addr < _res_pmp_is_match_T_213; // @[PMP.scala 210:14]
  wire  _res_pmp_is_match_T_229 = _res_pmp_is_match_T_224 & _res_pmp_is_match_T_228; // @[PMP.scala 228:56]
  wire  _res_pmp_is_match_T_230 = _res_pmp_is_match_T_219 & _res_pmp_is_match_T_229; // @[PMP.scala 200:10]
  wire  res_pmp_is_match_10 = io_check_env_pmp_10_cfg_a[1] ? _res_pmp_is_match_T_218 : _res_pmp_is_match_T_230; // @[PMP.scala 199:8]
  wire  res_pmp_ignore_10 = res_pmp_passThrough & ~io_check_env_pmp_10_cfg_l; // @[PMP.scala 434:32]
  wire  res_pmp_cur_10_cfg_r = io_check_env_pmp_10_cfg_r | res_pmp_ignore_10; // @[PMP.scala 438:42]
  wire  res_pmp_cur_10_cfg_w = io_check_env_pmp_10_cfg_w | res_pmp_ignore_10; // @[PMP.scala 439:42]
  wire  res_pmp_cur_10_cfg_x = io_check_env_pmp_10_cfg_x | res_pmp_ignore_10; // @[PMP.scala 440:42]
  wire [35:0] _res_pmp_is_match_T_232 = {io_check_env_pmp_11_addr, 2'h0}; // @[PMP.scala 190:35]
  wire [35:0] _res_pmp_is_match_T_234 = _res_pmp_is_match_T_232 & 36'hffffff000; // @[PMP.scala 190:50]
  wire [35:0] _res_pmp_is_match_T_235 = ~io_check_env_pmp_11_mask; // @[PMP.scala 232:10]
  wire [35:0] _res_pmp_is_match_T_236 = io_req_bits_addr & _res_pmp_is_match_T_235; // @[PMP.scala 232:8]
  wire [35:0] _res_pmp_is_match_T_238 = _res_pmp_is_match_T_234 & _res_pmp_is_match_T_235; // @[PMP.scala 232:21]
  wire  _res_pmp_is_match_T_239 = _res_pmp_is_match_T_236 == _res_pmp_is_match_T_238; // @[PMP.scala 232:14]
  wire  _res_pmp_is_match_T_240 = io_check_env_pmp_11_cfg_a == 2'h1; // @[PMP.scala 53:15]
  wire  _res_pmp_is_match_T_245 = ~_res_pmp_is_match_T_228; // @[PMP.scala 220:5]
  wire  _res_pmp_is_match_T_249 = io_req_bits_addr < _res_pmp_is_match_T_234; // @[PMP.scala 210:14]
  wire  _res_pmp_is_match_T_250 = _res_pmp_is_match_T_245 & _res_pmp_is_match_T_249; // @[PMP.scala 228:56]
  wire  _res_pmp_is_match_T_251 = _res_pmp_is_match_T_240 & _res_pmp_is_match_T_250; // @[PMP.scala 200:10]
  wire  res_pmp_is_match_11 = io_check_env_pmp_11_cfg_a[1] ? _res_pmp_is_match_T_239 : _res_pmp_is_match_T_251; // @[PMP.scala 199:8]
  wire  res_pmp_ignore_11 = res_pmp_passThrough & ~io_check_env_pmp_11_cfg_l; // @[PMP.scala 434:32]
  wire  res_pmp_cur_11_cfg_r = io_check_env_pmp_11_cfg_r | res_pmp_ignore_11; // @[PMP.scala 438:42]
  wire  res_pmp_cur_11_cfg_w = io_check_env_pmp_11_cfg_w | res_pmp_ignore_11; // @[PMP.scala 439:42]
  wire  res_pmp_cur_11_cfg_x = io_check_env_pmp_11_cfg_x | res_pmp_ignore_11; // @[PMP.scala 440:42]
  wire [35:0] _res_pmp_is_match_T_253 = {io_check_env_pmp_12_addr, 2'h0}; // @[PMP.scala 190:35]
  wire [35:0] _res_pmp_is_match_T_255 = _res_pmp_is_match_T_253 & 36'hffffff000; // @[PMP.scala 190:50]
  wire [35:0] _res_pmp_is_match_T_256 = ~io_check_env_pmp_12_mask; // @[PMP.scala 232:10]
  wire [35:0] _res_pmp_is_match_T_257 = io_req_bits_addr & _res_pmp_is_match_T_256; // @[PMP.scala 232:8]
  wire [35:0] _res_pmp_is_match_T_259 = _res_pmp_is_match_T_255 & _res_pmp_is_match_T_256; // @[PMP.scala 232:21]
  wire  _res_pmp_is_match_T_260 = _res_pmp_is_match_T_257 == _res_pmp_is_match_T_259; // @[PMP.scala 232:14]
  wire  _res_pmp_is_match_T_261 = io_check_env_pmp_12_cfg_a == 2'h1; // @[PMP.scala 53:15]
  wire  _res_pmp_is_match_T_266 = ~_res_pmp_is_match_T_249; // @[PMP.scala 220:5]
  wire  _res_pmp_is_match_T_270 = io_req_bits_addr < _res_pmp_is_match_T_255; // @[PMP.scala 210:14]
  wire  _res_pmp_is_match_T_271 = _res_pmp_is_match_T_266 & _res_pmp_is_match_T_270; // @[PMP.scala 228:56]
  wire  _res_pmp_is_match_T_272 = _res_pmp_is_match_T_261 & _res_pmp_is_match_T_271; // @[PMP.scala 200:10]
  wire  res_pmp_is_match_12 = io_check_env_pmp_12_cfg_a[1] ? _res_pmp_is_match_T_260 : _res_pmp_is_match_T_272; // @[PMP.scala 199:8]
  wire  res_pmp_ignore_12 = res_pmp_passThrough & ~io_check_env_pmp_12_cfg_l; // @[PMP.scala 434:32]
  wire  res_pmp_cur_12_cfg_r = io_check_env_pmp_12_cfg_r | res_pmp_ignore_12; // @[PMP.scala 438:42]
  wire  res_pmp_cur_12_cfg_w = io_check_env_pmp_12_cfg_w | res_pmp_ignore_12; // @[PMP.scala 439:42]
  wire  res_pmp_cur_12_cfg_x = io_check_env_pmp_12_cfg_x | res_pmp_ignore_12; // @[PMP.scala 440:42]
  wire [35:0] _res_pmp_is_match_T_274 = {io_check_env_pmp_13_addr, 2'h0}; // @[PMP.scala 190:35]
  wire [35:0] _res_pmp_is_match_T_276 = _res_pmp_is_match_T_274 & 36'hffffff000; // @[PMP.scala 190:50]
  wire [35:0] _res_pmp_is_match_T_277 = ~io_check_env_pmp_13_mask; // @[PMP.scala 232:10]
  wire [35:0] _res_pmp_is_match_T_278 = io_req_bits_addr & _res_pmp_is_match_T_277; // @[PMP.scala 232:8]
  wire [35:0] _res_pmp_is_match_T_280 = _res_pmp_is_match_T_276 & _res_pmp_is_match_T_277; // @[PMP.scala 232:21]
  wire  _res_pmp_is_match_T_281 = _res_pmp_is_match_T_278 == _res_pmp_is_match_T_280; // @[PMP.scala 232:14]
  wire  _res_pmp_is_match_T_282 = io_check_env_pmp_13_cfg_a == 2'h1; // @[PMP.scala 53:15]
  wire  _res_pmp_is_match_T_287 = ~_res_pmp_is_match_T_270; // @[PMP.scala 220:5]
  wire  _res_pmp_is_match_T_291 = io_req_bits_addr < _res_pmp_is_match_T_276; // @[PMP.scala 210:14]
  wire  _res_pmp_is_match_T_292 = _res_pmp_is_match_T_287 & _res_pmp_is_match_T_291; // @[PMP.scala 228:56]
  wire  _res_pmp_is_match_T_293 = _res_pmp_is_match_T_282 & _res_pmp_is_match_T_292; // @[PMP.scala 200:10]
  wire  res_pmp_is_match_13 = io_check_env_pmp_13_cfg_a[1] ? _res_pmp_is_match_T_281 : _res_pmp_is_match_T_293; // @[PMP.scala 199:8]
  wire  res_pmp_ignore_13 = res_pmp_passThrough & ~io_check_env_pmp_13_cfg_l; // @[PMP.scala 434:32]
  wire  res_pmp_cur_13_cfg_r = io_check_env_pmp_13_cfg_r | res_pmp_ignore_13; // @[PMP.scala 438:42]
  wire  res_pmp_cur_13_cfg_w = io_check_env_pmp_13_cfg_w | res_pmp_ignore_13; // @[PMP.scala 439:42]
  wire  res_pmp_cur_13_cfg_x = io_check_env_pmp_13_cfg_x | res_pmp_ignore_13; // @[PMP.scala 440:42]
  wire [35:0] _res_pmp_is_match_T_295 = {io_check_env_pmp_14_addr, 2'h0}; // @[PMP.scala 190:35]
  wire [35:0] _res_pmp_is_match_T_297 = _res_pmp_is_match_T_295 & 36'hffffff000; // @[PMP.scala 190:50]
  wire [35:0] _res_pmp_is_match_T_298 = ~io_check_env_pmp_14_mask; // @[PMP.scala 232:10]
  wire [35:0] _res_pmp_is_match_T_299 = io_req_bits_addr & _res_pmp_is_match_T_298; // @[PMP.scala 232:8]
  wire [35:0] _res_pmp_is_match_T_301 = _res_pmp_is_match_T_297 & _res_pmp_is_match_T_298; // @[PMP.scala 232:21]
  wire  _res_pmp_is_match_T_302 = _res_pmp_is_match_T_299 == _res_pmp_is_match_T_301; // @[PMP.scala 232:14]
  wire  _res_pmp_is_match_T_303 = io_check_env_pmp_14_cfg_a == 2'h1; // @[PMP.scala 53:15]
  wire  _res_pmp_is_match_T_308 = ~_res_pmp_is_match_T_291; // @[PMP.scala 220:5]
  wire  _res_pmp_is_match_T_312 = io_req_bits_addr < _res_pmp_is_match_T_297; // @[PMP.scala 210:14]
  wire  _res_pmp_is_match_T_313 = _res_pmp_is_match_T_308 & _res_pmp_is_match_T_312; // @[PMP.scala 228:56]
  wire  _res_pmp_is_match_T_314 = _res_pmp_is_match_T_303 & _res_pmp_is_match_T_313; // @[PMP.scala 200:10]
  wire  res_pmp_is_match_14 = io_check_env_pmp_14_cfg_a[1] ? _res_pmp_is_match_T_302 : _res_pmp_is_match_T_314; // @[PMP.scala 199:8]
  wire  res_pmp_ignore_14 = res_pmp_passThrough & ~io_check_env_pmp_14_cfg_l; // @[PMP.scala 434:32]
  wire  res_pmp_cur_14_cfg_r = io_check_env_pmp_14_cfg_r | res_pmp_ignore_14; // @[PMP.scala 438:42]
  wire  res_pmp_cur_14_cfg_w = io_check_env_pmp_14_cfg_w | res_pmp_ignore_14; // @[PMP.scala 439:42]
  wire  res_pmp_cur_14_cfg_x = io_check_env_pmp_14_cfg_x | res_pmp_ignore_14; // @[PMP.scala 440:42]
  wire [35:0] _res_pmp_is_match_T_316 = {io_check_env_pmp_15_addr, 2'h0}; // @[PMP.scala 190:35]
  wire [35:0] _res_pmp_is_match_T_318 = _res_pmp_is_match_T_316 & 36'hffffff000; // @[PMP.scala 190:50]
  wire [35:0] _res_pmp_is_match_T_319 = ~io_check_env_pmp_15_mask; // @[PMP.scala 232:10]
  wire [35:0] _res_pmp_is_match_T_320 = io_req_bits_addr & _res_pmp_is_match_T_319; // @[PMP.scala 232:8]
  wire [35:0] _res_pmp_is_match_T_322 = _res_pmp_is_match_T_318 & _res_pmp_is_match_T_319; // @[PMP.scala 232:21]
  wire  _res_pmp_is_match_T_323 = _res_pmp_is_match_T_320 == _res_pmp_is_match_T_322; // @[PMP.scala 232:14]
  wire  _res_pmp_is_match_T_324 = io_check_env_pmp_15_cfg_a == 2'h1; // @[PMP.scala 53:15]
  wire  _res_pmp_is_match_T_329 = ~_res_pmp_is_match_T_312; // @[PMP.scala 220:5]
  wire  _res_pmp_is_match_T_333 = io_req_bits_addr < _res_pmp_is_match_T_318; // @[PMP.scala 210:14]
  wire  _res_pmp_is_match_T_334 = _res_pmp_is_match_T_329 & _res_pmp_is_match_T_333; // @[PMP.scala 228:56]
  wire  _res_pmp_is_match_T_335 = _res_pmp_is_match_T_324 & _res_pmp_is_match_T_334; // @[PMP.scala 200:10]
  wire  res_pmp_is_match_15 = io_check_env_pmp_15_cfg_a[1] ? _res_pmp_is_match_T_323 : _res_pmp_is_match_T_335; // @[PMP.scala 199:8]
  wire  res_pmp_ignore_15 = res_pmp_passThrough & ~io_check_env_pmp_15_cfg_l; // @[PMP.scala 434:32]
  wire  res_pmp_cur_15_cfg_r = io_check_env_pmp_15_cfg_r | res_pmp_ignore_15; // @[PMP.scala 438:42]
  wire  res_pmp_cur_15_cfg_w = io_check_env_pmp_15_cfg_w | res_pmp_ignore_15; // @[PMP.scala 439:42]
  wire  res_pmp_cur_15_cfg_x = io_check_env_pmp_15_cfg_x | res_pmp_ignore_15; // @[PMP.scala 440:42]
  wire  _res_pmp_T_1_cfg_x = res_pmp_is_match ? res_pmp_cur_cfg_x : res_pmp_cur_1_cfg_x; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_1_cfg_w = res_pmp_is_match ? res_pmp_cur_cfg_w : res_pmp_cur_1_cfg_w; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_1_cfg_r = res_pmp_is_match ? res_pmp_cur_cfg_r : res_pmp_cur_1_cfg_r; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_3_cfg_x = res_pmp_is_match_2 ? res_pmp_cur_2_cfg_x : res_pmp_cur_3_cfg_x; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_3_cfg_w = res_pmp_is_match_2 ? res_pmp_cur_2_cfg_w : res_pmp_cur_3_cfg_w; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_3_cfg_r = res_pmp_is_match_2 ? res_pmp_cur_2_cfg_r : res_pmp_cur_3_cfg_r; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_5_cfg_x = res_pmp_is_match | res_pmp_is_match_1 ? _res_pmp_T_1_cfg_x : _res_pmp_T_3_cfg_x; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_5_cfg_w = res_pmp_is_match | res_pmp_is_match_1 ? _res_pmp_T_1_cfg_w : _res_pmp_T_3_cfg_w; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_5_cfg_r = res_pmp_is_match | res_pmp_is_match_1 ? _res_pmp_T_1_cfg_r : _res_pmp_T_3_cfg_r; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_7_cfg_x = res_pmp_is_match_4 ? res_pmp_cur_4_cfg_x : res_pmp_cur_5_cfg_x; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_7_cfg_w = res_pmp_is_match_4 ? res_pmp_cur_4_cfg_w : res_pmp_cur_5_cfg_w; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_7_cfg_r = res_pmp_is_match_4 ? res_pmp_cur_4_cfg_r : res_pmp_cur_5_cfg_r; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_9_cfg_x = res_pmp_is_match_6 ? res_pmp_cur_6_cfg_x : res_pmp_cur_7_cfg_x; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_9_cfg_w = res_pmp_is_match_6 ? res_pmp_cur_6_cfg_w : res_pmp_cur_7_cfg_w; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_9_cfg_r = res_pmp_is_match_6 ? res_pmp_cur_6_cfg_r : res_pmp_cur_7_cfg_r; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_11_cfg_x = res_pmp_is_match_4 | res_pmp_is_match_5 ? _res_pmp_T_7_cfg_x : _res_pmp_T_9_cfg_x; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_11_cfg_w = res_pmp_is_match_4 | res_pmp_is_match_5 ? _res_pmp_T_7_cfg_w : _res_pmp_T_9_cfg_w; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_11_cfg_r = res_pmp_is_match_4 | res_pmp_is_match_5 ? _res_pmp_T_7_cfg_r : _res_pmp_T_9_cfg_r; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_13_cfg_x = res_pmp_is_match | res_pmp_is_match_1 | (res_pmp_is_match_2 | res_pmp_is_match_3) ?
    _res_pmp_T_5_cfg_x : _res_pmp_T_11_cfg_x; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_13_cfg_w = res_pmp_is_match | res_pmp_is_match_1 | (res_pmp_is_match_2 | res_pmp_is_match_3) ?
    _res_pmp_T_5_cfg_w : _res_pmp_T_11_cfg_w; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_13_cfg_r = res_pmp_is_match | res_pmp_is_match_1 | (res_pmp_is_match_2 | res_pmp_is_match_3) ?
    _res_pmp_T_5_cfg_r : _res_pmp_T_11_cfg_r; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_15_cfg_x = res_pmp_is_match_8 ? res_pmp_cur_8_cfg_x : res_pmp_cur_9_cfg_x; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_15_cfg_w = res_pmp_is_match_8 ? res_pmp_cur_8_cfg_w : res_pmp_cur_9_cfg_w; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_15_cfg_r = res_pmp_is_match_8 ? res_pmp_cur_8_cfg_r : res_pmp_cur_9_cfg_r; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_17_cfg_x = res_pmp_is_match_10 ? res_pmp_cur_10_cfg_x : res_pmp_cur_11_cfg_x; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_17_cfg_w = res_pmp_is_match_10 ? res_pmp_cur_10_cfg_w : res_pmp_cur_11_cfg_w; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_17_cfg_r = res_pmp_is_match_10 ? res_pmp_cur_10_cfg_r : res_pmp_cur_11_cfg_r; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_19_cfg_x = res_pmp_is_match_8 | res_pmp_is_match_9 ? _res_pmp_T_15_cfg_x : _res_pmp_T_17_cfg_x; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_19_cfg_w = res_pmp_is_match_8 | res_pmp_is_match_9 ? _res_pmp_T_15_cfg_w : _res_pmp_T_17_cfg_w; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_19_cfg_r = res_pmp_is_match_8 | res_pmp_is_match_9 ? _res_pmp_T_15_cfg_r : _res_pmp_T_17_cfg_r; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_21_cfg_x = res_pmp_is_match_12 ? res_pmp_cur_12_cfg_x : res_pmp_cur_13_cfg_x; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_21_cfg_w = res_pmp_is_match_12 ? res_pmp_cur_12_cfg_w : res_pmp_cur_13_cfg_w; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_21_cfg_r = res_pmp_is_match_12 ? res_pmp_cur_12_cfg_r : res_pmp_cur_13_cfg_r; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_23_cfg_x = res_pmp_is_match_15 ? res_pmp_cur_15_cfg_x : res_pmp_passThrough; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_23_cfg_w = res_pmp_is_match_15 ? res_pmp_cur_15_cfg_w : res_pmp_passThrough; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_23_cfg_r = res_pmp_is_match_15 ? res_pmp_cur_15_cfg_r : res_pmp_passThrough; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_25_cfg_x = res_pmp_is_match_14 ? res_pmp_cur_14_cfg_x : _res_pmp_T_23_cfg_x; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_25_cfg_w = res_pmp_is_match_14 ? res_pmp_cur_14_cfg_w : _res_pmp_T_23_cfg_w; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_25_cfg_r = res_pmp_is_match_14 ? res_pmp_cur_14_cfg_r : _res_pmp_T_23_cfg_r; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_27_cfg_x = res_pmp_is_match_12 | res_pmp_is_match_13 ? _res_pmp_T_21_cfg_x : _res_pmp_T_25_cfg_x; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_27_cfg_w = res_pmp_is_match_12 | res_pmp_is_match_13 ? _res_pmp_T_21_cfg_w : _res_pmp_T_25_cfg_w; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_27_cfg_r = res_pmp_is_match_12 | res_pmp_is_match_13 ? _res_pmp_T_21_cfg_r : _res_pmp_T_25_cfg_r; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_29_cfg_x = res_pmp_is_match_8 | res_pmp_is_match_9 | (res_pmp_is_match_10 | res_pmp_is_match_11) ?
    _res_pmp_T_19_cfg_x : _res_pmp_T_27_cfg_x; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_29_cfg_w = res_pmp_is_match_8 | res_pmp_is_match_9 | (res_pmp_is_match_10 | res_pmp_is_match_11) ?
    _res_pmp_T_19_cfg_w : _res_pmp_T_27_cfg_w; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_29_cfg_r = res_pmp_is_match_8 | res_pmp_is_match_9 | (res_pmp_is_match_10 | res_pmp_is_match_11) ?
    _res_pmp_T_19_cfg_r : _res_pmp_T_27_cfg_r; // @[ParallelMux.scala 90:77]
  wire  res_pmp_cfg_x = res_pmp_is_match | res_pmp_is_match_1 | (res_pmp_is_match_2 | res_pmp_is_match_3) | (
    res_pmp_is_match_4 | res_pmp_is_match_5 | (res_pmp_is_match_6 | res_pmp_is_match_7)) ? _res_pmp_T_13_cfg_x :
    _res_pmp_T_29_cfg_x; // @[ParallelMux.scala 90:77]
  wire  res_pmp_cfg_w = res_pmp_is_match | res_pmp_is_match_1 | (res_pmp_is_match_2 | res_pmp_is_match_3) | (
    res_pmp_is_match_4 | res_pmp_is_match_5 | (res_pmp_is_match_6 | res_pmp_is_match_7)) ? _res_pmp_T_13_cfg_w :
    _res_pmp_T_29_cfg_w; // @[ParallelMux.scala 90:77]
  wire  res_pmp_cfg_r = res_pmp_is_match | res_pmp_is_match_1 | (res_pmp_is_match_2 | res_pmp_is_match_3) | (
    res_pmp_is_match_4 | res_pmp_is_match_5 | (res_pmp_is_match_6 | res_pmp_is_match_7)) ? _res_pmp_T_13_cfg_r :
    _res_pmp_T_29_cfg_r; // @[ParallelMux.scala 90:77]
  wire [35:0] _res_pma_is_match_T_1 = {io_check_env_pma_0_addr, 2'h0}; // @[PMP.scala 190:35]
  wire [35:0] _res_pma_is_match_T_3 = _res_pma_is_match_T_1 & 36'hffffff000; // @[PMP.scala 190:50]
  wire [35:0] _res_pma_is_match_T_4 = ~io_check_env_pma_0_mask; // @[PMP.scala 232:10]
  wire [35:0] _res_pma_is_match_T_5 = io_req_bits_addr & _res_pma_is_match_T_4; // @[PMP.scala 232:8]
  wire [35:0] _res_pma_is_match_T_7 = _res_pma_is_match_T_3 & _res_pma_is_match_T_4; // @[PMP.scala 232:21]
  wire  _res_pma_is_match_T_8 = _res_pma_is_match_T_5 == _res_pma_is_match_T_7; // @[PMP.scala 232:14]
  wire  _res_pma_is_match_T_9 = io_check_env_pma_0_cfg_a == 2'h1; // @[PMP.scala 53:15]
  wire  _res_pma_is_match_T_18 = io_req_bits_addr < _res_pma_is_match_T_3; // @[PMP.scala 210:14]
  wire  _res_pma_is_match_T_20 = _res_pma_is_match_T_9 & _res_pma_is_match_T_18; // @[PMP.scala 200:10]
  wire  res_pma_is_match = io_check_env_pma_0_cfg_a[1] ? _res_pma_is_match_T_8 : _res_pma_is_match_T_20; // @[PMP.scala 199:8]
  wire [35:0] _res_pma_is_match_T_22 = {io_check_env_pma_1_addr, 2'h0}; // @[PMP.scala 190:35]
  wire [35:0] _res_pma_is_match_T_24 = _res_pma_is_match_T_22 & 36'hffffff000; // @[PMP.scala 190:50]
  wire [35:0] _res_pma_is_match_T_25 = ~io_check_env_pma_1_mask; // @[PMP.scala 232:10]
  wire [35:0] _res_pma_is_match_T_26 = io_req_bits_addr & _res_pma_is_match_T_25; // @[PMP.scala 232:8]
  wire [35:0] _res_pma_is_match_T_28 = _res_pma_is_match_T_24 & _res_pma_is_match_T_25; // @[PMP.scala 232:21]
  wire  _res_pma_is_match_T_29 = _res_pma_is_match_T_26 == _res_pma_is_match_T_28; // @[PMP.scala 232:14]
  wire  _res_pma_is_match_T_30 = io_check_env_pma_1_cfg_a == 2'h1; // @[PMP.scala 53:15]
  wire  _res_pma_is_match_T_35 = ~_res_pma_is_match_T_18; // @[PMP.scala 220:5]
  wire  _res_pma_is_match_T_39 = io_req_bits_addr < _res_pma_is_match_T_24; // @[PMP.scala 210:14]
  wire  _res_pma_is_match_T_40 = _res_pma_is_match_T_35 & _res_pma_is_match_T_39; // @[PMP.scala 228:56]
  wire  _res_pma_is_match_T_41 = _res_pma_is_match_T_30 & _res_pma_is_match_T_40; // @[PMP.scala 200:10]
  wire  res_pma_is_match_1 = io_check_env_pma_1_cfg_a[1] ? _res_pma_is_match_T_29 : _res_pma_is_match_T_41; // @[PMP.scala 199:8]
  wire [35:0] _res_pma_is_match_T_43 = {io_check_env_pma_2_addr, 2'h0}; // @[PMP.scala 190:35]
  wire [35:0] _res_pma_is_match_T_45 = _res_pma_is_match_T_43 & 36'hffffff000; // @[PMP.scala 190:50]
  wire [35:0] _res_pma_is_match_T_46 = ~io_check_env_pma_2_mask; // @[PMP.scala 232:10]
  wire [35:0] _res_pma_is_match_T_47 = io_req_bits_addr & _res_pma_is_match_T_46; // @[PMP.scala 232:8]
  wire [35:0] _res_pma_is_match_T_49 = _res_pma_is_match_T_45 & _res_pma_is_match_T_46; // @[PMP.scala 232:21]
  wire  _res_pma_is_match_T_50 = _res_pma_is_match_T_47 == _res_pma_is_match_T_49; // @[PMP.scala 232:14]
  wire  _res_pma_is_match_T_51 = io_check_env_pma_2_cfg_a == 2'h1; // @[PMP.scala 53:15]
  wire  _res_pma_is_match_T_56 = ~_res_pma_is_match_T_39; // @[PMP.scala 220:5]
  wire  _res_pma_is_match_T_60 = io_req_bits_addr < _res_pma_is_match_T_45; // @[PMP.scala 210:14]
  wire  _res_pma_is_match_T_61 = _res_pma_is_match_T_56 & _res_pma_is_match_T_60; // @[PMP.scala 228:56]
  wire  _res_pma_is_match_T_62 = _res_pma_is_match_T_51 & _res_pma_is_match_T_61; // @[PMP.scala 200:10]
  wire  res_pma_is_match_2 = io_check_env_pma_2_cfg_a[1] ? _res_pma_is_match_T_50 : _res_pma_is_match_T_62; // @[PMP.scala 199:8]
  wire [35:0] _res_pma_is_match_T_64 = {io_check_env_pma_3_addr, 2'h0}; // @[PMP.scala 190:35]
  wire [35:0] _res_pma_is_match_T_66 = _res_pma_is_match_T_64 & 36'hffffff000; // @[PMP.scala 190:50]
  wire [35:0] _res_pma_is_match_T_67 = ~io_check_env_pma_3_mask; // @[PMP.scala 232:10]
  wire [35:0] _res_pma_is_match_T_68 = io_req_bits_addr & _res_pma_is_match_T_67; // @[PMP.scala 232:8]
  wire [35:0] _res_pma_is_match_T_70 = _res_pma_is_match_T_66 & _res_pma_is_match_T_67; // @[PMP.scala 232:21]
  wire  _res_pma_is_match_T_71 = _res_pma_is_match_T_68 == _res_pma_is_match_T_70; // @[PMP.scala 232:14]
  wire  _res_pma_is_match_T_72 = io_check_env_pma_3_cfg_a == 2'h1; // @[PMP.scala 53:15]
  wire  _res_pma_is_match_T_77 = ~_res_pma_is_match_T_60; // @[PMP.scala 220:5]
  wire  _res_pma_is_match_T_81 = io_req_bits_addr < _res_pma_is_match_T_66; // @[PMP.scala 210:14]
  wire  _res_pma_is_match_T_82 = _res_pma_is_match_T_77 & _res_pma_is_match_T_81; // @[PMP.scala 228:56]
  wire  _res_pma_is_match_T_83 = _res_pma_is_match_T_72 & _res_pma_is_match_T_82; // @[PMP.scala 200:10]
  wire  res_pma_is_match_3 = io_check_env_pma_3_cfg_a[1] ? _res_pma_is_match_T_71 : _res_pma_is_match_T_83; // @[PMP.scala 199:8]
  wire [35:0] _res_pma_is_match_T_85 = {io_check_env_pma_4_addr, 2'h0}; // @[PMP.scala 190:35]
  wire [35:0] _res_pma_is_match_T_87 = _res_pma_is_match_T_85 & 36'hffffff000; // @[PMP.scala 190:50]
  wire [35:0] _res_pma_is_match_T_88 = ~io_check_env_pma_4_mask; // @[PMP.scala 232:10]
  wire [35:0] _res_pma_is_match_T_89 = io_req_bits_addr & _res_pma_is_match_T_88; // @[PMP.scala 232:8]
  wire [35:0] _res_pma_is_match_T_91 = _res_pma_is_match_T_87 & _res_pma_is_match_T_88; // @[PMP.scala 232:21]
  wire  _res_pma_is_match_T_92 = _res_pma_is_match_T_89 == _res_pma_is_match_T_91; // @[PMP.scala 232:14]
  wire  _res_pma_is_match_T_93 = io_check_env_pma_4_cfg_a == 2'h1; // @[PMP.scala 53:15]
  wire  _res_pma_is_match_T_98 = ~_res_pma_is_match_T_81; // @[PMP.scala 220:5]
  wire  _res_pma_is_match_T_102 = io_req_bits_addr < _res_pma_is_match_T_87; // @[PMP.scala 210:14]
  wire  _res_pma_is_match_T_103 = _res_pma_is_match_T_98 & _res_pma_is_match_T_102; // @[PMP.scala 228:56]
  wire  _res_pma_is_match_T_104 = _res_pma_is_match_T_93 & _res_pma_is_match_T_103; // @[PMP.scala 200:10]
  wire  res_pma_is_match_4 = io_check_env_pma_4_cfg_a[1] ? _res_pma_is_match_T_92 : _res_pma_is_match_T_104; // @[PMP.scala 199:8]
  wire [35:0] _res_pma_is_match_T_106 = {io_check_env_pma_5_addr, 2'h0}; // @[PMP.scala 190:35]
  wire [35:0] _res_pma_is_match_T_108 = _res_pma_is_match_T_106 & 36'hffffff000; // @[PMP.scala 190:50]
  wire [35:0] _res_pma_is_match_T_109 = ~io_check_env_pma_5_mask; // @[PMP.scala 232:10]
  wire [35:0] _res_pma_is_match_T_110 = io_req_bits_addr & _res_pma_is_match_T_109; // @[PMP.scala 232:8]
  wire [35:0] _res_pma_is_match_T_112 = _res_pma_is_match_T_108 & _res_pma_is_match_T_109; // @[PMP.scala 232:21]
  wire  _res_pma_is_match_T_113 = _res_pma_is_match_T_110 == _res_pma_is_match_T_112; // @[PMP.scala 232:14]
  wire  _res_pma_is_match_T_114 = io_check_env_pma_5_cfg_a == 2'h1; // @[PMP.scala 53:15]
  wire  _res_pma_is_match_T_119 = ~_res_pma_is_match_T_102; // @[PMP.scala 220:5]
  wire  _res_pma_is_match_T_123 = io_req_bits_addr < _res_pma_is_match_T_108; // @[PMP.scala 210:14]
  wire  _res_pma_is_match_T_124 = _res_pma_is_match_T_119 & _res_pma_is_match_T_123; // @[PMP.scala 228:56]
  wire  _res_pma_is_match_T_125 = _res_pma_is_match_T_114 & _res_pma_is_match_T_124; // @[PMP.scala 200:10]
  wire  res_pma_is_match_5 = io_check_env_pma_5_cfg_a[1] ? _res_pma_is_match_T_113 : _res_pma_is_match_T_125; // @[PMP.scala 199:8]
  wire [35:0] _res_pma_is_match_T_127 = {io_check_env_pma_6_addr, 2'h0}; // @[PMP.scala 190:35]
  wire [35:0] _res_pma_is_match_T_129 = _res_pma_is_match_T_127 & 36'hffffff000; // @[PMP.scala 190:50]
  wire [35:0] _res_pma_is_match_T_130 = ~io_check_env_pma_6_mask; // @[PMP.scala 232:10]
  wire [35:0] _res_pma_is_match_T_131 = io_req_bits_addr & _res_pma_is_match_T_130; // @[PMP.scala 232:8]
  wire [35:0] _res_pma_is_match_T_133 = _res_pma_is_match_T_129 & _res_pma_is_match_T_130; // @[PMP.scala 232:21]
  wire  _res_pma_is_match_T_134 = _res_pma_is_match_T_131 == _res_pma_is_match_T_133; // @[PMP.scala 232:14]
  wire  _res_pma_is_match_T_135 = io_check_env_pma_6_cfg_a == 2'h1; // @[PMP.scala 53:15]
  wire  _res_pma_is_match_T_140 = ~_res_pma_is_match_T_123; // @[PMP.scala 220:5]
  wire  _res_pma_is_match_T_144 = io_req_bits_addr < _res_pma_is_match_T_129; // @[PMP.scala 210:14]
  wire  _res_pma_is_match_T_145 = _res_pma_is_match_T_140 & _res_pma_is_match_T_144; // @[PMP.scala 228:56]
  wire  _res_pma_is_match_T_146 = _res_pma_is_match_T_135 & _res_pma_is_match_T_145; // @[PMP.scala 200:10]
  wire  res_pma_is_match_6 = io_check_env_pma_6_cfg_a[1] ? _res_pma_is_match_T_134 : _res_pma_is_match_T_146; // @[PMP.scala 199:8]
  wire [35:0] _res_pma_is_match_T_148 = {io_check_env_pma_7_addr, 2'h0}; // @[PMP.scala 190:35]
  wire [35:0] _res_pma_is_match_T_150 = _res_pma_is_match_T_148 & 36'hffffff000; // @[PMP.scala 190:50]
  wire [35:0] _res_pma_is_match_T_151 = ~io_check_env_pma_7_mask; // @[PMP.scala 232:10]
  wire [35:0] _res_pma_is_match_T_152 = io_req_bits_addr & _res_pma_is_match_T_151; // @[PMP.scala 232:8]
  wire [35:0] _res_pma_is_match_T_154 = _res_pma_is_match_T_150 & _res_pma_is_match_T_151; // @[PMP.scala 232:21]
  wire  _res_pma_is_match_T_155 = _res_pma_is_match_T_152 == _res_pma_is_match_T_154; // @[PMP.scala 232:14]
  wire  _res_pma_is_match_T_156 = io_check_env_pma_7_cfg_a == 2'h1; // @[PMP.scala 53:15]
  wire  _res_pma_is_match_T_161 = ~_res_pma_is_match_T_144; // @[PMP.scala 220:5]
  wire  _res_pma_is_match_T_165 = io_req_bits_addr < _res_pma_is_match_T_150; // @[PMP.scala 210:14]
  wire  _res_pma_is_match_T_166 = _res_pma_is_match_T_161 & _res_pma_is_match_T_165; // @[PMP.scala 228:56]
  wire  _res_pma_is_match_T_167 = _res_pma_is_match_T_156 & _res_pma_is_match_T_166; // @[PMP.scala 200:10]
  wire  res_pma_is_match_7 = io_check_env_pma_7_cfg_a[1] ? _res_pma_is_match_T_155 : _res_pma_is_match_T_167; // @[PMP.scala 199:8]
  wire [35:0] _res_pma_is_match_T_169 = {io_check_env_pma_8_addr, 2'h0}; // @[PMP.scala 190:35]
  wire [35:0] _res_pma_is_match_T_171 = _res_pma_is_match_T_169 & 36'hffffff000; // @[PMP.scala 190:50]
  wire [35:0] _res_pma_is_match_T_172 = ~io_check_env_pma_8_mask; // @[PMP.scala 232:10]
  wire [35:0] _res_pma_is_match_T_173 = io_req_bits_addr & _res_pma_is_match_T_172; // @[PMP.scala 232:8]
  wire [35:0] _res_pma_is_match_T_175 = _res_pma_is_match_T_171 & _res_pma_is_match_T_172; // @[PMP.scala 232:21]
  wire  _res_pma_is_match_T_176 = _res_pma_is_match_T_173 == _res_pma_is_match_T_175; // @[PMP.scala 232:14]
  wire  _res_pma_is_match_T_177 = io_check_env_pma_8_cfg_a == 2'h1; // @[PMP.scala 53:15]
  wire  _res_pma_is_match_T_182 = ~_res_pma_is_match_T_165; // @[PMP.scala 220:5]
  wire  _res_pma_is_match_T_186 = io_req_bits_addr < _res_pma_is_match_T_171; // @[PMP.scala 210:14]
  wire  _res_pma_is_match_T_187 = _res_pma_is_match_T_182 & _res_pma_is_match_T_186; // @[PMP.scala 228:56]
  wire  _res_pma_is_match_T_188 = _res_pma_is_match_T_177 & _res_pma_is_match_T_187; // @[PMP.scala 200:10]
  wire  res_pma_is_match_8 = io_check_env_pma_8_cfg_a[1] ? _res_pma_is_match_T_176 : _res_pma_is_match_T_188; // @[PMP.scala 199:8]
  wire [35:0] _res_pma_is_match_T_190 = {io_check_env_pma_9_addr, 2'h0}; // @[PMP.scala 190:35]
  wire [35:0] _res_pma_is_match_T_192 = _res_pma_is_match_T_190 & 36'hffffff000; // @[PMP.scala 190:50]
  wire [35:0] _res_pma_is_match_T_193 = ~io_check_env_pma_9_mask; // @[PMP.scala 232:10]
  wire [35:0] _res_pma_is_match_T_194 = io_req_bits_addr & _res_pma_is_match_T_193; // @[PMP.scala 232:8]
  wire [35:0] _res_pma_is_match_T_196 = _res_pma_is_match_T_192 & _res_pma_is_match_T_193; // @[PMP.scala 232:21]
  wire  _res_pma_is_match_T_197 = _res_pma_is_match_T_194 == _res_pma_is_match_T_196; // @[PMP.scala 232:14]
  wire  _res_pma_is_match_T_198 = io_check_env_pma_9_cfg_a == 2'h1; // @[PMP.scala 53:15]
  wire  _res_pma_is_match_T_203 = ~_res_pma_is_match_T_186; // @[PMP.scala 220:5]
  wire  _res_pma_is_match_T_207 = io_req_bits_addr < _res_pma_is_match_T_192; // @[PMP.scala 210:14]
  wire  _res_pma_is_match_T_208 = _res_pma_is_match_T_203 & _res_pma_is_match_T_207; // @[PMP.scala 228:56]
  wire  _res_pma_is_match_T_209 = _res_pma_is_match_T_198 & _res_pma_is_match_T_208; // @[PMP.scala 200:10]
  wire  res_pma_is_match_9 = io_check_env_pma_9_cfg_a[1] ? _res_pma_is_match_T_197 : _res_pma_is_match_T_209; // @[PMP.scala 199:8]
  wire [35:0] _res_pma_is_match_T_211 = {io_check_env_pma_10_addr, 2'h0}; // @[PMP.scala 190:35]
  wire [35:0] _res_pma_is_match_T_213 = _res_pma_is_match_T_211 & 36'hffffff000; // @[PMP.scala 190:50]
  wire [35:0] _res_pma_is_match_T_214 = ~io_check_env_pma_10_mask; // @[PMP.scala 232:10]
  wire [35:0] _res_pma_is_match_T_215 = io_req_bits_addr & _res_pma_is_match_T_214; // @[PMP.scala 232:8]
  wire [35:0] _res_pma_is_match_T_217 = _res_pma_is_match_T_213 & _res_pma_is_match_T_214; // @[PMP.scala 232:21]
  wire  _res_pma_is_match_T_218 = _res_pma_is_match_T_215 == _res_pma_is_match_T_217; // @[PMP.scala 232:14]
  wire  _res_pma_is_match_T_219 = io_check_env_pma_10_cfg_a == 2'h1; // @[PMP.scala 53:15]
  wire  _res_pma_is_match_T_224 = ~_res_pma_is_match_T_207; // @[PMP.scala 220:5]
  wire  _res_pma_is_match_T_228 = io_req_bits_addr < _res_pma_is_match_T_213; // @[PMP.scala 210:14]
  wire  _res_pma_is_match_T_229 = _res_pma_is_match_T_224 & _res_pma_is_match_T_228; // @[PMP.scala 228:56]
  wire  _res_pma_is_match_T_230 = _res_pma_is_match_T_219 & _res_pma_is_match_T_229; // @[PMP.scala 200:10]
  wire  res_pma_is_match_10 = io_check_env_pma_10_cfg_a[1] ? _res_pma_is_match_T_218 : _res_pma_is_match_T_230; // @[PMP.scala 199:8]
  wire [35:0] _res_pma_is_match_T_232 = {io_check_env_pma_11_addr, 2'h0}; // @[PMP.scala 190:35]
  wire [35:0] _res_pma_is_match_T_234 = _res_pma_is_match_T_232 & 36'hffffff000; // @[PMP.scala 190:50]
  wire [35:0] _res_pma_is_match_T_235 = ~io_check_env_pma_11_mask; // @[PMP.scala 232:10]
  wire [35:0] _res_pma_is_match_T_236 = io_req_bits_addr & _res_pma_is_match_T_235; // @[PMP.scala 232:8]
  wire [35:0] _res_pma_is_match_T_238 = _res_pma_is_match_T_234 & _res_pma_is_match_T_235; // @[PMP.scala 232:21]
  wire  _res_pma_is_match_T_239 = _res_pma_is_match_T_236 == _res_pma_is_match_T_238; // @[PMP.scala 232:14]
  wire  _res_pma_is_match_T_240 = io_check_env_pma_11_cfg_a == 2'h1; // @[PMP.scala 53:15]
  wire  _res_pma_is_match_T_245 = ~_res_pma_is_match_T_228; // @[PMP.scala 220:5]
  wire  _res_pma_is_match_T_249 = io_req_bits_addr < _res_pma_is_match_T_234; // @[PMP.scala 210:14]
  wire  _res_pma_is_match_T_250 = _res_pma_is_match_T_245 & _res_pma_is_match_T_249; // @[PMP.scala 228:56]
  wire  _res_pma_is_match_T_251 = _res_pma_is_match_T_240 & _res_pma_is_match_T_250; // @[PMP.scala 200:10]
  wire  res_pma_is_match_11 = io_check_env_pma_11_cfg_a[1] ? _res_pma_is_match_T_239 : _res_pma_is_match_T_251; // @[PMP.scala 199:8]
  wire [35:0] _res_pma_is_match_T_253 = {io_check_env_pma_12_addr, 2'h0}; // @[PMP.scala 190:35]
  wire [35:0] _res_pma_is_match_T_255 = _res_pma_is_match_T_253 & 36'hffffff000; // @[PMP.scala 190:50]
  wire [35:0] _res_pma_is_match_T_256 = ~io_check_env_pma_12_mask; // @[PMP.scala 232:10]
  wire [35:0] _res_pma_is_match_T_257 = io_req_bits_addr & _res_pma_is_match_T_256; // @[PMP.scala 232:8]
  wire [35:0] _res_pma_is_match_T_259 = _res_pma_is_match_T_255 & _res_pma_is_match_T_256; // @[PMP.scala 232:21]
  wire  _res_pma_is_match_T_260 = _res_pma_is_match_T_257 == _res_pma_is_match_T_259; // @[PMP.scala 232:14]
  wire  _res_pma_is_match_T_261 = io_check_env_pma_12_cfg_a == 2'h1; // @[PMP.scala 53:15]
  wire  _res_pma_is_match_T_266 = ~_res_pma_is_match_T_249; // @[PMP.scala 220:5]
  wire  _res_pma_is_match_T_270 = io_req_bits_addr < _res_pma_is_match_T_255; // @[PMP.scala 210:14]
  wire  _res_pma_is_match_T_271 = _res_pma_is_match_T_266 & _res_pma_is_match_T_270; // @[PMP.scala 228:56]
  wire  _res_pma_is_match_T_272 = _res_pma_is_match_T_261 & _res_pma_is_match_T_271; // @[PMP.scala 200:10]
  wire  res_pma_is_match_12 = io_check_env_pma_12_cfg_a[1] ? _res_pma_is_match_T_260 : _res_pma_is_match_T_272; // @[PMP.scala 199:8]
  wire [35:0] _res_pma_is_match_T_274 = {io_check_env_pma_13_addr, 2'h0}; // @[PMP.scala 190:35]
  wire [35:0] _res_pma_is_match_T_276 = _res_pma_is_match_T_274 & 36'hffffff000; // @[PMP.scala 190:50]
  wire [35:0] _res_pma_is_match_T_277 = ~io_check_env_pma_13_mask; // @[PMP.scala 232:10]
  wire [35:0] _res_pma_is_match_T_278 = io_req_bits_addr & _res_pma_is_match_T_277; // @[PMP.scala 232:8]
  wire [35:0] _res_pma_is_match_T_280 = _res_pma_is_match_T_276 & _res_pma_is_match_T_277; // @[PMP.scala 232:21]
  wire  _res_pma_is_match_T_281 = _res_pma_is_match_T_278 == _res_pma_is_match_T_280; // @[PMP.scala 232:14]
  wire  _res_pma_is_match_T_282 = io_check_env_pma_13_cfg_a == 2'h1; // @[PMP.scala 53:15]
  wire  _res_pma_is_match_T_287 = ~_res_pma_is_match_T_270; // @[PMP.scala 220:5]
  wire  _res_pma_is_match_T_291 = io_req_bits_addr < _res_pma_is_match_T_276; // @[PMP.scala 210:14]
  wire  _res_pma_is_match_T_292 = _res_pma_is_match_T_287 & _res_pma_is_match_T_291; // @[PMP.scala 228:56]
  wire  _res_pma_is_match_T_293 = _res_pma_is_match_T_282 & _res_pma_is_match_T_292; // @[PMP.scala 200:10]
  wire  res_pma_is_match_13 = io_check_env_pma_13_cfg_a[1] ? _res_pma_is_match_T_281 : _res_pma_is_match_T_293; // @[PMP.scala 199:8]
  wire [35:0] _res_pma_is_match_T_295 = {io_check_env_pma_14_addr, 2'h0}; // @[PMP.scala 190:35]
  wire [35:0] _res_pma_is_match_T_297 = _res_pma_is_match_T_295 & 36'hffffff000; // @[PMP.scala 190:50]
  wire [35:0] _res_pma_is_match_T_298 = ~io_check_env_pma_14_mask; // @[PMP.scala 232:10]
  wire [35:0] _res_pma_is_match_T_299 = io_req_bits_addr & _res_pma_is_match_T_298; // @[PMP.scala 232:8]
  wire [35:0] _res_pma_is_match_T_301 = _res_pma_is_match_T_297 & _res_pma_is_match_T_298; // @[PMP.scala 232:21]
  wire  _res_pma_is_match_T_302 = _res_pma_is_match_T_299 == _res_pma_is_match_T_301; // @[PMP.scala 232:14]
  wire  _res_pma_is_match_T_303 = io_check_env_pma_14_cfg_a == 2'h1; // @[PMP.scala 53:15]
  wire  _res_pma_is_match_T_308 = ~_res_pma_is_match_T_291; // @[PMP.scala 220:5]
  wire  _res_pma_is_match_T_312 = io_req_bits_addr < _res_pma_is_match_T_297; // @[PMP.scala 210:14]
  wire  _res_pma_is_match_T_313 = _res_pma_is_match_T_308 & _res_pma_is_match_T_312; // @[PMP.scala 228:56]
  wire  _res_pma_is_match_T_314 = _res_pma_is_match_T_303 & _res_pma_is_match_T_313; // @[PMP.scala 200:10]
  wire  res_pma_is_match_14 = io_check_env_pma_14_cfg_a[1] ? _res_pma_is_match_T_302 : _res_pma_is_match_T_314; // @[PMP.scala 199:8]
  wire [35:0] _res_pma_is_match_T_316 = {io_check_env_pma_15_addr, 2'h0}; // @[PMP.scala 190:35]
  wire [35:0] _res_pma_is_match_T_318 = _res_pma_is_match_T_316 & 36'hffffff000; // @[PMP.scala 190:50]
  wire [35:0] _res_pma_is_match_T_319 = ~io_check_env_pma_15_mask; // @[PMP.scala 232:10]
  wire [35:0] _res_pma_is_match_T_320 = io_req_bits_addr & _res_pma_is_match_T_319; // @[PMP.scala 232:8]
  wire [35:0] _res_pma_is_match_T_322 = _res_pma_is_match_T_318 & _res_pma_is_match_T_319; // @[PMP.scala 232:21]
  wire  _res_pma_is_match_T_323 = _res_pma_is_match_T_320 == _res_pma_is_match_T_322; // @[PMP.scala 232:14]
  wire  _res_pma_is_match_T_324 = io_check_env_pma_15_cfg_a == 2'h1; // @[PMP.scala 53:15]
  wire  _res_pma_is_match_T_329 = ~_res_pma_is_match_T_312; // @[PMP.scala 220:5]
  wire  _res_pma_is_match_T_333 = io_req_bits_addr < _res_pma_is_match_T_318; // @[PMP.scala 210:14]
  wire  _res_pma_is_match_T_334 = _res_pma_is_match_T_329 & _res_pma_is_match_T_333; // @[PMP.scala 228:56]
  wire  _res_pma_is_match_T_335 = _res_pma_is_match_T_324 & _res_pma_is_match_T_334; // @[PMP.scala 200:10]
  wire  res_pma_is_match_15 = io_check_env_pma_15_cfg_a[1] ? _res_pma_is_match_T_323 : _res_pma_is_match_T_335; // @[PMP.scala 199:8]
  wire  _res_pma_T_1_cfg_c = res_pma_is_match ? io_check_env_pma_0_cfg_c : io_check_env_pma_1_cfg_c; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_1_cfg_atomic = res_pma_is_match ? io_check_env_pma_0_cfg_atomic : io_check_env_pma_1_cfg_atomic; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_1_cfg_x = res_pma_is_match ? io_check_env_pma_0_cfg_x : io_check_env_pma_1_cfg_x; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_1_cfg_w = res_pma_is_match ? io_check_env_pma_0_cfg_w : io_check_env_pma_1_cfg_w; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_1_cfg_r = res_pma_is_match ? io_check_env_pma_0_cfg_r : io_check_env_pma_1_cfg_r; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_3_cfg_c = res_pma_is_match_2 ? io_check_env_pma_2_cfg_c : io_check_env_pma_3_cfg_c; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_3_cfg_atomic = res_pma_is_match_2 ? io_check_env_pma_2_cfg_atomic : io_check_env_pma_3_cfg_atomic; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_3_cfg_x = res_pma_is_match_2 ? io_check_env_pma_2_cfg_x : io_check_env_pma_3_cfg_x; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_3_cfg_w = res_pma_is_match_2 ? io_check_env_pma_2_cfg_w : io_check_env_pma_3_cfg_w; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_3_cfg_r = res_pma_is_match_2 ? io_check_env_pma_2_cfg_r : io_check_env_pma_3_cfg_r; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_5_cfg_c = res_pma_is_match | res_pma_is_match_1 ? _res_pma_T_1_cfg_c : _res_pma_T_3_cfg_c; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_5_cfg_atomic = res_pma_is_match | res_pma_is_match_1 ? _res_pma_T_1_cfg_atomic :
    _res_pma_T_3_cfg_atomic; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_5_cfg_x = res_pma_is_match | res_pma_is_match_1 ? _res_pma_T_1_cfg_x : _res_pma_T_3_cfg_x; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_5_cfg_w = res_pma_is_match | res_pma_is_match_1 ? _res_pma_T_1_cfg_w : _res_pma_T_3_cfg_w; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_5_cfg_r = res_pma_is_match | res_pma_is_match_1 ? _res_pma_T_1_cfg_r : _res_pma_T_3_cfg_r; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_7_cfg_c = res_pma_is_match_4 ? io_check_env_pma_4_cfg_c : io_check_env_pma_5_cfg_c; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_7_cfg_atomic = res_pma_is_match_4 ? io_check_env_pma_4_cfg_atomic : io_check_env_pma_5_cfg_atomic; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_7_cfg_x = res_pma_is_match_4 ? io_check_env_pma_4_cfg_x : io_check_env_pma_5_cfg_x; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_7_cfg_w = res_pma_is_match_4 ? io_check_env_pma_4_cfg_w : io_check_env_pma_5_cfg_w; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_7_cfg_r = res_pma_is_match_4 ? io_check_env_pma_4_cfg_r : io_check_env_pma_5_cfg_r; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_9_cfg_c = res_pma_is_match_6 ? io_check_env_pma_6_cfg_c : io_check_env_pma_7_cfg_c; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_9_cfg_atomic = res_pma_is_match_6 ? io_check_env_pma_6_cfg_atomic : io_check_env_pma_7_cfg_atomic; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_9_cfg_x = res_pma_is_match_6 ? io_check_env_pma_6_cfg_x : io_check_env_pma_7_cfg_x; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_9_cfg_w = res_pma_is_match_6 ? io_check_env_pma_6_cfg_w : io_check_env_pma_7_cfg_w; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_9_cfg_r = res_pma_is_match_6 ? io_check_env_pma_6_cfg_r : io_check_env_pma_7_cfg_r; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_11_cfg_c = res_pma_is_match_4 | res_pma_is_match_5 ? _res_pma_T_7_cfg_c : _res_pma_T_9_cfg_c; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_11_cfg_atomic = res_pma_is_match_4 | res_pma_is_match_5 ? _res_pma_T_7_cfg_atomic :
    _res_pma_T_9_cfg_atomic; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_11_cfg_x = res_pma_is_match_4 | res_pma_is_match_5 ? _res_pma_T_7_cfg_x : _res_pma_T_9_cfg_x; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_11_cfg_w = res_pma_is_match_4 | res_pma_is_match_5 ? _res_pma_T_7_cfg_w : _res_pma_T_9_cfg_w; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_11_cfg_r = res_pma_is_match_4 | res_pma_is_match_5 ? _res_pma_T_7_cfg_r : _res_pma_T_9_cfg_r; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_13_cfg_c = res_pma_is_match | res_pma_is_match_1 | (res_pma_is_match_2 | res_pma_is_match_3) ?
    _res_pma_T_5_cfg_c : _res_pma_T_11_cfg_c; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_13_cfg_atomic = res_pma_is_match | res_pma_is_match_1 | (res_pma_is_match_2 | res_pma_is_match_3) ?
    _res_pma_T_5_cfg_atomic : _res_pma_T_11_cfg_atomic; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_13_cfg_x = res_pma_is_match | res_pma_is_match_1 | (res_pma_is_match_2 | res_pma_is_match_3) ?
    _res_pma_T_5_cfg_x : _res_pma_T_11_cfg_x; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_13_cfg_w = res_pma_is_match | res_pma_is_match_1 | (res_pma_is_match_2 | res_pma_is_match_3) ?
    _res_pma_T_5_cfg_w : _res_pma_T_11_cfg_w; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_13_cfg_r = res_pma_is_match | res_pma_is_match_1 | (res_pma_is_match_2 | res_pma_is_match_3) ?
    _res_pma_T_5_cfg_r : _res_pma_T_11_cfg_r; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_15_cfg_c = res_pma_is_match_8 ? io_check_env_pma_8_cfg_c : io_check_env_pma_9_cfg_c; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_15_cfg_atomic = res_pma_is_match_8 ? io_check_env_pma_8_cfg_atomic : io_check_env_pma_9_cfg_atomic; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_15_cfg_x = res_pma_is_match_8 ? io_check_env_pma_8_cfg_x : io_check_env_pma_9_cfg_x; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_15_cfg_w = res_pma_is_match_8 ? io_check_env_pma_8_cfg_w : io_check_env_pma_9_cfg_w; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_15_cfg_r = res_pma_is_match_8 ? io_check_env_pma_8_cfg_r : io_check_env_pma_9_cfg_r; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_17_cfg_c = res_pma_is_match_10 ? io_check_env_pma_10_cfg_c : io_check_env_pma_11_cfg_c; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_17_cfg_atomic = res_pma_is_match_10 ? io_check_env_pma_10_cfg_atomic : io_check_env_pma_11_cfg_atomic
    ; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_17_cfg_x = res_pma_is_match_10 ? io_check_env_pma_10_cfg_x : io_check_env_pma_11_cfg_x; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_17_cfg_w = res_pma_is_match_10 ? io_check_env_pma_10_cfg_w : io_check_env_pma_11_cfg_w; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_17_cfg_r = res_pma_is_match_10 ? io_check_env_pma_10_cfg_r : io_check_env_pma_11_cfg_r; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_19_cfg_c = res_pma_is_match_8 | res_pma_is_match_9 ? _res_pma_T_15_cfg_c : _res_pma_T_17_cfg_c; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_19_cfg_atomic = res_pma_is_match_8 | res_pma_is_match_9 ? _res_pma_T_15_cfg_atomic :
    _res_pma_T_17_cfg_atomic; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_19_cfg_x = res_pma_is_match_8 | res_pma_is_match_9 ? _res_pma_T_15_cfg_x : _res_pma_T_17_cfg_x; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_19_cfg_w = res_pma_is_match_8 | res_pma_is_match_9 ? _res_pma_T_15_cfg_w : _res_pma_T_17_cfg_w; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_19_cfg_r = res_pma_is_match_8 | res_pma_is_match_9 ? _res_pma_T_15_cfg_r : _res_pma_T_17_cfg_r; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_21_cfg_c = res_pma_is_match_12 ? io_check_env_pma_12_cfg_c : io_check_env_pma_13_cfg_c; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_21_cfg_atomic = res_pma_is_match_12 ? io_check_env_pma_12_cfg_atomic : io_check_env_pma_13_cfg_atomic
    ; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_21_cfg_x = res_pma_is_match_12 ? io_check_env_pma_12_cfg_x : io_check_env_pma_13_cfg_x; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_21_cfg_w = res_pma_is_match_12 ? io_check_env_pma_12_cfg_w : io_check_env_pma_13_cfg_w; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_21_cfg_r = res_pma_is_match_12 ? io_check_env_pma_12_cfg_r : io_check_env_pma_13_cfg_r; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_25_cfg_c = res_pma_is_match_14 ? io_check_env_pma_14_cfg_c : res_pma_is_match_15 &
    io_check_env_pma_15_cfg_c; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_25_cfg_atomic = res_pma_is_match_14 ? io_check_env_pma_14_cfg_atomic : res_pma_is_match_15 &
    io_check_env_pma_15_cfg_atomic; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_25_cfg_x = res_pma_is_match_14 ? io_check_env_pma_14_cfg_x : res_pma_is_match_15 &
    io_check_env_pma_15_cfg_x; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_25_cfg_w = res_pma_is_match_14 ? io_check_env_pma_14_cfg_w : res_pma_is_match_15 &
    io_check_env_pma_15_cfg_w; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_25_cfg_r = res_pma_is_match_14 ? io_check_env_pma_14_cfg_r : res_pma_is_match_15 &
    io_check_env_pma_15_cfg_r; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_27_cfg_c = res_pma_is_match_12 | res_pma_is_match_13 ? _res_pma_T_21_cfg_c : _res_pma_T_25_cfg_c; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_27_cfg_atomic = res_pma_is_match_12 | res_pma_is_match_13 ? _res_pma_T_21_cfg_atomic :
    _res_pma_T_25_cfg_atomic; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_27_cfg_x = res_pma_is_match_12 | res_pma_is_match_13 ? _res_pma_T_21_cfg_x : _res_pma_T_25_cfg_x; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_27_cfg_w = res_pma_is_match_12 | res_pma_is_match_13 ? _res_pma_T_21_cfg_w : _res_pma_T_25_cfg_w; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_27_cfg_r = res_pma_is_match_12 | res_pma_is_match_13 ? _res_pma_T_21_cfg_r : _res_pma_T_25_cfg_r; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_29_cfg_c = res_pma_is_match_8 | res_pma_is_match_9 | (res_pma_is_match_10 | res_pma_is_match_11) ?
    _res_pma_T_19_cfg_c : _res_pma_T_27_cfg_c; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_29_cfg_atomic = res_pma_is_match_8 | res_pma_is_match_9 | (res_pma_is_match_10 | res_pma_is_match_11)
     ? _res_pma_T_19_cfg_atomic : _res_pma_T_27_cfg_atomic; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_29_cfg_x = res_pma_is_match_8 | res_pma_is_match_9 | (res_pma_is_match_10 | res_pma_is_match_11) ?
    _res_pma_T_19_cfg_x : _res_pma_T_27_cfg_x; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_29_cfg_w = res_pma_is_match_8 | res_pma_is_match_9 | (res_pma_is_match_10 | res_pma_is_match_11) ?
    _res_pma_T_19_cfg_w : _res_pma_T_27_cfg_w; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_29_cfg_r = res_pma_is_match_8 | res_pma_is_match_9 | (res_pma_is_match_10 | res_pma_is_match_11) ?
    _res_pma_T_19_cfg_r : _res_pma_T_27_cfg_r; // @[ParallelMux.scala 90:77]
  wire  res_pma_cfg_c = res_pma_is_match | res_pma_is_match_1 | (res_pma_is_match_2 | res_pma_is_match_3) | (
    res_pma_is_match_4 | res_pma_is_match_5 | (res_pma_is_match_6 | res_pma_is_match_7)) ? _res_pma_T_13_cfg_c :
    _res_pma_T_29_cfg_c; // @[ParallelMux.scala 90:77]
  wire  res_pma_cfg_atomic = res_pma_is_match | res_pma_is_match_1 | (res_pma_is_match_2 | res_pma_is_match_3) | (
    res_pma_is_match_4 | res_pma_is_match_5 | (res_pma_is_match_6 | res_pma_is_match_7)) ? _res_pma_T_13_cfg_atomic :
    _res_pma_T_29_cfg_atomic; // @[ParallelMux.scala 90:77]
  wire  res_pma_cfg_x = res_pma_is_match | res_pma_is_match_1 | (res_pma_is_match_2 | res_pma_is_match_3) | (
    res_pma_is_match_4 | res_pma_is_match_5 | (res_pma_is_match_6 | res_pma_is_match_7)) ? _res_pma_T_13_cfg_x :
    _res_pma_T_29_cfg_x; // @[ParallelMux.scala 90:77]
  wire  res_pma_cfg_w = res_pma_is_match | res_pma_is_match_1 | (res_pma_is_match_2 | res_pma_is_match_3) | (
    res_pma_is_match_4 | res_pma_is_match_5 | (res_pma_is_match_6 | res_pma_is_match_7)) ? _res_pma_T_13_cfg_w :
    _res_pma_T_29_cfg_w; // @[ParallelMux.scala 90:77]
  wire  res_pma_cfg_r = res_pma_is_match | res_pma_is_match_1 | (res_pma_is_match_2 | res_pma_is_match_3) | (
    res_pma_is_match_4 | res_pma_is_match_5 | (res_pma_is_match_6 | res_pma_is_match_7)) ? _res_pma_T_13_cfg_r :
    _res_pma_T_29_cfg_r; // @[ParallelMux.scala 90:77]
  wire  _resp_pmp_resp_ld_T_1 = io_req_bits_cmd[1:0] == 2'h0; // @[MMUBundle.scala 234:31]
  wire  _resp_pmp_resp_ld_T_2 = io_req_bits_cmd == 3'h5; // @[MMUBundle.scala 239:25]
  wire  resp_pmp_ld = _resp_pmp_resp_ld_T_1 & ~_resp_pmp_resp_ld_T_2 & ~res_pmp_cfg_r; // @[PMP.scala 405:57]
  wire  _resp_pmp_resp_st_T_1 = io_req_bits_cmd[1:0] == 2'h1; // @[MMUBundle.scala 235:32]
  wire  resp_pmp_st = (_resp_pmp_resp_st_T_1 | _resp_pmp_resp_ld_T_2) & ~res_pmp_cfg_w; // @[PMP.scala 406:59]
  wire  _resp_pmp_resp_instr_T_1 = io_req_bits_cmd[1:0] == 2'h2; // @[MMUBundle.scala 236:31]
  wire  resp_pmp_instr = _resp_pmp_resp_instr_T_1 & ~res_pmp_cfg_x; // @[PMP.scala 407:38]
  wire  resp_pma_ld = _resp_pmp_resp_ld_T_1 & ~io_req_bits_cmd[2] & ~res_pma_cfg_r; // @[PMA.scala 212:58]
  wire  resp_pma_st = (_resp_pmp_resp_st_T_1 | io_req_bits_cmd[2] & res_pma_cfg_atomic) & ~res_pma_cfg_w; // @[PMA.scala 213:74]
  wire  resp_pma_instr = _resp_pmp_resp_instr_T_1 & ~res_pma_cfg_x; // @[PMA.scala 214:38]
  assign io_resp_ld = resp_pmp_ld | resp_pma_ld; // @[PMP.scala 393:23]
  assign io_resp_st = resp_pmp_st | resp_pma_st; // @[PMP.scala 394:23]
  assign io_resp_instr = resp_pmp_instr | resp_pma_instr; // @[PMP.scala 395:29]
  assign io_resp_mmio = ~res_pma_cfg_c; // @[PMA.scala 215:18]
  assign io_resp_atomic = res_pma_is_match | res_pma_is_match_1 | (res_pma_is_match_2 | res_pma_is_match_3) | (
    res_pma_is_match_4 | res_pma_is_match_5 | (res_pma_is_match_6 | res_pma_is_match_7)) ? _res_pma_T_13_cfg_atomic :
    _res_pma_T_29_cfg_atomic; // @[ParallelMux.scala 90:77]
endmodule

