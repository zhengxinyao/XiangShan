module TLPMA(
  input         clock,
  input         reset,
  output        auto_in_a_ready,
  input         auto_in_a_valid,
  input  [2:0]  auto_in_a_bits_opcode,
  input  [1:0]  auto_in_a_bits_size,
  input  [2:0]  auto_in_a_bits_source,
  input  [29:0] auto_in_a_bits_address,
  input  [7:0]  auto_in_a_bits_mask,
  input  [63:0] auto_in_a_bits_data,
  input         auto_in_d_ready,
  output        auto_in_d_valid,
  output [2:0]  auto_in_d_bits_opcode,
  output [1:0]  auto_in_d_bits_size,
  output [2:0]  auto_in_d_bits_source,
  output [63:0] auto_in_d_bits_data,
  input  [35:0] io_req_0_bits_addr,
  input  [35:0] io_req_1_bits_addr,
  output        io_resp_0_ld,
  output        io_resp_0_st,
  output        io_resp_0_instr,
  output        io_resp_0_mmio,
  output        io_resp_0_atomic,
  output        io_resp_1_ld,
  output        io_resp_1_st,
  output        io_resp_1_instr,
  output        io_resp_1_mmio,
  output        io_resp_1_atomic
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [63:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
`endif // RANDOMIZE_REG_INIT
  wire  out_back_clock; // @[Decoupled.scala 361:21]
  wire  out_back_reset; // @[Decoupled.scala 361:21]
  wire  out_back_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  out_back_io_enq_valid; // @[Decoupled.scala 361:21]
  wire  out_back_io_enq_bits_read; // @[Decoupled.scala 361:21]
  wire [8:0] out_back_io_enq_bits_index; // @[Decoupled.scala 361:21]
  wire [63:0] out_back_io_enq_bits_data; // @[Decoupled.scala 361:21]
  wire [7:0] out_back_io_enq_bits_mask; // @[Decoupled.scala 361:21]
  wire [2:0] out_back_io_enq_bits_extra_tlrr_extra_source; // @[Decoupled.scala 361:21]
  wire [1:0] out_back_io_enq_bits_extra_tlrr_extra_size; // @[Decoupled.scala 361:21]
  wire  out_back_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  out_back_io_deq_valid; // @[Decoupled.scala 361:21]
  wire  out_back_io_deq_bits_read; // @[Decoupled.scala 361:21]
  wire [8:0] out_back_io_deq_bits_index; // @[Decoupled.scala 361:21]
  wire [63:0] out_back_io_deq_bits_data; // @[Decoupled.scala 361:21]
  wire [7:0] out_back_io_deq_bits_mask; // @[Decoupled.scala 361:21]
  wire [2:0] out_back_io_deq_bits_extra_tlrr_extra_source; // @[Decoupled.scala 361:21]
  wire [1:0] out_back_io_deq_bits_extra_tlrr_extra_size; // @[Decoupled.scala 361:21]
  wire [1:0] PMPChecker_io_check_env_mode; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pmp_0_cfg_l; // @[TLPMA.scala 47:13]
  wire [1:0] PMPChecker_io_check_env_pmp_0_cfg_a; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pmp_0_cfg_x; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pmp_0_cfg_w; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pmp_0_cfg_r; // @[TLPMA.scala 47:13]
  wire [33:0] PMPChecker_io_check_env_pmp_0_addr; // @[TLPMA.scala 47:13]
  wire [35:0] PMPChecker_io_check_env_pmp_0_mask; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pmp_1_cfg_l; // @[TLPMA.scala 47:13]
  wire [1:0] PMPChecker_io_check_env_pmp_1_cfg_a; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pmp_1_cfg_x; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pmp_1_cfg_w; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pmp_1_cfg_r; // @[TLPMA.scala 47:13]
  wire [33:0] PMPChecker_io_check_env_pmp_1_addr; // @[TLPMA.scala 47:13]
  wire [35:0] PMPChecker_io_check_env_pmp_1_mask; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pmp_2_cfg_l; // @[TLPMA.scala 47:13]
  wire [1:0] PMPChecker_io_check_env_pmp_2_cfg_a; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pmp_2_cfg_x; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pmp_2_cfg_w; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pmp_2_cfg_r; // @[TLPMA.scala 47:13]
  wire [33:0] PMPChecker_io_check_env_pmp_2_addr; // @[TLPMA.scala 47:13]
  wire [35:0] PMPChecker_io_check_env_pmp_2_mask; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pmp_3_cfg_l; // @[TLPMA.scala 47:13]
  wire [1:0] PMPChecker_io_check_env_pmp_3_cfg_a; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pmp_3_cfg_x; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pmp_3_cfg_w; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pmp_3_cfg_r; // @[TLPMA.scala 47:13]
  wire [33:0] PMPChecker_io_check_env_pmp_3_addr; // @[TLPMA.scala 47:13]
  wire [35:0] PMPChecker_io_check_env_pmp_3_mask; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pmp_4_cfg_l; // @[TLPMA.scala 47:13]
  wire [1:0] PMPChecker_io_check_env_pmp_4_cfg_a; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pmp_4_cfg_x; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pmp_4_cfg_w; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pmp_4_cfg_r; // @[TLPMA.scala 47:13]
  wire [33:0] PMPChecker_io_check_env_pmp_4_addr; // @[TLPMA.scala 47:13]
  wire [35:0] PMPChecker_io_check_env_pmp_4_mask; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pmp_5_cfg_l; // @[TLPMA.scala 47:13]
  wire [1:0] PMPChecker_io_check_env_pmp_5_cfg_a; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pmp_5_cfg_x; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pmp_5_cfg_w; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pmp_5_cfg_r; // @[TLPMA.scala 47:13]
  wire [33:0] PMPChecker_io_check_env_pmp_5_addr; // @[TLPMA.scala 47:13]
  wire [35:0] PMPChecker_io_check_env_pmp_5_mask; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pmp_6_cfg_l; // @[TLPMA.scala 47:13]
  wire [1:0] PMPChecker_io_check_env_pmp_6_cfg_a; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pmp_6_cfg_x; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pmp_6_cfg_w; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pmp_6_cfg_r; // @[TLPMA.scala 47:13]
  wire [33:0] PMPChecker_io_check_env_pmp_6_addr; // @[TLPMA.scala 47:13]
  wire [35:0] PMPChecker_io_check_env_pmp_6_mask; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pmp_7_cfg_l; // @[TLPMA.scala 47:13]
  wire [1:0] PMPChecker_io_check_env_pmp_7_cfg_a; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pmp_7_cfg_x; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pmp_7_cfg_w; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pmp_7_cfg_r; // @[TLPMA.scala 47:13]
  wire [33:0] PMPChecker_io_check_env_pmp_7_addr; // @[TLPMA.scala 47:13]
  wire [35:0] PMPChecker_io_check_env_pmp_7_mask; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pmp_8_cfg_l; // @[TLPMA.scala 47:13]
  wire [1:0] PMPChecker_io_check_env_pmp_8_cfg_a; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pmp_8_cfg_x; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pmp_8_cfg_w; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pmp_8_cfg_r; // @[TLPMA.scala 47:13]
  wire [33:0] PMPChecker_io_check_env_pmp_8_addr; // @[TLPMA.scala 47:13]
  wire [35:0] PMPChecker_io_check_env_pmp_8_mask; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pmp_9_cfg_l; // @[TLPMA.scala 47:13]
  wire [1:0] PMPChecker_io_check_env_pmp_9_cfg_a; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pmp_9_cfg_x; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pmp_9_cfg_w; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pmp_9_cfg_r; // @[TLPMA.scala 47:13]
  wire [33:0] PMPChecker_io_check_env_pmp_9_addr; // @[TLPMA.scala 47:13]
  wire [35:0] PMPChecker_io_check_env_pmp_9_mask; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pmp_10_cfg_l; // @[TLPMA.scala 47:13]
  wire [1:0] PMPChecker_io_check_env_pmp_10_cfg_a; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pmp_10_cfg_x; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pmp_10_cfg_w; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pmp_10_cfg_r; // @[TLPMA.scala 47:13]
  wire [33:0] PMPChecker_io_check_env_pmp_10_addr; // @[TLPMA.scala 47:13]
  wire [35:0] PMPChecker_io_check_env_pmp_10_mask; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pmp_11_cfg_l; // @[TLPMA.scala 47:13]
  wire [1:0] PMPChecker_io_check_env_pmp_11_cfg_a; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pmp_11_cfg_x; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pmp_11_cfg_w; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pmp_11_cfg_r; // @[TLPMA.scala 47:13]
  wire [33:0] PMPChecker_io_check_env_pmp_11_addr; // @[TLPMA.scala 47:13]
  wire [35:0] PMPChecker_io_check_env_pmp_11_mask; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pmp_12_cfg_l; // @[TLPMA.scala 47:13]
  wire [1:0] PMPChecker_io_check_env_pmp_12_cfg_a; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pmp_12_cfg_x; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pmp_12_cfg_w; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pmp_12_cfg_r; // @[TLPMA.scala 47:13]
  wire [33:0] PMPChecker_io_check_env_pmp_12_addr; // @[TLPMA.scala 47:13]
  wire [35:0] PMPChecker_io_check_env_pmp_12_mask; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pmp_13_cfg_l; // @[TLPMA.scala 47:13]
  wire [1:0] PMPChecker_io_check_env_pmp_13_cfg_a; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pmp_13_cfg_x; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pmp_13_cfg_w; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pmp_13_cfg_r; // @[TLPMA.scala 47:13]
  wire [33:0] PMPChecker_io_check_env_pmp_13_addr; // @[TLPMA.scala 47:13]
  wire [35:0] PMPChecker_io_check_env_pmp_13_mask; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pmp_14_cfg_l; // @[TLPMA.scala 47:13]
  wire [1:0] PMPChecker_io_check_env_pmp_14_cfg_a; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pmp_14_cfg_x; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pmp_14_cfg_w; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pmp_14_cfg_r; // @[TLPMA.scala 47:13]
  wire [33:0] PMPChecker_io_check_env_pmp_14_addr; // @[TLPMA.scala 47:13]
  wire [35:0] PMPChecker_io_check_env_pmp_14_mask; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pmp_15_cfg_l; // @[TLPMA.scala 47:13]
  wire [1:0] PMPChecker_io_check_env_pmp_15_cfg_a; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pmp_15_cfg_x; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pmp_15_cfg_w; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pmp_15_cfg_r; // @[TLPMA.scala 47:13]
  wire [33:0] PMPChecker_io_check_env_pmp_15_addr; // @[TLPMA.scala 47:13]
  wire [35:0] PMPChecker_io_check_env_pmp_15_mask; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_0_cfg_c; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_0_cfg_atomic; // @[TLPMA.scala 47:13]
  wire [1:0] PMPChecker_io_check_env_pma_0_cfg_a; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_0_cfg_x; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_0_cfg_w; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_0_cfg_r; // @[TLPMA.scala 47:13]
  wire [33:0] PMPChecker_io_check_env_pma_0_addr; // @[TLPMA.scala 47:13]
  wire [35:0] PMPChecker_io_check_env_pma_0_mask; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_1_cfg_c; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_1_cfg_atomic; // @[TLPMA.scala 47:13]
  wire [1:0] PMPChecker_io_check_env_pma_1_cfg_a; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_1_cfg_x; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_1_cfg_w; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_1_cfg_r; // @[TLPMA.scala 47:13]
  wire [33:0] PMPChecker_io_check_env_pma_1_addr; // @[TLPMA.scala 47:13]
  wire [35:0] PMPChecker_io_check_env_pma_1_mask; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_2_cfg_c; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_2_cfg_atomic; // @[TLPMA.scala 47:13]
  wire [1:0] PMPChecker_io_check_env_pma_2_cfg_a; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_2_cfg_x; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_2_cfg_w; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_2_cfg_r; // @[TLPMA.scala 47:13]
  wire [33:0] PMPChecker_io_check_env_pma_2_addr; // @[TLPMA.scala 47:13]
  wire [35:0] PMPChecker_io_check_env_pma_2_mask; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_3_cfg_c; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_3_cfg_atomic; // @[TLPMA.scala 47:13]
  wire [1:0] PMPChecker_io_check_env_pma_3_cfg_a; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_3_cfg_x; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_3_cfg_w; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_3_cfg_r; // @[TLPMA.scala 47:13]
  wire [33:0] PMPChecker_io_check_env_pma_3_addr; // @[TLPMA.scala 47:13]
  wire [35:0] PMPChecker_io_check_env_pma_3_mask; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_4_cfg_c; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_4_cfg_atomic; // @[TLPMA.scala 47:13]
  wire [1:0] PMPChecker_io_check_env_pma_4_cfg_a; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_4_cfg_x; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_4_cfg_w; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_4_cfg_r; // @[TLPMA.scala 47:13]
  wire [33:0] PMPChecker_io_check_env_pma_4_addr; // @[TLPMA.scala 47:13]
  wire [35:0] PMPChecker_io_check_env_pma_4_mask; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_5_cfg_c; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_5_cfg_atomic; // @[TLPMA.scala 47:13]
  wire [1:0] PMPChecker_io_check_env_pma_5_cfg_a; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_5_cfg_x; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_5_cfg_w; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_5_cfg_r; // @[TLPMA.scala 47:13]
  wire [33:0] PMPChecker_io_check_env_pma_5_addr; // @[TLPMA.scala 47:13]
  wire [35:0] PMPChecker_io_check_env_pma_5_mask; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_6_cfg_c; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_6_cfg_atomic; // @[TLPMA.scala 47:13]
  wire [1:0] PMPChecker_io_check_env_pma_6_cfg_a; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_6_cfg_x; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_6_cfg_w; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_6_cfg_r; // @[TLPMA.scala 47:13]
  wire [33:0] PMPChecker_io_check_env_pma_6_addr; // @[TLPMA.scala 47:13]
  wire [35:0] PMPChecker_io_check_env_pma_6_mask; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_7_cfg_c; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_7_cfg_atomic; // @[TLPMA.scala 47:13]
  wire [1:0] PMPChecker_io_check_env_pma_7_cfg_a; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_7_cfg_x; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_7_cfg_w; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_7_cfg_r; // @[TLPMA.scala 47:13]
  wire [33:0] PMPChecker_io_check_env_pma_7_addr; // @[TLPMA.scala 47:13]
  wire [35:0] PMPChecker_io_check_env_pma_7_mask; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_8_cfg_c; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_8_cfg_atomic; // @[TLPMA.scala 47:13]
  wire [1:0] PMPChecker_io_check_env_pma_8_cfg_a; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_8_cfg_x; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_8_cfg_w; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_8_cfg_r; // @[TLPMA.scala 47:13]
  wire [33:0] PMPChecker_io_check_env_pma_8_addr; // @[TLPMA.scala 47:13]
  wire [35:0] PMPChecker_io_check_env_pma_8_mask; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_9_cfg_c; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_9_cfg_atomic; // @[TLPMA.scala 47:13]
  wire [1:0] PMPChecker_io_check_env_pma_9_cfg_a; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_9_cfg_x; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_9_cfg_w; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_9_cfg_r; // @[TLPMA.scala 47:13]
  wire [33:0] PMPChecker_io_check_env_pma_9_addr; // @[TLPMA.scala 47:13]
  wire [35:0] PMPChecker_io_check_env_pma_9_mask; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_10_cfg_c; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_10_cfg_atomic; // @[TLPMA.scala 47:13]
  wire [1:0] PMPChecker_io_check_env_pma_10_cfg_a; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_10_cfg_x; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_10_cfg_w; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_10_cfg_r; // @[TLPMA.scala 47:13]
  wire [33:0] PMPChecker_io_check_env_pma_10_addr; // @[TLPMA.scala 47:13]
  wire [35:0] PMPChecker_io_check_env_pma_10_mask; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_11_cfg_c; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_11_cfg_atomic; // @[TLPMA.scala 47:13]
  wire [1:0] PMPChecker_io_check_env_pma_11_cfg_a; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_11_cfg_x; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_11_cfg_w; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_11_cfg_r; // @[TLPMA.scala 47:13]
  wire [33:0] PMPChecker_io_check_env_pma_11_addr; // @[TLPMA.scala 47:13]
  wire [35:0] PMPChecker_io_check_env_pma_11_mask; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_12_cfg_c; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_12_cfg_atomic; // @[TLPMA.scala 47:13]
  wire [1:0] PMPChecker_io_check_env_pma_12_cfg_a; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_12_cfg_x; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_12_cfg_w; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_12_cfg_r; // @[TLPMA.scala 47:13]
  wire [33:0] PMPChecker_io_check_env_pma_12_addr; // @[TLPMA.scala 47:13]
  wire [35:0] PMPChecker_io_check_env_pma_12_mask; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_13_cfg_c; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_13_cfg_atomic; // @[TLPMA.scala 47:13]
  wire [1:0] PMPChecker_io_check_env_pma_13_cfg_a; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_13_cfg_x; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_13_cfg_w; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_13_cfg_r; // @[TLPMA.scala 47:13]
  wire [33:0] PMPChecker_io_check_env_pma_13_addr; // @[TLPMA.scala 47:13]
  wire [35:0] PMPChecker_io_check_env_pma_13_mask; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_14_cfg_c; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_14_cfg_atomic; // @[TLPMA.scala 47:13]
  wire [1:0] PMPChecker_io_check_env_pma_14_cfg_a; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_14_cfg_x; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_14_cfg_w; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_14_cfg_r; // @[TLPMA.scala 47:13]
  wire [33:0] PMPChecker_io_check_env_pma_14_addr; // @[TLPMA.scala 47:13]
  wire [35:0] PMPChecker_io_check_env_pma_14_mask; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_15_cfg_c; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_15_cfg_atomic; // @[TLPMA.scala 47:13]
  wire [1:0] PMPChecker_io_check_env_pma_15_cfg_a; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_15_cfg_x; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_15_cfg_w; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_check_env_pma_15_cfg_r; // @[TLPMA.scala 47:13]
  wire [33:0] PMPChecker_io_check_env_pma_15_addr; // @[TLPMA.scala 47:13]
  wire [35:0] PMPChecker_io_check_env_pma_15_mask; // @[TLPMA.scala 47:13]
  wire [35:0] PMPChecker_io_req_bits_addr; // @[TLPMA.scala 47:13]
  wire [2:0] PMPChecker_io_req_bits_cmd; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_resp_ld; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_resp_st; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_resp_instr; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_resp_mmio; // @[TLPMA.scala 47:13]
  wire  PMPChecker_io_resp_atomic; // @[TLPMA.scala 47:13]
  wire [1:0] PMPChecker_1_io_check_env_mode; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pmp_0_cfg_l; // @[TLPMA.scala 47:13]
  wire [1:0] PMPChecker_1_io_check_env_pmp_0_cfg_a; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pmp_0_cfg_x; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pmp_0_cfg_w; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pmp_0_cfg_r; // @[TLPMA.scala 47:13]
  wire [33:0] PMPChecker_1_io_check_env_pmp_0_addr; // @[TLPMA.scala 47:13]
  wire [35:0] PMPChecker_1_io_check_env_pmp_0_mask; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pmp_1_cfg_l; // @[TLPMA.scala 47:13]
  wire [1:0] PMPChecker_1_io_check_env_pmp_1_cfg_a; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pmp_1_cfg_x; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pmp_1_cfg_w; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pmp_1_cfg_r; // @[TLPMA.scala 47:13]
  wire [33:0] PMPChecker_1_io_check_env_pmp_1_addr; // @[TLPMA.scala 47:13]
  wire [35:0] PMPChecker_1_io_check_env_pmp_1_mask; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pmp_2_cfg_l; // @[TLPMA.scala 47:13]
  wire [1:0] PMPChecker_1_io_check_env_pmp_2_cfg_a; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pmp_2_cfg_x; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pmp_2_cfg_w; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pmp_2_cfg_r; // @[TLPMA.scala 47:13]
  wire [33:0] PMPChecker_1_io_check_env_pmp_2_addr; // @[TLPMA.scala 47:13]
  wire [35:0] PMPChecker_1_io_check_env_pmp_2_mask; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pmp_3_cfg_l; // @[TLPMA.scala 47:13]
  wire [1:0] PMPChecker_1_io_check_env_pmp_3_cfg_a; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pmp_3_cfg_x; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pmp_3_cfg_w; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pmp_3_cfg_r; // @[TLPMA.scala 47:13]
  wire [33:0] PMPChecker_1_io_check_env_pmp_3_addr; // @[TLPMA.scala 47:13]
  wire [35:0] PMPChecker_1_io_check_env_pmp_3_mask; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pmp_4_cfg_l; // @[TLPMA.scala 47:13]
  wire [1:0] PMPChecker_1_io_check_env_pmp_4_cfg_a; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pmp_4_cfg_x; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pmp_4_cfg_w; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pmp_4_cfg_r; // @[TLPMA.scala 47:13]
  wire [33:0] PMPChecker_1_io_check_env_pmp_4_addr; // @[TLPMA.scala 47:13]
  wire [35:0] PMPChecker_1_io_check_env_pmp_4_mask; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pmp_5_cfg_l; // @[TLPMA.scala 47:13]
  wire [1:0] PMPChecker_1_io_check_env_pmp_5_cfg_a; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pmp_5_cfg_x; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pmp_5_cfg_w; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pmp_5_cfg_r; // @[TLPMA.scala 47:13]
  wire [33:0] PMPChecker_1_io_check_env_pmp_5_addr; // @[TLPMA.scala 47:13]
  wire [35:0] PMPChecker_1_io_check_env_pmp_5_mask; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pmp_6_cfg_l; // @[TLPMA.scala 47:13]
  wire [1:0] PMPChecker_1_io_check_env_pmp_6_cfg_a; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pmp_6_cfg_x; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pmp_6_cfg_w; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pmp_6_cfg_r; // @[TLPMA.scala 47:13]
  wire [33:0] PMPChecker_1_io_check_env_pmp_6_addr; // @[TLPMA.scala 47:13]
  wire [35:0] PMPChecker_1_io_check_env_pmp_6_mask; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pmp_7_cfg_l; // @[TLPMA.scala 47:13]
  wire [1:0] PMPChecker_1_io_check_env_pmp_7_cfg_a; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pmp_7_cfg_x; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pmp_7_cfg_w; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pmp_7_cfg_r; // @[TLPMA.scala 47:13]
  wire [33:0] PMPChecker_1_io_check_env_pmp_7_addr; // @[TLPMA.scala 47:13]
  wire [35:0] PMPChecker_1_io_check_env_pmp_7_mask; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pmp_8_cfg_l; // @[TLPMA.scala 47:13]
  wire [1:0] PMPChecker_1_io_check_env_pmp_8_cfg_a; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pmp_8_cfg_x; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pmp_8_cfg_w; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pmp_8_cfg_r; // @[TLPMA.scala 47:13]
  wire [33:0] PMPChecker_1_io_check_env_pmp_8_addr; // @[TLPMA.scala 47:13]
  wire [35:0] PMPChecker_1_io_check_env_pmp_8_mask; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pmp_9_cfg_l; // @[TLPMA.scala 47:13]
  wire [1:0] PMPChecker_1_io_check_env_pmp_9_cfg_a; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pmp_9_cfg_x; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pmp_9_cfg_w; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pmp_9_cfg_r; // @[TLPMA.scala 47:13]
  wire [33:0] PMPChecker_1_io_check_env_pmp_9_addr; // @[TLPMA.scala 47:13]
  wire [35:0] PMPChecker_1_io_check_env_pmp_9_mask; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pmp_10_cfg_l; // @[TLPMA.scala 47:13]
  wire [1:0] PMPChecker_1_io_check_env_pmp_10_cfg_a; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pmp_10_cfg_x; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pmp_10_cfg_w; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pmp_10_cfg_r; // @[TLPMA.scala 47:13]
  wire [33:0] PMPChecker_1_io_check_env_pmp_10_addr; // @[TLPMA.scala 47:13]
  wire [35:0] PMPChecker_1_io_check_env_pmp_10_mask; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pmp_11_cfg_l; // @[TLPMA.scala 47:13]
  wire [1:0] PMPChecker_1_io_check_env_pmp_11_cfg_a; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pmp_11_cfg_x; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pmp_11_cfg_w; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pmp_11_cfg_r; // @[TLPMA.scala 47:13]
  wire [33:0] PMPChecker_1_io_check_env_pmp_11_addr; // @[TLPMA.scala 47:13]
  wire [35:0] PMPChecker_1_io_check_env_pmp_11_mask; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pmp_12_cfg_l; // @[TLPMA.scala 47:13]
  wire [1:0] PMPChecker_1_io_check_env_pmp_12_cfg_a; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pmp_12_cfg_x; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pmp_12_cfg_w; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pmp_12_cfg_r; // @[TLPMA.scala 47:13]
  wire [33:0] PMPChecker_1_io_check_env_pmp_12_addr; // @[TLPMA.scala 47:13]
  wire [35:0] PMPChecker_1_io_check_env_pmp_12_mask; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pmp_13_cfg_l; // @[TLPMA.scala 47:13]
  wire [1:0] PMPChecker_1_io_check_env_pmp_13_cfg_a; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pmp_13_cfg_x; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pmp_13_cfg_w; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pmp_13_cfg_r; // @[TLPMA.scala 47:13]
  wire [33:0] PMPChecker_1_io_check_env_pmp_13_addr; // @[TLPMA.scala 47:13]
  wire [35:0] PMPChecker_1_io_check_env_pmp_13_mask; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pmp_14_cfg_l; // @[TLPMA.scala 47:13]
  wire [1:0] PMPChecker_1_io_check_env_pmp_14_cfg_a; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pmp_14_cfg_x; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pmp_14_cfg_w; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pmp_14_cfg_r; // @[TLPMA.scala 47:13]
  wire [33:0] PMPChecker_1_io_check_env_pmp_14_addr; // @[TLPMA.scala 47:13]
  wire [35:0] PMPChecker_1_io_check_env_pmp_14_mask; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pmp_15_cfg_l; // @[TLPMA.scala 47:13]
  wire [1:0] PMPChecker_1_io_check_env_pmp_15_cfg_a; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pmp_15_cfg_x; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pmp_15_cfg_w; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pmp_15_cfg_r; // @[TLPMA.scala 47:13]
  wire [33:0] PMPChecker_1_io_check_env_pmp_15_addr; // @[TLPMA.scala 47:13]
  wire [35:0] PMPChecker_1_io_check_env_pmp_15_mask; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_0_cfg_c; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_0_cfg_atomic; // @[TLPMA.scala 47:13]
  wire [1:0] PMPChecker_1_io_check_env_pma_0_cfg_a; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_0_cfg_x; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_0_cfg_w; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_0_cfg_r; // @[TLPMA.scala 47:13]
  wire [33:0] PMPChecker_1_io_check_env_pma_0_addr; // @[TLPMA.scala 47:13]
  wire [35:0] PMPChecker_1_io_check_env_pma_0_mask; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_1_cfg_c; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_1_cfg_atomic; // @[TLPMA.scala 47:13]
  wire [1:0] PMPChecker_1_io_check_env_pma_1_cfg_a; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_1_cfg_x; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_1_cfg_w; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_1_cfg_r; // @[TLPMA.scala 47:13]
  wire [33:0] PMPChecker_1_io_check_env_pma_1_addr; // @[TLPMA.scala 47:13]
  wire [35:0] PMPChecker_1_io_check_env_pma_1_mask; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_2_cfg_c; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_2_cfg_atomic; // @[TLPMA.scala 47:13]
  wire [1:0] PMPChecker_1_io_check_env_pma_2_cfg_a; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_2_cfg_x; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_2_cfg_w; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_2_cfg_r; // @[TLPMA.scala 47:13]
  wire [33:0] PMPChecker_1_io_check_env_pma_2_addr; // @[TLPMA.scala 47:13]
  wire [35:0] PMPChecker_1_io_check_env_pma_2_mask; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_3_cfg_c; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_3_cfg_atomic; // @[TLPMA.scala 47:13]
  wire [1:0] PMPChecker_1_io_check_env_pma_3_cfg_a; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_3_cfg_x; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_3_cfg_w; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_3_cfg_r; // @[TLPMA.scala 47:13]
  wire [33:0] PMPChecker_1_io_check_env_pma_3_addr; // @[TLPMA.scala 47:13]
  wire [35:0] PMPChecker_1_io_check_env_pma_3_mask; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_4_cfg_c; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_4_cfg_atomic; // @[TLPMA.scala 47:13]
  wire [1:0] PMPChecker_1_io_check_env_pma_4_cfg_a; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_4_cfg_x; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_4_cfg_w; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_4_cfg_r; // @[TLPMA.scala 47:13]
  wire [33:0] PMPChecker_1_io_check_env_pma_4_addr; // @[TLPMA.scala 47:13]
  wire [35:0] PMPChecker_1_io_check_env_pma_4_mask; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_5_cfg_c; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_5_cfg_atomic; // @[TLPMA.scala 47:13]
  wire [1:0] PMPChecker_1_io_check_env_pma_5_cfg_a; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_5_cfg_x; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_5_cfg_w; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_5_cfg_r; // @[TLPMA.scala 47:13]
  wire [33:0] PMPChecker_1_io_check_env_pma_5_addr; // @[TLPMA.scala 47:13]
  wire [35:0] PMPChecker_1_io_check_env_pma_5_mask; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_6_cfg_c; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_6_cfg_atomic; // @[TLPMA.scala 47:13]
  wire [1:0] PMPChecker_1_io_check_env_pma_6_cfg_a; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_6_cfg_x; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_6_cfg_w; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_6_cfg_r; // @[TLPMA.scala 47:13]
  wire [33:0] PMPChecker_1_io_check_env_pma_6_addr; // @[TLPMA.scala 47:13]
  wire [35:0] PMPChecker_1_io_check_env_pma_6_mask; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_7_cfg_c; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_7_cfg_atomic; // @[TLPMA.scala 47:13]
  wire [1:0] PMPChecker_1_io_check_env_pma_7_cfg_a; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_7_cfg_x; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_7_cfg_w; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_7_cfg_r; // @[TLPMA.scala 47:13]
  wire [33:0] PMPChecker_1_io_check_env_pma_7_addr; // @[TLPMA.scala 47:13]
  wire [35:0] PMPChecker_1_io_check_env_pma_7_mask; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_8_cfg_c; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_8_cfg_atomic; // @[TLPMA.scala 47:13]
  wire [1:0] PMPChecker_1_io_check_env_pma_8_cfg_a; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_8_cfg_x; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_8_cfg_w; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_8_cfg_r; // @[TLPMA.scala 47:13]
  wire [33:0] PMPChecker_1_io_check_env_pma_8_addr; // @[TLPMA.scala 47:13]
  wire [35:0] PMPChecker_1_io_check_env_pma_8_mask; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_9_cfg_c; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_9_cfg_atomic; // @[TLPMA.scala 47:13]
  wire [1:0] PMPChecker_1_io_check_env_pma_9_cfg_a; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_9_cfg_x; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_9_cfg_w; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_9_cfg_r; // @[TLPMA.scala 47:13]
  wire [33:0] PMPChecker_1_io_check_env_pma_9_addr; // @[TLPMA.scala 47:13]
  wire [35:0] PMPChecker_1_io_check_env_pma_9_mask; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_10_cfg_c; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_10_cfg_atomic; // @[TLPMA.scala 47:13]
  wire [1:0] PMPChecker_1_io_check_env_pma_10_cfg_a; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_10_cfg_x; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_10_cfg_w; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_10_cfg_r; // @[TLPMA.scala 47:13]
  wire [33:0] PMPChecker_1_io_check_env_pma_10_addr; // @[TLPMA.scala 47:13]
  wire [35:0] PMPChecker_1_io_check_env_pma_10_mask; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_11_cfg_c; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_11_cfg_atomic; // @[TLPMA.scala 47:13]
  wire [1:0] PMPChecker_1_io_check_env_pma_11_cfg_a; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_11_cfg_x; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_11_cfg_w; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_11_cfg_r; // @[TLPMA.scala 47:13]
  wire [33:0] PMPChecker_1_io_check_env_pma_11_addr; // @[TLPMA.scala 47:13]
  wire [35:0] PMPChecker_1_io_check_env_pma_11_mask; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_12_cfg_c; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_12_cfg_atomic; // @[TLPMA.scala 47:13]
  wire [1:0] PMPChecker_1_io_check_env_pma_12_cfg_a; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_12_cfg_x; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_12_cfg_w; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_12_cfg_r; // @[TLPMA.scala 47:13]
  wire [33:0] PMPChecker_1_io_check_env_pma_12_addr; // @[TLPMA.scala 47:13]
  wire [35:0] PMPChecker_1_io_check_env_pma_12_mask; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_13_cfg_c; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_13_cfg_atomic; // @[TLPMA.scala 47:13]
  wire [1:0] PMPChecker_1_io_check_env_pma_13_cfg_a; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_13_cfg_x; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_13_cfg_w; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_13_cfg_r; // @[TLPMA.scala 47:13]
  wire [33:0] PMPChecker_1_io_check_env_pma_13_addr; // @[TLPMA.scala 47:13]
  wire [35:0] PMPChecker_1_io_check_env_pma_13_mask; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_14_cfg_c; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_14_cfg_atomic; // @[TLPMA.scala 47:13]
  wire [1:0] PMPChecker_1_io_check_env_pma_14_cfg_a; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_14_cfg_x; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_14_cfg_w; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_14_cfg_r; // @[TLPMA.scala 47:13]
  wire [33:0] PMPChecker_1_io_check_env_pma_14_addr; // @[TLPMA.scala 47:13]
  wire [35:0] PMPChecker_1_io_check_env_pma_14_mask; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_15_cfg_c; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_15_cfg_atomic; // @[TLPMA.scala 47:13]
  wire [1:0] PMPChecker_1_io_check_env_pma_15_cfg_a; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_15_cfg_x; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_15_cfg_w; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_check_env_pma_15_cfg_r; // @[TLPMA.scala 47:13]
  wire [33:0] PMPChecker_1_io_check_env_pma_15_addr; // @[TLPMA.scala 47:13]
  wire [35:0] PMPChecker_1_io_check_env_pma_15_mask; // @[TLPMA.scala 47:13]
  wire [35:0] PMPChecker_1_io_req_bits_addr; // @[TLPMA.scala 47:13]
  wire [2:0] PMPChecker_1_io_req_bits_cmd; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_resp_ld; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_resp_st; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_resp_instr; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_resp_mmio; // @[TLPMA.scala 47:13]
  wire  PMPChecker_1_io_resp_atomic; // @[TLPMA.scala 47:13]
  reg [63:0] pmaCfgMerged_0; // @[PMA.scala 50:31]
  reg [63:0] pmaCfgMerged_1; // @[PMA.scala 50:31]
  reg [33:0] addr_0; // @[PMA.scala 51:23]
  reg [33:0] addr_1; // @[PMA.scala 51:23]
  reg [33:0] addr_2; // @[PMA.scala 51:23]
  reg [33:0] addr_3; // @[PMA.scala 51:23]
  reg [33:0] addr_4; // @[PMA.scala 51:23]
  reg [33:0] addr_5; // @[PMA.scala 51:23]
  reg [33:0] addr_6; // @[PMA.scala 51:23]
  reg [33:0] addr_7; // @[PMA.scala 51:23]
  reg [33:0] addr_8; // @[PMA.scala 51:23]
  reg [33:0] addr_9; // @[PMA.scala 51:23]
  reg [33:0] addr_10; // @[PMA.scala 51:23]
  reg [33:0] addr_11; // @[PMA.scala 51:23]
  reg [33:0] addr_12; // @[PMA.scala 51:23]
  reg [33:0] addr_13; // @[PMA.scala 51:23]
  reg [33:0] addr_14; // @[PMA.scala 51:23]
  reg [33:0] addr_15; // @[PMA.scala 51:23]
  reg [35:0] mask_0; // @[PMA.scala 52:23]
  reg [35:0] mask_1; // @[PMA.scala 52:23]
  reg [35:0] mask_2; // @[PMA.scala 52:23]
  reg [35:0] mask_3; // @[PMA.scala 52:23]
  reg [35:0] mask_4; // @[PMA.scala 52:23]
  reg [35:0] mask_5; // @[PMA.scala 52:23]
  reg [35:0] mask_6; // @[PMA.scala 52:23]
  reg [35:0] mask_7; // @[PMA.scala 52:23]
  reg [35:0] mask_8; // @[PMA.scala 52:23]
  reg [35:0] mask_9; // @[PMA.scala 52:23]
  reg [35:0] mask_10; // @[PMA.scala 52:23]
  reg [35:0] mask_11; // @[PMA.scala 52:23]
  reg [35:0] mask_12; // @[PMA.scala 52:23]
  reg [35:0] mask_13; // @[PMA.scala 52:23]
  reg [35:0] mask_14; // @[PMA.scala 52:23]
  reg [35:0] mask_15; // @[PMA.scala 52:23]
  wire [127:0] _cfg_T = {pmaCfgMerged_1,pmaCfgMerged_0}; // @[PMA.scala 53:46]
  wire [1:0] cfg_0_a = _cfg_T[4:3]; // @[PMA.scala 53:46]
  wire  cfg_0_l = _cfg_T[7]; // @[PMA.scala 53:46]
  wire [1:0] cfg_1_a = _cfg_T[12:11]; // @[PMA.scala 53:46]
  wire  cfg_1_l = _cfg_T[15]; // @[PMA.scala 53:46]
  wire [1:0] cfg_2_a = _cfg_T[20:19]; // @[PMA.scala 53:46]
  wire  cfg_2_l = _cfg_T[23]; // @[PMA.scala 53:46]
  wire [1:0] cfg_3_a = _cfg_T[28:27]; // @[PMA.scala 53:46]
  wire  cfg_3_l = _cfg_T[31]; // @[PMA.scala 53:46]
  wire [1:0] cfg_4_a = _cfg_T[36:35]; // @[PMA.scala 53:46]
  wire  cfg_4_l = _cfg_T[39]; // @[PMA.scala 53:46]
  wire [1:0] cfg_5_a = _cfg_T[44:43]; // @[PMA.scala 53:46]
  wire  cfg_5_l = _cfg_T[47]; // @[PMA.scala 53:46]
  wire [1:0] cfg_6_a = _cfg_T[52:51]; // @[PMA.scala 53:46]
  wire  cfg_6_l = _cfg_T[55]; // @[PMA.scala 53:46]
  wire [1:0] cfg_7_a = _cfg_T[60:59]; // @[PMA.scala 53:46]
  wire  cfg_7_l = _cfg_T[63]; // @[PMA.scala 53:46]
  wire [1:0] cfg_8_a = _cfg_T[68:67]; // @[PMA.scala 53:46]
  wire  cfg_8_l = _cfg_T[71]; // @[PMA.scala 53:46]
  wire [1:0] cfg_9_a = _cfg_T[76:75]; // @[PMA.scala 53:46]
  wire  cfg_9_l = _cfg_T[79]; // @[PMA.scala 53:46]
  wire [1:0] cfg_10_a = _cfg_T[84:83]; // @[PMA.scala 53:46]
  wire  cfg_10_l = _cfg_T[87]; // @[PMA.scala 53:46]
  wire [1:0] cfg_11_a = _cfg_T[92:91]; // @[PMA.scala 53:46]
  wire  cfg_11_l = _cfg_T[95]; // @[PMA.scala 53:46]
  wire [1:0] cfg_12_a = _cfg_T[100:99]; // @[PMA.scala 53:46]
  wire  cfg_12_l = _cfg_T[103]; // @[PMA.scala 53:46]
  wire [1:0] cfg_13_a = _cfg_T[108:107]; // @[PMA.scala 53:46]
  wire  cfg_13_l = _cfg_T[111]; // @[PMA.scala 53:46]
  wire [1:0] cfg_14_a = _cfg_T[116:115]; // @[PMA.scala 53:46]
  wire  cfg_14_l = _cfg_T[119]; // @[PMA.scala 53:46]
  wire [1:0] cfg_15_a = _cfg_T[124:123]; // @[PMA.scala 53:46]
  wire  cfg_15_l = _cfg_T[127]; // @[PMA.scala 53:46]
  wire [33:0] _T_1 = addr_0 | 34'h1ff; // @[PMP.scala 126:10]
  wire [33:0] _T_3 = {addr_0[33:10],10'h0}; // @[Cat.scala 31:58]
  wire [33:0] _T_4 = cfg_0_a[1] ? _T_1 : _T_3; // @[PMP.scala 112:10]
  wire [63:0] _T_5 = {30'h0,_T_4}; // @[Cat.scala 31:58]
  wire [33:0] _T_7 = addr_1 | 34'h1ff; // @[PMP.scala 126:10]
  wire [33:0] _T_9 = {addr_1[33:10],10'h0}; // @[Cat.scala 31:58]
  wire [33:0] _T_10 = cfg_1_a[1] ? _T_7 : _T_9; // @[PMP.scala 112:10]
  wire [63:0] _T_11 = {30'h0,_T_10}; // @[Cat.scala 31:58]
  wire [33:0] _T_13 = addr_2 | 34'h1ff; // @[PMP.scala 126:10]
  wire [33:0] _T_15 = {addr_2[33:10],10'h0}; // @[Cat.scala 31:58]
  wire [33:0] _T_16 = cfg_2_a[1] ? _T_13 : _T_15; // @[PMP.scala 112:10]
  wire [63:0] _T_17 = {30'h0,_T_16}; // @[Cat.scala 31:58]
  wire [33:0] _T_19 = addr_3 | 34'h1ff; // @[PMP.scala 126:10]
  wire [33:0] _T_21 = {addr_3[33:10],10'h0}; // @[Cat.scala 31:58]
  wire [33:0] _T_22 = cfg_3_a[1] ? _T_19 : _T_21; // @[PMP.scala 112:10]
  wire [63:0] _T_23 = {30'h0,_T_22}; // @[Cat.scala 31:58]
  wire [33:0] _T_25 = addr_4 | 34'h1ff; // @[PMP.scala 126:10]
  wire [33:0] _T_27 = {addr_4[33:10],10'h0}; // @[Cat.scala 31:58]
  wire [33:0] _T_28 = cfg_4_a[1] ? _T_25 : _T_27; // @[PMP.scala 112:10]
  wire [63:0] _T_29 = {30'h0,_T_28}; // @[Cat.scala 31:58]
  wire [33:0] _T_31 = addr_5 | 34'h1ff; // @[PMP.scala 126:10]
  wire [33:0] _T_33 = {addr_5[33:10],10'h0}; // @[Cat.scala 31:58]
  wire [33:0] _T_34 = cfg_5_a[1] ? _T_31 : _T_33; // @[PMP.scala 112:10]
  wire [63:0] _T_35 = {30'h0,_T_34}; // @[Cat.scala 31:58]
  wire [33:0] _T_37 = addr_6 | 34'h1ff; // @[PMP.scala 126:10]
  wire [33:0] _T_39 = {addr_6[33:10],10'h0}; // @[Cat.scala 31:58]
  wire [33:0] _T_40 = cfg_6_a[1] ? _T_37 : _T_39; // @[PMP.scala 112:10]
  wire [63:0] _T_41 = {30'h0,_T_40}; // @[Cat.scala 31:58]
  wire [33:0] _T_43 = addr_7 | 34'h1ff; // @[PMP.scala 126:10]
  wire [33:0] _T_45 = {addr_7[33:10],10'h0}; // @[Cat.scala 31:58]
  wire [33:0] _T_46 = cfg_7_a[1] ? _T_43 : _T_45; // @[PMP.scala 112:10]
  wire [63:0] _T_47 = {30'h0,_T_46}; // @[Cat.scala 31:58]
  wire [33:0] _T_49 = addr_8 | 34'h1ff; // @[PMP.scala 126:10]
  wire [33:0] _T_51 = {addr_8[33:10],10'h0}; // @[Cat.scala 31:58]
  wire [33:0] _T_52 = cfg_8_a[1] ? _T_49 : _T_51; // @[PMP.scala 112:10]
  wire [63:0] _T_53 = {30'h0,_T_52}; // @[Cat.scala 31:58]
  wire [33:0] _T_55 = addr_9 | 34'h1ff; // @[PMP.scala 126:10]
  wire [33:0] _T_57 = {addr_9[33:10],10'h0}; // @[Cat.scala 31:58]
  wire [33:0] _T_58 = cfg_9_a[1] ? _T_55 : _T_57; // @[PMP.scala 112:10]
  wire [63:0] _T_59 = {30'h0,_T_58}; // @[Cat.scala 31:58]
  wire [33:0] _T_61 = addr_10 | 34'h1ff; // @[PMP.scala 126:10]
  wire [33:0] _T_63 = {addr_10[33:10],10'h0}; // @[Cat.scala 31:58]
  wire [33:0] _T_64 = cfg_10_a[1] ? _T_61 : _T_63; // @[PMP.scala 112:10]
  wire [63:0] _T_65 = {30'h0,_T_64}; // @[Cat.scala 31:58]
  wire [33:0] _T_67 = addr_11 | 34'h1ff; // @[PMP.scala 126:10]
  wire [33:0] _T_69 = {addr_11[33:10],10'h0}; // @[Cat.scala 31:58]
  wire [33:0] _T_70 = cfg_11_a[1] ? _T_67 : _T_69; // @[PMP.scala 112:10]
  wire [63:0] _T_71 = {30'h0,_T_70}; // @[Cat.scala 31:58]
  wire [33:0] _T_73 = addr_12 | 34'h1ff; // @[PMP.scala 126:10]
  wire [33:0] _T_75 = {addr_12[33:10],10'h0}; // @[Cat.scala 31:58]
  wire [33:0] _T_76 = cfg_12_a[1] ? _T_73 : _T_75; // @[PMP.scala 112:10]
  wire [63:0] _T_77 = {30'h0,_T_76}; // @[Cat.scala 31:58]
  wire [33:0] _T_79 = addr_13 | 34'h1ff; // @[PMP.scala 126:10]
  wire [33:0] _T_81 = {addr_13[33:10],10'h0}; // @[Cat.scala 31:58]
  wire [33:0] _T_82 = cfg_13_a[1] ? _T_79 : _T_81; // @[PMP.scala 112:10]
  wire [63:0] _T_83 = {30'h0,_T_82}; // @[Cat.scala 31:58]
  wire [33:0] _T_85 = addr_14 | 34'h1ff; // @[PMP.scala 126:10]
  wire [33:0] _T_87 = {addr_14[33:10],10'h0}; // @[Cat.scala 31:58]
  wire [33:0] _T_88 = cfg_14_a[1] ? _T_85 : _T_87; // @[PMP.scala 112:10]
  wire [63:0] _T_89 = {30'h0,_T_88}; // @[Cat.scala 31:58]
  wire [33:0] _T_91 = addr_15 | 34'h1ff; // @[PMP.scala 126:10]
  wire [33:0] _T_93 = {addr_15[33:10],10'h0}; // @[Cat.scala 31:58]
  wire [33:0] _T_94 = cfg_15_a[1] ? _T_91 : _T_93; // @[PMP.scala 112:10]
  wire [63:0] _T_95 = {30'h0,_T_94}; // @[Cat.scala 31:58]
  wire  in_bits_read = auto_in_a_bits_opcode == 3'h4; // @[RegisterRouter.scala 71:36]
  wire [8:0] in_bits_index = auto_in_a_bits_address[11:3]; // @[RegisterRouter.scala 70:18 72:19]
  wire [8:0] out_findex = in_bits_index & 9'h1d0; // @[RegisterRouter.scala 82:24]
  wire [8:0] out_bindex = out_back_io_deq_bits_index & 9'h1d0; // @[RegisterRouter.scala 82:24]
  wire  _out_T_1 = out_bindex == 9'h0; // @[RegisterRouter.scala 82:24]
  wire [7:0] _out_frontMask_T_9 = auto_in_a_bits_mask[0] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _out_frontMask_T_11 = auto_in_a_bits_mask[1] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _out_frontMask_T_13 = auto_in_a_bits_mask[2] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _out_frontMask_T_15 = auto_in_a_bits_mask[3] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _out_frontMask_T_17 = auto_in_a_bits_mask[4] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _out_frontMask_T_19 = auto_in_a_bits_mask[5] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _out_frontMask_T_21 = auto_in_a_bits_mask[6] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _out_frontMask_T_23 = auto_in_a_bits_mask[7] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [63:0] out_frontMask = {_out_frontMask_T_23,_out_frontMask_T_21,_out_frontMask_T_19,_out_frontMask_T_17,
    _out_frontMask_T_15,_out_frontMask_T_13,_out_frontMask_T_11,_out_frontMask_T_9}; // @[Cat.scala 31:58]
  wire [7:0] _out_backMask_T_9 = out_back_io_deq_bits_mask[0] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _out_backMask_T_11 = out_back_io_deq_bits_mask[1] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _out_backMask_T_13 = out_back_io_deq_bits_mask[2] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _out_backMask_T_15 = out_back_io_deq_bits_mask[3] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _out_backMask_T_17 = out_back_io_deq_bits_mask[4] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _out_backMask_T_19 = out_back_io_deq_bits_mask[5] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _out_backMask_T_21 = out_back_io_deq_bits_mask[6] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _out_backMask_T_23 = out_back_io_deq_bits_mask[7] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [63:0] out_backMask = {_out_backMask_T_23,_out_backMask_T_21,_out_backMask_T_19,_out_backMask_T_17,
    _out_backMask_T_15,_out_backMask_T_13,_out_backMask_T_11,_out_backMask_T_9}; // @[Cat.scala 31:58]
  wire  out_rimask = |out_frontMask; // @[RegisterRouter.scala 82:24]
  wire  out_romask = |out_backMask; // @[RegisterRouter.scala 82:24]
  wire  out_womask = &out_backMask; // @[RegisterRouter.scala 82:24]
  wire  out_front_ready = out_back_io_enq_ready; // @[Decoupled.scala 365:17 RegisterRouter.scala 82:24]
  wire [4:0] out_iindex = {in_bits_index[5],in_bits_index[3],in_bits_index[2],in_bits_index[1],in_bits_index[0]}; // @[Cat.scala 31:58]
  wire [31:0] _out_frontSel_T = 32'h1 << out_iindex; // @[OneHot.scala 57:35]
  wire  out_frontSel_0 = _out_frontSel_T[0]; // @[RegisterRouter.scala 82:24]
  wire  out_rivalid_0 = auto_in_a_valid & out_front_ready & in_bits_read & out_frontSel_0 & out_findex == 9'h0; // @[RegisterRouter.scala 82:24]
  wire  out_f_rivalid = out_rivalid_0 & out_rimask; // @[RegisterRouter.scala 82:24]
  wire [4:0] out_oindex = {out_back_io_deq_bits_index[5],out_back_io_deq_bits_index[3],out_back_io_deq_bits_index[2],
    out_back_io_deq_bits_index[1],out_back_io_deq_bits_index[0]}; // @[Cat.scala 31:58]
  wire [31:0] _out_backSel_T = 32'h1 << out_oindex; // @[OneHot.scala 57:35]
  wire  out_backSel_0 = _out_backSel_T[0]; // @[RegisterRouter.scala 82:24]
  wire  out_roready_0 = out_back_io_deq_valid & auto_in_d_ready & out_back_io_deq_bits_read & out_backSel_0 & out_bindex
     == 9'h0; // @[RegisterRouter.scala 82:24]
  wire  out_f_roready = out_roready_0 & out_romask; // @[RegisterRouter.scala 82:24]
  wire  out_woready_0 = out_back_io_deq_valid & auto_in_d_ready & ~out_back_io_deq_bits_read & out_backSel_0 &
    out_bindex == 9'h0; // @[RegisterRouter.scala 82:24]
  wire  out_f_woready = out_woready_0 & out_womask; // @[RegisterRouter.scala 82:24]
  reg  out_v_reg; // @[Hold.scala 40:24]
  wire  out_f_riready = ~out_v_reg; // @[PMA.scala 67:20]
  wire  _out_v_reg_T = out_f_riready & out_f_rivalid; // @[PMA.scala 66:39]
  wire  _out_v_reg_T_1 = out_v_reg & out_f_roready; // @[PMA.scala 66:58]
  wire  _GEN_0 = _out_v_reg_T_1 ? 1'h0 : out_v_reg; // @[Hold.scala 41:20 40:24 41:28]
  wire [63:0] _out_T_40 = out_back_io_deq_bits_data; // @[RegisterRouter.scala 82:24]
  wire  out_pmaCfgMerged_0_cfg_wm_tmp_r = _out_T_40[0]; // @[PMP.scala 93:61]
  wire  out_pmaCfgMerged_0_cfg_wm_tmp_w = _out_T_40[1]; // @[PMP.scala 93:61]
  wire  out_pmaCfgMerged_0_cfg_wm_tmp_x = _out_T_40[2]; // @[PMP.scala 93:61]
  wire [1:0] out_pmaCfgMerged_0_cfg_wm_tmp_a = _out_T_40[4:3]; // @[PMP.scala 93:61]
  wire  out_pmaCfgMerged_0_cfg_wm_tmp_atomic = _out_T_40[5]; // @[PMP.scala 93:61]
  wire  out_pmaCfgMerged_0_cfg_wm_tmp_c = _out_T_40[6]; // @[PMP.scala 93:61]
  wire  out_pmaCfgMerged_0_cfg_wm_tmp_l = _out_T_40[7]; // @[PMP.scala 93:61]
  wire  _out_pmaCfgMerged_0_cfgVec_0_a_T_1 = |out_pmaCfgMerged_0_cfg_wm_tmp_a; // @[PMP.scala 97:80]
  wire [1:0] _out_pmaCfgMerged_0_cfgVec_0_a_T_2 = {out_pmaCfgMerged_0_cfg_wm_tmp_a[1],
    _out_pmaCfgMerged_0_cfgVec_0_a_T_1}; // @[Cat.scala 31:58]
  wire [1:0] out_pmaCfgMerged_0_cfgVec_0_a = ~out_pmaCfgMerged_0_cfg_wm_tmp_l ? _out_pmaCfgMerged_0_cfgVec_0_a_T_2 :
    out_pmaCfgMerged_0_cfg_wm_tmp_a; // @[PMP.scala 94:17 95:29 97:41]
  wire [34:0] _out_pmaCfgMerged_0_mask_0_match_mask_c_addr_T_1 = {addr_0,out_pmaCfgMerged_0_cfgVec_0_a[0]}; // @[Cat.scala 31:58]
  wire [34:0] out_pmaCfgMerged_0_mask_0_match_mask_c_addr = _out_pmaCfgMerged_0_mask_0_match_mask_c_addr_T_1 | 35'h3ff; // @[PMP.scala 86:50]
  wire [34:0] _out_pmaCfgMerged_0_mask_0_T_1 = out_pmaCfgMerged_0_mask_0_match_mask_c_addr + 35'h1; // @[PMP.scala 87:49]
  wire [34:0] _out_pmaCfgMerged_0_mask_0_T_2 = ~_out_pmaCfgMerged_0_mask_0_T_1; // @[PMP.scala 87:29]
  wire [34:0] _out_pmaCfgMerged_0_mask_0_T_3 = out_pmaCfgMerged_0_mask_0_match_mask_c_addr &
    _out_pmaCfgMerged_0_mask_0_T_2; // @[PMP.scala 87:27]
  wire [36:0] _out_pmaCfgMerged_0_mask_0_T_4 = {_out_pmaCfgMerged_0_mask_0_T_3,2'h3}; // @[Cat.scala 31:58]
  wire [36:0] _GEN_3 = out_pmaCfgMerged_0_cfgVec_0_a[1] ? _out_pmaCfgMerged_0_mask_0_T_4 : {{1'd0}, mask_0}; // @[PMA.scala 52:23 PMP.scala 98:36 99:27]
  wire  out_pmaCfgMerged_0_cfgVec_0_w = ~out_pmaCfgMerged_0_cfg_wm_tmp_l ? out_pmaCfgMerged_0_cfg_wm_tmp_w &
    out_pmaCfgMerged_0_cfg_wm_tmp_r : out_pmaCfgMerged_0_cfg_wm_tmp_w; // @[PMP.scala 94:17 95:29 96:21]
  wire [36:0] _GEN_6 = ~out_pmaCfgMerged_0_cfg_wm_tmp_l ? _GEN_3 : {{1'd0}, mask_0}; // @[PMA.scala 52:23 PMP.scala 95:29]
  wire  out_pmaCfgMerged_0_cfg_wm_tmp_1_r = _out_T_40[8]; // @[PMP.scala 93:61]
  wire  out_pmaCfgMerged_0_cfg_wm_tmp_1_w = _out_T_40[9]; // @[PMP.scala 93:61]
  wire  out_pmaCfgMerged_0_cfg_wm_tmp_1_x = _out_T_40[10]; // @[PMP.scala 93:61]
  wire [1:0] out_pmaCfgMerged_0_cfg_wm_tmp_1_a = _out_T_40[12:11]; // @[PMP.scala 93:61]
  wire  out_pmaCfgMerged_0_cfg_wm_tmp_1_atomic = _out_T_40[13]; // @[PMP.scala 93:61]
  wire  out_pmaCfgMerged_0_cfg_wm_tmp_1_c = _out_T_40[14]; // @[PMP.scala 93:61]
  wire  out_pmaCfgMerged_0_cfg_wm_tmp_1_l = _out_T_40[15]; // @[PMP.scala 93:61]
  wire  _out_pmaCfgMerged_0_cfgVec_1_a_T_1 = |out_pmaCfgMerged_0_cfg_wm_tmp_1_a; // @[PMP.scala 97:80]
  wire [1:0] _out_pmaCfgMerged_0_cfgVec_1_a_T_2 = {out_pmaCfgMerged_0_cfg_wm_tmp_1_a[1],
    _out_pmaCfgMerged_0_cfgVec_1_a_T_1}; // @[Cat.scala 31:58]
  wire [1:0] out_pmaCfgMerged_0_cfgVec_1_a = ~out_pmaCfgMerged_0_cfg_wm_tmp_1_l ? _out_pmaCfgMerged_0_cfgVec_1_a_T_2 :
    out_pmaCfgMerged_0_cfg_wm_tmp_1_a; // @[PMP.scala 94:17 95:29 97:41]
  wire [34:0] _out_pmaCfgMerged_0_mask_1_match_mask_c_addr_T_1 = {addr_1,out_pmaCfgMerged_0_cfgVec_1_a[0]}; // @[Cat.scala 31:58]
  wire [34:0] out_pmaCfgMerged_0_mask_1_match_mask_c_addr = _out_pmaCfgMerged_0_mask_1_match_mask_c_addr_T_1 | 35'h3ff; // @[PMP.scala 86:50]
  wire [34:0] _out_pmaCfgMerged_0_mask_1_T_1 = out_pmaCfgMerged_0_mask_1_match_mask_c_addr + 35'h1; // @[PMP.scala 87:49]
  wire [34:0] _out_pmaCfgMerged_0_mask_1_T_2 = ~_out_pmaCfgMerged_0_mask_1_T_1; // @[PMP.scala 87:29]
  wire [34:0] _out_pmaCfgMerged_0_mask_1_T_3 = out_pmaCfgMerged_0_mask_1_match_mask_c_addr &
    _out_pmaCfgMerged_0_mask_1_T_2; // @[PMP.scala 87:27]
  wire [36:0] _out_pmaCfgMerged_0_mask_1_T_4 = {_out_pmaCfgMerged_0_mask_1_T_3,2'h3}; // @[Cat.scala 31:58]
  wire [36:0] _GEN_7 = out_pmaCfgMerged_0_cfgVec_1_a[1] ? _out_pmaCfgMerged_0_mask_1_T_4 : {{1'd0}, mask_1}; // @[PMA.scala 52:23 PMP.scala 98:36 99:27]
  wire  out_pmaCfgMerged_0_cfgVec_1_w = ~out_pmaCfgMerged_0_cfg_wm_tmp_1_l ? out_pmaCfgMerged_0_cfg_wm_tmp_1_w &
    out_pmaCfgMerged_0_cfg_wm_tmp_1_r : out_pmaCfgMerged_0_cfg_wm_tmp_1_w; // @[PMP.scala 94:17 95:29 96:21]
  wire [36:0] _GEN_10 = ~out_pmaCfgMerged_0_cfg_wm_tmp_1_l ? _GEN_7 : {{1'd0}, mask_1}; // @[PMA.scala 52:23 PMP.scala 95:29]
  wire  out_pmaCfgMerged_0_cfg_wm_tmp_2_r = _out_T_40[16]; // @[PMP.scala 93:61]
  wire  out_pmaCfgMerged_0_cfg_wm_tmp_2_w = _out_T_40[17]; // @[PMP.scala 93:61]
  wire  out_pmaCfgMerged_0_cfg_wm_tmp_2_x = _out_T_40[18]; // @[PMP.scala 93:61]
  wire [1:0] out_pmaCfgMerged_0_cfg_wm_tmp_2_a = _out_T_40[20:19]; // @[PMP.scala 93:61]
  wire  out_pmaCfgMerged_0_cfg_wm_tmp_2_atomic = _out_T_40[21]; // @[PMP.scala 93:61]
  wire  out_pmaCfgMerged_0_cfg_wm_tmp_2_c = _out_T_40[22]; // @[PMP.scala 93:61]
  wire  out_pmaCfgMerged_0_cfg_wm_tmp_2_l = _out_T_40[23]; // @[PMP.scala 93:61]
  wire  _out_pmaCfgMerged_0_cfgVec_2_a_T_1 = |out_pmaCfgMerged_0_cfg_wm_tmp_2_a; // @[PMP.scala 97:80]
  wire [1:0] _out_pmaCfgMerged_0_cfgVec_2_a_T_2 = {out_pmaCfgMerged_0_cfg_wm_tmp_2_a[1],
    _out_pmaCfgMerged_0_cfgVec_2_a_T_1}; // @[Cat.scala 31:58]
  wire [1:0] out_pmaCfgMerged_0_cfgVec_2_a = ~out_pmaCfgMerged_0_cfg_wm_tmp_2_l ? _out_pmaCfgMerged_0_cfgVec_2_a_T_2 :
    out_pmaCfgMerged_0_cfg_wm_tmp_2_a; // @[PMP.scala 94:17 95:29 97:41]
  wire [34:0] _out_pmaCfgMerged_0_mask_2_match_mask_c_addr_T_1 = {addr_2,out_pmaCfgMerged_0_cfgVec_2_a[0]}; // @[Cat.scala 31:58]
  wire [34:0] out_pmaCfgMerged_0_mask_2_match_mask_c_addr = _out_pmaCfgMerged_0_mask_2_match_mask_c_addr_T_1 | 35'h3ff; // @[PMP.scala 86:50]
  wire [34:0] _out_pmaCfgMerged_0_mask_2_T_1 = out_pmaCfgMerged_0_mask_2_match_mask_c_addr + 35'h1; // @[PMP.scala 87:49]
  wire [34:0] _out_pmaCfgMerged_0_mask_2_T_2 = ~_out_pmaCfgMerged_0_mask_2_T_1; // @[PMP.scala 87:29]
  wire [34:0] _out_pmaCfgMerged_0_mask_2_T_3 = out_pmaCfgMerged_0_mask_2_match_mask_c_addr &
    _out_pmaCfgMerged_0_mask_2_T_2; // @[PMP.scala 87:27]
  wire [36:0] _out_pmaCfgMerged_0_mask_2_T_4 = {_out_pmaCfgMerged_0_mask_2_T_3,2'h3}; // @[Cat.scala 31:58]
  wire [36:0] _GEN_11 = out_pmaCfgMerged_0_cfgVec_2_a[1] ? _out_pmaCfgMerged_0_mask_2_T_4 : {{1'd0}, mask_2}; // @[PMA.scala 52:23 PMP.scala 98:36 99:27]
  wire  out_pmaCfgMerged_0_cfgVec_2_w = ~out_pmaCfgMerged_0_cfg_wm_tmp_2_l ? out_pmaCfgMerged_0_cfg_wm_tmp_2_w &
    out_pmaCfgMerged_0_cfg_wm_tmp_2_r : out_pmaCfgMerged_0_cfg_wm_tmp_2_w; // @[PMP.scala 94:17 95:29 96:21]
  wire [36:0] _GEN_14 = ~out_pmaCfgMerged_0_cfg_wm_tmp_2_l ? _GEN_11 : {{1'd0}, mask_2}; // @[PMA.scala 52:23 PMP.scala 95:29]
  wire  out_pmaCfgMerged_0_cfg_wm_tmp_3_r = _out_T_40[24]; // @[PMP.scala 93:61]
  wire  out_pmaCfgMerged_0_cfg_wm_tmp_3_w = _out_T_40[25]; // @[PMP.scala 93:61]
  wire  out_pmaCfgMerged_0_cfg_wm_tmp_3_x = _out_T_40[26]; // @[PMP.scala 93:61]
  wire [1:0] out_pmaCfgMerged_0_cfg_wm_tmp_3_a = _out_T_40[28:27]; // @[PMP.scala 93:61]
  wire  out_pmaCfgMerged_0_cfg_wm_tmp_3_atomic = _out_T_40[29]; // @[PMP.scala 93:61]
  wire  out_pmaCfgMerged_0_cfg_wm_tmp_3_c = _out_T_40[30]; // @[PMP.scala 93:61]
  wire  out_pmaCfgMerged_0_cfg_wm_tmp_3_l = _out_T_40[31]; // @[PMP.scala 93:61]
  wire  _out_pmaCfgMerged_0_cfgVec_3_a_T_1 = |out_pmaCfgMerged_0_cfg_wm_tmp_3_a; // @[PMP.scala 97:80]
  wire [1:0] _out_pmaCfgMerged_0_cfgVec_3_a_T_2 = {out_pmaCfgMerged_0_cfg_wm_tmp_3_a[1],
    _out_pmaCfgMerged_0_cfgVec_3_a_T_1}; // @[Cat.scala 31:58]
  wire [1:0] out_pmaCfgMerged_0_cfgVec_3_a = ~out_pmaCfgMerged_0_cfg_wm_tmp_3_l ? _out_pmaCfgMerged_0_cfgVec_3_a_T_2 :
    out_pmaCfgMerged_0_cfg_wm_tmp_3_a; // @[PMP.scala 94:17 95:29 97:41]
  wire [34:0] _out_pmaCfgMerged_0_mask_3_match_mask_c_addr_T_1 = {addr_3,out_pmaCfgMerged_0_cfgVec_3_a[0]}; // @[Cat.scala 31:58]
  wire [34:0] out_pmaCfgMerged_0_mask_3_match_mask_c_addr = _out_pmaCfgMerged_0_mask_3_match_mask_c_addr_T_1 | 35'h3ff; // @[PMP.scala 86:50]
  wire [34:0] _out_pmaCfgMerged_0_mask_3_T_1 = out_pmaCfgMerged_0_mask_3_match_mask_c_addr + 35'h1; // @[PMP.scala 87:49]
  wire [34:0] _out_pmaCfgMerged_0_mask_3_T_2 = ~_out_pmaCfgMerged_0_mask_3_T_1; // @[PMP.scala 87:29]
  wire [34:0] _out_pmaCfgMerged_0_mask_3_T_3 = out_pmaCfgMerged_0_mask_3_match_mask_c_addr &
    _out_pmaCfgMerged_0_mask_3_T_2; // @[PMP.scala 87:27]
  wire [36:0] _out_pmaCfgMerged_0_mask_3_T_4 = {_out_pmaCfgMerged_0_mask_3_T_3,2'h3}; // @[Cat.scala 31:58]
  wire [36:0] _GEN_15 = out_pmaCfgMerged_0_cfgVec_3_a[1] ? _out_pmaCfgMerged_0_mask_3_T_4 : {{1'd0}, mask_3}; // @[PMA.scala 52:23 PMP.scala 98:36 99:27]
  wire  out_pmaCfgMerged_0_cfgVec_3_w = ~out_pmaCfgMerged_0_cfg_wm_tmp_3_l ? out_pmaCfgMerged_0_cfg_wm_tmp_3_w &
    out_pmaCfgMerged_0_cfg_wm_tmp_3_r : out_pmaCfgMerged_0_cfg_wm_tmp_3_w; // @[PMP.scala 94:17 95:29 96:21]
  wire [36:0] _GEN_18 = ~out_pmaCfgMerged_0_cfg_wm_tmp_3_l ? _GEN_15 : {{1'd0}, mask_3}; // @[PMA.scala 52:23 PMP.scala 95:29]
  wire  out_pmaCfgMerged_0_cfg_wm_tmp_4_r = _out_T_40[32]; // @[PMP.scala 93:61]
  wire  out_pmaCfgMerged_0_cfg_wm_tmp_4_w = _out_T_40[33]; // @[PMP.scala 93:61]
  wire  out_pmaCfgMerged_0_cfg_wm_tmp_4_x = _out_T_40[34]; // @[PMP.scala 93:61]
  wire [1:0] out_pmaCfgMerged_0_cfg_wm_tmp_4_a = _out_T_40[36:35]; // @[PMP.scala 93:61]
  wire  out_pmaCfgMerged_0_cfg_wm_tmp_4_atomic = _out_T_40[37]; // @[PMP.scala 93:61]
  wire  out_pmaCfgMerged_0_cfg_wm_tmp_4_c = _out_T_40[38]; // @[PMP.scala 93:61]
  wire  out_pmaCfgMerged_0_cfg_wm_tmp_4_l = _out_T_40[39]; // @[PMP.scala 93:61]
  wire  _out_pmaCfgMerged_0_cfgVec_4_a_T_1 = |out_pmaCfgMerged_0_cfg_wm_tmp_4_a; // @[PMP.scala 97:80]
  wire [1:0] _out_pmaCfgMerged_0_cfgVec_4_a_T_2 = {out_pmaCfgMerged_0_cfg_wm_tmp_4_a[1],
    _out_pmaCfgMerged_0_cfgVec_4_a_T_1}; // @[Cat.scala 31:58]
  wire [1:0] out_pmaCfgMerged_0_cfgVec_4_a = ~out_pmaCfgMerged_0_cfg_wm_tmp_4_l ? _out_pmaCfgMerged_0_cfgVec_4_a_T_2 :
    out_pmaCfgMerged_0_cfg_wm_tmp_4_a; // @[PMP.scala 94:17 95:29 97:41]
  wire [34:0] _out_pmaCfgMerged_0_mask_4_match_mask_c_addr_T_1 = {addr_4,out_pmaCfgMerged_0_cfgVec_4_a[0]}; // @[Cat.scala 31:58]
  wire [34:0] out_pmaCfgMerged_0_mask_4_match_mask_c_addr = _out_pmaCfgMerged_0_mask_4_match_mask_c_addr_T_1 | 35'h3ff; // @[PMP.scala 86:50]
  wire [34:0] _out_pmaCfgMerged_0_mask_4_T_1 = out_pmaCfgMerged_0_mask_4_match_mask_c_addr + 35'h1; // @[PMP.scala 87:49]
  wire [34:0] _out_pmaCfgMerged_0_mask_4_T_2 = ~_out_pmaCfgMerged_0_mask_4_T_1; // @[PMP.scala 87:29]
  wire [34:0] _out_pmaCfgMerged_0_mask_4_T_3 = out_pmaCfgMerged_0_mask_4_match_mask_c_addr &
    _out_pmaCfgMerged_0_mask_4_T_2; // @[PMP.scala 87:27]
  wire [36:0] _out_pmaCfgMerged_0_mask_4_T_4 = {_out_pmaCfgMerged_0_mask_4_T_3,2'h3}; // @[Cat.scala 31:58]
  wire [36:0] _GEN_19 = out_pmaCfgMerged_0_cfgVec_4_a[1] ? _out_pmaCfgMerged_0_mask_4_T_4 : {{1'd0}, mask_4}; // @[PMA.scala 52:23 PMP.scala 98:36 99:27]
  wire  out_pmaCfgMerged_0_cfgVec_4_w = ~out_pmaCfgMerged_0_cfg_wm_tmp_4_l ? out_pmaCfgMerged_0_cfg_wm_tmp_4_w &
    out_pmaCfgMerged_0_cfg_wm_tmp_4_r : out_pmaCfgMerged_0_cfg_wm_tmp_4_w; // @[PMP.scala 94:17 95:29 96:21]
  wire [36:0] _GEN_22 = ~out_pmaCfgMerged_0_cfg_wm_tmp_4_l ? _GEN_19 : {{1'd0}, mask_4}; // @[PMA.scala 52:23 PMP.scala 95:29]
  wire  out_pmaCfgMerged_0_cfg_wm_tmp_5_r = _out_T_40[40]; // @[PMP.scala 93:61]
  wire  out_pmaCfgMerged_0_cfg_wm_tmp_5_w = _out_T_40[41]; // @[PMP.scala 93:61]
  wire  out_pmaCfgMerged_0_cfg_wm_tmp_5_x = _out_T_40[42]; // @[PMP.scala 93:61]
  wire [1:0] out_pmaCfgMerged_0_cfg_wm_tmp_5_a = _out_T_40[44:43]; // @[PMP.scala 93:61]
  wire  out_pmaCfgMerged_0_cfg_wm_tmp_5_atomic = _out_T_40[45]; // @[PMP.scala 93:61]
  wire  out_pmaCfgMerged_0_cfg_wm_tmp_5_c = _out_T_40[46]; // @[PMP.scala 93:61]
  wire  out_pmaCfgMerged_0_cfg_wm_tmp_5_l = _out_T_40[47]; // @[PMP.scala 93:61]
  wire  _out_pmaCfgMerged_0_cfgVec_5_a_T_1 = |out_pmaCfgMerged_0_cfg_wm_tmp_5_a; // @[PMP.scala 97:80]
  wire [1:0] _out_pmaCfgMerged_0_cfgVec_5_a_T_2 = {out_pmaCfgMerged_0_cfg_wm_tmp_5_a[1],
    _out_pmaCfgMerged_0_cfgVec_5_a_T_1}; // @[Cat.scala 31:58]
  wire [1:0] out_pmaCfgMerged_0_cfgVec_5_a = ~out_pmaCfgMerged_0_cfg_wm_tmp_5_l ? _out_pmaCfgMerged_0_cfgVec_5_a_T_2 :
    out_pmaCfgMerged_0_cfg_wm_tmp_5_a; // @[PMP.scala 94:17 95:29 97:41]
  wire [34:0] _out_pmaCfgMerged_0_mask_5_match_mask_c_addr_T_1 = {addr_5,out_pmaCfgMerged_0_cfgVec_5_a[0]}; // @[Cat.scala 31:58]
  wire [34:0] out_pmaCfgMerged_0_mask_5_match_mask_c_addr = _out_pmaCfgMerged_0_mask_5_match_mask_c_addr_T_1 | 35'h3ff; // @[PMP.scala 86:50]
  wire [34:0] _out_pmaCfgMerged_0_mask_5_T_1 = out_pmaCfgMerged_0_mask_5_match_mask_c_addr + 35'h1; // @[PMP.scala 87:49]
  wire [34:0] _out_pmaCfgMerged_0_mask_5_T_2 = ~_out_pmaCfgMerged_0_mask_5_T_1; // @[PMP.scala 87:29]
  wire [34:0] _out_pmaCfgMerged_0_mask_5_T_3 = out_pmaCfgMerged_0_mask_5_match_mask_c_addr &
    _out_pmaCfgMerged_0_mask_5_T_2; // @[PMP.scala 87:27]
  wire [36:0] _out_pmaCfgMerged_0_mask_5_T_4 = {_out_pmaCfgMerged_0_mask_5_T_3,2'h3}; // @[Cat.scala 31:58]
  wire [36:0] _GEN_23 = out_pmaCfgMerged_0_cfgVec_5_a[1] ? _out_pmaCfgMerged_0_mask_5_T_4 : {{1'd0}, mask_5}; // @[PMA.scala 52:23 PMP.scala 98:36 99:27]
  wire  out_pmaCfgMerged_0_cfgVec_5_w = ~out_pmaCfgMerged_0_cfg_wm_tmp_5_l ? out_pmaCfgMerged_0_cfg_wm_tmp_5_w &
    out_pmaCfgMerged_0_cfg_wm_tmp_5_r : out_pmaCfgMerged_0_cfg_wm_tmp_5_w; // @[PMP.scala 94:17 95:29 96:21]
  wire [36:0] _GEN_26 = ~out_pmaCfgMerged_0_cfg_wm_tmp_5_l ? _GEN_23 : {{1'd0}, mask_5}; // @[PMA.scala 52:23 PMP.scala 95:29]
  wire  out_pmaCfgMerged_0_cfg_wm_tmp_6_r = _out_T_40[48]; // @[PMP.scala 93:61]
  wire  out_pmaCfgMerged_0_cfg_wm_tmp_6_w = _out_T_40[49]; // @[PMP.scala 93:61]
  wire  out_pmaCfgMerged_0_cfg_wm_tmp_6_x = _out_T_40[50]; // @[PMP.scala 93:61]
  wire [1:0] out_pmaCfgMerged_0_cfg_wm_tmp_6_a = _out_T_40[52:51]; // @[PMP.scala 93:61]
  wire  out_pmaCfgMerged_0_cfg_wm_tmp_6_atomic = _out_T_40[53]; // @[PMP.scala 93:61]
  wire  out_pmaCfgMerged_0_cfg_wm_tmp_6_c = _out_T_40[54]; // @[PMP.scala 93:61]
  wire  out_pmaCfgMerged_0_cfg_wm_tmp_6_l = _out_T_40[55]; // @[PMP.scala 93:61]
  wire  _out_pmaCfgMerged_0_cfgVec_6_a_T_1 = |out_pmaCfgMerged_0_cfg_wm_tmp_6_a; // @[PMP.scala 97:80]
  wire [1:0] _out_pmaCfgMerged_0_cfgVec_6_a_T_2 = {out_pmaCfgMerged_0_cfg_wm_tmp_6_a[1],
    _out_pmaCfgMerged_0_cfgVec_6_a_T_1}; // @[Cat.scala 31:58]
  wire [1:0] out_pmaCfgMerged_0_cfgVec_6_a = ~out_pmaCfgMerged_0_cfg_wm_tmp_6_l ? _out_pmaCfgMerged_0_cfgVec_6_a_T_2 :
    out_pmaCfgMerged_0_cfg_wm_tmp_6_a; // @[PMP.scala 94:17 95:29 97:41]
  wire [34:0] _out_pmaCfgMerged_0_mask_6_match_mask_c_addr_T_1 = {addr_6,out_pmaCfgMerged_0_cfgVec_6_a[0]}; // @[Cat.scala 31:58]
  wire [34:0] out_pmaCfgMerged_0_mask_6_match_mask_c_addr = _out_pmaCfgMerged_0_mask_6_match_mask_c_addr_T_1 | 35'h3ff; // @[PMP.scala 86:50]
  wire [34:0] _out_pmaCfgMerged_0_mask_6_T_1 = out_pmaCfgMerged_0_mask_6_match_mask_c_addr + 35'h1; // @[PMP.scala 87:49]
  wire [34:0] _out_pmaCfgMerged_0_mask_6_T_2 = ~_out_pmaCfgMerged_0_mask_6_T_1; // @[PMP.scala 87:29]
  wire [34:0] _out_pmaCfgMerged_0_mask_6_T_3 = out_pmaCfgMerged_0_mask_6_match_mask_c_addr &
    _out_pmaCfgMerged_0_mask_6_T_2; // @[PMP.scala 87:27]
  wire [36:0] _out_pmaCfgMerged_0_mask_6_T_4 = {_out_pmaCfgMerged_0_mask_6_T_3,2'h3}; // @[Cat.scala 31:58]
  wire [36:0] _GEN_27 = out_pmaCfgMerged_0_cfgVec_6_a[1] ? _out_pmaCfgMerged_0_mask_6_T_4 : {{1'd0}, mask_6}; // @[PMA.scala 52:23 PMP.scala 98:36 99:27]
  wire  out_pmaCfgMerged_0_cfgVec_6_w = ~out_pmaCfgMerged_0_cfg_wm_tmp_6_l ? out_pmaCfgMerged_0_cfg_wm_tmp_6_w &
    out_pmaCfgMerged_0_cfg_wm_tmp_6_r : out_pmaCfgMerged_0_cfg_wm_tmp_6_w; // @[PMP.scala 94:17 95:29 96:21]
  wire [36:0] _GEN_30 = ~out_pmaCfgMerged_0_cfg_wm_tmp_6_l ? _GEN_27 : {{1'd0}, mask_6}; // @[PMA.scala 52:23 PMP.scala 95:29]
  wire  out_pmaCfgMerged_0_cfg_wm_tmp_7_r = _out_T_40[56]; // @[PMP.scala 93:61]
  wire  out_pmaCfgMerged_0_cfg_wm_tmp_7_w = _out_T_40[57]; // @[PMP.scala 93:61]
  wire  out_pmaCfgMerged_0_cfg_wm_tmp_7_x = _out_T_40[58]; // @[PMP.scala 93:61]
  wire [1:0] out_pmaCfgMerged_0_cfg_wm_tmp_7_a = _out_T_40[60:59]; // @[PMP.scala 93:61]
  wire  out_pmaCfgMerged_0_cfg_wm_tmp_7_atomic = _out_T_40[61]; // @[PMP.scala 93:61]
  wire  out_pmaCfgMerged_0_cfg_wm_tmp_7_c = _out_T_40[62]; // @[PMP.scala 93:61]
  wire  out_pmaCfgMerged_0_cfg_wm_tmp_7_l = _out_T_40[63]; // @[PMP.scala 93:61]
  wire  _out_pmaCfgMerged_0_cfgVec_7_a_T_1 = |out_pmaCfgMerged_0_cfg_wm_tmp_7_a; // @[PMP.scala 97:80]
  wire [1:0] _out_pmaCfgMerged_0_cfgVec_7_a_T_2 = {out_pmaCfgMerged_0_cfg_wm_tmp_7_a[1],
    _out_pmaCfgMerged_0_cfgVec_7_a_T_1}; // @[Cat.scala 31:58]
  wire [1:0] out_pmaCfgMerged_0_cfgVec_7_a = ~out_pmaCfgMerged_0_cfg_wm_tmp_7_l ? _out_pmaCfgMerged_0_cfgVec_7_a_T_2 :
    out_pmaCfgMerged_0_cfg_wm_tmp_7_a; // @[PMP.scala 94:17 95:29 97:41]
  wire [34:0] _out_pmaCfgMerged_0_mask_7_match_mask_c_addr_T_1 = {addr_7,out_pmaCfgMerged_0_cfgVec_7_a[0]}; // @[Cat.scala 31:58]
  wire [34:0] out_pmaCfgMerged_0_mask_7_match_mask_c_addr = _out_pmaCfgMerged_0_mask_7_match_mask_c_addr_T_1 | 35'h3ff; // @[PMP.scala 86:50]
  wire [34:0] _out_pmaCfgMerged_0_mask_7_T_1 = out_pmaCfgMerged_0_mask_7_match_mask_c_addr + 35'h1; // @[PMP.scala 87:49]
  wire [34:0] _out_pmaCfgMerged_0_mask_7_T_2 = ~_out_pmaCfgMerged_0_mask_7_T_1; // @[PMP.scala 87:29]
  wire [34:0] _out_pmaCfgMerged_0_mask_7_T_3 = out_pmaCfgMerged_0_mask_7_match_mask_c_addr &
    _out_pmaCfgMerged_0_mask_7_T_2; // @[PMP.scala 87:27]
  wire [36:0] _out_pmaCfgMerged_0_mask_7_T_4 = {_out_pmaCfgMerged_0_mask_7_T_3,2'h3}; // @[Cat.scala 31:58]
  wire [36:0] _GEN_31 = out_pmaCfgMerged_0_cfgVec_7_a[1] ? _out_pmaCfgMerged_0_mask_7_T_4 : {{1'd0}, mask_7}; // @[PMA.scala 52:23 PMP.scala 98:36 99:27]
  wire  out_pmaCfgMerged_0_cfgVec_7_w = ~out_pmaCfgMerged_0_cfg_wm_tmp_7_l ? out_pmaCfgMerged_0_cfg_wm_tmp_7_w &
    out_pmaCfgMerged_0_cfg_wm_tmp_7_r : out_pmaCfgMerged_0_cfg_wm_tmp_7_w; // @[PMP.scala 94:17 95:29 96:21]
  wire [36:0] _GEN_34 = ~out_pmaCfgMerged_0_cfg_wm_tmp_7_l ? _GEN_31 : {{1'd0}, mask_7}; // @[PMA.scala 52:23 PMP.scala 95:29]
  wire [7:0] out_pmaCfgMerged_0_lo_lo_lo = {out_pmaCfgMerged_0_cfg_wm_tmp_l,out_pmaCfgMerged_0_cfg_wm_tmp_c,
    out_pmaCfgMerged_0_cfg_wm_tmp_atomic,out_pmaCfgMerged_0_cfgVec_0_a,out_pmaCfgMerged_0_cfg_wm_tmp_x,
    out_pmaCfgMerged_0_cfgVec_0_w,out_pmaCfgMerged_0_cfg_wm_tmp_r}; // @[PMP.scala 103:12]
  wire [15:0] out_pmaCfgMerged_0_lo_lo = {out_pmaCfgMerged_0_cfg_wm_tmp_1_l,out_pmaCfgMerged_0_cfg_wm_tmp_1_c,
    out_pmaCfgMerged_0_cfg_wm_tmp_1_atomic,out_pmaCfgMerged_0_cfgVec_1_a,out_pmaCfgMerged_0_cfg_wm_tmp_1_x,
    out_pmaCfgMerged_0_cfgVec_1_w,out_pmaCfgMerged_0_cfg_wm_tmp_1_r,out_pmaCfgMerged_0_lo_lo_lo}; // @[PMP.scala 103:12]
  wire [7:0] out_pmaCfgMerged_0_lo_hi_lo = {out_pmaCfgMerged_0_cfg_wm_tmp_2_l,out_pmaCfgMerged_0_cfg_wm_tmp_2_c,
    out_pmaCfgMerged_0_cfg_wm_tmp_2_atomic,out_pmaCfgMerged_0_cfgVec_2_a,out_pmaCfgMerged_0_cfg_wm_tmp_2_x,
    out_pmaCfgMerged_0_cfgVec_2_w,out_pmaCfgMerged_0_cfg_wm_tmp_2_r}; // @[PMP.scala 103:12]
  wire [31:0] out_pmaCfgMerged_0_lo = {out_pmaCfgMerged_0_cfg_wm_tmp_3_l,out_pmaCfgMerged_0_cfg_wm_tmp_3_c,
    out_pmaCfgMerged_0_cfg_wm_tmp_3_atomic,out_pmaCfgMerged_0_cfgVec_3_a,out_pmaCfgMerged_0_cfg_wm_tmp_3_x,
    out_pmaCfgMerged_0_cfgVec_3_w,out_pmaCfgMerged_0_cfg_wm_tmp_3_r,out_pmaCfgMerged_0_lo_hi_lo,
    out_pmaCfgMerged_0_lo_lo}; // @[PMP.scala 103:12]
  wire [7:0] out_pmaCfgMerged_0_hi_lo_lo = {out_pmaCfgMerged_0_cfg_wm_tmp_4_l,out_pmaCfgMerged_0_cfg_wm_tmp_4_c,
    out_pmaCfgMerged_0_cfg_wm_tmp_4_atomic,out_pmaCfgMerged_0_cfgVec_4_a,out_pmaCfgMerged_0_cfg_wm_tmp_4_x,
    out_pmaCfgMerged_0_cfgVec_4_w,out_pmaCfgMerged_0_cfg_wm_tmp_4_r}; // @[PMP.scala 103:12]
  wire [15:0] out_pmaCfgMerged_0_hi_lo = {out_pmaCfgMerged_0_cfg_wm_tmp_5_l,out_pmaCfgMerged_0_cfg_wm_tmp_5_c,
    out_pmaCfgMerged_0_cfg_wm_tmp_5_atomic,out_pmaCfgMerged_0_cfgVec_5_a,out_pmaCfgMerged_0_cfg_wm_tmp_5_x,
    out_pmaCfgMerged_0_cfgVec_5_w,out_pmaCfgMerged_0_cfg_wm_tmp_5_r,out_pmaCfgMerged_0_hi_lo_lo}; // @[PMP.scala 103:12]
  wire [7:0] out_pmaCfgMerged_0_hi_hi_lo = {out_pmaCfgMerged_0_cfg_wm_tmp_6_l,out_pmaCfgMerged_0_cfg_wm_tmp_6_c,
    out_pmaCfgMerged_0_cfg_wm_tmp_6_atomic,out_pmaCfgMerged_0_cfgVec_6_a,out_pmaCfgMerged_0_cfg_wm_tmp_6_x,
    out_pmaCfgMerged_0_cfgVec_6_w,out_pmaCfgMerged_0_cfg_wm_tmp_6_r}; // @[PMP.scala 103:12]
  wire [63:0] _out_pmaCfgMerged_0_T_16 = {out_pmaCfgMerged_0_cfg_wm_tmp_7_l,out_pmaCfgMerged_0_cfg_wm_tmp_7_c,
    out_pmaCfgMerged_0_cfg_wm_tmp_7_atomic,out_pmaCfgMerged_0_cfgVec_7_a,out_pmaCfgMerged_0_cfg_wm_tmp_7_x,
    out_pmaCfgMerged_0_cfgVec_7_w,out_pmaCfgMerged_0_cfg_wm_tmp_7_r,out_pmaCfgMerged_0_hi_hi_lo,
    out_pmaCfgMerged_0_hi_lo,out_pmaCfgMerged_0_lo}; // @[PMP.scala 103:12]
  wire [36:0] _GEN_35 = out_f_woready ? _GEN_6 : {{1'd0}, mask_0}; // @[PMA.scala 52:23 73:38]
  wire [36:0] _GEN_36 = out_f_woready ? _GEN_10 : {{1'd0}, mask_1}; // @[PMA.scala 52:23 73:38]
  wire [36:0] _GEN_37 = out_f_woready ? _GEN_14 : {{1'd0}, mask_2}; // @[PMA.scala 52:23 73:38]
  wire [36:0] _GEN_38 = out_f_woready ? _GEN_18 : {{1'd0}, mask_3}; // @[PMA.scala 52:23 73:38]
  wire [36:0] _GEN_39 = out_f_woready ? _GEN_22 : {{1'd0}, mask_4}; // @[PMA.scala 52:23 73:38]
  wire [36:0] _GEN_40 = out_f_woready ? _GEN_26 : {{1'd0}, mask_5}; // @[PMA.scala 52:23 73:38]
  wire [36:0] _GEN_41 = out_f_woready ? _GEN_30 : {{1'd0}, mask_6}; // @[PMA.scala 52:23 73:38]
  wire [36:0] _GEN_42 = out_f_woready ? _GEN_34 : {{1'd0}, mask_7}; // @[PMA.scala 52:23 73:38]
  wire  out_rifireMux_out = out_f_riready | ~out_rimask; // @[RegisterRouter.scala 82:24]
  wire  out_rofireMux_out = out_v_reg | ~out_romask; // @[RegisterRouter.scala 82:24]
  wire  out_backSel_26 = _out_backSel_T[26]; // @[RegisterRouter.scala 82:24]
  wire  out_woready_1 = out_back_io_deq_valid & auto_in_d_ready & ~out_back_io_deq_bits_read & out_backSel_26 &
    out_bindex == 9'h0; // @[RegisterRouter.scala 82:24]
  wire  out_f_woready_1 = out_woready_1 & out_womask; // @[RegisterRouter.scala 82:24]
  wire  _out_addr_10_locked_T = cfg_9_a == 2'h1; // @[PMP.scala 53:15]
  wire  out_addr_10_locked = cfg_10_l | cfg_9_l & _out_addr_10_locked_T; // @[PMP.scala 61:51]
  wire  _out_addr_10_mask_10_T = ~out_addr_10_locked; // @[PMP.scala 120:17]
  wire [34:0] _out_addr_10_mask_10_match_mask_c_addr_T_1 = {_out_T_40[33:0],cfg_10_a[0]}; // @[Cat.scala 31:58]
  wire [34:0] out_addr_10_mask_10_match_mask_c_addr = _out_addr_10_mask_10_match_mask_c_addr_T_1 | 35'h3ff; // @[PMP.scala 86:50]
  wire [34:0] _out_addr_10_mask_10_T_2 = out_addr_10_mask_10_match_mask_c_addr + 35'h1; // @[PMP.scala 87:49]
  wire [34:0] _out_addr_10_mask_10_T_3 = ~_out_addr_10_mask_10_T_2; // @[PMP.scala 87:29]
  wire [34:0] _out_addr_10_mask_10_T_4 = out_addr_10_mask_10_match_mask_c_addr & _out_addr_10_mask_10_T_3; // @[PMP.scala 87:27]
  wire [36:0] _out_addr_10_mask_10_T_5 = {_out_addr_10_mask_10_T_4,2'h3}; // @[Cat.scala 31:58]
  wire [36:0] _out_addr_10_mask_10_T_6 = ~out_addr_10_locked ? _out_addr_10_mask_10_T_5 : {{1'd0}, mask_10}; // @[PMP.scala 120:16]
  wire [36:0] _GEN_44 = out_f_woready_1 ? _out_addr_10_mask_10_T_6 : {{1'd0}, mask_10}; // @[PMA.scala 84:24 PMP.scala 120:10 PMA.scala 52:23]
  wire  out_backSel_21 = _out_backSel_T[21]; // @[RegisterRouter.scala 82:24]
  wire  out_woready_2 = out_back_io_deq_valid & auto_in_d_ready & ~out_back_io_deq_bits_read & out_backSel_21 &
    out_bindex == 9'h0; // @[RegisterRouter.scala 82:24]
  wire  out_f_woready_2 = out_woready_2 & out_womask; // @[RegisterRouter.scala 82:24]
  wire  _out_addr_5_locked_T = cfg_4_a == 2'h1; // @[PMP.scala 53:15]
  wire  out_addr_5_locked = cfg_5_l | cfg_4_l & _out_addr_5_locked_T; // @[PMP.scala 61:51]
  wire  _out_addr_5_mask_5_T = ~out_addr_5_locked; // @[PMP.scala 120:17]
  wire [34:0] _out_addr_5_mask_5_match_mask_c_addr_T_1 = {_out_T_40[33:0],cfg_5_a[0]}; // @[Cat.scala 31:58]
  wire [34:0] out_addr_5_mask_5_match_mask_c_addr = _out_addr_5_mask_5_match_mask_c_addr_T_1 | 35'h3ff; // @[PMP.scala 86:50]
  wire [34:0] _out_addr_5_mask_5_T_2 = out_addr_5_mask_5_match_mask_c_addr + 35'h1; // @[PMP.scala 87:49]
  wire [34:0] _out_addr_5_mask_5_T_3 = ~_out_addr_5_mask_5_T_2; // @[PMP.scala 87:29]
  wire [34:0] _out_addr_5_mask_5_T_4 = out_addr_5_mask_5_match_mask_c_addr & _out_addr_5_mask_5_T_3; // @[PMP.scala 87:27]
  wire [36:0] _out_addr_5_mask_5_T_5 = {_out_addr_5_mask_5_T_4,2'h3}; // @[Cat.scala 31:58]
  wire [36:0] _out_addr_5_mask_5_T_6 = ~out_addr_5_locked ? _out_addr_5_mask_5_T_5 : {{1'd0}, mask_5}; // @[PMP.scala 120:16]
  wire [36:0] _GEN_46 = out_f_woready_2 ? _out_addr_5_mask_5_T_6 : _GEN_40; // @[PMA.scala 84:24 PMP.scala 120:10]
  wire  out_backSel_30 = _out_backSel_T[30]; // @[RegisterRouter.scala 82:24]
  wire  out_woready_3 = out_back_io_deq_valid & auto_in_d_ready & ~out_back_io_deq_bits_read & out_backSel_30 &
    out_bindex == 9'h0; // @[RegisterRouter.scala 82:24]
  wire  out_f_woready_3 = out_woready_3 & out_womask; // @[RegisterRouter.scala 82:24]
  wire  _out_addr_14_locked_T = cfg_13_a == 2'h1; // @[PMP.scala 53:15]
  wire  out_addr_14_locked = cfg_14_l | cfg_13_l & _out_addr_14_locked_T; // @[PMP.scala 61:51]
  wire  _out_addr_14_mask_14_T = ~out_addr_14_locked; // @[PMP.scala 120:17]
  wire [34:0] _out_addr_14_mask_14_match_mask_c_addr_T_1 = {_out_T_40[33:0],cfg_14_a[0]}; // @[Cat.scala 31:58]
  wire [34:0] out_addr_14_mask_14_match_mask_c_addr = _out_addr_14_mask_14_match_mask_c_addr_T_1 | 35'h3ff; // @[PMP.scala 86:50]
  wire [34:0] _out_addr_14_mask_14_T_2 = out_addr_14_mask_14_match_mask_c_addr + 35'h1; // @[PMP.scala 87:49]
  wire [34:0] _out_addr_14_mask_14_T_3 = ~_out_addr_14_mask_14_T_2; // @[PMP.scala 87:29]
  wire [34:0] _out_addr_14_mask_14_T_4 = out_addr_14_mask_14_match_mask_c_addr & _out_addr_14_mask_14_T_3; // @[PMP.scala 87:27]
  wire [36:0] _out_addr_14_mask_14_T_5 = {_out_addr_14_mask_14_T_4,2'h3}; // @[Cat.scala 31:58]
  wire [36:0] _out_addr_14_mask_14_T_6 = ~out_addr_14_locked ? _out_addr_14_mask_14_T_5 : {{1'd0}, mask_14}; // @[PMP.scala 120:16]
  wire [36:0] _GEN_48 = out_f_woready_3 ? _out_addr_14_mask_14_T_6 : {{1'd0}, mask_14}; // @[PMA.scala 84:24 PMP.scala 120:10 PMA.scala 52:23]
  wire  out_frontSel_1 = _out_frontSel_T[1]; // @[RegisterRouter.scala 82:24]
  wire  out_rivalid_4 = auto_in_a_valid & out_front_ready & in_bits_read & out_frontSel_1 & out_findex == 9'h0; // @[RegisterRouter.scala 82:24]
  wire  out_f_rivalid_4 = out_rivalid_4 & out_rimask; // @[RegisterRouter.scala 82:24]
  wire  out_backSel_1 = _out_backSel_T[1]; // @[RegisterRouter.scala 82:24]
  wire  out_roready_4 = out_back_io_deq_valid & auto_in_d_ready & out_back_io_deq_bits_read & out_backSel_1 & out_bindex
     == 9'h0; // @[RegisterRouter.scala 82:24]
  wire  out_f_roready_4 = out_roready_4 & out_romask; // @[RegisterRouter.scala 82:24]
  reg  out_v_reg_1; // @[Hold.scala 40:24]
  wire  out_f_riready_1 = ~out_v_reg_1; // @[PMA.scala 67:20]
  wire  _out_v_reg_T_2 = out_f_riready_1 & out_f_rivalid_4; // @[PMA.scala 66:39]
  wire  _out_v_reg_T_3 = out_v_reg_1 & out_f_roready_4; // @[PMA.scala 66:58]
  wire  _GEN_50 = _out_v_reg_T_3 ? 1'h0 : out_v_reg_1; // @[Hold.scala 41:20 40:24 41:28]
  wire  out_rifireMux_out_1 = out_f_riready_1 | ~out_rimask; // @[RegisterRouter.scala 82:24]
  wire  out_rofireMux_out_1 = out_v_reg_1 | ~out_romask; // @[RegisterRouter.scala 82:24]
  wire  out_backSel_22 = _out_backSel_T[22]; // @[RegisterRouter.scala 82:24]
  wire  out_woready_5 = out_back_io_deq_valid & auto_in_d_ready & ~out_back_io_deq_bits_read & out_backSel_22 &
    out_bindex == 9'h0; // @[RegisterRouter.scala 82:24]
  wire  out_f_woready_5 = out_woready_5 & out_womask; // @[RegisterRouter.scala 82:24]
  wire  _out_addr_6_locked_T = cfg_5_a == 2'h1; // @[PMP.scala 53:15]
  wire  out_addr_6_locked = cfg_6_l | cfg_5_l & _out_addr_6_locked_T; // @[PMP.scala 61:51]
  wire  _out_addr_6_mask_6_T = ~out_addr_6_locked; // @[PMP.scala 120:17]
  wire [34:0] _out_addr_6_mask_6_match_mask_c_addr_T_1 = {_out_T_40[33:0],cfg_6_a[0]}; // @[Cat.scala 31:58]
  wire [34:0] out_addr_6_mask_6_match_mask_c_addr = _out_addr_6_mask_6_match_mask_c_addr_T_1 | 35'h3ff; // @[PMP.scala 86:50]
  wire [34:0] _out_addr_6_mask_6_T_2 = out_addr_6_mask_6_match_mask_c_addr + 35'h1; // @[PMP.scala 87:49]
  wire [34:0] _out_addr_6_mask_6_T_3 = ~_out_addr_6_mask_6_T_2; // @[PMP.scala 87:29]
  wire [34:0] _out_addr_6_mask_6_T_4 = out_addr_6_mask_6_match_mask_c_addr & _out_addr_6_mask_6_T_3; // @[PMP.scala 87:27]
  wire [36:0] _out_addr_6_mask_6_T_5 = {_out_addr_6_mask_6_T_4,2'h3}; // @[Cat.scala 31:58]
  wire [36:0] _out_addr_6_mask_6_T_6 = ~out_addr_6_locked ? _out_addr_6_mask_6_T_5 : {{1'd0}, mask_6}; // @[PMP.scala 120:16]
  wire [36:0] _GEN_53 = out_f_woready_5 ? _out_addr_6_mask_6_T_6 : _GEN_41; // @[PMA.scala 84:24 PMP.scala 120:10]
  wire  out_backSel_17 = _out_backSel_T[17]; // @[RegisterRouter.scala 82:24]
  wire  out_woready_6 = out_back_io_deq_valid & auto_in_d_ready & ~out_back_io_deq_bits_read & out_backSel_17 &
    out_bindex == 9'h0; // @[RegisterRouter.scala 82:24]
  wire  out_f_woready_6 = out_woready_6 & out_womask; // @[RegisterRouter.scala 82:24]
  wire  _out_addr_1_locked_T = cfg_0_a == 2'h1; // @[PMP.scala 53:15]
  wire  out_addr_1_locked = cfg_1_l | cfg_0_l & _out_addr_1_locked_T; // @[PMP.scala 61:51]
  wire  _out_addr_1_mask_1_T = ~out_addr_1_locked; // @[PMP.scala 120:17]
  wire [34:0] _out_addr_1_mask_1_match_mask_c_addr_T_1 = {_out_T_40[33:0],cfg_1_a[0]}; // @[Cat.scala 31:58]
  wire [34:0] out_addr_1_mask_1_match_mask_c_addr = _out_addr_1_mask_1_match_mask_c_addr_T_1 | 35'h3ff; // @[PMP.scala 86:50]
  wire [34:0] _out_addr_1_mask_1_T_2 = out_addr_1_mask_1_match_mask_c_addr + 35'h1; // @[PMP.scala 87:49]
  wire [34:0] _out_addr_1_mask_1_T_3 = ~_out_addr_1_mask_1_T_2; // @[PMP.scala 87:29]
  wire [34:0] _out_addr_1_mask_1_T_4 = out_addr_1_mask_1_match_mask_c_addr & _out_addr_1_mask_1_T_3; // @[PMP.scala 87:27]
  wire [36:0] _out_addr_1_mask_1_T_5 = {_out_addr_1_mask_1_T_4,2'h3}; // @[Cat.scala 31:58]
  wire [36:0] _out_addr_1_mask_1_T_6 = ~out_addr_1_locked ? _out_addr_1_mask_1_T_5 : {{1'd0}, mask_1}; // @[PMP.scala 120:16]
  wire [36:0] _GEN_55 = out_f_woready_6 ? _out_addr_1_mask_1_T_6 : _GEN_36; // @[PMA.scala 84:24 PMP.scala 120:10]
  wire  out_backSel_25 = _out_backSel_T[25]; // @[RegisterRouter.scala 82:24]
  wire  out_woready_7 = out_back_io_deq_valid & auto_in_d_ready & ~out_back_io_deq_bits_read & out_backSel_25 &
    out_bindex == 9'h0; // @[RegisterRouter.scala 82:24]
  wire  out_f_woready_7 = out_woready_7 & out_womask; // @[RegisterRouter.scala 82:24]
  wire  _out_addr_9_locked_T = cfg_8_a == 2'h1; // @[PMP.scala 53:15]
  wire  out_addr_9_locked = cfg_9_l | cfg_8_l & _out_addr_9_locked_T; // @[PMP.scala 61:51]
  wire  _out_addr_9_mask_9_T = ~out_addr_9_locked; // @[PMP.scala 120:17]
  wire [34:0] _out_addr_9_mask_9_match_mask_c_addr_T_1 = {_out_T_40[33:0],cfg_9_a[0]}; // @[Cat.scala 31:58]
  wire [34:0] out_addr_9_mask_9_match_mask_c_addr = _out_addr_9_mask_9_match_mask_c_addr_T_1 | 35'h3ff; // @[PMP.scala 86:50]
  wire [34:0] _out_addr_9_mask_9_T_2 = out_addr_9_mask_9_match_mask_c_addr + 35'h1; // @[PMP.scala 87:49]
  wire [34:0] _out_addr_9_mask_9_T_3 = ~_out_addr_9_mask_9_T_2; // @[PMP.scala 87:29]
  wire [34:0] _out_addr_9_mask_9_T_4 = out_addr_9_mask_9_match_mask_c_addr & _out_addr_9_mask_9_T_3; // @[PMP.scala 87:27]
  wire [36:0] _out_addr_9_mask_9_T_5 = {_out_addr_9_mask_9_T_4,2'h3}; // @[Cat.scala 31:58]
  wire [36:0] _out_addr_9_mask_9_T_6 = ~out_addr_9_locked ? _out_addr_9_mask_9_T_5 : {{1'd0}, mask_9}; // @[PMP.scala 120:16]
  wire [36:0] _GEN_57 = out_f_woready_7 ? _out_addr_9_mask_9_T_6 : {{1'd0}, mask_9}; // @[PMA.scala 84:24 PMP.scala 120:10 PMA.scala 52:23]
  wire  out_frontSel_2 = _out_frontSel_T[2]; // @[RegisterRouter.scala 82:24]
  wire  out_rivalid_8 = auto_in_a_valid & out_front_ready & in_bits_read & out_frontSel_2 & out_findex == 9'h0; // @[RegisterRouter.scala 82:24]
  wire  out_f_rivalid_8 = out_rivalid_8 & out_rimask; // @[RegisterRouter.scala 82:24]
  wire  out_backSel_2 = _out_backSel_T[2]; // @[RegisterRouter.scala 82:24]
  wire  out_roready_8 = out_back_io_deq_valid & auto_in_d_ready & out_back_io_deq_bits_read & out_backSel_2 & out_bindex
     == 9'h0; // @[RegisterRouter.scala 82:24]
  wire  out_f_roready_8 = out_roready_8 & out_romask; // @[RegisterRouter.scala 82:24]
  wire  out_woready_8 = out_back_io_deq_valid & auto_in_d_ready & ~out_back_io_deq_bits_read & out_backSel_2 &
    out_bindex == 9'h0; // @[RegisterRouter.scala 82:24]
  wire  out_f_woready_8 = out_woready_8 & out_womask; // @[RegisterRouter.scala 82:24]
  reg  out_v_reg_2; // @[Hold.scala 40:24]
  wire  out_f_riready_2 = ~out_v_reg_2; // @[PMA.scala 67:20]
  wire  _out_v_reg_T_4 = out_f_riready_2 & out_f_rivalid_8; // @[PMA.scala 66:39]
  wire  _out_v_reg_T_5 = out_v_reg_2 & out_f_roready_8; // @[PMA.scala 66:58]
  wire  _GEN_59 = _out_v_reg_T_5 ? 1'h0 : out_v_reg_2; // @[Hold.scala 41:20 40:24 41:28]
  wire [34:0] _out_pmaCfgMerged_1_mask_8_match_mask_c_addr_T_1 = {addr_8,out_pmaCfgMerged_0_cfgVec_0_a[0]}; // @[Cat.scala 31:58]
  wire [34:0] out_pmaCfgMerged_1_mask_8_match_mask_c_addr = _out_pmaCfgMerged_1_mask_8_match_mask_c_addr_T_1 | 35'h3ff; // @[PMP.scala 86:50]
  wire [34:0] _out_pmaCfgMerged_1_mask_8_T_1 = out_pmaCfgMerged_1_mask_8_match_mask_c_addr + 35'h1; // @[PMP.scala 87:49]
  wire [34:0] _out_pmaCfgMerged_1_mask_8_T_2 = ~_out_pmaCfgMerged_1_mask_8_T_1; // @[PMP.scala 87:29]
  wire [34:0] _out_pmaCfgMerged_1_mask_8_T_3 = out_pmaCfgMerged_1_mask_8_match_mask_c_addr &
    _out_pmaCfgMerged_1_mask_8_T_2; // @[PMP.scala 87:27]
  wire [36:0] _out_pmaCfgMerged_1_mask_8_T_4 = {_out_pmaCfgMerged_1_mask_8_T_3,2'h3}; // @[Cat.scala 31:58]
  wire [36:0] _GEN_62 = out_pmaCfgMerged_0_cfgVec_0_a[1] ? _out_pmaCfgMerged_1_mask_8_T_4 : {{1'd0}, mask_8}; // @[PMA.scala 52:23 PMP.scala 98:36 99:27]
  wire [36:0] _GEN_65 = ~out_pmaCfgMerged_0_cfg_wm_tmp_l ? _GEN_62 : {{1'd0}, mask_8}; // @[PMA.scala 52:23 PMP.scala 95:29]
  wire [34:0] _out_pmaCfgMerged_1_mask_9_match_mask_c_addr_T_1 = {addr_9,out_pmaCfgMerged_0_cfgVec_1_a[0]}; // @[Cat.scala 31:58]
  wire [34:0] out_pmaCfgMerged_1_mask_9_match_mask_c_addr = _out_pmaCfgMerged_1_mask_9_match_mask_c_addr_T_1 | 35'h3ff; // @[PMP.scala 86:50]
  wire [34:0] _out_pmaCfgMerged_1_mask_9_T_1 = out_pmaCfgMerged_1_mask_9_match_mask_c_addr + 35'h1; // @[PMP.scala 87:49]
  wire [34:0] _out_pmaCfgMerged_1_mask_9_T_2 = ~_out_pmaCfgMerged_1_mask_9_T_1; // @[PMP.scala 87:29]
  wire [34:0] _out_pmaCfgMerged_1_mask_9_T_3 = out_pmaCfgMerged_1_mask_9_match_mask_c_addr &
    _out_pmaCfgMerged_1_mask_9_T_2; // @[PMP.scala 87:27]
  wire [36:0] _out_pmaCfgMerged_1_mask_9_T_4 = {_out_pmaCfgMerged_1_mask_9_T_3,2'h3}; // @[Cat.scala 31:58]
  wire [36:0] _GEN_66 = out_pmaCfgMerged_0_cfgVec_1_a[1] ? _out_pmaCfgMerged_1_mask_9_T_4 : _GEN_57; // @[PMP.scala 98:36 99:27]
  wire [36:0] _GEN_69 = ~out_pmaCfgMerged_0_cfg_wm_tmp_1_l ? _GEN_66 : _GEN_57; // @[PMP.scala 95:29]
  wire [34:0] _out_pmaCfgMerged_1_mask_10_match_mask_c_addr_T_1 = {addr_10,out_pmaCfgMerged_0_cfgVec_2_a[0]}; // @[Cat.scala 31:58]
  wire [34:0] out_pmaCfgMerged_1_mask_10_match_mask_c_addr = _out_pmaCfgMerged_1_mask_10_match_mask_c_addr_T_1 | 35'h3ff
    ; // @[PMP.scala 86:50]
  wire [34:0] _out_pmaCfgMerged_1_mask_10_T_1 = out_pmaCfgMerged_1_mask_10_match_mask_c_addr + 35'h1; // @[PMP.scala 87:49]
  wire [34:0] _out_pmaCfgMerged_1_mask_10_T_2 = ~_out_pmaCfgMerged_1_mask_10_T_1; // @[PMP.scala 87:29]
  wire [34:0] _out_pmaCfgMerged_1_mask_10_T_3 = out_pmaCfgMerged_1_mask_10_match_mask_c_addr &
    _out_pmaCfgMerged_1_mask_10_T_2; // @[PMP.scala 87:27]
  wire [36:0] _out_pmaCfgMerged_1_mask_10_T_4 = {_out_pmaCfgMerged_1_mask_10_T_3,2'h3}; // @[Cat.scala 31:58]
  wire [36:0] _GEN_70 = out_pmaCfgMerged_0_cfgVec_2_a[1] ? _out_pmaCfgMerged_1_mask_10_T_4 : _GEN_44; // @[PMP.scala 98:36 99:27]
  wire [36:0] _GEN_73 = ~out_pmaCfgMerged_0_cfg_wm_tmp_2_l ? _GEN_70 : _GEN_44; // @[PMP.scala 95:29]
  wire [34:0] _out_pmaCfgMerged_1_mask_11_match_mask_c_addr_T_1 = {addr_11,out_pmaCfgMerged_0_cfgVec_3_a[0]}; // @[Cat.scala 31:58]
  wire [34:0] out_pmaCfgMerged_1_mask_11_match_mask_c_addr = _out_pmaCfgMerged_1_mask_11_match_mask_c_addr_T_1 | 35'h3ff
    ; // @[PMP.scala 86:50]
  wire [34:0] _out_pmaCfgMerged_1_mask_11_T_1 = out_pmaCfgMerged_1_mask_11_match_mask_c_addr + 35'h1; // @[PMP.scala 87:49]
  wire [34:0] _out_pmaCfgMerged_1_mask_11_T_2 = ~_out_pmaCfgMerged_1_mask_11_T_1; // @[PMP.scala 87:29]
  wire [34:0] _out_pmaCfgMerged_1_mask_11_T_3 = out_pmaCfgMerged_1_mask_11_match_mask_c_addr &
    _out_pmaCfgMerged_1_mask_11_T_2; // @[PMP.scala 87:27]
  wire [36:0] _out_pmaCfgMerged_1_mask_11_T_4 = {_out_pmaCfgMerged_1_mask_11_T_3,2'h3}; // @[Cat.scala 31:58]
  wire [36:0] _GEN_74 = out_pmaCfgMerged_0_cfgVec_3_a[1] ? _out_pmaCfgMerged_1_mask_11_T_4 : {{1'd0}, mask_11}; // @[PMA.scala 52:23 PMP.scala 98:36 99:27]
  wire [36:0] _GEN_77 = ~out_pmaCfgMerged_0_cfg_wm_tmp_3_l ? _GEN_74 : {{1'd0}, mask_11}; // @[PMA.scala 52:23 PMP.scala 95:29]
  wire [34:0] _out_pmaCfgMerged_1_mask_12_match_mask_c_addr_T_1 = {addr_12,out_pmaCfgMerged_0_cfgVec_4_a[0]}; // @[Cat.scala 31:58]
  wire [34:0] out_pmaCfgMerged_1_mask_12_match_mask_c_addr = _out_pmaCfgMerged_1_mask_12_match_mask_c_addr_T_1 | 35'h3ff
    ; // @[PMP.scala 86:50]
  wire [34:0] _out_pmaCfgMerged_1_mask_12_T_1 = out_pmaCfgMerged_1_mask_12_match_mask_c_addr + 35'h1; // @[PMP.scala 87:49]
  wire [34:0] _out_pmaCfgMerged_1_mask_12_T_2 = ~_out_pmaCfgMerged_1_mask_12_T_1; // @[PMP.scala 87:29]
  wire [34:0] _out_pmaCfgMerged_1_mask_12_T_3 = out_pmaCfgMerged_1_mask_12_match_mask_c_addr &
    _out_pmaCfgMerged_1_mask_12_T_2; // @[PMP.scala 87:27]
  wire [36:0] _out_pmaCfgMerged_1_mask_12_T_4 = {_out_pmaCfgMerged_1_mask_12_T_3,2'h3}; // @[Cat.scala 31:58]
  wire [36:0] _GEN_78 = out_pmaCfgMerged_0_cfgVec_4_a[1] ? _out_pmaCfgMerged_1_mask_12_T_4 : {{1'd0}, mask_12}; // @[PMA.scala 52:23 PMP.scala 98:36 99:27]
  wire [36:0] _GEN_81 = ~out_pmaCfgMerged_0_cfg_wm_tmp_4_l ? _GEN_78 : {{1'd0}, mask_12}; // @[PMA.scala 52:23 PMP.scala 95:29]
  wire [34:0] _out_pmaCfgMerged_1_mask_13_match_mask_c_addr_T_1 = {addr_13,out_pmaCfgMerged_0_cfgVec_5_a[0]}; // @[Cat.scala 31:58]
  wire [34:0] out_pmaCfgMerged_1_mask_13_match_mask_c_addr = _out_pmaCfgMerged_1_mask_13_match_mask_c_addr_T_1 | 35'h3ff
    ; // @[PMP.scala 86:50]
  wire [34:0] _out_pmaCfgMerged_1_mask_13_T_1 = out_pmaCfgMerged_1_mask_13_match_mask_c_addr + 35'h1; // @[PMP.scala 87:49]
  wire [34:0] _out_pmaCfgMerged_1_mask_13_T_2 = ~_out_pmaCfgMerged_1_mask_13_T_1; // @[PMP.scala 87:29]
  wire [34:0] _out_pmaCfgMerged_1_mask_13_T_3 = out_pmaCfgMerged_1_mask_13_match_mask_c_addr &
    _out_pmaCfgMerged_1_mask_13_T_2; // @[PMP.scala 87:27]
  wire [36:0] _out_pmaCfgMerged_1_mask_13_T_4 = {_out_pmaCfgMerged_1_mask_13_T_3,2'h3}; // @[Cat.scala 31:58]
  wire [36:0] _GEN_82 = out_pmaCfgMerged_0_cfgVec_5_a[1] ? _out_pmaCfgMerged_1_mask_13_T_4 : {{1'd0}, mask_13}; // @[PMA.scala 52:23 PMP.scala 98:36 99:27]
  wire [36:0] _GEN_85 = ~out_pmaCfgMerged_0_cfg_wm_tmp_5_l ? _GEN_82 : {{1'd0}, mask_13}; // @[PMA.scala 52:23 PMP.scala 95:29]
  wire [34:0] _out_pmaCfgMerged_1_mask_14_match_mask_c_addr_T_1 = {addr_14,out_pmaCfgMerged_0_cfgVec_6_a[0]}; // @[Cat.scala 31:58]
  wire [34:0] out_pmaCfgMerged_1_mask_14_match_mask_c_addr = _out_pmaCfgMerged_1_mask_14_match_mask_c_addr_T_1 | 35'h3ff
    ; // @[PMP.scala 86:50]
  wire [34:0] _out_pmaCfgMerged_1_mask_14_T_1 = out_pmaCfgMerged_1_mask_14_match_mask_c_addr + 35'h1; // @[PMP.scala 87:49]
  wire [34:0] _out_pmaCfgMerged_1_mask_14_T_2 = ~_out_pmaCfgMerged_1_mask_14_T_1; // @[PMP.scala 87:29]
  wire [34:0] _out_pmaCfgMerged_1_mask_14_T_3 = out_pmaCfgMerged_1_mask_14_match_mask_c_addr &
    _out_pmaCfgMerged_1_mask_14_T_2; // @[PMP.scala 87:27]
  wire [36:0] _out_pmaCfgMerged_1_mask_14_T_4 = {_out_pmaCfgMerged_1_mask_14_T_3,2'h3}; // @[Cat.scala 31:58]
  wire [36:0] _GEN_86 = out_pmaCfgMerged_0_cfgVec_6_a[1] ? _out_pmaCfgMerged_1_mask_14_T_4 : _GEN_48; // @[PMP.scala 98:36 99:27]
  wire [36:0] _GEN_89 = ~out_pmaCfgMerged_0_cfg_wm_tmp_6_l ? _GEN_86 : _GEN_48; // @[PMP.scala 95:29]
  wire [34:0] _out_pmaCfgMerged_1_mask_15_match_mask_c_addr_T_1 = {addr_15,out_pmaCfgMerged_0_cfgVec_7_a[0]}; // @[Cat.scala 31:58]
  wire [34:0] out_pmaCfgMerged_1_mask_15_match_mask_c_addr = _out_pmaCfgMerged_1_mask_15_match_mask_c_addr_T_1 | 35'h3ff
    ; // @[PMP.scala 86:50]
  wire [34:0] _out_pmaCfgMerged_1_mask_15_T_1 = out_pmaCfgMerged_1_mask_15_match_mask_c_addr + 35'h1; // @[PMP.scala 87:49]
  wire [34:0] _out_pmaCfgMerged_1_mask_15_T_2 = ~_out_pmaCfgMerged_1_mask_15_T_1; // @[PMP.scala 87:29]
  wire [34:0] _out_pmaCfgMerged_1_mask_15_T_3 = out_pmaCfgMerged_1_mask_15_match_mask_c_addr &
    _out_pmaCfgMerged_1_mask_15_T_2; // @[PMP.scala 87:27]
  wire [36:0] _out_pmaCfgMerged_1_mask_15_T_4 = {_out_pmaCfgMerged_1_mask_15_T_3,2'h3}; // @[Cat.scala 31:58]
  wire [36:0] _GEN_90 = out_pmaCfgMerged_0_cfgVec_7_a[1] ? _out_pmaCfgMerged_1_mask_15_T_4 : {{1'd0}, mask_15}; // @[PMA.scala 52:23 PMP.scala 98:36 99:27]
  wire [36:0] _GEN_93 = ~out_pmaCfgMerged_0_cfg_wm_tmp_7_l ? _GEN_90 : {{1'd0}, mask_15}; // @[PMA.scala 52:23 PMP.scala 95:29]
  wire [36:0] _GEN_94 = out_f_woready_8 ? _GEN_65 : {{1'd0}, mask_8}; // @[PMA.scala 52:23 73:38]
  wire [36:0] _GEN_95 = out_f_woready_8 ? _GEN_69 : _GEN_57; // @[PMA.scala 73:38]
  wire [36:0] _GEN_96 = out_f_woready_8 ? _GEN_73 : _GEN_44; // @[PMA.scala 73:38]
  wire [36:0] _GEN_97 = out_f_woready_8 ? _GEN_77 : {{1'd0}, mask_11}; // @[PMA.scala 52:23 73:38]
  wire [36:0] _GEN_98 = out_f_woready_8 ? _GEN_81 : {{1'd0}, mask_12}; // @[PMA.scala 52:23 73:38]
  wire [36:0] _GEN_99 = out_f_woready_8 ? _GEN_85 : {{1'd0}, mask_13}; // @[PMA.scala 52:23 73:38]
  wire [36:0] _GEN_100 = out_f_woready_8 ? _GEN_89 : _GEN_48; // @[PMA.scala 73:38]
  wire [36:0] _GEN_101 = out_f_woready_8 ? _GEN_93 : {{1'd0}, mask_15}; // @[PMA.scala 52:23 73:38]
  wire  out_rifireMux_out_2 = out_f_riready_2 | ~out_rimask; // @[RegisterRouter.scala 82:24]
  wire  out_rofireMux_out_2 = out_v_reg_2 | ~out_romask; // @[RegisterRouter.scala 82:24]
  wire  out_backSel_16 = _out_backSel_T[16]; // @[RegisterRouter.scala 82:24]
  wire  out_woready_9 = out_back_io_deq_valid & auto_in_d_ready & ~out_back_io_deq_bits_read & out_backSel_16 &
    out_bindex == 9'h0; // @[RegisterRouter.scala 82:24]
  wire  out_f_woready_9 = out_woready_9 & out_womask; // @[RegisterRouter.scala 82:24]
  wire  _out_addr_0_mask_0_T = ~cfg_0_l; // @[PMP.scala 120:17]
  wire [34:0] _out_addr_0_mask_0_match_mask_c_addr_T_1 = {_out_T_40[33:0],cfg_0_a[0]}; // @[Cat.scala 31:58]
  wire [34:0] out_addr_0_mask_0_match_mask_c_addr = _out_addr_0_mask_0_match_mask_c_addr_T_1 | 35'h3ff; // @[PMP.scala 86:50]
  wire [34:0] _out_addr_0_mask_0_T_2 = out_addr_0_mask_0_match_mask_c_addr + 35'h1; // @[PMP.scala 87:49]
  wire [34:0] _out_addr_0_mask_0_T_3 = ~_out_addr_0_mask_0_T_2; // @[PMP.scala 87:29]
  wire [34:0] _out_addr_0_mask_0_T_4 = out_addr_0_mask_0_match_mask_c_addr & _out_addr_0_mask_0_T_3; // @[PMP.scala 87:27]
  wire [36:0] _out_addr_0_mask_0_T_5 = {_out_addr_0_mask_0_T_4,2'h3}; // @[Cat.scala 31:58]
  wire [36:0] _out_addr_0_mask_0_T_6 = ~cfg_0_l ? _out_addr_0_mask_0_T_5 : {{1'd0}, mask_0}; // @[PMP.scala 120:16]
  wire [36:0] _GEN_103 = out_f_woready_9 ? _out_addr_0_mask_0_T_6 : _GEN_35; // @[PMA.scala 84:24 PMP.scala 120:10]
  wire  out_backSel_18 = _out_backSel_T[18]; // @[RegisterRouter.scala 82:24]
  wire  out_woready_10 = out_back_io_deq_valid & auto_in_d_ready & ~out_back_io_deq_bits_read & out_backSel_18 &
    out_bindex == 9'h0; // @[RegisterRouter.scala 82:24]
  wire  out_f_woready_10 = out_woready_10 & out_womask; // @[RegisterRouter.scala 82:24]
  wire  _out_addr_2_locked_T = cfg_1_a == 2'h1; // @[PMP.scala 53:15]
  wire  out_addr_2_locked = cfg_2_l | cfg_1_l & _out_addr_2_locked_T; // @[PMP.scala 61:51]
  wire  _out_addr_2_mask_2_T = ~out_addr_2_locked; // @[PMP.scala 120:17]
  wire [34:0] _out_addr_2_mask_2_match_mask_c_addr_T_1 = {_out_T_40[33:0],cfg_2_a[0]}; // @[Cat.scala 31:58]
  wire [34:0] out_addr_2_mask_2_match_mask_c_addr = _out_addr_2_mask_2_match_mask_c_addr_T_1 | 35'h3ff; // @[PMP.scala 86:50]
  wire [34:0] _out_addr_2_mask_2_T_2 = out_addr_2_mask_2_match_mask_c_addr + 35'h1; // @[PMP.scala 87:49]
  wire [34:0] _out_addr_2_mask_2_T_3 = ~_out_addr_2_mask_2_T_2; // @[PMP.scala 87:29]
  wire [34:0] _out_addr_2_mask_2_T_4 = out_addr_2_mask_2_match_mask_c_addr & _out_addr_2_mask_2_T_3; // @[PMP.scala 87:27]
  wire [36:0] _out_addr_2_mask_2_T_5 = {_out_addr_2_mask_2_T_4,2'h3}; // @[Cat.scala 31:58]
  wire [36:0] _out_addr_2_mask_2_T_6 = ~out_addr_2_locked ? _out_addr_2_mask_2_T_5 : {{1'd0}, mask_2}; // @[PMP.scala 120:16]
  wire [36:0] _GEN_105 = out_f_woready_10 ? _out_addr_2_mask_2_T_6 : _GEN_37; // @[PMA.scala 84:24 PMP.scala 120:10]
  wire  out_backSel_29 = _out_backSel_T[29]; // @[RegisterRouter.scala 82:24]
  wire  out_woready_11 = out_back_io_deq_valid & auto_in_d_ready & ~out_back_io_deq_bits_read & out_backSel_29 &
    out_bindex == 9'h0; // @[RegisterRouter.scala 82:24]
  wire  out_f_woready_11 = out_woready_11 & out_womask; // @[RegisterRouter.scala 82:24]
  wire  _out_addr_13_locked_T = cfg_12_a == 2'h1; // @[PMP.scala 53:15]
  wire  out_addr_13_locked = cfg_13_l | cfg_12_l & _out_addr_13_locked_T; // @[PMP.scala 61:51]
  wire  _out_addr_13_mask_13_T = ~out_addr_13_locked; // @[PMP.scala 120:17]
  wire [34:0] _out_addr_13_mask_13_match_mask_c_addr_T_1 = {_out_T_40[33:0],cfg_13_a[0]}; // @[Cat.scala 31:58]
  wire [34:0] out_addr_13_mask_13_match_mask_c_addr = _out_addr_13_mask_13_match_mask_c_addr_T_1 | 35'h3ff; // @[PMP.scala 86:50]
  wire [34:0] _out_addr_13_mask_13_T_2 = out_addr_13_mask_13_match_mask_c_addr + 35'h1; // @[PMP.scala 87:49]
  wire [34:0] _out_addr_13_mask_13_T_3 = ~_out_addr_13_mask_13_T_2; // @[PMP.scala 87:29]
  wire [34:0] _out_addr_13_mask_13_T_4 = out_addr_13_mask_13_match_mask_c_addr & _out_addr_13_mask_13_T_3; // @[PMP.scala 87:27]
  wire [36:0] _out_addr_13_mask_13_T_5 = {_out_addr_13_mask_13_T_4,2'h3}; // @[Cat.scala 31:58]
  wire [36:0] _out_addr_13_mask_13_T_6 = ~out_addr_13_locked ? _out_addr_13_mask_13_T_5 : {{1'd0}, mask_13}; // @[PMP.scala 120:16]
  wire [36:0] _GEN_107 = out_f_woready_11 ? _out_addr_13_mask_13_T_6 : _GEN_99; // @[PMA.scala 84:24 PMP.scala 120:10]
  wire  out_backSel_28 = _out_backSel_T[28]; // @[RegisterRouter.scala 82:24]
  wire  out_woready_12 = out_back_io_deq_valid & auto_in_d_ready & ~out_back_io_deq_bits_read & out_backSel_28 &
    out_bindex == 9'h0; // @[RegisterRouter.scala 82:24]
  wire  out_f_woready_12 = out_woready_12 & out_womask; // @[RegisterRouter.scala 82:24]
  wire  _out_addr_12_locked_T = cfg_11_a == 2'h1; // @[PMP.scala 53:15]
  wire  out_addr_12_locked = cfg_12_l | cfg_11_l & _out_addr_12_locked_T; // @[PMP.scala 61:51]
  wire  _out_addr_12_mask_12_T = ~out_addr_12_locked; // @[PMP.scala 120:17]
  wire [34:0] _out_addr_12_mask_12_match_mask_c_addr_T_1 = {_out_T_40[33:0],cfg_12_a[0]}; // @[Cat.scala 31:58]
  wire [34:0] out_addr_12_mask_12_match_mask_c_addr = _out_addr_12_mask_12_match_mask_c_addr_T_1 | 35'h3ff; // @[PMP.scala 86:50]
  wire [34:0] _out_addr_12_mask_12_T_2 = out_addr_12_mask_12_match_mask_c_addr + 35'h1; // @[PMP.scala 87:49]
  wire [34:0] _out_addr_12_mask_12_T_3 = ~_out_addr_12_mask_12_T_2; // @[PMP.scala 87:29]
  wire [34:0] _out_addr_12_mask_12_T_4 = out_addr_12_mask_12_match_mask_c_addr & _out_addr_12_mask_12_T_3; // @[PMP.scala 87:27]
  wire [36:0] _out_addr_12_mask_12_T_5 = {_out_addr_12_mask_12_T_4,2'h3}; // @[Cat.scala 31:58]
  wire [36:0] _out_addr_12_mask_12_T_6 = ~out_addr_12_locked ? _out_addr_12_mask_12_T_5 : {{1'd0}, mask_12}; // @[PMP.scala 120:16]
  wire [36:0] _GEN_109 = out_f_woready_12 ? _out_addr_12_mask_12_T_6 : _GEN_98; // @[PMA.scala 84:24 PMP.scala 120:10]
  wire  out_backSel_23 = _out_backSel_T[23]; // @[RegisterRouter.scala 82:24]
  wire  out_woready_13 = out_back_io_deq_valid & auto_in_d_ready & ~out_back_io_deq_bits_read & out_backSel_23 &
    out_bindex == 9'h0; // @[RegisterRouter.scala 82:24]
  wire  out_f_woready_13 = out_woready_13 & out_womask; // @[RegisterRouter.scala 82:24]
  wire  _out_addr_7_locked_T = cfg_6_a == 2'h1; // @[PMP.scala 53:15]
  wire  out_addr_7_locked = cfg_7_l | cfg_6_l & _out_addr_7_locked_T; // @[PMP.scala 61:51]
  wire  _out_addr_7_mask_7_T = ~out_addr_7_locked; // @[PMP.scala 120:17]
  wire [34:0] _out_addr_7_mask_7_match_mask_c_addr_T_1 = {_out_T_40[33:0],cfg_7_a[0]}; // @[Cat.scala 31:58]
  wire [34:0] out_addr_7_mask_7_match_mask_c_addr = _out_addr_7_mask_7_match_mask_c_addr_T_1 | 35'h3ff; // @[PMP.scala 86:50]
  wire [34:0] _out_addr_7_mask_7_T_2 = out_addr_7_mask_7_match_mask_c_addr + 35'h1; // @[PMP.scala 87:49]
  wire [34:0] _out_addr_7_mask_7_T_3 = ~_out_addr_7_mask_7_T_2; // @[PMP.scala 87:29]
  wire [34:0] _out_addr_7_mask_7_T_4 = out_addr_7_mask_7_match_mask_c_addr & _out_addr_7_mask_7_T_3; // @[PMP.scala 87:27]
  wire [36:0] _out_addr_7_mask_7_T_5 = {_out_addr_7_mask_7_T_4,2'h3}; // @[Cat.scala 31:58]
  wire [36:0] _out_addr_7_mask_7_T_6 = ~out_addr_7_locked ? _out_addr_7_mask_7_T_5 : {{1'd0}, mask_7}; // @[PMP.scala 120:16]
  wire [36:0] _GEN_111 = out_f_woready_13 ? _out_addr_7_mask_7_T_6 : _GEN_42; // @[PMA.scala 84:24 PMP.scala 120:10]
  wire  out_frontSel_3 = _out_frontSel_T[3]; // @[RegisterRouter.scala 82:24]
  wire  out_rivalid_14 = auto_in_a_valid & out_front_ready & in_bits_read & out_frontSel_3 & out_findex == 9'h0; // @[RegisterRouter.scala 82:24]
  wire  out_f_rivalid_14 = out_rivalid_14 & out_rimask; // @[RegisterRouter.scala 82:24]
  wire  out_backSel_3 = _out_backSel_T[3]; // @[RegisterRouter.scala 82:24]
  wire  out_roready_14 = out_back_io_deq_valid & auto_in_d_ready & out_back_io_deq_bits_read & out_backSel_3 &
    out_bindex == 9'h0; // @[RegisterRouter.scala 82:24]
  wire  out_f_roready_14 = out_roready_14 & out_romask; // @[RegisterRouter.scala 82:24]
  reg  out_v_reg_3; // @[Hold.scala 40:24]
  wire  out_f_riready_3 = ~out_v_reg_3; // @[PMA.scala 67:20]
  wire  _out_v_reg_T_6 = out_f_riready_3 & out_f_rivalid_14; // @[PMA.scala 66:39]
  wire  _out_v_reg_T_7 = out_v_reg_3 & out_f_roready_14; // @[PMA.scala 66:58]
  wire  _GEN_113 = _out_v_reg_T_7 ? 1'h0 : out_v_reg_3; // @[Hold.scala 41:20 40:24 41:28]
  wire  out_rifireMux_out_3 = out_f_riready_3 | ~out_rimask; // @[RegisterRouter.scala 82:24]
  wire  out_rofireMux_out_3 = out_v_reg_3 | ~out_romask; // @[RegisterRouter.scala 82:24]
  wire  out_backSel_19 = _out_backSel_T[19]; // @[RegisterRouter.scala 82:24]
  wire  out_woready_15 = out_back_io_deq_valid & auto_in_d_ready & ~out_back_io_deq_bits_read & out_backSel_19 &
    out_bindex == 9'h0; // @[RegisterRouter.scala 82:24]
  wire  out_f_woready_15 = out_woready_15 & out_womask; // @[RegisterRouter.scala 82:24]
  wire  _out_addr_3_locked_T = cfg_2_a == 2'h1; // @[PMP.scala 53:15]
  wire  out_addr_3_locked = cfg_3_l | cfg_2_l & _out_addr_3_locked_T; // @[PMP.scala 61:51]
  wire  _out_addr_3_mask_3_T = ~out_addr_3_locked; // @[PMP.scala 120:17]
  wire [34:0] _out_addr_3_mask_3_match_mask_c_addr_T_1 = {_out_T_40[33:0],cfg_3_a[0]}; // @[Cat.scala 31:58]
  wire [34:0] out_addr_3_mask_3_match_mask_c_addr = _out_addr_3_mask_3_match_mask_c_addr_T_1 | 35'h3ff; // @[PMP.scala 86:50]
  wire [34:0] _out_addr_3_mask_3_T_2 = out_addr_3_mask_3_match_mask_c_addr + 35'h1; // @[PMP.scala 87:49]
  wire [34:0] _out_addr_3_mask_3_T_3 = ~_out_addr_3_mask_3_T_2; // @[PMP.scala 87:29]
  wire [34:0] _out_addr_3_mask_3_T_4 = out_addr_3_mask_3_match_mask_c_addr & _out_addr_3_mask_3_T_3; // @[PMP.scala 87:27]
  wire [36:0] _out_addr_3_mask_3_T_5 = {_out_addr_3_mask_3_T_4,2'h3}; // @[Cat.scala 31:58]
  wire [36:0] _out_addr_3_mask_3_T_6 = ~out_addr_3_locked ? _out_addr_3_mask_3_T_5 : {{1'd0}, mask_3}; // @[PMP.scala 120:16]
  wire [36:0] _GEN_116 = out_f_woready_15 ? _out_addr_3_mask_3_T_6 : _GEN_38; // @[PMA.scala 84:24 PMP.scala 120:10]
  wire  out_backSel_27 = _out_backSel_T[27]; // @[RegisterRouter.scala 82:24]
  wire  out_woready_16 = out_back_io_deq_valid & auto_in_d_ready & ~out_back_io_deq_bits_read & out_backSel_27 &
    out_bindex == 9'h0; // @[RegisterRouter.scala 82:24]
  wire  out_f_woready_16 = out_woready_16 & out_womask; // @[RegisterRouter.scala 82:24]
  wire  _out_addr_11_locked_T = cfg_10_a == 2'h1; // @[PMP.scala 53:15]
  wire  out_addr_11_locked = cfg_11_l | cfg_10_l & _out_addr_11_locked_T; // @[PMP.scala 61:51]
  wire  _out_addr_11_mask_11_T = ~out_addr_11_locked; // @[PMP.scala 120:17]
  wire [34:0] _out_addr_11_mask_11_match_mask_c_addr_T_1 = {_out_T_40[33:0],cfg_11_a[0]}; // @[Cat.scala 31:58]
  wire [34:0] out_addr_11_mask_11_match_mask_c_addr = _out_addr_11_mask_11_match_mask_c_addr_T_1 | 35'h3ff; // @[PMP.scala 86:50]
  wire [34:0] _out_addr_11_mask_11_T_2 = out_addr_11_mask_11_match_mask_c_addr + 35'h1; // @[PMP.scala 87:49]
  wire [34:0] _out_addr_11_mask_11_T_3 = ~_out_addr_11_mask_11_T_2; // @[PMP.scala 87:29]
  wire [34:0] _out_addr_11_mask_11_T_4 = out_addr_11_mask_11_match_mask_c_addr & _out_addr_11_mask_11_T_3; // @[PMP.scala 87:27]
  wire [36:0] _out_addr_11_mask_11_T_5 = {_out_addr_11_mask_11_T_4,2'h3}; // @[Cat.scala 31:58]
  wire [36:0] _out_addr_11_mask_11_T_6 = ~out_addr_11_locked ? _out_addr_11_mask_11_T_5 : {{1'd0}, mask_11}; // @[PMP.scala 120:16]
  wire [36:0] _GEN_118 = out_f_woready_16 ? _out_addr_11_mask_11_T_6 : _GEN_97; // @[PMA.scala 84:24 PMP.scala 120:10]
  wire  out_backSel_24 = _out_backSel_T[24]; // @[RegisterRouter.scala 82:24]
  wire  out_woready_17 = out_back_io_deq_valid & auto_in_d_ready & ~out_back_io_deq_bits_read & out_backSel_24 &
    out_bindex == 9'h0; // @[RegisterRouter.scala 82:24]
  wire  out_f_woready_17 = out_woready_17 & out_womask; // @[RegisterRouter.scala 82:24]
  wire  _out_addr_8_locked_T = cfg_7_a == 2'h1; // @[PMP.scala 53:15]
  wire  out_addr_8_locked = cfg_8_l | cfg_7_l & _out_addr_8_locked_T; // @[PMP.scala 61:51]
  wire  _out_addr_8_mask_8_T = ~out_addr_8_locked; // @[PMP.scala 120:17]
  wire [34:0] _out_addr_8_mask_8_match_mask_c_addr_T_1 = {_out_T_40[33:0],cfg_8_a[0]}; // @[Cat.scala 31:58]
  wire [34:0] out_addr_8_mask_8_match_mask_c_addr = _out_addr_8_mask_8_match_mask_c_addr_T_1 | 35'h3ff; // @[PMP.scala 86:50]
  wire [34:0] _out_addr_8_mask_8_T_2 = out_addr_8_mask_8_match_mask_c_addr + 35'h1; // @[PMP.scala 87:49]
  wire [34:0] _out_addr_8_mask_8_T_3 = ~_out_addr_8_mask_8_T_2; // @[PMP.scala 87:29]
  wire [34:0] _out_addr_8_mask_8_T_4 = out_addr_8_mask_8_match_mask_c_addr & _out_addr_8_mask_8_T_3; // @[PMP.scala 87:27]
  wire [36:0] _out_addr_8_mask_8_T_5 = {_out_addr_8_mask_8_T_4,2'h3}; // @[Cat.scala 31:58]
  wire [36:0] _out_addr_8_mask_8_T_6 = ~out_addr_8_locked ? _out_addr_8_mask_8_T_5 : {{1'd0}, mask_8}; // @[PMP.scala 120:16]
  wire [36:0] _GEN_120 = out_f_woready_17 ? _out_addr_8_mask_8_T_6 : _GEN_94; // @[PMA.scala 84:24 PMP.scala 120:10]
  wire  out_backSel_20 = _out_backSel_T[20]; // @[RegisterRouter.scala 82:24]
  wire  out_woready_18 = out_back_io_deq_valid & auto_in_d_ready & ~out_back_io_deq_bits_read & out_backSel_20 &
    out_bindex == 9'h0; // @[RegisterRouter.scala 82:24]
  wire  out_f_woready_18 = out_woready_18 & out_womask; // @[RegisterRouter.scala 82:24]
  wire  _out_addr_4_locked_T = cfg_3_a == 2'h1; // @[PMP.scala 53:15]
  wire  out_addr_4_locked = cfg_4_l | cfg_3_l & _out_addr_4_locked_T; // @[PMP.scala 61:51]
  wire  _out_addr_4_mask_4_T = ~out_addr_4_locked; // @[PMP.scala 120:17]
  wire [34:0] _out_addr_4_mask_4_match_mask_c_addr_T_1 = {_out_T_40[33:0],cfg_4_a[0]}; // @[Cat.scala 31:58]
  wire [34:0] out_addr_4_mask_4_match_mask_c_addr = _out_addr_4_mask_4_match_mask_c_addr_T_1 | 35'h3ff; // @[PMP.scala 86:50]
  wire [34:0] _out_addr_4_mask_4_T_2 = out_addr_4_mask_4_match_mask_c_addr + 35'h1; // @[PMP.scala 87:49]
  wire [34:0] _out_addr_4_mask_4_T_3 = ~_out_addr_4_mask_4_T_2; // @[PMP.scala 87:29]
  wire [34:0] _out_addr_4_mask_4_T_4 = out_addr_4_mask_4_match_mask_c_addr & _out_addr_4_mask_4_T_3; // @[PMP.scala 87:27]
  wire [36:0] _out_addr_4_mask_4_T_5 = {_out_addr_4_mask_4_T_4,2'h3}; // @[Cat.scala 31:58]
  wire [36:0] _out_addr_4_mask_4_T_6 = ~out_addr_4_locked ? _out_addr_4_mask_4_T_5 : {{1'd0}, mask_4}; // @[PMP.scala 120:16]
  wire [36:0] _GEN_122 = out_f_woready_18 ? _out_addr_4_mask_4_T_6 : _GEN_39; // @[PMA.scala 84:24 PMP.scala 120:10]
  wire  out_backSel_31 = _out_backSel_T[31]; // @[RegisterRouter.scala 82:24]
  wire  out_woready_19 = out_back_io_deq_valid & auto_in_d_ready & ~out_back_io_deq_bits_read & out_backSel_31 &
    out_bindex == 9'h0; // @[RegisterRouter.scala 82:24]
  wire  out_f_woready_19 = out_woready_19 & out_womask; // @[RegisterRouter.scala 82:24]
  wire  _out_addr_15_locked_T = cfg_14_a == 2'h1; // @[PMP.scala 53:15]
  wire  out_addr_15_locked = cfg_15_l | cfg_14_l & _out_addr_15_locked_T; // @[PMP.scala 61:51]
  wire  _out_addr_15_mask_15_T = ~out_addr_15_locked; // @[PMP.scala 120:17]
  wire [34:0] _out_addr_15_mask_15_match_mask_c_addr_T_1 = {_out_T_40[33:0],cfg_15_a[0]}; // @[Cat.scala 31:58]
  wire [34:0] out_addr_15_mask_15_match_mask_c_addr = _out_addr_15_mask_15_match_mask_c_addr_T_1 | 35'h3ff; // @[PMP.scala 86:50]
  wire [34:0] _out_addr_15_mask_15_T_2 = out_addr_15_mask_15_match_mask_c_addr + 35'h1; // @[PMP.scala 87:49]
  wire [34:0] _out_addr_15_mask_15_T_3 = ~_out_addr_15_mask_15_T_2; // @[PMP.scala 87:29]
  wire [34:0] _out_addr_15_mask_15_T_4 = out_addr_15_mask_15_match_mask_c_addr & _out_addr_15_mask_15_T_3; // @[PMP.scala 87:27]
  wire [36:0] _out_addr_15_mask_15_T_5 = {_out_addr_15_mask_15_T_4,2'h3}; // @[Cat.scala 31:58]
  wire [36:0] _out_addr_15_mask_15_T_6 = ~out_addr_15_locked ? _out_addr_15_mask_15_T_5 : {{1'd0}, mask_15}; // @[PMP.scala 120:16]
  wire [36:0] _GEN_124 = out_f_woready_19 ? _out_addr_15_mask_15_T_6 : _GEN_101; // @[PMA.scala 84:24 PMP.scala 120:10]
  wire  _out_rifireMux_T_5 = out_rifireMux_out | ~(out_findex == 9'h0); // @[RegisterRouter.scala 82:24]
  wire  _out_rifireMux_T_9 = out_rifireMux_out_1 | ~(out_findex == 9'h0); // @[RegisterRouter.scala 82:24]
  wire  _out_rifireMux_T_13 = out_rifireMux_out_2 | ~(out_findex == 9'h0); // @[RegisterRouter.scala 82:24]
  wire  _out_rifireMux_T_17 = out_rifireMux_out_3 | ~(out_findex == 9'h0); // @[RegisterRouter.scala 82:24]
  wire  _GEN_127 = 5'h1 == out_iindex ? _out_rifireMux_T_9 : _out_rifireMux_T_5; // @[MuxLiteral.scala 48:{10,10}]
  wire  _GEN_128 = 5'h2 == out_iindex ? _out_rifireMux_T_13 : _GEN_127; // @[MuxLiteral.scala 48:{10,10}]
  wire  _GEN_129 = 5'h3 == out_iindex ? _out_rifireMux_T_17 : _GEN_128; // @[MuxLiteral.scala 48:{10,10}]
  wire  _GEN_144 = 5'h12 == out_iindex | (5'h11 == out_iindex | (5'h10 == out_iindex | (5'hf == out_iindex | (5'he ==
    out_iindex | (5'hd == out_iindex | (5'hc == out_iindex | (5'hb == out_iindex | (5'ha == out_iindex | (5'h9 ==
    out_iindex | (5'h8 == out_iindex | (5'h7 == out_iindex | (5'h6 == out_iindex | (5'h5 == out_iindex | (5'h4 ==
    out_iindex | _GEN_129)))))))))))))); // @[MuxLiteral.scala 48:{10,10}]
  wire  out_rifireMux = 5'h1f == out_iindex | (5'h1e == out_iindex | (5'h1d == out_iindex | (5'h1c == out_iindex | (5'h1b
     == out_iindex | (5'h1a == out_iindex | (5'h19 == out_iindex | (5'h18 == out_iindex | (5'h17 == out_iindex | (5'h16
     == out_iindex | (5'h15 == out_iindex | (5'h14 == out_iindex | (5'h13 == out_iindex | _GEN_144)))))))))))); // @[MuxLiteral.scala 48:{10,10}]
  wire  _out_rofireMux_T_5 = out_rofireMux_out | ~(out_bindex == 9'h0); // @[RegisterRouter.scala 82:24]
  wire  _out_rofireMux_T_9 = out_rofireMux_out_1 | ~(out_bindex == 9'h0); // @[RegisterRouter.scala 82:24]
  wire  _out_rofireMux_T_13 = out_rofireMux_out_2 | ~(out_bindex == 9'h0); // @[RegisterRouter.scala 82:24]
  wire  _out_rofireMux_T_17 = out_rofireMux_out_3 | ~(out_bindex == 9'h0); // @[RegisterRouter.scala 82:24]
  wire  _GEN_191 = 5'h1 == out_oindex ? _out_rofireMux_T_9 : _out_rofireMux_T_5; // @[MuxLiteral.scala 48:{10,10}]
  wire  _GEN_192 = 5'h2 == out_oindex ? _out_rofireMux_T_13 : _GEN_191; // @[MuxLiteral.scala 48:{10,10}]
  wire  _GEN_193 = 5'h3 == out_oindex ? _out_rofireMux_T_17 : _GEN_192; // @[MuxLiteral.scala 48:{10,10}]
  wire  _GEN_208 = 5'h12 == out_oindex | (5'h11 == out_oindex | (5'h10 == out_oindex | (5'hf == out_oindex | (5'he ==
    out_oindex | (5'hd == out_oindex | (5'hc == out_oindex | (5'hb == out_oindex | (5'ha == out_oindex | (5'h9 ==
    out_oindex | (5'h8 == out_oindex | (5'h7 == out_oindex | (5'h6 == out_oindex | (5'h5 == out_oindex | (5'h4 ==
    out_oindex | _GEN_193)))))))))))))); // @[MuxLiteral.scala 48:{10,10}]
  wire  out_rofireMux = 5'h1f == out_oindex | (5'h1e == out_oindex | (5'h1d == out_oindex | (5'h1c == out_oindex | (5'h1b
     == out_oindex | (5'h1a == out_oindex | (5'h19 == out_oindex | (5'h18 == out_oindex | (5'h17 == out_oindex | (5'h16
     == out_oindex | (5'h15 == out_oindex | (5'h14 == out_oindex | (5'h13 == out_oindex | _GEN_208)))))))))))); // @[MuxLiteral.scala 48:{10,10}]
  wire  out_iready = in_bits_read ? out_rifireMux : 1'h1; // @[RegisterRouter.scala 82:24]
  wire  out_oready = out_back_io_deq_bits_read ? out_rofireMux : 1'h1; // @[RegisterRouter.scala 82:24]
  wire  _GEN_255 = 5'h1 == out_oindex ? _out_T_1 : _out_T_1; // @[MuxLiteral.scala 48:{10,10}]
  wire  _GEN_256 = 5'h2 == out_oindex ? _out_T_1 : _GEN_255; // @[MuxLiteral.scala 48:{10,10}]
  wire  _GEN_257 = 5'h3 == out_oindex ? _out_T_1 : _GEN_256; // @[MuxLiteral.scala 48:{10,10}]
  wire  _GEN_270 = 5'h10 == out_oindex ? _out_T_1 : 5'hf == out_oindex | (5'he == out_oindex | (5'hd == out_oindex | (5'hc
     == out_oindex | (5'hb == out_oindex | (5'ha == out_oindex | (5'h9 == out_oindex | (5'h8 == out_oindex | (5'h7 ==
    out_oindex | (5'h6 == out_oindex | (5'h5 == out_oindex | (5'h4 == out_oindex | _GEN_257))))))))))); // @[MuxLiteral.scala 48:{10,10}]
  wire  _GEN_271 = 5'h11 == out_oindex ? _out_T_1 : _GEN_270; // @[MuxLiteral.scala 48:{10,10}]
  wire  _GEN_272 = 5'h12 == out_oindex ? _out_T_1 : _GEN_271; // @[MuxLiteral.scala 48:{10,10}]
  wire  _GEN_273 = 5'h13 == out_oindex ? _out_T_1 : _GEN_272; // @[MuxLiteral.scala 48:{10,10}]
  wire  _GEN_274 = 5'h14 == out_oindex ? _out_T_1 : _GEN_273; // @[MuxLiteral.scala 48:{10,10}]
  wire  _GEN_275 = 5'h15 == out_oindex ? _out_T_1 : _GEN_274; // @[MuxLiteral.scala 48:{10,10}]
  wire  _GEN_276 = 5'h16 == out_oindex ? _out_T_1 : _GEN_275; // @[MuxLiteral.scala 48:{10,10}]
  wire  _GEN_277 = 5'h17 == out_oindex ? _out_T_1 : _GEN_276; // @[MuxLiteral.scala 48:{10,10}]
  wire  _GEN_278 = 5'h18 == out_oindex ? _out_T_1 : _GEN_277; // @[MuxLiteral.scala 48:{10,10}]
  wire  _GEN_279 = 5'h19 == out_oindex ? _out_T_1 : _GEN_278; // @[MuxLiteral.scala 48:{10,10}]
  wire  _GEN_280 = 5'h1a == out_oindex ? _out_T_1 : _GEN_279; // @[MuxLiteral.scala 48:{10,10}]
  wire  _GEN_281 = 5'h1b == out_oindex ? _out_T_1 : _GEN_280; // @[MuxLiteral.scala 48:{10,10}]
  wire  _GEN_282 = 5'h1c == out_oindex ? _out_T_1 : _GEN_281; // @[MuxLiteral.scala 48:{10,10}]
  wire  _GEN_283 = 5'h1d == out_oindex ? _out_T_1 : _GEN_282; // @[MuxLiteral.scala 48:{10,10}]
  wire  _GEN_284 = 5'h1e == out_oindex ? _out_T_1 : _GEN_283; // @[MuxLiteral.scala 48:{10,10}]
  wire  _GEN_285 = 5'h1f == out_oindex ? _out_T_1 : _GEN_284; // @[MuxLiteral.scala 48:{10,10}]
  wire [63:0] _GEN_287 = 5'h1 == out_oindex ? 64'h0 : pmaCfgMerged_0; // @[MuxLiteral.scala 48:{10,10}]
  wire [63:0] _GEN_288 = 5'h2 == out_oindex ? pmaCfgMerged_1 : _GEN_287; // @[MuxLiteral.scala 48:{10,10}]
  wire [63:0] _GEN_289 = 5'h3 == out_oindex ? 64'h0 : _GEN_288; // @[MuxLiteral.scala 48:{10,10}]
  wire [63:0] _GEN_290 = 5'h4 == out_oindex ? 64'h0 : _GEN_289; // @[MuxLiteral.scala 48:{10,10}]
  wire [63:0] _GEN_291 = 5'h5 == out_oindex ? 64'h0 : _GEN_290; // @[MuxLiteral.scala 48:{10,10}]
  wire [63:0] _GEN_292 = 5'h6 == out_oindex ? 64'h0 : _GEN_291; // @[MuxLiteral.scala 48:{10,10}]
  wire [63:0] _GEN_293 = 5'h7 == out_oindex ? 64'h0 : _GEN_292; // @[MuxLiteral.scala 48:{10,10}]
  wire [63:0] _GEN_294 = 5'h8 == out_oindex ? 64'h0 : _GEN_293; // @[MuxLiteral.scala 48:{10,10}]
  wire [63:0] _GEN_295 = 5'h9 == out_oindex ? 64'h0 : _GEN_294; // @[MuxLiteral.scala 48:{10,10}]
  wire [63:0] _GEN_296 = 5'ha == out_oindex ? 64'h0 : _GEN_295; // @[MuxLiteral.scala 48:{10,10}]
  wire [63:0] _GEN_297 = 5'hb == out_oindex ? 64'h0 : _GEN_296; // @[MuxLiteral.scala 48:{10,10}]
  wire [63:0] _GEN_298 = 5'hc == out_oindex ? 64'h0 : _GEN_297; // @[MuxLiteral.scala 48:{10,10}]
  wire [63:0] _GEN_299 = 5'hd == out_oindex ? 64'h0 : _GEN_298; // @[MuxLiteral.scala 48:{10,10}]
  wire [63:0] _GEN_300 = 5'he == out_oindex ? 64'h0 : _GEN_299; // @[MuxLiteral.scala 48:{10,10}]
  wire [63:0] _GEN_301 = 5'hf == out_oindex ? 64'h0 : _GEN_300; // @[MuxLiteral.scala 48:{10,10}]
  wire [63:0] _GEN_302 = 5'h10 == out_oindex ? _T_5 : _GEN_301; // @[MuxLiteral.scala 48:{10,10}]
  wire [63:0] _GEN_303 = 5'h11 == out_oindex ? _T_11 : _GEN_302; // @[MuxLiteral.scala 48:{10,10}]
  wire [63:0] _GEN_304 = 5'h12 == out_oindex ? _T_17 : _GEN_303; // @[MuxLiteral.scala 48:{10,10}]
  wire [63:0] _GEN_305 = 5'h13 == out_oindex ? _T_23 : _GEN_304; // @[MuxLiteral.scala 48:{10,10}]
  wire [63:0] _GEN_306 = 5'h14 == out_oindex ? _T_29 : _GEN_305; // @[MuxLiteral.scala 48:{10,10}]
  wire [63:0] _GEN_307 = 5'h15 == out_oindex ? _T_35 : _GEN_306; // @[MuxLiteral.scala 48:{10,10}]
  wire [63:0] _GEN_308 = 5'h16 == out_oindex ? _T_41 : _GEN_307; // @[MuxLiteral.scala 48:{10,10}]
  wire [63:0] _GEN_309 = 5'h17 == out_oindex ? _T_47 : _GEN_308; // @[MuxLiteral.scala 48:{10,10}]
  wire [63:0] _GEN_310 = 5'h18 == out_oindex ? _T_53 : _GEN_309; // @[MuxLiteral.scala 48:{10,10}]
  wire [63:0] _GEN_311 = 5'h19 == out_oindex ? _T_59 : _GEN_310; // @[MuxLiteral.scala 48:{10,10}]
  wire [63:0] _GEN_312 = 5'h1a == out_oindex ? _T_65 : _GEN_311; // @[MuxLiteral.scala 48:{10,10}]
  wire [63:0] _GEN_313 = 5'h1b == out_oindex ? _T_71 : _GEN_312; // @[MuxLiteral.scala 48:{10,10}]
  wire [63:0] _GEN_314 = 5'h1c == out_oindex ? _T_77 : _GEN_313; // @[MuxLiteral.scala 48:{10,10}]
  wire [63:0] _GEN_315 = 5'h1d == out_oindex ? _T_83 : _GEN_314; // @[MuxLiteral.scala 48:{10,10}]
  wire [63:0] _GEN_316 = 5'h1e == out_oindex ? _T_89 : _GEN_315; // @[MuxLiteral.scala 48:{10,10}]
  wire [63:0] _GEN_317 = 5'h1f == out_oindex ? _T_95 : _GEN_316; // @[MuxLiteral.scala 48:{10,10}]
  wire  out_bits_read = out_back_io_deq_bits_read; // @[RegisterRouter.scala 82:{24,24}]
  Queue_132 out_back ( // @[Decoupled.scala 361:21]
    .clock(out_back_clock),
    .reset(out_back_reset),
    .io_enq_ready(out_back_io_enq_ready),
    .io_enq_valid(out_back_io_enq_valid),
    .io_enq_bits_read(out_back_io_enq_bits_read),
    .io_enq_bits_index(out_back_io_enq_bits_index),
    .io_enq_bits_data(out_back_io_enq_bits_data),
    .io_enq_bits_mask(out_back_io_enq_bits_mask),
    .io_enq_bits_extra_tlrr_extra_source(out_back_io_enq_bits_extra_tlrr_extra_source),
    .io_enq_bits_extra_tlrr_extra_size(out_back_io_enq_bits_extra_tlrr_extra_size),
    .io_deq_ready(out_back_io_deq_ready),
    .io_deq_valid(out_back_io_deq_valid),
    .io_deq_bits_read(out_back_io_deq_bits_read),
    .io_deq_bits_index(out_back_io_deq_bits_index),
    .io_deq_bits_data(out_back_io_deq_bits_data),
    .io_deq_bits_mask(out_back_io_deq_bits_mask),
    .io_deq_bits_extra_tlrr_extra_source(out_back_io_deq_bits_extra_tlrr_extra_source),
    .io_deq_bits_extra_tlrr_extra_size(out_back_io_deq_bits_extra_tlrr_extra_size)
  );
  PMPChecker PMPChecker ( // @[TLPMA.scala 47:13]
    .io_check_env_mode(PMPChecker_io_check_env_mode),
    .io_check_env_pmp_0_cfg_l(PMPChecker_io_check_env_pmp_0_cfg_l),
    .io_check_env_pmp_0_cfg_a(PMPChecker_io_check_env_pmp_0_cfg_a),
    .io_check_env_pmp_0_cfg_x(PMPChecker_io_check_env_pmp_0_cfg_x),
    .io_check_env_pmp_0_cfg_w(PMPChecker_io_check_env_pmp_0_cfg_w),
    .io_check_env_pmp_0_cfg_r(PMPChecker_io_check_env_pmp_0_cfg_r),
    .io_check_env_pmp_0_addr(PMPChecker_io_check_env_pmp_0_addr),
    .io_check_env_pmp_0_mask(PMPChecker_io_check_env_pmp_0_mask),
    .io_check_env_pmp_1_cfg_l(PMPChecker_io_check_env_pmp_1_cfg_l),
    .io_check_env_pmp_1_cfg_a(PMPChecker_io_check_env_pmp_1_cfg_a),
    .io_check_env_pmp_1_cfg_x(PMPChecker_io_check_env_pmp_1_cfg_x),
    .io_check_env_pmp_1_cfg_w(PMPChecker_io_check_env_pmp_1_cfg_w),
    .io_check_env_pmp_1_cfg_r(PMPChecker_io_check_env_pmp_1_cfg_r),
    .io_check_env_pmp_1_addr(PMPChecker_io_check_env_pmp_1_addr),
    .io_check_env_pmp_1_mask(PMPChecker_io_check_env_pmp_1_mask),
    .io_check_env_pmp_2_cfg_l(PMPChecker_io_check_env_pmp_2_cfg_l),
    .io_check_env_pmp_2_cfg_a(PMPChecker_io_check_env_pmp_2_cfg_a),
    .io_check_env_pmp_2_cfg_x(PMPChecker_io_check_env_pmp_2_cfg_x),
    .io_check_env_pmp_2_cfg_w(PMPChecker_io_check_env_pmp_2_cfg_w),
    .io_check_env_pmp_2_cfg_r(PMPChecker_io_check_env_pmp_2_cfg_r),
    .io_check_env_pmp_2_addr(PMPChecker_io_check_env_pmp_2_addr),
    .io_check_env_pmp_2_mask(PMPChecker_io_check_env_pmp_2_mask),
    .io_check_env_pmp_3_cfg_l(PMPChecker_io_check_env_pmp_3_cfg_l),
    .io_check_env_pmp_3_cfg_a(PMPChecker_io_check_env_pmp_3_cfg_a),
    .io_check_env_pmp_3_cfg_x(PMPChecker_io_check_env_pmp_3_cfg_x),
    .io_check_env_pmp_3_cfg_w(PMPChecker_io_check_env_pmp_3_cfg_w),
    .io_check_env_pmp_3_cfg_r(PMPChecker_io_check_env_pmp_3_cfg_r),
    .io_check_env_pmp_3_addr(PMPChecker_io_check_env_pmp_3_addr),
    .io_check_env_pmp_3_mask(PMPChecker_io_check_env_pmp_3_mask),
    .io_check_env_pmp_4_cfg_l(PMPChecker_io_check_env_pmp_4_cfg_l),
    .io_check_env_pmp_4_cfg_a(PMPChecker_io_check_env_pmp_4_cfg_a),
    .io_check_env_pmp_4_cfg_x(PMPChecker_io_check_env_pmp_4_cfg_x),
    .io_check_env_pmp_4_cfg_w(PMPChecker_io_check_env_pmp_4_cfg_w),
    .io_check_env_pmp_4_cfg_r(PMPChecker_io_check_env_pmp_4_cfg_r),
    .io_check_env_pmp_4_addr(PMPChecker_io_check_env_pmp_4_addr),
    .io_check_env_pmp_4_mask(PMPChecker_io_check_env_pmp_4_mask),
    .io_check_env_pmp_5_cfg_l(PMPChecker_io_check_env_pmp_5_cfg_l),
    .io_check_env_pmp_5_cfg_a(PMPChecker_io_check_env_pmp_5_cfg_a),
    .io_check_env_pmp_5_cfg_x(PMPChecker_io_check_env_pmp_5_cfg_x),
    .io_check_env_pmp_5_cfg_w(PMPChecker_io_check_env_pmp_5_cfg_w),
    .io_check_env_pmp_5_cfg_r(PMPChecker_io_check_env_pmp_5_cfg_r),
    .io_check_env_pmp_5_addr(PMPChecker_io_check_env_pmp_5_addr),
    .io_check_env_pmp_5_mask(PMPChecker_io_check_env_pmp_5_mask),
    .io_check_env_pmp_6_cfg_l(PMPChecker_io_check_env_pmp_6_cfg_l),
    .io_check_env_pmp_6_cfg_a(PMPChecker_io_check_env_pmp_6_cfg_a),
    .io_check_env_pmp_6_cfg_x(PMPChecker_io_check_env_pmp_6_cfg_x),
    .io_check_env_pmp_6_cfg_w(PMPChecker_io_check_env_pmp_6_cfg_w),
    .io_check_env_pmp_6_cfg_r(PMPChecker_io_check_env_pmp_6_cfg_r),
    .io_check_env_pmp_6_addr(PMPChecker_io_check_env_pmp_6_addr),
    .io_check_env_pmp_6_mask(PMPChecker_io_check_env_pmp_6_mask),
    .io_check_env_pmp_7_cfg_l(PMPChecker_io_check_env_pmp_7_cfg_l),
    .io_check_env_pmp_7_cfg_a(PMPChecker_io_check_env_pmp_7_cfg_a),
    .io_check_env_pmp_7_cfg_x(PMPChecker_io_check_env_pmp_7_cfg_x),
    .io_check_env_pmp_7_cfg_w(PMPChecker_io_check_env_pmp_7_cfg_w),
    .io_check_env_pmp_7_cfg_r(PMPChecker_io_check_env_pmp_7_cfg_r),
    .io_check_env_pmp_7_addr(PMPChecker_io_check_env_pmp_7_addr),
    .io_check_env_pmp_7_mask(PMPChecker_io_check_env_pmp_7_mask),
    .io_check_env_pmp_8_cfg_l(PMPChecker_io_check_env_pmp_8_cfg_l),
    .io_check_env_pmp_8_cfg_a(PMPChecker_io_check_env_pmp_8_cfg_a),
    .io_check_env_pmp_8_cfg_x(PMPChecker_io_check_env_pmp_8_cfg_x),
    .io_check_env_pmp_8_cfg_w(PMPChecker_io_check_env_pmp_8_cfg_w),
    .io_check_env_pmp_8_cfg_r(PMPChecker_io_check_env_pmp_8_cfg_r),
    .io_check_env_pmp_8_addr(PMPChecker_io_check_env_pmp_8_addr),
    .io_check_env_pmp_8_mask(PMPChecker_io_check_env_pmp_8_mask),
    .io_check_env_pmp_9_cfg_l(PMPChecker_io_check_env_pmp_9_cfg_l),
    .io_check_env_pmp_9_cfg_a(PMPChecker_io_check_env_pmp_9_cfg_a),
    .io_check_env_pmp_9_cfg_x(PMPChecker_io_check_env_pmp_9_cfg_x),
    .io_check_env_pmp_9_cfg_w(PMPChecker_io_check_env_pmp_9_cfg_w),
    .io_check_env_pmp_9_cfg_r(PMPChecker_io_check_env_pmp_9_cfg_r),
    .io_check_env_pmp_9_addr(PMPChecker_io_check_env_pmp_9_addr),
    .io_check_env_pmp_9_mask(PMPChecker_io_check_env_pmp_9_mask),
    .io_check_env_pmp_10_cfg_l(PMPChecker_io_check_env_pmp_10_cfg_l),
    .io_check_env_pmp_10_cfg_a(PMPChecker_io_check_env_pmp_10_cfg_a),
    .io_check_env_pmp_10_cfg_x(PMPChecker_io_check_env_pmp_10_cfg_x),
    .io_check_env_pmp_10_cfg_w(PMPChecker_io_check_env_pmp_10_cfg_w),
    .io_check_env_pmp_10_cfg_r(PMPChecker_io_check_env_pmp_10_cfg_r),
    .io_check_env_pmp_10_addr(PMPChecker_io_check_env_pmp_10_addr),
    .io_check_env_pmp_10_mask(PMPChecker_io_check_env_pmp_10_mask),
    .io_check_env_pmp_11_cfg_l(PMPChecker_io_check_env_pmp_11_cfg_l),
    .io_check_env_pmp_11_cfg_a(PMPChecker_io_check_env_pmp_11_cfg_a),
    .io_check_env_pmp_11_cfg_x(PMPChecker_io_check_env_pmp_11_cfg_x),
    .io_check_env_pmp_11_cfg_w(PMPChecker_io_check_env_pmp_11_cfg_w),
    .io_check_env_pmp_11_cfg_r(PMPChecker_io_check_env_pmp_11_cfg_r),
    .io_check_env_pmp_11_addr(PMPChecker_io_check_env_pmp_11_addr),
    .io_check_env_pmp_11_mask(PMPChecker_io_check_env_pmp_11_mask),
    .io_check_env_pmp_12_cfg_l(PMPChecker_io_check_env_pmp_12_cfg_l),
    .io_check_env_pmp_12_cfg_a(PMPChecker_io_check_env_pmp_12_cfg_a),
    .io_check_env_pmp_12_cfg_x(PMPChecker_io_check_env_pmp_12_cfg_x),
    .io_check_env_pmp_12_cfg_w(PMPChecker_io_check_env_pmp_12_cfg_w),
    .io_check_env_pmp_12_cfg_r(PMPChecker_io_check_env_pmp_12_cfg_r),
    .io_check_env_pmp_12_addr(PMPChecker_io_check_env_pmp_12_addr),
    .io_check_env_pmp_12_mask(PMPChecker_io_check_env_pmp_12_mask),
    .io_check_env_pmp_13_cfg_l(PMPChecker_io_check_env_pmp_13_cfg_l),
    .io_check_env_pmp_13_cfg_a(PMPChecker_io_check_env_pmp_13_cfg_a),
    .io_check_env_pmp_13_cfg_x(PMPChecker_io_check_env_pmp_13_cfg_x),
    .io_check_env_pmp_13_cfg_w(PMPChecker_io_check_env_pmp_13_cfg_w),
    .io_check_env_pmp_13_cfg_r(PMPChecker_io_check_env_pmp_13_cfg_r),
    .io_check_env_pmp_13_addr(PMPChecker_io_check_env_pmp_13_addr),
    .io_check_env_pmp_13_mask(PMPChecker_io_check_env_pmp_13_mask),
    .io_check_env_pmp_14_cfg_l(PMPChecker_io_check_env_pmp_14_cfg_l),
    .io_check_env_pmp_14_cfg_a(PMPChecker_io_check_env_pmp_14_cfg_a),
    .io_check_env_pmp_14_cfg_x(PMPChecker_io_check_env_pmp_14_cfg_x),
    .io_check_env_pmp_14_cfg_w(PMPChecker_io_check_env_pmp_14_cfg_w),
    .io_check_env_pmp_14_cfg_r(PMPChecker_io_check_env_pmp_14_cfg_r),
    .io_check_env_pmp_14_addr(PMPChecker_io_check_env_pmp_14_addr),
    .io_check_env_pmp_14_mask(PMPChecker_io_check_env_pmp_14_mask),
    .io_check_env_pmp_15_cfg_l(PMPChecker_io_check_env_pmp_15_cfg_l),
    .io_check_env_pmp_15_cfg_a(PMPChecker_io_check_env_pmp_15_cfg_a),
    .io_check_env_pmp_15_cfg_x(PMPChecker_io_check_env_pmp_15_cfg_x),
    .io_check_env_pmp_15_cfg_w(PMPChecker_io_check_env_pmp_15_cfg_w),
    .io_check_env_pmp_15_cfg_r(PMPChecker_io_check_env_pmp_15_cfg_r),
    .io_check_env_pmp_15_addr(PMPChecker_io_check_env_pmp_15_addr),
    .io_check_env_pmp_15_mask(PMPChecker_io_check_env_pmp_15_mask),
    .io_check_env_pma_0_cfg_c(PMPChecker_io_check_env_pma_0_cfg_c),
    .io_check_env_pma_0_cfg_atomic(PMPChecker_io_check_env_pma_0_cfg_atomic),
    .io_check_env_pma_0_cfg_a(PMPChecker_io_check_env_pma_0_cfg_a),
    .io_check_env_pma_0_cfg_x(PMPChecker_io_check_env_pma_0_cfg_x),
    .io_check_env_pma_0_cfg_w(PMPChecker_io_check_env_pma_0_cfg_w),
    .io_check_env_pma_0_cfg_r(PMPChecker_io_check_env_pma_0_cfg_r),
    .io_check_env_pma_0_addr(PMPChecker_io_check_env_pma_0_addr),
    .io_check_env_pma_0_mask(PMPChecker_io_check_env_pma_0_mask),
    .io_check_env_pma_1_cfg_c(PMPChecker_io_check_env_pma_1_cfg_c),
    .io_check_env_pma_1_cfg_atomic(PMPChecker_io_check_env_pma_1_cfg_atomic),
    .io_check_env_pma_1_cfg_a(PMPChecker_io_check_env_pma_1_cfg_a),
    .io_check_env_pma_1_cfg_x(PMPChecker_io_check_env_pma_1_cfg_x),
    .io_check_env_pma_1_cfg_w(PMPChecker_io_check_env_pma_1_cfg_w),
    .io_check_env_pma_1_cfg_r(PMPChecker_io_check_env_pma_1_cfg_r),
    .io_check_env_pma_1_addr(PMPChecker_io_check_env_pma_1_addr),
    .io_check_env_pma_1_mask(PMPChecker_io_check_env_pma_1_mask),
    .io_check_env_pma_2_cfg_c(PMPChecker_io_check_env_pma_2_cfg_c),
    .io_check_env_pma_2_cfg_atomic(PMPChecker_io_check_env_pma_2_cfg_atomic),
    .io_check_env_pma_2_cfg_a(PMPChecker_io_check_env_pma_2_cfg_a),
    .io_check_env_pma_2_cfg_x(PMPChecker_io_check_env_pma_2_cfg_x),
    .io_check_env_pma_2_cfg_w(PMPChecker_io_check_env_pma_2_cfg_w),
    .io_check_env_pma_2_cfg_r(PMPChecker_io_check_env_pma_2_cfg_r),
    .io_check_env_pma_2_addr(PMPChecker_io_check_env_pma_2_addr),
    .io_check_env_pma_2_mask(PMPChecker_io_check_env_pma_2_mask),
    .io_check_env_pma_3_cfg_c(PMPChecker_io_check_env_pma_3_cfg_c),
    .io_check_env_pma_3_cfg_atomic(PMPChecker_io_check_env_pma_3_cfg_atomic),
    .io_check_env_pma_3_cfg_a(PMPChecker_io_check_env_pma_3_cfg_a),
    .io_check_env_pma_3_cfg_x(PMPChecker_io_check_env_pma_3_cfg_x),
    .io_check_env_pma_3_cfg_w(PMPChecker_io_check_env_pma_3_cfg_w),
    .io_check_env_pma_3_cfg_r(PMPChecker_io_check_env_pma_3_cfg_r),
    .io_check_env_pma_3_addr(PMPChecker_io_check_env_pma_3_addr),
    .io_check_env_pma_3_mask(PMPChecker_io_check_env_pma_3_mask),
    .io_check_env_pma_4_cfg_c(PMPChecker_io_check_env_pma_4_cfg_c),
    .io_check_env_pma_4_cfg_atomic(PMPChecker_io_check_env_pma_4_cfg_atomic),
    .io_check_env_pma_4_cfg_a(PMPChecker_io_check_env_pma_4_cfg_a),
    .io_check_env_pma_4_cfg_x(PMPChecker_io_check_env_pma_4_cfg_x),
    .io_check_env_pma_4_cfg_w(PMPChecker_io_check_env_pma_4_cfg_w),
    .io_check_env_pma_4_cfg_r(PMPChecker_io_check_env_pma_4_cfg_r),
    .io_check_env_pma_4_addr(PMPChecker_io_check_env_pma_4_addr),
    .io_check_env_pma_4_mask(PMPChecker_io_check_env_pma_4_mask),
    .io_check_env_pma_5_cfg_c(PMPChecker_io_check_env_pma_5_cfg_c),
    .io_check_env_pma_5_cfg_atomic(PMPChecker_io_check_env_pma_5_cfg_atomic),
    .io_check_env_pma_5_cfg_a(PMPChecker_io_check_env_pma_5_cfg_a),
    .io_check_env_pma_5_cfg_x(PMPChecker_io_check_env_pma_5_cfg_x),
    .io_check_env_pma_5_cfg_w(PMPChecker_io_check_env_pma_5_cfg_w),
    .io_check_env_pma_5_cfg_r(PMPChecker_io_check_env_pma_5_cfg_r),
    .io_check_env_pma_5_addr(PMPChecker_io_check_env_pma_5_addr),
    .io_check_env_pma_5_mask(PMPChecker_io_check_env_pma_5_mask),
    .io_check_env_pma_6_cfg_c(PMPChecker_io_check_env_pma_6_cfg_c),
    .io_check_env_pma_6_cfg_atomic(PMPChecker_io_check_env_pma_6_cfg_atomic),
    .io_check_env_pma_6_cfg_a(PMPChecker_io_check_env_pma_6_cfg_a),
    .io_check_env_pma_6_cfg_x(PMPChecker_io_check_env_pma_6_cfg_x),
    .io_check_env_pma_6_cfg_w(PMPChecker_io_check_env_pma_6_cfg_w),
    .io_check_env_pma_6_cfg_r(PMPChecker_io_check_env_pma_6_cfg_r),
    .io_check_env_pma_6_addr(PMPChecker_io_check_env_pma_6_addr),
    .io_check_env_pma_6_mask(PMPChecker_io_check_env_pma_6_mask),
    .io_check_env_pma_7_cfg_c(PMPChecker_io_check_env_pma_7_cfg_c),
    .io_check_env_pma_7_cfg_atomic(PMPChecker_io_check_env_pma_7_cfg_atomic),
    .io_check_env_pma_7_cfg_a(PMPChecker_io_check_env_pma_7_cfg_a),
    .io_check_env_pma_7_cfg_x(PMPChecker_io_check_env_pma_7_cfg_x),
    .io_check_env_pma_7_cfg_w(PMPChecker_io_check_env_pma_7_cfg_w),
    .io_check_env_pma_7_cfg_r(PMPChecker_io_check_env_pma_7_cfg_r),
    .io_check_env_pma_7_addr(PMPChecker_io_check_env_pma_7_addr),
    .io_check_env_pma_7_mask(PMPChecker_io_check_env_pma_7_mask),
    .io_check_env_pma_8_cfg_c(PMPChecker_io_check_env_pma_8_cfg_c),
    .io_check_env_pma_8_cfg_atomic(PMPChecker_io_check_env_pma_8_cfg_atomic),
    .io_check_env_pma_8_cfg_a(PMPChecker_io_check_env_pma_8_cfg_a),
    .io_check_env_pma_8_cfg_x(PMPChecker_io_check_env_pma_8_cfg_x),
    .io_check_env_pma_8_cfg_w(PMPChecker_io_check_env_pma_8_cfg_w),
    .io_check_env_pma_8_cfg_r(PMPChecker_io_check_env_pma_8_cfg_r),
    .io_check_env_pma_8_addr(PMPChecker_io_check_env_pma_8_addr),
    .io_check_env_pma_8_mask(PMPChecker_io_check_env_pma_8_mask),
    .io_check_env_pma_9_cfg_c(PMPChecker_io_check_env_pma_9_cfg_c),
    .io_check_env_pma_9_cfg_atomic(PMPChecker_io_check_env_pma_9_cfg_atomic),
    .io_check_env_pma_9_cfg_a(PMPChecker_io_check_env_pma_9_cfg_a),
    .io_check_env_pma_9_cfg_x(PMPChecker_io_check_env_pma_9_cfg_x),
    .io_check_env_pma_9_cfg_w(PMPChecker_io_check_env_pma_9_cfg_w),
    .io_check_env_pma_9_cfg_r(PMPChecker_io_check_env_pma_9_cfg_r),
    .io_check_env_pma_9_addr(PMPChecker_io_check_env_pma_9_addr),
    .io_check_env_pma_9_mask(PMPChecker_io_check_env_pma_9_mask),
    .io_check_env_pma_10_cfg_c(PMPChecker_io_check_env_pma_10_cfg_c),
    .io_check_env_pma_10_cfg_atomic(PMPChecker_io_check_env_pma_10_cfg_atomic),
    .io_check_env_pma_10_cfg_a(PMPChecker_io_check_env_pma_10_cfg_a),
    .io_check_env_pma_10_cfg_x(PMPChecker_io_check_env_pma_10_cfg_x),
    .io_check_env_pma_10_cfg_w(PMPChecker_io_check_env_pma_10_cfg_w),
    .io_check_env_pma_10_cfg_r(PMPChecker_io_check_env_pma_10_cfg_r),
    .io_check_env_pma_10_addr(PMPChecker_io_check_env_pma_10_addr),
    .io_check_env_pma_10_mask(PMPChecker_io_check_env_pma_10_mask),
    .io_check_env_pma_11_cfg_c(PMPChecker_io_check_env_pma_11_cfg_c),
    .io_check_env_pma_11_cfg_atomic(PMPChecker_io_check_env_pma_11_cfg_atomic),
    .io_check_env_pma_11_cfg_a(PMPChecker_io_check_env_pma_11_cfg_a),
    .io_check_env_pma_11_cfg_x(PMPChecker_io_check_env_pma_11_cfg_x),
    .io_check_env_pma_11_cfg_w(PMPChecker_io_check_env_pma_11_cfg_w),
    .io_check_env_pma_11_cfg_r(PMPChecker_io_check_env_pma_11_cfg_r),
    .io_check_env_pma_11_addr(PMPChecker_io_check_env_pma_11_addr),
    .io_check_env_pma_11_mask(PMPChecker_io_check_env_pma_11_mask),
    .io_check_env_pma_12_cfg_c(PMPChecker_io_check_env_pma_12_cfg_c),
    .io_check_env_pma_12_cfg_atomic(PMPChecker_io_check_env_pma_12_cfg_atomic),
    .io_check_env_pma_12_cfg_a(PMPChecker_io_check_env_pma_12_cfg_a),
    .io_check_env_pma_12_cfg_x(PMPChecker_io_check_env_pma_12_cfg_x),
    .io_check_env_pma_12_cfg_w(PMPChecker_io_check_env_pma_12_cfg_w),
    .io_check_env_pma_12_cfg_r(PMPChecker_io_check_env_pma_12_cfg_r),
    .io_check_env_pma_12_addr(PMPChecker_io_check_env_pma_12_addr),
    .io_check_env_pma_12_mask(PMPChecker_io_check_env_pma_12_mask),
    .io_check_env_pma_13_cfg_c(PMPChecker_io_check_env_pma_13_cfg_c),
    .io_check_env_pma_13_cfg_atomic(PMPChecker_io_check_env_pma_13_cfg_atomic),
    .io_check_env_pma_13_cfg_a(PMPChecker_io_check_env_pma_13_cfg_a),
    .io_check_env_pma_13_cfg_x(PMPChecker_io_check_env_pma_13_cfg_x),
    .io_check_env_pma_13_cfg_w(PMPChecker_io_check_env_pma_13_cfg_w),
    .io_check_env_pma_13_cfg_r(PMPChecker_io_check_env_pma_13_cfg_r),
    .io_check_env_pma_13_addr(PMPChecker_io_check_env_pma_13_addr),
    .io_check_env_pma_13_mask(PMPChecker_io_check_env_pma_13_mask),
    .io_check_env_pma_14_cfg_c(PMPChecker_io_check_env_pma_14_cfg_c),
    .io_check_env_pma_14_cfg_atomic(PMPChecker_io_check_env_pma_14_cfg_atomic),
    .io_check_env_pma_14_cfg_a(PMPChecker_io_check_env_pma_14_cfg_a),
    .io_check_env_pma_14_cfg_x(PMPChecker_io_check_env_pma_14_cfg_x),
    .io_check_env_pma_14_cfg_w(PMPChecker_io_check_env_pma_14_cfg_w),
    .io_check_env_pma_14_cfg_r(PMPChecker_io_check_env_pma_14_cfg_r),
    .io_check_env_pma_14_addr(PMPChecker_io_check_env_pma_14_addr),
    .io_check_env_pma_14_mask(PMPChecker_io_check_env_pma_14_mask),
    .io_check_env_pma_15_cfg_c(PMPChecker_io_check_env_pma_15_cfg_c),
    .io_check_env_pma_15_cfg_atomic(PMPChecker_io_check_env_pma_15_cfg_atomic),
    .io_check_env_pma_15_cfg_a(PMPChecker_io_check_env_pma_15_cfg_a),
    .io_check_env_pma_15_cfg_x(PMPChecker_io_check_env_pma_15_cfg_x),
    .io_check_env_pma_15_cfg_w(PMPChecker_io_check_env_pma_15_cfg_w),
    .io_check_env_pma_15_cfg_r(PMPChecker_io_check_env_pma_15_cfg_r),
    .io_check_env_pma_15_addr(PMPChecker_io_check_env_pma_15_addr),
    .io_check_env_pma_15_mask(PMPChecker_io_check_env_pma_15_mask),
    .io_req_bits_addr(PMPChecker_io_req_bits_addr),
    .io_req_bits_cmd(PMPChecker_io_req_bits_cmd),
    .io_resp_ld(PMPChecker_io_resp_ld),
    .io_resp_st(PMPChecker_io_resp_st),
    .io_resp_instr(PMPChecker_io_resp_instr),
    .io_resp_mmio(PMPChecker_io_resp_mmio),
    .io_resp_atomic(PMPChecker_io_resp_atomic)
  );
  PMPChecker PMPChecker_1 ( // @[TLPMA.scala 47:13]
    .io_check_env_mode(PMPChecker_1_io_check_env_mode),
    .io_check_env_pmp_0_cfg_l(PMPChecker_1_io_check_env_pmp_0_cfg_l),
    .io_check_env_pmp_0_cfg_a(PMPChecker_1_io_check_env_pmp_0_cfg_a),
    .io_check_env_pmp_0_cfg_x(PMPChecker_1_io_check_env_pmp_0_cfg_x),
    .io_check_env_pmp_0_cfg_w(PMPChecker_1_io_check_env_pmp_0_cfg_w),
    .io_check_env_pmp_0_cfg_r(PMPChecker_1_io_check_env_pmp_0_cfg_r),
    .io_check_env_pmp_0_addr(PMPChecker_1_io_check_env_pmp_0_addr),
    .io_check_env_pmp_0_mask(PMPChecker_1_io_check_env_pmp_0_mask),
    .io_check_env_pmp_1_cfg_l(PMPChecker_1_io_check_env_pmp_1_cfg_l),
    .io_check_env_pmp_1_cfg_a(PMPChecker_1_io_check_env_pmp_1_cfg_a),
    .io_check_env_pmp_1_cfg_x(PMPChecker_1_io_check_env_pmp_1_cfg_x),
    .io_check_env_pmp_1_cfg_w(PMPChecker_1_io_check_env_pmp_1_cfg_w),
    .io_check_env_pmp_1_cfg_r(PMPChecker_1_io_check_env_pmp_1_cfg_r),
    .io_check_env_pmp_1_addr(PMPChecker_1_io_check_env_pmp_1_addr),
    .io_check_env_pmp_1_mask(PMPChecker_1_io_check_env_pmp_1_mask),
    .io_check_env_pmp_2_cfg_l(PMPChecker_1_io_check_env_pmp_2_cfg_l),
    .io_check_env_pmp_2_cfg_a(PMPChecker_1_io_check_env_pmp_2_cfg_a),
    .io_check_env_pmp_2_cfg_x(PMPChecker_1_io_check_env_pmp_2_cfg_x),
    .io_check_env_pmp_2_cfg_w(PMPChecker_1_io_check_env_pmp_2_cfg_w),
    .io_check_env_pmp_2_cfg_r(PMPChecker_1_io_check_env_pmp_2_cfg_r),
    .io_check_env_pmp_2_addr(PMPChecker_1_io_check_env_pmp_2_addr),
    .io_check_env_pmp_2_mask(PMPChecker_1_io_check_env_pmp_2_mask),
    .io_check_env_pmp_3_cfg_l(PMPChecker_1_io_check_env_pmp_3_cfg_l),
    .io_check_env_pmp_3_cfg_a(PMPChecker_1_io_check_env_pmp_3_cfg_a),
    .io_check_env_pmp_3_cfg_x(PMPChecker_1_io_check_env_pmp_3_cfg_x),
    .io_check_env_pmp_3_cfg_w(PMPChecker_1_io_check_env_pmp_3_cfg_w),
    .io_check_env_pmp_3_cfg_r(PMPChecker_1_io_check_env_pmp_3_cfg_r),
    .io_check_env_pmp_3_addr(PMPChecker_1_io_check_env_pmp_3_addr),
    .io_check_env_pmp_3_mask(PMPChecker_1_io_check_env_pmp_3_mask),
    .io_check_env_pmp_4_cfg_l(PMPChecker_1_io_check_env_pmp_4_cfg_l),
    .io_check_env_pmp_4_cfg_a(PMPChecker_1_io_check_env_pmp_4_cfg_a),
    .io_check_env_pmp_4_cfg_x(PMPChecker_1_io_check_env_pmp_4_cfg_x),
    .io_check_env_pmp_4_cfg_w(PMPChecker_1_io_check_env_pmp_4_cfg_w),
    .io_check_env_pmp_4_cfg_r(PMPChecker_1_io_check_env_pmp_4_cfg_r),
    .io_check_env_pmp_4_addr(PMPChecker_1_io_check_env_pmp_4_addr),
    .io_check_env_pmp_4_mask(PMPChecker_1_io_check_env_pmp_4_mask),
    .io_check_env_pmp_5_cfg_l(PMPChecker_1_io_check_env_pmp_5_cfg_l),
    .io_check_env_pmp_5_cfg_a(PMPChecker_1_io_check_env_pmp_5_cfg_a),
    .io_check_env_pmp_5_cfg_x(PMPChecker_1_io_check_env_pmp_5_cfg_x),
    .io_check_env_pmp_5_cfg_w(PMPChecker_1_io_check_env_pmp_5_cfg_w),
    .io_check_env_pmp_5_cfg_r(PMPChecker_1_io_check_env_pmp_5_cfg_r),
    .io_check_env_pmp_5_addr(PMPChecker_1_io_check_env_pmp_5_addr),
    .io_check_env_pmp_5_mask(PMPChecker_1_io_check_env_pmp_5_mask),
    .io_check_env_pmp_6_cfg_l(PMPChecker_1_io_check_env_pmp_6_cfg_l),
    .io_check_env_pmp_6_cfg_a(PMPChecker_1_io_check_env_pmp_6_cfg_a),
    .io_check_env_pmp_6_cfg_x(PMPChecker_1_io_check_env_pmp_6_cfg_x),
    .io_check_env_pmp_6_cfg_w(PMPChecker_1_io_check_env_pmp_6_cfg_w),
    .io_check_env_pmp_6_cfg_r(PMPChecker_1_io_check_env_pmp_6_cfg_r),
    .io_check_env_pmp_6_addr(PMPChecker_1_io_check_env_pmp_6_addr),
    .io_check_env_pmp_6_mask(PMPChecker_1_io_check_env_pmp_6_mask),
    .io_check_env_pmp_7_cfg_l(PMPChecker_1_io_check_env_pmp_7_cfg_l),
    .io_check_env_pmp_7_cfg_a(PMPChecker_1_io_check_env_pmp_7_cfg_a),
    .io_check_env_pmp_7_cfg_x(PMPChecker_1_io_check_env_pmp_7_cfg_x),
    .io_check_env_pmp_7_cfg_w(PMPChecker_1_io_check_env_pmp_7_cfg_w),
    .io_check_env_pmp_7_cfg_r(PMPChecker_1_io_check_env_pmp_7_cfg_r),
    .io_check_env_pmp_7_addr(PMPChecker_1_io_check_env_pmp_7_addr),
    .io_check_env_pmp_7_mask(PMPChecker_1_io_check_env_pmp_7_mask),
    .io_check_env_pmp_8_cfg_l(PMPChecker_1_io_check_env_pmp_8_cfg_l),
    .io_check_env_pmp_8_cfg_a(PMPChecker_1_io_check_env_pmp_8_cfg_a),
    .io_check_env_pmp_8_cfg_x(PMPChecker_1_io_check_env_pmp_8_cfg_x),
    .io_check_env_pmp_8_cfg_w(PMPChecker_1_io_check_env_pmp_8_cfg_w),
    .io_check_env_pmp_8_cfg_r(PMPChecker_1_io_check_env_pmp_8_cfg_r),
    .io_check_env_pmp_8_addr(PMPChecker_1_io_check_env_pmp_8_addr),
    .io_check_env_pmp_8_mask(PMPChecker_1_io_check_env_pmp_8_mask),
    .io_check_env_pmp_9_cfg_l(PMPChecker_1_io_check_env_pmp_9_cfg_l),
    .io_check_env_pmp_9_cfg_a(PMPChecker_1_io_check_env_pmp_9_cfg_a),
    .io_check_env_pmp_9_cfg_x(PMPChecker_1_io_check_env_pmp_9_cfg_x),
    .io_check_env_pmp_9_cfg_w(PMPChecker_1_io_check_env_pmp_9_cfg_w),
    .io_check_env_pmp_9_cfg_r(PMPChecker_1_io_check_env_pmp_9_cfg_r),
    .io_check_env_pmp_9_addr(PMPChecker_1_io_check_env_pmp_9_addr),
    .io_check_env_pmp_9_mask(PMPChecker_1_io_check_env_pmp_9_mask),
    .io_check_env_pmp_10_cfg_l(PMPChecker_1_io_check_env_pmp_10_cfg_l),
    .io_check_env_pmp_10_cfg_a(PMPChecker_1_io_check_env_pmp_10_cfg_a),
    .io_check_env_pmp_10_cfg_x(PMPChecker_1_io_check_env_pmp_10_cfg_x),
    .io_check_env_pmp_10_cfg_w(PMPChecker_1_io_check_env_pmp_10_cfg_w),
    .io_check_env_pmp_10_cfg_r(PMPChecker_1_io_check_env_pmp_10_cfg_r),
    .io_check_env_pmp_10_addr(PMPChecker_1_io_check_env_pmp_10_addr),
    .io_check_env_pmp_10_mask(PMPChecker_1_io_check_env_pmp_10_mask),
    .io_check_env_pmp_11_cfg_l(PMPChecker_1_io_check_env_pmp_11_cfg_l),
    .io_check_env_pmp_11_cfg_a(PMPChecker_1_io_check_env_pmp_11_cfg_a),
    .io_check_env_pmp_11_cfg_x(PMPChecker_1_io_check_env_pmp_11_cfg_x),
    .io_check_env_pmp_11_cfg_w(PMPChecker_1_io_check_env_pmp_11_cfg_w),
    .io_check_env_pmp_11_cfg_r(PMPChecker_1_io_check_env_pmp_11_cfg_r),
    .io_check_env_pmp_11_addr(PMPChecker_1_io_check_env_pmp_11_addr),
    .io_check_env_pmp_11_mask(PMPChecker_1_io_check_env_pmp_11_mask),
    .io_check_env_pmp_12_cfg_l(PMPChecker_1_io_check_env_pmp_12_cfg_l),
    .io_check_env_pmp_12_cfg_a(PMPChecker_1_io_check_env_pmp_12_cfg_a),
    .io_check_env_pmp_12_cfg_x(PMPChecker_1_io_check_env_pmp_12_cfg_x),
    .io_check_env_pmp_12_cfg_w(PMPChecker_1_io_check_env_pmp_12_cfg_w),
    .io_check_env_pmp_12_cfg_r(PMPChecker_1_io_check_env_pmp_12_cfg_r),
    .io_check_env_pmp_12_addr(PMPChecker_1_io_check_env_pmp_12_addr),
    .io_check_env_pmp_12_mask(PMPChecker_1_io_check_env_pmp_12_mask),
    .io_check_env_pmp_13_cfg_l(PMPChecker_1_io_check_env_pmp_13_cfg_l),
    .io_check_env_pmp_13_cfg_a(PMPChecker_1_io_check_env_pmp_13_cfg_a),
    .io_check_env_pmp_13_cfg_x(PMPChecker_1_io_check_env_pmp_13_cfg_x),
    .io_check_env_pmp_13_cfg_w(PMPChecker_1_io_check_env_pmp_13_cfg_w),
    .io_check_env_pmp_13_cfg_r(PMPChecker_1_io_check_env_pmp_13_cfg_r),
    .io_check_env_pmp_13_addr(PMPChecker_1_io_check_env_pmp_13_addr),
    .io_check_env_pmp_13_mask(PMPChecker_1_io_check_env_pmp_13_mask),
    .io_check_env_pmp_14_cfg_l(PMPChecker_1_io_check_env_pmp_14_cfg_l),
    .io_check_env_pmp_14_cfg_a(PMPChecker_1_io_check_env_pmp_14_cfg_a),
    .io_check_env_pmp_14_cfg_x(PMPChecker_1_io_check_env_pmp_14_cfg_x),
    .io_check_env_pmp_14_cfg_w(PMPChecker_1_io_check_env_pmp_14_cfg_w),
    .io_check_env_pmp_14_cfg_r(PMPChecker_1_io_check_env_pmp_14_cfg_r),
    .io_check_env_pmp_14_addr(PMPChecker_1_io_check_env_pmp_14_addr),
    .io_check_env_pmp_14_mask(PMPChecker_1_io_check_env_pmp_14_mask),
    .io_check_env_pmp_15_cfg_l(PMPChecker_1_io_check_env_pmp_15_cfg_l),
    .io_check_env_pmp_15_cfg_a(PMPChecker_1_io_check_env_pmp_15_cfg_a),
    .io_check_env_pmp_15_cfg_x(PMPChecker_1_io_check_env_pmp_15_cfg_x),
    .io_check_env_pmp_15_cfg_w(PMPChecker_1_io_check_env_pmp_15_cfg_w),
    .io_check_env_pmp_15_cfg_r(PMPChecker_1_io_check_env_pmp_15_cfg_r),
    .io_check_env_pmp_15_addr(PMPChecker_1_io_check_env_pmp_15_addr),
    .io_check_env_pmp_15_mask(PMPChecker_1_io_check_env_pmp_15_mask),
    .io_check_env_pma_0_cfg_c(PMPChecker_1_io_check_env_pma_0_cfg_c),
    .io_check_env_pma_0_cfg_atomic(PMPChecker_1_io_check_env_pma_0_cfg_atomic),
    .io_check_env_pma_0_cfg_a(PMPChecker_1_io_check_env_pma_0_cfg_a),
    .io_check_env_pma_0_cfg_x(PMPChecker_1_io_check_env_pma_0_cfg_x),
    .io_check_env_pma_0_cfg_w(PMPChecker_1_io_check_env_pma_0_cfg_w),
    .io_check_env_pma_0_cfg_r(PMPChecker_1_io_check_env_pma_0_cfg_r),
    .io_check_env_pma_0_addr(PMPChecker_1_io_check_env_pma_0_addr),
    .io_check_env_pma_0_mask(PMPChecker_1_io_check_env_pma_0_mask),
    .io_check_env_pma_1_cfg_c(PMPChecker_1_io_check_env_pma_1_cfg_c),
    .io_check_env_pma_1_cfg_atomic(PMPChecker_1_io_check_env_pma_1_cfg_atomic),
    .io_check_env_pma_1_cfg_a(PMPChecker_1_io_check_env_pma_1_cfg_a),
    .io_check_env_pma_1_cfg_x(PMPChecker_1_io_check_env_pma_1_cfg_x),
    .io_check_env_pma_1_cfg_w(PMPChecker_1_io_check_env_pma_1_cfg_w),
    .io_check_env_pma_1_cfg_r(PMPChecker_1_io_check_env_pma_1_cfg_r),
    .io_check_env_pma_1_addr(PMPChecker_1_io_check_env_pma_1_addr),
    .io_check_env_pma_1_mask(PMPChecker_1_io_check_env_pma_1_mask),
    .io_check_env_pma_2_cfg_c(PMPChecker_1_io_check_env_pma_2_cfg_c),
    .io_check_env_pma_2_cfg_atomic(PMPChecker_1_io_check_env_pma_2_cfg_atomic),
    .io_check_env_pma_2_cfg_a(PMPChecker_1_io_check_env_pma_2_cfg_a),
    .io_check_env_pma_2_cfg_x(PMPChecker_1_io_check_env_pma_2_cfg_x),
    .io_check_env_pma_2_cfg_w(PMPChecker_1_io_check_env_pma_2_cfg_w),
    .io_check_env_pma_2_cfg_r(PMPChecker_1_io_check_env_pma_2_cfg_r),
    .io_check_env_pma_2_addr(PMPChecker_1_io_check_env_pma_2_addr),
    .io_check_env_pma_2_mask(PMPChecker_1_io_check_env_pma_2_mask),
    .io_check_env_pma_3_cfg_c(PMPChecker_1_io_check_env_pma_3_cfg_c),
    .io_check_env_pma_3_cfg_atomic(PMPChecker_1_io_check_env_pma_3_cfg_atomic),
    .io_check_env_pma_3_cfg_a(PMPChecker_1_io_check_env_pma_3_cfg_a),
    .io_check_env_pma_3_cfg_x(PMPChecker_1_io_check_env_pma_3_cfg_x),
    .io_check_env_pma_3_cfg_w(PMPChecker_1_io_check_env_pma_3_cfg_w),
    .io_check_env_pma_3_cfg_r(PMPChecker_1_io_check_env_pma_3_cfg_r),
    .io_check_env_pma_3_addr(PMPChecker_1_io_check_env_pma_3_addr),
    .io_check_env_pma_3_mask(PMPChecker_1_io_check_env_pma_3_mask),
    .io_check_env_pma_4_cfg_c(PMPChecker_1_io_check_env_pma_4_cfg_c),
    .io_check_env_pma_4_cfg_atomic(PMPChecker_1_io_check_env_pma_4_cfg_atomic),
    .io_check_env_pma_4_cfg_a(PMPChecker_1_io_check_env_pma_4_cfg_a),
    .io_check_env_pma_4_cfg_x(PMPChecker_1_io_check_env_pma_4_cfg_x),
    .io_check_env_pma_4_cfg_w(PMPChecker_1_io_check_env_pma_4_cfg_w),
    .io_check_env_pma_4_cfg_r(PMPChecker_1_io_check_env_pma_4_cfg_r),
    .io_check_env_pma_4_addr(PMPChecker_1_io_check_env_pma_4_addr),
    .io_check_env_pma_4_mask(PMPChecker_1_io_check_env_pma_4_mask),
    .io_check_env_pma_5_cfg_c(PMPChecker_1_io_check_env_pma_5_cfg_c),
    .io_check_env_pma_5_cfg_atomic(PMPChecker_1_io_check_env_pma_5_cfg_atomic),
    .io_check_env_pma_5_cfg_a(PMPChecker_1_io_check_env_pma_5_cfg_a),
    .io_check_env_pma_5_cfg_x(PMPChecker_1_io_check_env_pma_5_cfg_x),
    .io_check_env_pma_5_cfg_w(PMPChecker_1_io_check_env_pma_5_cfg_w),
    .io_check_env_pma_5_cfg_r(PMPChecker_1_io_check_env_pma_5_cfg_r),
    .io_check_env_pma_5_addr(PMPChecker_1_io_check_env_pma_5_addr),
    .io_check_env_pma_5_mask(PMPChecker_1_io_check_env_pma_5_mask),
    .io_check_env_pma_6_cfg_c(PMPChecker_1_io_check_env_pma_6_cfg_c),
    .io_check_env_pma_6_cfg_atomic(PMPChecker_1_io_check_env_pma_6_cfg_atomic),
    .io_check_env_pma_6_cfg_a(PMPChecker_1_io_check_env_pma_6_cfg_a),
    .io_check_env_pma_6_cfg_x(PMPChecker_1_io_check_env_pma_6_cfg_x),
    .io_check_env_pma_6_cfg_w(PMPChecker_1_io_check_env_pma_6_cfg_w),
    .io_check_env_pma_6_cfg_r(PMPChecker_1_io_check_env_pma_6_cfg_r),
    .io_check_env_pma_6_addr(PMPChecker_1_io_check_env_pma_6_addr),
    .io_check_env_pma_6_mask(PMPChecker_1_io_check_env_pma_6_mask),
    .io_check_env_pma_7_cfg_c(PMPChecker_1_io_check_env_pma_7_cfg_c),
    .io_check_env_pma_7_cfg_atomic(PMPChecker_1_io_check_env_pma_7_cfg_atomic),
    .io_check_env_pma_7_cfg_a(PMPChecker_1_io_check_env_pma_7_cfg_a),
    .io_check_env_pma_7_cfg_x(PMPChecker_1_io_check_env_pma_7_cfg_x),
    .io_check_env_pma_7_cfg_w(PMPChecker_1_io_check_env_pma_7_cfg_w),
    .io_check_env_pma_7_cfg_r(PMPChecker_1_io_check_env_pma_7_cfg_r),
    .io_check_env_pma_7_addr(PMPChecker_1_io_check_env_pma_7_addr),
    .io_check_env_pma_7_mask(PMPChecker_1_io_check_env_pma_7_mask),
    .io_check_env_pma_8_cfg_c(PMPChecker_1_io_check_env_pma_8_cfg_c),
    .io_check_env_pma_8_cfg_atomic(PMPChecker_1_io_check_env_pma_8_cfg_atomic),
    .io_check_env_pma_8_cfg_a(PMPChecker_1_io_check_env_pma_8_cfg_a),
    .io_check_env_pma_8_cfg_x(PMPChecker_1_io_check_env_pma_8_cfg_x),
    .io_check_env_pma_8_cfg_w(PMPChecker_1_io_check_env_pma_8_cfg_w),
    .io_check_env_pma_8_cfg_r(PMPChecker_1_io_check_env_pma_8_cfg_r),
    .io_check_env_pma_8_addr(PMPChecker_1_io_check_env_pma_8_addr),
    .io_check_env_pma_8_mask(PMPChecker_1_io_check_env_pma_8_mask),
    .io_check_env_pma_9_cfg_c(PMPChecker_1_io_check_env_pma_9_cfg_c),
    .io_check_env_pma_9_cfg_atomic(PMPChecker_1_io_check_env_pma_9_cfg_atomic),
    .io_check_env_pma_9_cfg_a(PMPChecker_1_io_check_env_pma_9_cfg_a),
    .io_check_env_pma_9_cfg_x(PMPChecker_1_io_check_env_pma_9_cfg_x),
    .io_check_env_pma_9_cfg_w(PMPChecker_1_io_check_env_pma_9_cfg_w),
    .io_check_env_pma_9_cfg_r(PMPChecker_1_io_check_env_pma_9_cfg_r),
    .io_check_env_pma_9_addr(PMPChecker_1_io_check_env_pma_9_addr),
    .io_check_env_pma_9_mask(PMPChecker_1_io_check_env_pma_9_mask),
    .io_check_env_pma_10_cfg_c(PMPChecker_1_io_check_env_pma_10_cfg_c),
    .io_check_env_pma_10_cfg_atomic(PMPChecker_1_io_check_env_pma_10_cfg_atomic),
    .io_check_env_pma_10_cfg_a(PMPChecker_1_io_check_env_pma_10_cfg_a),
    .io_check_env_pma_10_cfg_x(PMPChecker_1_io_check_env_pma_10_cfg_x),
    .io_check_env_pma_10_cfg_w(PMPChecker_1_io_check_env_pma_10_cfg_w),
    .io_check_env_pma_10_cfg_r(PMPChecker_1_io_check_env_pma_10_cfg_r),
    .io_check_env_pma_10_addr(PMPChecker_1_io_check_env_pma_10_addr),
    .io_check_env_pma_10_mask(PMPChecker_1_io_check_env_pma_10_mask),
    .io_check_env_pma_11_cfg_c(PMPChecker_1_io_check_env_pma_11_cfg_c),
    .io_check_env_pma_11_cfg_atomic(PMPChecker_1_io_check_env_pma_11_cfg_atomic),
    .io_check_env_pma_11_cfg_a(PMPChecker_1_io_check_env_pma_11_cfg_a),
    .io_check_env_pma_11_cfg_x(PMPChecker_1_io_check_env_pma_11_cfg_x),
    .io_check_env_pma_11_cfg_w(PMPChecker_1_io_check_env_pma_11_cfg_w),
    .io_check_env_pma_11_cfg_r(PMPChecker_1_io_check_env_pma_11_cfg_r),
    .io_check_env_pma_11_addr(PMPChecker_1_io_check_env_pma_11_addr),
    .io_check_env_pma_11_mask(PMPChecker_1_io_check_env_pma_11_mask),
    .io_check_env_pma_12_cfg_c(PMPChecker_1_io_check_env_pma_12_cfg_c),
    .io_check_env_pma_12_cfg_atomic(PMPChecker_1_io_check_env_pma_12_cfg_atomic),
    .io_check_env_pma_12_cfg_a(PMPChecker_1_io_check_env_pma_12_cfg_a),
    .io_check_env_pma_12_cfg_x(PMPChecker_1_io_check_env_pma_12_cfg_x),
    .io_check_env_pma_12_cfg_w(PMPChecker_1_io_check_env_pma_12_cfg_w),
    .io_check_env_pma_12_cfg_r(PMPChecker_1_io_check_env_pma_12_cfg_r),
    .io_check_env_pma_12_addr(PMPChecker_1_io_check_env_pma_12_addr),
    .io_check_env_pma_12_mask(PMPChecker_1_io_check_env_pma_12_mask),
    .io_check_env_pma_13_cfg_c(PMPChecker_1_io_check_env_pma_13_cfg_c),
    .io_check_env_pma_13_cfg_atomic(PMPChecker_1_io_check_env_pma_13_cfg_atomic),
    .io_check_env_pma_13_cfg_a(PMPChecker_1_io_check_env_pma_13_cfg_a),
    .io_check_env_pma_13_cfg_x(PMPChecker_1_io_check_env_pma_13_cfg_x),
    .io_check_env_pma_13_cfg_w(PMPChecker_1_io_check_env_pma_13_cfg_w),
    .io_check_env_pma_13_cfg_r(PMPChecker_1_io_check_env_pma_13_cfg_r),
    .io_check_env_pma_13_addr(PMPChecker_1_io_check_env_pma_13_addr),
    .io_check_env_pma_13_mask(PMPChecker_1_io_check_env_pma_13_mask),
    .io_check_env_pma_14_cfg_c(PMPChecker_1_io_check_env_pma_14_cfg_c),
    .io_check_env_pma_14_cfg_atomic(PMPChecker_1_io_check_env_pma_14_cfg_atomic),
    .io_check_env_pma_14_cfg_a(PMPChecker_1_io_check_env_pma_14_cfg_a),
    .io_check_env_pma_14_cfg_x(PMPChecker_1_io_check_env_pma_14_cfg_x),
    .io_check_env_pma_14_cfg_w(PMPChecker_1_io_check_env_pma_14_cfg_w),
    .io_check_env_pma_14_cfg_r(PMPChecker_1_io_check_env_pma_14_cfg_r),
    .io_check_env_pma_14_addr(PMPChecker_1_io_check_env_pma_14_addr),
    .io_check_env_pma_14_mask(PMPChecker_1_io_check_env_pma_14_mask),
    .io_check_env_pma_15_cfg_c(PMPChecker_1_io_check_env_pma_15_cfg_c),
    .io_check_env_pma_15_cfg_atomic(PMPChecker_1_io_check_env_pma_15_cfg_atomic),
    .io_check_env_pma_15_cfg_a(PMPChecker_1_io_check_env_pma_15_cfg_a),
    .io_check_env_pma_15_cfg_x(PMPChecker_1_io_check_env_pma_15_cfg_x),
    .io_check_env_pma_15_cfg_w(PMPChecker_1_io_check_env_pma_15_cfg_w),
    .io_check_env_pma_15_cfg_r(PMPChecker_1_io_check_env_pma_15_cfg_r),
    .io_check_env_pma_15_addr(PMPChecker_1_io_check_env_pma_15_addr),
    .io_check_env_pma_15_mask(PMPChecker_1_io_check_env_pma_15_mask),
    .io_req_bits_addr(PMPChecker_1_io_req_bits_addr),
    .io_req_bits_cmd(PMPChecker_1_io_req_bits_cmd),
    .io_resp_ld(PMPChecker_1_io_resp_ld),
    .io_resp_st(PMPChecker_1_io_resp_st),
    .io_resp_instr(PMPChecker_1_io_resp_instr),
    .io_resp_mmio(PMPChecker_1_io_resp_mmio),
    .io_resp_atomic(PMPChecker_1_io_resp_atomic)
  );
  assign auto_in_a_ready = out_front_ready & out_iready; // @[RegisterRouter.scala 82:24]
  assign auto_in_d_valid = out_back_io_deq_valid & out_oready; // @[RegisterRouter.scala 82:24]
  assign auto_in_d_bits_opcode = {{2'd0}, out_bits_read}; // @[Nodes.scala 1210:84 RegisterRouter.scala 97:19]
  assign auto_in_d_bits_size = out_back_io_deq_bits_extra_tlrr_extra_size; // @[RegisterRouter.scala 82:{24,24}]
  assign auto_in_d_bits_source = out_back_io_deq_bits_extra_tlrr_extra_source; // @[RegisterRouter.scala 82:{24,24}]
  assign auto_in_d_bits_data = _GEN_285 ? _GEN_317 : 64'h0; // @[RegisterRouter.scala 82:24]
  assign io_resp_0_ld = PMPChecker_io_resp_ld; // @[TLPMA.scala 46:{28,28}]
  assign io_resp_0_st = PMPChecker_io_resp_st; // @[TLPMA.scala 46:{28,28}]
  assign io_resp_0_instr = PMPChecker_io_resp_instr; // @[TLPMA.scala 46:{28,28}]
  assign io_resp_0_mmio = PMPChecker_io_resp_mmio; // @[TLPMA.scala 46:{28,28}]
  assign io_resp_0_atomic = PMPChecker_io_resp_atomic; // @[TLPMA.scala 46:{28,28}]
  assign io_resp_1_ld = PMPChecker_1_io_resp_ld; // @[TLPMA.scala 46:{28,28}]
  assign io_resp_1_st = PMPChecker_1_io_resp_st; // @[TLPMA.scala 46:{28,28}]
  assign io_resp_1_instr = PMPChecker_1_io_resp_instr; // @[TLPMA.scala 46:{28,28}]
  assign io_resp_1_mmio = PMPChecker_1_io_resp_mmio; // @[TLPMA.scala 46:{28,28}]
  assign io_resp_1_atomic = PMPChecker_1_io_resp_atomic; // @[TLPMA.scala 46:{28,28}]
  assign out_back_clock = clock;
  assign out_back_reset = reset;
  assign out_back_io_enq_valid = auto_in_a_valid & out_iready; // @[RegisterRouter.scala 82:24]
  assign out_back_io_enq_bits_read = auto_in_a_bits_opcode == 3'h4; // @[RegisterRouter.scala 71:36]
  assign out_back_io_enq_bits_index = auto_in_a_bits_address[11:3]; // @[RegisterRouter.scala 70:18 72:19]
  assign out_back_io_enq_bits_data = auto_in_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign out_back_io_enq_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign out_back_io_enq_bits_extra_tlrr_extra_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign out_back_io_enq_bits_extra_tlrr_extra_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign out_back_io_deq_ready = auto_in_d_ready & out_oready; // @[RegisterRouter.scala 82:24]
  assign PMPChecker_io_check_env_mode = 2'h3; // @[TLPMA.scala 46:28 PMP.scala 465:15]
  assign PMPChecker_io_check_env_pmp_0_cfg_l = _cfg_T[7]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_0_cfg_a = _cfg_T[4:3]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_0_cfg_x = _cfg_T[2]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_0_cfg_w = _cfg_T[1]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_0_cfg_r = _cfg_T[0]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_0_addr = addr_0; // @[PMA.scala 45:19 PMP.scala 283:15]
  assign PMPChecker_io_check_env_pmp_0_mask = mask_0; // @[PMA.scala 45:19 PMP.scala 284:15]
  assign PMPChecker_io_check_env_pmp_1_cfg_l = _cfg_T[15]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_1_cfg_a = _cfg_T[12:11]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_1_cfg_x = _cfg_T[10]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_1_cfg_w = _cfg_T[9]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_1_cfg_r = _cfg_T[8]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_1_addr = addr_1; // @[PMA.scala 45:19 PMP.scala 283:15]
  assign PMPChecker_io_check_env_pmp_1_mask = mask_1; // @[PMA.scala 45:19 PMP.scala 284:15]
  assign PMPChecker_io_check_env_pmp_2_cfg_l = _cfg_T[23]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_2_cfg_a = _cfg_T[20:19]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_2_cfg_x = _cfg_T[18]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_2_cfg_w = _cfg_T[17]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_2_cfg_r = _cfg_T[16]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_2_addr = addr_2; // @[PMA.scala 45:19 PMP.scala 283:15]
  assign PMPChecker_io_check_env_pmp_2_mask = mask_2; // @[PMA.scala 45:19 PMP.scala 284:15]
  assign PMPChecker_io_check_env_pmp_3_cfg_l = _cfg_T[31]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_3_cfg_a = _cfg_T[28:27]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_3_cfg_x = _cfg_T[26]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_3_cfg_w = _cfg_T[25]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_3_cfg_r = _cfg_T[24]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_3_addr = addr_3; // @[PMA.scala 45:19 PMP.scala 283:15]
  assign PMPChecker_io_check_env_pmp_3_mask = mask_3; // @[PMA.scala 45:19 PMP.scala 284:15]
  assign PMPChecker_io_check_env_pmp_4_cfg_l = _cfg_T[39]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_4_cfg_a = _cfg_T[36:35]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_4_cfg_x = _cfg_T[34]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_4_cfg_w = _cfg_T[33]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_4_cfg_r = _cfg_T[32]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_4_addr = addr_4; // @[PMA.scala 45:19 PMP.scala 283:15]
  assign PMPChecker_io_check_env_pmp_4_mask = mask_4; // @[PMA.scala 45:19 PMP.scala 284:15]
  assign PMPChecker_io_check_env_pmp_5_cfg_l = _cfg_T[47]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_5_cfg_a = _cfg_T[44:43]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_5_cfg_x = _cfg_T[42]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_5_cfg_w = _cfg_T[41]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_5_cfg_r = _cfg_T[40]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_5_addr = addr_5; // @[PMA.scala 45:19 PMP.scala 283:15]
  assign PMPChecker_io_check_env_pmp_5_mask = mask_5; // @[PMA.scala 45:19 PMP.scala 284:15]
  assign PMPChecker_io_check_env_pmp_6_cfg_l = _cfg_T[55]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_6_cfg_a = _cfg_T[52:51]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_6_cfg_x = _cfg_T[50]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_6_cfg_w = _cfg_T[49]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_6_cfg_r = _cfg_T[48]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_6_addr = addr_6; // @[PMA.scala 45:19 PMP.scala 283:15]
  assign PMPChecker_io_check_env_pmp_6_mask = mask_6; // @[PMA.scala 45:19 PMP.scala 284:15]
  assign PMPChecker_io_check_env_pmp_7_cfg_l = _cfg_T[63]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_7_cfg_a = _cfg_T[60:59]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_7_cfg_x = _cfg_T[58]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_7_cfg_w = _cfg_T[57]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_7_cfg_r = _cfg_T[56]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_7_addr = addr_7; // @[PMA.scala 45:19 PMP.scala 283:15]
  assign PMPChecker_io_check_env_pmp_7_mask = mask_7; // @[PMA.scala 45:19 PMP.scala 284:15]
  assign PMPChecker_io_check_env_pmp_8_cfg_l = _cfg_T[71]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_8_cfg_a = _cfg_T[68:67]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_8_cfg_x = _cfg_T[66]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_8_cfg_w = _cfg_T[65]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_8_cfg_r = _cfg_T[64]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_8_addr = addr_8; // @[PMA.scala 45:19 PMP.scala 283:15]
  assign PMPChecker_io_check_env_pmp_8_mask = mask_8; // @[PMA.scala 45:19 PMP.scala 284:15]
  assign PMPChecker_io_check_env_pmp_9_cfg_l = _cfg_T[79]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_9_cfg_a = _cfg_T[76:75]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_9_cfg_x = _cfg_T[74]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_9_cfg_w = _cfg_T[73]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_9_cfg_r = _cfg_T[72]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_9_addr = addr_9; // @[PMA.scala 45:19 PMP.scala 283:15]
  assign PMPChecker_io_check_env_pmp_9_mask = mask_9; // @[PMA.scala 45:19 PMP.scala 284:15]
  assign PMPChecker_io_check_env_pmp_10_cfg_l = _cfg_T[87]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_10_cfg_a = _cfg_T[84:83]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_10_cfg_x = _cfg_T[82]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_10_cfg_w = _cfg_T[81]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_10_cfg_r = _cfg_T[80]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_10_addr = addr_10; // @[PMA.scala 45:19 PMP.scala 283:15]
  assign PMPChecker_io_check_env_pmp_10_mask = mask_10; // @[PMA.scala 45:19 PMP.scala 284:15]
  assign PMPChecker_io_check_env_pmp_11_cfg_l = _cfg_T[95]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_11_cfg_a = _cfg_T[92:91]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_11_cfg_x = _cfg_T[90]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_11_cfg_w = _cfg_T[89]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_11_cfg_r = _cfg_T[88]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_11_addr = addr_11; // @[PMA.scala 45:19 PMP.scala 283:15]
  assign PMPChecker_io_check_env_pmp_11_mask = mask_11; // @[PMA.scala 45:19 PMP.scala 284:15]
  assign PMPChecker_io_check_env_pmp_12_cfg_l = _cfg_T[103]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_12_cfg_a = _cfg_T[100:99]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_12_cfg_x = _cfg_T[98]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_12_cfg_w = _cfg_T[97]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_12_cfg_r = _cfg_T[96]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_12_addr = addr_12; // @[PMA.scala 45:19 PMP.scala 283:15]
  assign PMPChecker_io_check_env_pmp_12_mask = mask_12; // @[PMA.scala 45:19 PMP.scala 284:15]
  assign PMPChecker_io_check_env_pmp_13_cfg_l = _cfg_T[111]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_13_cfg_a = _cfg_T[108:107]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_13_cfg_x = _cfg_T[106]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_13_cfg_w = _cfg_T[105]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_13_cfg_r = _cfg_T[104]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_13_addr = addr_13; // @[PMA.scala 45:19 PMP.scala 283:15]
  assign PMPChecker_io_check_env_pmp_13_mask = mask_13; // @[PMA.scala 45:19 PMP.scala 284:15]
  assign PMPChecker_io_check_env_pmp_14_cfg_l = _cfg_T[119]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_14_cfg_a = _cfg_T[116:115]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_14_cfg_x = _cfg_T[114]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_14_cfg_w = _cfg_T[113]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_14_cfg_r = _cfg_T[112]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_14_addr = addr_14; // @[PMA.scala 45:19 PMP.scala 283:15]
  assign PMPChecker_io_check_env_pmp_14_mask = mask_14; // @[PMA.scala 45:19 PMP.scala 284:15]
  assign PMPChecker_io_check_env_pmp_15_cfg_l = _cfg_T[127]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_15_cfg_a = _cfg_T[124:123]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_15_cfg_x = _cfg_T[122]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_15_cfg_w = _cfg_T[121]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_15_cfg_r = _cfg_T[120]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pmp_15_addr = addr_15; // @[PMA.scala 45:19 PMP.scala 283:15]
  assign PMPChecker_io_check_env_pmp_15_mask = mask_15; // @[PMA.scala 45:19 PMP.scala 284:15]
  assign PMPChecker_io_check_env_pma_0_cfg_c = _cfg_T[6]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_0_cfg_atomic = _cfg_T[5]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_0_cfg_a = _cfg_T[4:3]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_0_cfg_x = _cfg_T[2]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_0_cfg_w = _cfg_T[1]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_0_cfg_r = _cfg_T[0]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_0_addr = addr_0; // @[PMA.scala 45:19 PMP.scala 283:15]
  assign PMPChecker_io_check_env_pma_0_mask = mask_0; // @[PMA.scala 45:19 PMP.scala 284:15]
  assign PMPChecker_io_check_env_pma_1_cfg_c = _cfg_T[14]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_1_cfg_atomic = _cfg_T[13]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_1_cfg_a = _cfg_T[12:11]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_1_cfg_x = _cfg_T[10]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_1_cfg_w = _cfg_T[9]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_1_cfg_r = _cfg_T[8]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_1_addr = addr_1; // @[PMA.scala 45:19 PMP.scala 283:15]
  assign PMPChecker_io_check_env_pma_1_mask = mask_1; // @[PMA.scala 45:19 PMP.scala 284:15]
  assign PMPChecker_io_check_env_pma_2_cfg_c = _cfg_T[22]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_2_cfg_atomic = _cfg_T[21]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_2_cfg_a = _cfg_T[20:19]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_2_cfg_x = _cfg_T[18]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_2_cfg_w = _cfg_T[17]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_2_cfg_r = _cfg_T[16]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_2_addr = addr_2; // @[PMA.scala 45:19 PMP.scala 283:15]
  assign PMPChecker_io_check_env_pma_2_mask = mask_2; // @[PMA.scala 45:19 PMP.scala 284:15]
  assign PMPChecker_io_check_env_pma_3_cfg_c = _cfg_T[30]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_3_cfg_atomic = _cfg_T[29]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_3_cfg_a = _cfg_T[28:27]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_3_cfg_x = _cfg_T[26]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_3_cfg_w = _cfg_T[25]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_3_cfg_r = _cfg_T[24]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_3_addr = addr_3; // @[PMA.scala 45:19 PMP.scala 283:15]
  assign PMPChecker_io_check_env_pma_3_mask = mask_3; // @[PMA.scala 45:19 PMP.scala 284:15]
  assign PMPChecker_io_check_env_pma_4_cfg_c = _cfg_T[38]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_4_cfg_atomic = _cfg_T[37]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_4_cfg_a = _cfg_T[36:35]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_4_cfg_x = _cfg_T[34]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_4_cfg_w = _cfg_T[33]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_4_cfg_r = _cfg_T[32]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_4_addr = addr_4; // @[PMA.scala 45:19 PMP.scala 283:15]
  assign PMPChecker_io_check_env_pma_4_mask = mask_4; // @[PMA.scala 45:19 PMP.scala 284:15]
  assign PMPChecker_io_check_env_pma_5_cfg_c = _cfg_T[46]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_5_cfg_atomic = _cfg_T[45]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_5_cfg_a = _cfg_T[44:43]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_5_cfg_x = _cfg_T[42]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_5_cfg_w = _cfg_T[41]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_5_cfg_r = _cfg_T[40]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_5_addr = addr_5; // @[PMA.scala 45:19 PMP.scala 283:15]
  assign PMPChecker_io_check_env_pma_5_mask = mask_5; // @[PMA.scala 45:19 PMP.scala 284:15]
  assign PMPChecker_io_check_env_pma_6_cfg_c = _cfg_T[54]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_6_cfg_atomic = _cfg_T[53]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_6_cfg_a = _cfg_T[52:51]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_6_cfg_x = _cfg_T[50]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_6_cfg_w = _cfg_T[49]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_6_cfg_r = _cfg_T[48]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_6_addr = addr_6; // @[PMA.scala 45:19 PMP.scala 283:15]
  assign PMPChecker_io_check_env_pma_6_mask = mask_6; // @[PMA.scala 45:19 PMP.scala 284:15]
  assign PMPChecker_io_check_env_pma_7_cfg_c = _cfg_T[62]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_7_cfg_atomic = _cfg_T[61]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_7_cfg_a = _cfg_T[60:59]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_7_cfg_x = _cfg_T[58]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_7_cfg_w = _cfg_T[57]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_7_cfg_r = _cfg_T[56]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_7_addr = addr_7; // @[PMA.scala 45:19 PMP.scala 283:15]
  assign PMPChecker_io_check_env_pma_7_mask = mask_7; // @[PMA.scala 45:19 PMP.scala 284:15]
  assign PMPChecker_io_check_env_pma_8_cfg_c = _cfg_T[70]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_8_cfg_atomic = _cfg_T[69]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_8_cfg_a = _cfg_T[68:67]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_8_cfg_x = _cfg_T[66]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_8_cfg_w = _cfg_T[65]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_8_cfg_r = _cfg_T[64]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_8_addr = addr_8; // @[PMA.scala 45:19 PMP.scala 283:15]
  assign PMPChecker_io_check_env_pma_8_mask = mask_8; // @[PMA.scala 45:19 PMP.scala 284:15]
  assign PMPChecker_io_check_env_pma_9_cfg_c = _cfg_T[78]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_9_cfg_atomic = _cfg_T[77]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_9_cfg_a = _cfg_T[76:75]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_9_cfg_x = _cfg_T[74]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_9_cfg_w = _cfg_T[73]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_9_cfg_r = _cfg_T[72]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_9_addr = addr_9; // @[PMA.scala 45:19 PMP.scala 283:15]
  assign PMPChecker_io_check_env_pma_9_mask = mask_9; // @[PMA.scala 45:19 PMP.scala 284:15]
  assign PMPChecker_io_check_env_pma_10_cfg_c = _cfg_T[86]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_10_cfg_atomic = _cfg_T[85]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_10_cfg_a = _cfg_T[84:83]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_10_cfg_x = _cfg_T[82]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_10_cfg_w = _cfg_T[81]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_10_cfg_r = _cfg_T[80]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_10_addr = addr_10; // @[PMA.scala 45:19 PMP.scala 283:15]
  assign PMPChecker_io_check_env_pma_10_mask = mask_10; // @[PMA.scala 45:19 PMP.scala 284:15]
  assign PMPChecker_io_check_env_pma_11_cfg_c = _cfg_T[94]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_11_cfg_atomic = _cfg_T[93]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_11_cfg_a = _cfg_T[92:91]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_11_cfg_x = _cfg_T[90]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_11_cfg_w = _cfg_T[89]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_11_cfg_r = _cfg_T[88]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_11_addr = addr_11; // @[PMA.scala 45:19 PMP.scala 283:15]
  assign PMPChecker_io_check_env_pma_11_mask = mask_11; // @[PMA.scala 45:19 PMP.scala 284:15]
  assign PMPChecker_io_check_env_pma_12_cfg_c = _cfg_T[102]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_12_cfg_atomic = _cfg_T[101]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_12_cfg_a = _cfg_T[100:99]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_12_cfg_x = _cfg_T[98]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_12_cfg_w = _cfg_T[97]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_12_cfg_r = _cfg_T[96]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_12_addr = addr_12; // @[PMA.scala 45:19 PMP.scala 283:15]
  assign PMPChecker_io_check_env_pma_12_mask = mask_12; // @[PMA.scala 45:19 PMP.scala 284:15]
  assign PMPChecker_io_check_env_pma_13_cfg_c = _cfg_T[110]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_13_cfg_atomic = _cfg_T[109]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_13_cfg_a = _cfg_T[108:107]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_13_cfg_x = _cfg_T[106]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_13_cfg_w = _cfg_T[105]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_13_cfg_r = _cfg_T[104]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_13_addr = addr_13; // @[PMA.scala 45:19 PMP.scala 283:15]
  assign PMPChecker_io_check_env_pma_13_mask = mask_13; // @[PMA.scala 45:19 PMP.scala 284:15]
  assign PMPChecker_io_check_env_pma_14_cfg_c = _cfg_T[118]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_14_cfg_atomic = _cfg_T[117]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_14_cfg_a = _cfg_T[116:115]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_14_cfg_x = _cfg_T[114]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_14_cfg_w = _cfg_T[113]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_14_cfg_r = _cfg_T[112]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_14_addr = addr_14; // @[PMA.scala 45:19 PMP.scala 283:15]
  assign PMPChecker_io_check_env_pma_14_mask = mask_14; // @[PMA.scala 45:19 PMP.scala 284:15]
  assign PMPChecker_io_check_env_pma_15_cfg_c = _cfg_T[126]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_15_cfg_atomic = _cfg_T[125]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_15_cfg_a = _cfg_T[124:123]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_15_cfg_x = _cfg_T[122]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_15_cfg_w = _cfg_T[121]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_15_cfg_r = _cfg_T[120]; // @[PMA.scala 53:46]
  assign PMPChecker_io_check_env_pma_15_addr = addr_15; // @[PMA.scala 45:19 PMP.scala 283:15]
  assign PMPChecker_io_check_env_pma_15_mask = mask_15; // @[PMA.scala 45:19 PMP.scala 284:15]
  assign PMPChecker_io_req_bits_addr = io_req_0_bits_addr; // @[PMP.scala 373:15 TLPMA.scala 46:28]
  assign PMPChecker_io_req_bits_cmd = 3'h0; // @[PMP.scala 375:14 TLPMA.scala 46:28]
  assign PMPChecker_1_io_check_env_mode = 2'h3; // @[TLPMA.scala 46:28 PMP.scala 465:15]
  assign PMPChecker_1_io_check_env_pmp_0_cfg_l = _cfg_T[7]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_0_cfg_a = _cfg_T[4:3]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_0_cfg_x = _cfg_T[2]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_0_cfg_w = _cfg_T[1]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_0_cfg_r = _cfg_T[0]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_0_addr = addr_0; // @[PMA.scala 45:19 PMP.scala 283:15]
  assign PMPChecker_1_io_check_env_pmp_0_mask = mask_0; // @[PMA.scala 45:19 PMP.scala 284:15]
  assign PMPChecker_1_io_check_env_pmp_1_cfg_l = _cfg_T[15]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_1_cfg_a = _cfg_T[12:11]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_1_cfg_x = _cfg_T[10]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_1_cfg_w = _cfg_T[9]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_1_cfg_r = _cfg_T[8]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_1_addr = addr_1; // @[PMA.scala 45:19 PMP.scala 283:15]
  assign PMPChecker_1_io_check_env_pmp_1_mask = mask_1; // @[PMA.scala 45:19 PMP.scala 284:15]
  assign PMPChecker_1_io_check_env_pmp_2_cfg_l = _cfg_T[23]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_2_cfg_a = _cfg_T[20:19]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_2_cfg_x = _cfg_T[18]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_2_cfg_w = _cfg_T[17]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_2_cfg_r = _cfg_T[16]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_2_addr = addr_2; // @[PMA.scala 45:19 PMP.scala 283:15]
  assign PMPChecker_1_io_check_env_pmp_2_mask = mask_2; // @[PMA.scala 45:19 PMP.scala 284:15]
  assign PMPChecker_1_io_check_env_pmp_3_cfg_l = _cfg_T[31]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_3_cfg_a = _cfg_T[28:27]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_3_cfg_x = _cfg_T[26]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_3_cfg_w = _cfg_T[25]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_3_cfg_r = _cfg_T[24]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_3_addr = addr_3; // @[PMA.scala 45:19 PMP.scala 283:15]
  assign PMPChecker_1_io_check_env_pmp_3_mask = mask_3; // @[PMA.scala 45:19 PMP.scala 284:15]
  assign PMPChecker_1_io_check_env_pmp_4_cfg_l = _cfg_T[39]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_4_cfg_a = _cfg_T[36:35]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_4_cfg_x = _cfg_T[34]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_4_cfg_w = _cfg_T[33]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_4_cfg_r = _cfg_T[32]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_4_addr = addr_4; // @[PMA.scala 45:19 PMP.scala 283:15]
  assign PMPChecker_1_io_check_env_pmp_4_mask = mask_4; // @[PMA.scala 45:19 PMP.scala 284:15]
  assign PMPChecker_1_io_check_env_pmp_5_cfg_l = _cfg_T[47]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_5_cfg_a = _cfg_T[44:43]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_5_cfg_x = _cfg_T[42]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_5_cfg_w = _cfg_T[41]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_5_cfg_r = _cfg_T[40]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_5_addr = addr_5; // @[PMA.scala 45:19 PMP.scala 283:15]
  assign PMPChecker_1_io_check_env_pmp_5_mask = mask_5; // @[PMA.scala 45:19 PMP.scala 284:15]
  assign PMPChecker_1_io_check_env_pmp_6_cfg_l = _cfg_T[55]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_6_cfg_a = _cfg_T[52:51]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_6_cfg_x = _cfg_T[50]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_6_cfg_w = _cfg_T[49]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_6_cfg_r = _cfg_T[48]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_6_addr = addr_6; // @[PMA.scala 45:19 PMP.scala 283:15]
  assign PMPChecker_1_io_check_env_pmp_6_mask = mask_6; // @[PMA.scala 45:19 PMP.scala 284:15]
  assign PMPChecker_1_io_check_env_pmp_7_cfg_l = _cfg_T[63]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_7_cfg_a = _cfg_T[60:59]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_7_cfg_x = _cfg_T[58]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_7_cfg_w = _cfg_T[57]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_7_cfg_r = _cfg_T[56]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_7_addr = addr_7; // @[PMA.scala 45:19 PMP.scala 283:15]
  assign PMPChecker_1_io_check_env_pmp_7_mask = mask_7; // @[PMA.scala 45:19 PMP.scala 284:15]
  assign PMPChecker_1_io_check_env_pmp_8_cfg_l = _cfg_T[71]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_8_cfg_a = _cfg_T[68:67]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_8_cfg_x = _cfg_T[66]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_8_cfg_w = _cfg_T[65]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_8_cfg_r = _cfg_T[64]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_8_addr = addr_8; // @[PMA.scala 45:19 PMP.scala 283:15]
  assign PMPChecker_1_io_check_env_pmp_8_mask = mask_8; // @[PMA.scala 45:19 PMP.scala 284:15]
  assign PMPChecker_1_io_check_env_pmp_9_cfg_l = _cfg_T[79]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_9_cfg_a = _cfg_T[76:75]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_9_cfg_x = _cfg_T[74]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_9_cfg_w = _cfg_T[73]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_9_cfg_r = _cfg_T[72]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_9_addr = addr_9; // @[PMA.scala 45:19 PMP.scala 283:15]
  assign PMPChecker_1_io_check_env_pmp_9_mask = mask_9; // @[PMA.scala 45:19 PMP.scala 284:15]
  assign PMPChecker_1_io_check_env_pmp_10_cfg_l = _cfg_T[87]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_10_cfg_a = _cfg_T[84:83]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_10_cfg_x = _cfg_T[82]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_10_cfg_w = _cfg_T[81]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_10_cfg_r = _cfg_T[80]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_10_addr = addr_10; // @[PMA.scala 45:19 PMP.scala 283:15]
  assign PMPChecker_1_io_check_env_pmp_10_mask = mask_10; // @[PMA.scala 45:19 PMP.scala 284:15]
  assign PMPChecker_1_io_check_env_pmp_11_cfg_l = _cfg_T[95]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_11_cfg_a = _cfg_T[92:91]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_11_cfg_x = _cfg_T[90]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_11_cfg_w = _cfg_T[89]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_11_cfg_r = _cfg_T[88]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_11_addr = addr_11; // @[PMA.scala 45:19 PMP.scala 283:15]
  assign PMPChecker_1_io_check_env_pmp_11_mask = mask_11; // @[PMA.scala 45:19 PMP.scala 284:15]
  assign PMPChecker_1_io_check_env_pmp_12_cfg_l = _cfg_T[103]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_12_cfg_a = _cfg_T[100:99]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_12_cfg_x = _cfg_T[98]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_12_cfg_w = _cfg_T[97]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_12_cfg_r = _cfg_T[96]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_12_addr = addr_12; // @[PMA.scala 45:19 PMP.scala 283:15]
  assign PMPChecker_1_io_check_env_pmp_12_mask = mask_12; // @[PMA.scala 45:19 PMP.scala 284:15]
  assign PMPChecker_1_io_check_env_pmp_13_cfg_l = _cfg_T[111]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_13_cfg_a = _cfg_T[108:107]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_13_cfg_x = _cfg_T[106]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_13_cfg_w = _cfg_T[105]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_13_cfg_r = _cfg_T[104]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_13_addr = addr_13; // @[PMA.scala 45:19 PMP.scala 283:15]
  assign PMPChecker_1_io_check_env_pmp_13_mask = mask_13; // @[PMA.scala 45:19 PMP.scala 284:15]
  assign PMPChecker_1_io_check_env_pmp_14_cfg_l = _cfg_T[119]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_14_cfg_a = _cfg_T[116:115]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_14_cfg_x = _cfg_T[114]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_14_cfg_w = _cfg_T[113]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_14_cfg_r = _cfg_T[112]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_14_addr = addr_14; // @[PMA.scala 45:19 PMP.scala 283:15]
  assign PMPChecker_1_io_check_env_pmp_14_mask = mask_14; // @[PMA.scala 45:19 PMP.scala 284:15]
  assign PMPChecker_1_io_check_env_pmp_15_cfg_l = _cfg_T[127]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_15_cfg_a = _cfg_T[124:123]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_15_cfg_x = _cfg_T[122]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_15_cfg_w = _cfg_T[121]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_15_cfg_r = _cfg_T[120]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pmp_15_addr = addr_15; // @[PMA.scala 45:19 PMP.scala 283:15]
  assign PMPChecker_1_io_check_env_pmp_15_mask = mask_15; // @[PMA.scala 45:19 PMP.scala 284:15]
  assign PMPChecker_1_io_check_env_pma_0_cfg_c = _cfg_T[6]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_0_cfg_atomic = _cfg_T[5]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_0_cfg_a = _cfg_T[4:3]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_0_cfg_x = _cfg_T[2]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_0_cfg_w = _cfg_T[1]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_0_cfg_r = _cfg_T[0]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_0_addr = addr_0; // @[PMA.scala 45:19 PMP.scala 283:15]
  assign PMPChecker_1_io_check_env_pma_0_mask = mask_0; // @[PMA.scala 45:19 PMP.scala 284:15]
  assign PMPChecker_1_io_check_env_pma_1_cfg_c = _cfg_T[14]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_1_cfg_atomic = _cfg_T[13]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_1_cfg_a = _cfg_T[12:11]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_1_cfg_x = _cfg_T[10]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_1_cfg_w = _cfg_T[9]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_1_cfg_r = _cfg_T[8]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_1_addr = addr_1; // @[PMA.scala 45:19 PMP.scala 283:15]
  assign PMPChecker_1_io_check_env_pma_1_mask = mask_1; // @[PMA.scala 45:19 PMP.scala 284:15]
  assign PMPChecker_1_io_check_env_pma_2_cfg_c = _cfg_T[22]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_2_cfg_atomic = _cfg_T[21]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_2_cfg_a = _cfg_T[20:19]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_2_cfg_x = _cfg_T[18]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_2_cfg_w = _cfg_T[17]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_2_cfg_r = _cfg_T[16]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_2_addr = addr_2; // @[PMA.scala 45:19 PMP.scala 283:15]
  assign PMPChecker_1_io_check_env_pma_2_mask = mask_2; // @[PMA.scala 45:19 PMP.scala 284:15]
  assign PMPChecker_1_io_check_env_pma_3_cfg_c = _cfg_T[30]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_3_cfg_atomic = _cfg_T[29]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_3_cfg_a = _cfg_T[28:27]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_3_cfg_x = _cfg_T[26]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_3_cfg_w = _cfg_T[25]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_3_cfg_r = _cfg_T[24]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_3_addr = addr_3; // @[PMA.scala 45:19 PMP.scala 283:15]
  assign PMPChecker_1_io_check_env_pma_3_mask = mask_3; // @[PMA.scala 45:19 PMP.scala 284:15]
  assign PMPChecker_1_io_check_env_pma_4_cfg_c = _cfg_T[38]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_4_cfg_atomic = _cfg_T[37]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_4_cfg_a = _cfg_T[36:35]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_4_cfg_x = _cfg_T[34]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_4_cfg_w = _cfg_T[33]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_4_cfg_r = _cfg_T[32]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_4_addr = addr_4; // @[PMA.scala 45:19 PMP.scala 283:15]
  assign PMPChecker_1_io_check_env_pma_4_mask = mask_4; // @[PMA.scala 45:19 PMP.scala 284:15]
  assign PMPChecker_1_io_check_env_pma_5_cfg_c = _cfg_T[46]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_5_cfg_atomic = _cfg_T[45]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_5_cfg_a = _cfg_T[44:43]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_5_cfg_x = _cfg_T[42]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_5_cfg_w = _cfg_T[41]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_5_cfg_r = _cfg_T[40]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_5_addr = addr_5; // @[PMA.scala 45:19 PMP.scala 283:15]
  assign PMPChecker_1_io_check_env_pma_5_mask = mask_5; // @[PMA.scala 45:19 PMP.scala 284:15]
  assign PMPChecker_1_io_check_env_pma_6_cfg_c = _cfg_T[54]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_6_cfg_atomic = _cfg_T[53]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_6_cfg_a = _cfg_T[52:51]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_6_cfg_x = _cfg_T[50]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_6_cfg_w = _cfg_T[49]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_6_cfg_r = _cfg_T[48]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_6_addr = addr_6; // @[PMA.scala 45:19 PMP.scala 283:15]
  assign PMPChecker_1_io_check_env_pma_6_mask = mask_6; // @[PMA.scala 45:19 PMP.scala 284:15]
  assign PMPChecker_1_io_check_env_pma_7_cfg_c = _cfg_T[62]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_7_cfg_atomic = _cfg_T[61]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_7_cfg_a = _cfg_T[60:59]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_7_cfg_x = _cfg_T[58]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_7_cfg_w = _cfg_T[57]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_7_cfg_r = _cfg_T[56]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_7_addr = addr_7; // @[PMA.scala 45:19 PMP.scala 283:15]
  assign PMPChecker_1_io_check_env_pma_7_mask = mask_7; // @[PMA.scala 45:19 PMP.scala 284:15]
  assign PMPChecker_1_io_check_env_pma_8_cfg_c = _cfg_T[70]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_8_cfg_atomic = _cfg_T[69]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_8_cfg_a = _cfg_T[68:67]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_8_cfg_x = _cfg_T[66]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_8_cfg_w = _cfg_T[65]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_8_cfg_r = _cfg_T[64]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_8_addr = addr_8; // @[PMA.scala 45:19 PMP.scala 283:15]
  assign PMPChecker_1_io_check_env_pma_8_mask = mask_8; // @[PMA.scala 45:19 PMP.scala 284:15]
  assign PMPChecker_1_io_check_env_pma_9_cfg_c = _cfg_T[78]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_9_cfg_atomic = _cfg_T[77]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_9_cfg_a = _cfg_T[76:75]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_9_cfg_x = _cfg_T[74]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_9_cfg_w = _cfg_T[73]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_9_cfg_r = _cfg_T[72]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_9_addr = addr_9; // @[PMA.scala 45:19 PMP.scala 283:15]
  assign PMPChecker_1_io_check_env_pma_9_mask = mask_9; // @[PMA.scala 45:19 PMP.scala 284:15]
  assign PMPChecker_1_io_check_env_pma_10_cfg_c = _cfg_T[86]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_10_cfg_atomic = _cfg_T[85]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_10_cfg_a = _cfg_T[84:83]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_10_cfg_x = _cfg_T[82]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_10_cfg_w = _cfg_T[81]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_10_cfg_r = _cfg_T[80]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_10_addr = addr_10; // @[PMA.scala 45:19 PMP.scala 283:15]
  assign PMPChecker_1_io_check_env_pma_10_mask = mask_10; // @[PMA.scala 45:19 PMP.scala 284:15]
  assign PMPChecker_1_io_check_env_pma_11_cfg_c = _cfg_T[94]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_11_cfg_atomic = _cfg_T[93]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_11_cfg_a = _cfg_T[92:91]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_11_cfg_x = _cfg_T[90]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_11_cfg_w = _cfg_T[89]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_11_cfg_r = _cfg_T[88]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_11_addr = addr_11; // @[PMA.scala 45:19 PMP.scala 283:15]
  assign PMPChecker_1_io_check_env_pma_11_mask = mask_11; // @[PMA.scala 45:19 PMP.scala 284:15]
  assign PMPChecker_1_io_check_env_pma_12_cfg_c = _cfg_T[102]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_12_cfg_atomic = _cfg_T[101]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_12_cfg_a = _cfg_T[100:99]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_12_cfg_x = _cfg_T[98]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_12_cfg_w = _cfg_T[97]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_12_cfg_r = _cfg_T[96]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_12_addr = addr_12; // @[PMA.scala 45:19 PMP.scala 283:15]
  assign PMPChecker_1_io_check_env_pma_12_mask = mask_12; // @[PMA.scala 45:19 PMP.scala 284:15]
  assign PMPChecker_1_io_check_env_pma_13_cfg_c = _cfg_T[110]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_13_cfg_atomic = _cfg_T[109]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_13_cfg_a = _cfg_T[108:107]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_13_cfg_x = _cfg_T[106]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_13_cfg_w = _cfg_T[105]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_13_cfg_r = _cfg_T[104]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_13_addr = addr_13; // @[PMA.scala 45:19 PMP.scala 283:15]
  assign PMPChecker_1_io_check_env_pma_13_mask = mask_13; // @[PMA.scala 45:19 PMP.scala 284:15]
  assign PMPChecker_1_io_check_env_pma_14_cfg_c = _cfg_T[118]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_14_cfg_atomic = _cfg_T[117]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_14_cfg_a = _cfg_T[116:115]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_14_cfg_x = _cfg_T[114]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_14_cfg_w = _cfg_T[113]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_14_cfg_r = _cfg_T[112]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_14_addr = addr_14; // @[PMA.scala 45:19 PMP.scala 283:15]
  assign PMPChecker_1_io_check_env_pma_14_mask = mask_14; // @[PMA.scala 45:19 PMP.scala 284:15]
  assign PMPChecker_1_io_check_env_pma_15_cfg_c = _cfg_T[126]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_15_cfg_atomic = _cfg_T[125]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_15_cfg_a = _cfg_T[124:123]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_15_cfg_x = _cfg_T[122]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_15_cfg_w = _cfg_T[121]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_15_cfg_r = _cfg_T[120]; // @[PMA.scala 53:46]
  assign PMPChecker_1_io_check_env_pma_15_addr = addr_15; // @[PMA.scala 45:19 PMP.scala 283:15]
  assign PMPChecker_1_io_check_env_pma_15_mask = mask_15; // @[PMA.scala 45:19 PMP.scala 284:15]
  assign PMPChecker_1_io_req_bits_addr = io_req_1_bits_addr; // @[PMP.scala 373:15 TLPMA.scala 46:28]
  assign PMPChecker_1_io_req_bits_cmd = 3'h0; // @[PMP.scala 375:14 TLPMA.scala 46:28]
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PMA.scala 73:38]
      pmaCfgMerged_0 <= 64'hf0b0b0b0f0b0000; // @[PMA.scala 73:69]
    end else if (out_f_woready) begin // @[PMA.scala 50:31]
      pmaCfgMerged_0 <= _out_pmaCfgMerged_0_T_16;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PMA.scala 73:38]
      pmaCfgMerged_1 <= 64'h7f1b080b080b080b; // @[PMA.scala 73:69]
    end else if (out_f_woready_8) begin // @[PMA.scala 50:31]
      pmaCfgMerged_1 <= _out_pmaCfgMerged_0_T_16;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PMA.scala 84:24]
      addr_0 <= 34'h0; // @[PMP.scala 121:8]
    end else if (out_f_woready_9) begin // @[PMA.scala 51:23]
      if (_out_addr_0_mask_0_T) begin
        addr_0 <= _out_T_40[33:0];
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PMA.scala 84:24]
      addr_1 <= 34'h0; // @[PMP.scala 121:8]
    end else if (out_f_woready_6) begin // @[PMA.scala 51:23]
      if (_out_addr_1_mask_1_T) begin
        addr_1 <= _out_T_40[33:0];
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PMA.scala 84:24]
      addr_2 <= 34'h4000000; // @[PMP.scala 121:8]
    end else if (out_f_woready_10) begin // @[PMA.scala 51:23]
      if (_out_addr_2_mask_2_T) begin
        addr_2 <= _out_T_40[33:0];
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PMA.scala 84:24]
      addr_3 <= 34'h8000000; // @[PMP.scala 121:8]
    end else if (out_f_woready_15) begin // @[PMA.scala 51:23]
      if (_out_addr_3_mask_3_T) begin
        addr_3 <= _out_T_40[33:0];
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PMA.scala 84:24]
      addr_4 <= 34'hc004000; // @[PMP.scala 121:8]
    end else if (out_f_woready_18) begin // @[PMA.scala 51:23]
      if (_out_addr_4_mask_4_T) begin
        addr_4 <= _out_T_40[33:0];
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PMA.scala 84:24]
      addr_5 <= 34'hc014000; // @[PMP.scala 121:8]
    end else if (out_f_woready_2) begin // @[PMA.scala 51:23]
      if (_out_addr_5_mask_5_T) begin
        addr_5 <= _out_T_40[33:0];
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PMA.scala 84:24]
      addr_6 <= 34'he008000; // @[PMP.scala 121:8]
    end else if (out_f_woready_5) begin // @[PMA.scala 51:23]
      if (_out_addr_6_mask_6_T) begin
        addr_6 <= _out_T_40[33:0];
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PMA.scala 84:24]
      addr_7 <= 34'he008400; // @[PMP.scala 121:8]
    end else if (out_f_woready_13) begin // @[PMA.scala 51:23]
      if (_out_addr_7_mask_7_T) begin
        addr_7 <= _out_T_40[33:0];
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PMA.scala 84:24]
      addr_8 <= 34'he008800; // @[PMP.scala 121:8]
    end else if (out_f_woready_17) begin // @[PMA.scala 51:23]
      if (_out_addr_8_mask_8_T) begin
        addr_8 <= _out_T_40[33:0];
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PMA.scala 84:24]
      addr_9 <= 34'he400000; // @[PMP.scala 121:8]
    end else if (out_f_woready_7) begin // @[PMA.scala 51:23]
      if (_out_addr_9_mask_9_T) begin
        addr_9 <= _out_T_40[33:0];
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PMA.scala 84:24]
      addr_10 <= 34'he400800; // @[PMP.scala 121:8]
    end else if (out_f_woready_1) begin // @[PMA.scala 51:23]
      if (_out_addr_10_mask_10_T) begin
        addr_10 <= _out_T_40[33:0];
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PMA.scala 84:24]
      addr_11 <= 34'he800000; // @[PMP.scala 121:8]
    end else if (out_f_woready_16) begin // @[PMA.scala 51:23]
      if (_out_addr_11_mask_11_T) begin
        addr_11 <= _out_T_40[33:0];
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PMA.scala 84:24]
      addr_12 <= 34'he800400; // @[PMP.scala 121:8]
    end else if (out_f_woready_12) begin // @[PMA.scala 51:23]
      if (_out_addr_12_mask_12_T) begin
        addr_12 <= _out_T_40[33:0];
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PMA.scala 84:24]
      addr_13 <= 34'hf000000; // @[PMP.scala 121:8]
    end else if (out_f_woready_11) begin // @[PMA.scala 51:23]
      if (_out_addr_13_mask_13_T) begin
        addr_13 <= _out_T_40[33:0];
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PMA.scala 84:24]
      addr_14 <= 34'hfffffff; // @[PMP.scala 121:8]
    end else if (out_f_woready_3) begin // @[PMA.scala 51:23]
      if (_out_addr_14_mask_14_T) begin
        addr_14 <= _out_T_40[33:0];
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PMA.scala 84:24]
      addr_15 <= 34'h1ffffffff; // @[PMP.scala 121:8]
    end else if (out_f_woready_19) begin // @[PMA.scala 51:23]
      if (_out_addr_15_mask_15_T) begin
        addr_15 <= _out_T_40[33:0];
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PMA.scala 52:23]
      mask_0 <= 36'hfff; // @[PMA.scala 52:23]
    end else begin
      mask_0 <= _GEN_103[35:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PMA.scala 52:23]
      mask_1 <= 36'hfff; // @[PMA.scala 52:23]
    end else begin
      mask_1 <= _GEN_55[35:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PMA.scala 52:23]
      mask_2 <= 36'hfff; // @[PMA.scala 52:23]
    end else begin
      mask_2 <= _GEN_105[35:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PMA.scala 52:23]
      mask_3 <= 36'hfff; // @[PMA.scala 52:23]
    end else begin
      mask_3 <= _GEN_116[35:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PMA.scala 52:23]
      mask_4 <= 36'hfff; // @[PMA.scala 52:23]
    end else begin
      mask_4 <= _GEN_122[35:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PMA.scala 52:23]
      mask_5 <= 36'hfff; // @[PMA.scala 52:23]
    end else begin
      mask_5 <= _GEN_46[35:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PMA.scala 52:23]
      mask_6 <= 36'hfff; // @[PMA.scala 52:23]
    end else begin
      mask_6 <= _GEN_53[35:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PMA.scala 52:23]
      mask_7 <= 36'hfff; // @[PMA.scala 52:23]
    end else begin
      mask_7 <= _GEN_111[35:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PMA.scala 52:23]
      mask_8 <= 36'hfff; // @[PMA.scala 52:23]
    end else begin
      mask_8 <= _GEN_120[35:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PMA.scala 52:23]
      mask_9 <= 36'hfff; // @[PMA.scala 52:23]
    end else begin
      mask_9 <= _GEN_95[35:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PMA.scala 52:23]
      mask_10 <= 36'hfff; // @[PMA.scala 52:23]
    end else begin
      mask_10 <= _GEN_96[35:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PMA.scala 52:23]
      mask_11 <= 36'hfff; // @[PMA.scala 52:23]
    end else begin
      mask_11 <= _GEN_118[35:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PMA.scala 52:23]
      mask_12 <= 36'hfff; // @[PMA.scala 52:23]
    end else begin
      mask_12 <= _GEN_109[35:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PMA.scala 52:23]
      mask_13 <= 36'hfff; // @[PMA.scala 52:23]
    end else begin
      mask_13 <= _GEN_107[35:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PMA.scala 52:23]
      mask_14 <= 36'h7fffffff; // @[PMA.scala 52:23]
    end else begin
      mask_14 <= _GEN_100[35:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PMA.scala 52:23]
      mask_15 <= 36'hfffffffff; // @[PMA.scala 52:23]
    end else begin
      mask_15 <= _GEN_124[35:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Hold.scala 42:19]
      out_v_reg <= 1'h0; // @[Hold.scala 42:27]
    end else begin
      out_v_reg <= _out_v_reg_T | _GEN_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Hold.scala 42:19]
      out_v_reg_1 <= 1'h0; // @[Hold.scala 42:27]
    end else begin
      out_v_reg_1 <= _out_v_reg_T_2 | _GEN_50;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Hold.scala 42:19]
      out_v_reg_2 <= 1'h0; // @[Hold.scala 42:27]
    end else begin
      out_v_reg_2 <= _out_v_reg_T_4 | _GEN_59;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Hold.scala 42:19]
      out_v_reg_3 <= 1'h0; // @[Hold.scala 42:27]
    end else begin
      out_v_reg_3 <= _out_v_reg_T_6 | _GEN_113;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  pmaCfgMerged_0 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  pmaCfgMerged_1 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  addr_0 = _RAND_2[33:0];
  _RAND_3 = {2{`RANDOM}};
  addr_1 = _RAND_3[33:0];
  _RAND_4 = {2{`RANDOM}};
  addr_2 = _RAND_4[33:0];
  _RAND_5 = {2{`RANDOM}};
  addr_3 = _RAND_5[33:0];
  _RAND_6 = {2{`RANDOM}};
  addr_4 = _RAND_6[33:0];
  _RAND_7 = {2{`RANDOM}};
  addr_5 = _RAND_7[33:0];
  _RAND_8 = {2{`RANDOM}};
  addr_6 = _RAND_8[33:0];
  _RAND_9 = {2{`RANDOM}};
  addr_7 = _RAND_9[33:0];
  _RAND_10 = {2{`RANDOM}};
  addr_8 = _RAND_10[33:0];
  _RAND_11 = {2{`RANDOM}};
  addr_9 = _RAND_11[33:0];
  _RAND_12 = {2{`RANDOM}};
  addr_10 = _RAND_12[33:0];
  _RAND_13 = {2{`RANDOM}};
  addr_11 = _RAND_13[33:0];
  _RAND_14 = {2{`RANDOM}};
  addr_12 = _RAND_14[33:0];
  _RAND_15 = {2{`RANDOM}};
  addr_13 = _RAND_15[33:0];
  _RAND_16 = {2{`RANDOM}};
  addr_14 = _RAND_16[33:0];
  _RAND_17 = {2{`RANDOM}};
  addr_15 = _RAND_17[33:0];
  _RAND_18 = {2{`RANDOM}};
  mask_0 = _RAND_18[35:0];
  _RAND_19 = {2{`RANDOM}};
  mask_1 = _RAND_19[35:0];
  _RAND_20 = {2{`RANDOM}};
  mask_2 = _RAND_20[35:0];
  _RAND_21 = {2{`RANDOM}};
  mask_3 = _RAND_21[35:0];
  _RAND_22 = {2{`RANDOM}};
  mask_4 = _RAND_22[35:0];
  _RAND_23 = {2{`RANDOM}};
  mask_5 = _RAND_23[35:0];
  _RAND_24 = {2{`RANDOM}};
  mask_6 = _RAND_24[35:0];
  _RAND_25 = {2{`RANDOM}};
  mask_7 = _RAND_25[35:0];
  _RAND_26 = {2{`RANDOM}};
  mask_8 = _RAND_26[35:0];
  _RAND_27 = {2{`RANDOM}};
  mask_9 = _RAND_27[35:0];
  _RAND_28 = {2{`RANDOM}};
  mask_10 = _RAND_28[35:0];
  _RAND_29 = {2{`RANDOM}};
  mask_11 = _RAND_29[35:0];
  _RAND_30 = {2{`RANDOM}};
  mask_12 = _RAND_30[35:0];
  _RAND_31 = {2{`RANDOM}};
  mask_13 = _RAND_31[35:0];
  _RAND_32 = {2{`RANDOM}};
  mask_14 = _RAND_32[35:0];
  _RAND_33 = {2{`RANDOM}};
  mask_15 = _RAND_33[35:0];
  _RAND_34 = {1{`RANDOM}};
  out_v_reg = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  out_v_reg_1 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  out_v_reg_2 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  out_v_reg_3 = _RAND_37[0:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    pmaCfgMerged_0 = 64'hf0b0b0b0f0b0000;
  end
  if (reset) begin
    pmaCfgMerged_1 = 64'h7f1b080b080b080b;
  end
  if (reset) begin
    addr_0 = 34'h0;
  end
  if (reset) begin
    addr_1 = 34'h0;
  end
  if (reset) begin
    addr_2 = 34'h4000000;
  end
  if (reset) begin
    addr_3 = 34'h8000000;
  end
  if (reset) begin
    addr_4 = 34'hc004000;
  end
  if (reset) begin
    addr_5 = 34'hc014000;
  end
  if (reset) begin
    addr_6 = 34'he008000;
  end
  if (reset) begin
    addr_7 = 34'he008400;
  end
  if (reset) begin
    addr_8 = 34'he008800;
  end
  if (reset) begin
    addr_9 = 34'he400000;
  end
  if (reset) begin
    addr_10 = 34'he400800;
  end
  if (reset) begin
    addr_11 = 34'he800000;
  end
  if (reset) begin
    addr_12 = 34'he800400;
  end
  if (reset) begin
    addr_13 = 34'hf000000;
  end
  if (reset) begin
    addr_14 = 34'hfffffff;
  end
  if (reset) begin
    addr_15 = 34'h1ffffffff;
  end
  if (reset) begin
    mask_0 = 36'hfff;
  end
  if (reset) begin
    mask_1 = 36'hfff;
  end
  if (reset) begin
    mask_2 = 36'hfff;
  end
  if (reset) begin
    mask_3 = 36'hfff;
  end
  if (reset) begin
    mask_4 = 36'hfff;
  end
  if (reset) begin
    mask_5 = 36'hfff;
  end
  if (reset) begin
    mask_6 = 36'hfff;
  end
  if (reset) begin
    mask_7 = 36'hfff;
  end
  if (reset) begin
    mask_8 = 36'hfff;
  end
  if (reset) begin
    mask_9 = 36'hfff;
  end
  if (reset) begin
    mask_10 = 36'hfff;
  end
  if (reset) begin
    mask_11 = 36'hfff;
  end
  if (reset) begin
    mask_12 = 36'hfff;
  end
  if (reset) begin
    mask_13 = 36'hfff;
  end
  if (reset) begin
    mask_14 = 36'h7fffffff;
  end
  if (reset) begin
    mask_15 = 36'hfffffffff;
  end
  if (reset) begin
    out_v_reg = 1'h0;
  end
  if (reset) begin
    out_v_reg_1 = 1'h0;
  end
  if (reset) begin
    out_v_reg_2 = 1'h0;
  end
  if (reset) begin
    out_v_reg_3 = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule

