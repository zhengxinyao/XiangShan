module PtwCache(
  input          clock,
  input          reset,
  output         io_req_ready,
  input          io_req_valid,
  input  [26:0]  io_req_bits_req_info_vpn,
  input  [1:0]   io_req_bits_req_info_source,
  input          io_req_bits_isFirst,
  input          io_resp_ready,
  output         io_resp_valid,
  output [26:0]  io_resp_bits_req_info_vpn,
  output [1:0]   io_resp_bits_req_info_source,
  output         io_resp_bits_isFirst,
  output         io_resp_bits_hit,
  output         io_resp_bits_prefetch,
  output         io_resp_bits_bypassed,
  output         io_resp_bits_toFsm_l1Hit,
  output         io_resp_bits_toFsm_l2Hit,
  output [23:0]  io_resp_bits_toFsm_ppn,
  output [26:0]  io_resp_bits_toTlb_tag,
  output [15:0]  io_resp_bits_toTlb_asid,
  output [23:0]  io_resp_bits_toTlb_ppn,
  output         io_resp_bits_toTlb_perm_d,
  output         io_resp_bits_toTlb_perm_a,
  output         io_resp_bits_toTlb_perm_g,
  output         io_resp_bits_toTlb_perm_u,
  output         io_resp_bits_toTlb_perm_x,
  output         io_resp_bits_toTlb_perm_w,
  output         io_resp_bits_toTlb_perm_r,
  output [1:0]   io_resp_bits_toTlb_level,
  output         io_resp_bits_toTlb_prefetch,
  output         io_resp_bits_toTlb_v,
  input          io_refill_valid,
  input  [511:0] io_refill_bits_ptes,
  input          io_refill_bits_levelOH_sp,
  input          io_refill_bits_levelOH_l3,
  input          io_refill_bits_levelOH_l2,
  input          io_refill_bits_levelOH_l1,
  input  [26:0]  io_refill_bits_req_info_dup_0_vpn,
  input  [1:0]   io_refill_bits_req_info_dup_0_source,
  input  [26:0]  io_refill_bits_req_info_dup_1_vpn,
  input  [1:0]   io_refill_bits_req_info_dup_1_source,
  input  [26:0]  io_refill_bits_req_info_dup_2_vpn,
  input  [1:0]   io_refill_bits_req_info_dup_2_source,
  input  [1:0]   io_refill_bits_level_dup_0,
  input  [1:0]   io_refill_bits_level_dup_1,
  input  [1:0]   io_refill_bits_level_dup_2,
  input  [63:0]  io_refill_bits_sel_pte_dup_0,
  input  [63:0]  io_refill_bits_sel_pte_dup_1,
  input  [63:0]  io_refill_bits_sel_pte_dup_2,
  input          io_sfence_dup_0_valid,
  input          io_sfence_dup_0_bits_rs1,
  input          io_sfence_dup_0_bits_rs2,
  input  [38:0]  io_sfence_dup_0_bits_addr,
  input  [15:0]  io_sfence_dup_0_bits_asid,
  input          io_sfence_dup_1_valid,
  input          io_sfence_dup_2_valid,
  input          io_sfence_dup_3_valid,
  input          io_sfence_dup_3_bits_rs1,
  input          io_sfence_dup_3_bits_rs2,
  input  [38:0]  io_sfence_dup_3_bits_addr,
  input  [15:0]  io_csr_dup_0_satp_asid,
  input          io_csr_dup_0_satp_changed,
  input  [15:0]  io_csr_dup_1_satp_asid,
  input          io_csr_dup_1_satp_changed,
  input  [15:0]  io_csr_dup_2_satp_asid,
  input          io_csr_dup_2_satp_changed,
  output [5:0]   io_perf_0_value,
  output [5:0]   io_perf_1_value,
  output [5:0]   io_perf_2_value,
  output [5:0]   io_perf_3_value,
  output [5:0]   io_perf_4_value,
  output [5:0]   io_perf_5_value,
  output [5:0]   io_perf_6_value,
  output [5:0]   io_perf_7_value
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [63:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [63:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [63:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [63:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [63:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [63:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_786;
  reg [63:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_789;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_793;
  reg [31:0] _RAND_794;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [31:0] _RAND_798;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_801;
  reg [31:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_804;
  reg [31:0] _RAND_805;
  reg [31:0] _RAND_806;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [31:0] _RAND_810;
  reg [31:0] _RAND_811;
  reg [31:0] _RAND_812;
  reg [31:0] _RAND_813;
  reg [31:0] _RAND_814;
  reg [31:0] _RAND_815;
  reg [31:0] _RAND_816;
  reg [31:0] _RAND_817;
  reg [31:0] _RAND_818;
  reg [31:0] _RAND_819;
  reg [31:0] _RAND_820;
  reg [31:0] _RAND_821;
  reg [31:0] _RAND_822;
  reg [31:0] _RAND_823;
  reg [31:0] _RAND_824;
  reg [31:0] _RAND_825;
  reg [31:0] _RAND_826;
  reg [31:0] _RAND_827;
  reg [31:0] _RAND_828;
  reg [31:0] _RAND_829;
  reg [31:0] _RAND_830;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
  reg [31:0] _RAND_834;
  reg [31:0] _RAND_835;
  reg [31:0] _RAND_836;
  reg [31:0] _RAND_837;
  reg [31:0] _RAND_838;
  reg [31:0] _RAND_839;
  reg [31:0] _RAND_840;
  reg [31:0] _RAND_841;
  reg [31:0] _RAND_842;
  reg [31:0] _RAND_843;
  reg [31:0] _RAND_844;
  reg [31:0] _RAND_845;
  reg [31:0] _RAND_846;
  reg [31:0] _RAND_847;
  reg [31:0] _RAND_848;
  reg [31:0] _RAND_849;
  reg [31:0] _RAND_850;
  reg [31:0] _RAND_851;
  reg [31:0] _RAND_852;
  reg [31:0] _RAND_853;
  reg [31:0] _RAND_854;
  reg [31:0] _RAND_855;
  reg [31:0] _RAND_856;
  reg [31:0] _RAND_857;
  reg [31:0] _RAND_858;
  reg [31:0] _RAND_859;
  reg [31:0] _RAND_860;
  reg [31:0] _RAND_861;
  reg [31:0] _RAND_862;
  reg [63:0] _RAND_863;
  reg [31:0] _RAND_864;
  reg [31:0] _RAND_865;
  reg [31:0] _RAND_866;
  reg [31:0] _RAND_867;
  reg [31:0] _RAND_868;
  reg [31:0] _RAND_869;
  reg [31:0] _RAND_870;
  reg [31:0] _RAND_871;
  reg [31:0] _RAND_872;
  reg [31:0] _RAND_873;
  reg [31:0] _RAND_874;
  reg [31:0] _RAND_875;
  reg [31:0] _RAND_876;
  reg [31:0] _RAND_877;
  reg [31:0] _RAND_878;
  reg [31:0] _RAND_879;
  reg [31:0] _RAND_880;
  reg [31:0] _RAND_881;
  reg [31:0] _RAND_882;
  reg [31:0] _RAND_883;
  reg [31:0] _RAND_884;
  reg [31:0] _RAND_885;
  reg [31:0] _RAND_886;
  reg [31:0] _RAND_887;
  reg [31:0] _RAND_888;
  reg [31:0] _RAND_889;
  reg [31:0] _RAND_890;
  reg [31:0] _RAND_891;
  reg [31:0] _RAND_892;
  reg [31:0] _RAND_893;
  reg [31:0] _RAND_894;
  reg [31:0] _RAND_895;
  reg [31:0] _RAND_896;
  reg [31:0] _RAND_897;
  reg [31:0] _RAND_898;
  reg [31:0] _RAND_899;
  reg [31:0] _RAND_900;
  reg [31:0] _RAND_901;
  reg [31:0] _RAND_902;
  reg [31:0] _RAND_903;
  reg [31:0] _RAND_904;
  reg [31:0] _RAND_905;
  reg [31:0] _RAND_906;
  reg [31:0] _RAND_907;
  reg [31:0] _RAND_908;
  reg [31:0] _RAND_909;
  reg [31:0] _RAND_910;
  reg [31:0] _RAND_911;
  reg [31:0] _RAND_912;
  reg [31:0] _RAND_913;
  reg [31:0] _RAND_914;
  reg [31:0] _RAND_915;
  reg [31:0] _RAND_916;
  reg [31:0] _RAND_917;
  reg [31:0] _RAND_918;
  reg [31:0] _RAND_919;
  reg [31:0] _RAND_920;
  reg [31:0] _RAND_921;
  reg [31:0] _RAND_922;
  reg [31:0] _RAND_923;
  reg [31:0] _RAND_924;
  reg [31:0] _RAND_925;
  reg [31:0] _RAND_926;
  reg [31:0] _RAND_927;
  reg [31:0] _RAND_928;
  reg [31:0] _RAND_929;
  reg [31:0] _RAND_930;
  reg [31:0] _RAND_931;
  reg [31:0] _RAND_932;
  reg [31:0] _RAND_933;
  reg [31:0] _RAND_934;
  reg [31:0] _RAND_935;
  reg [31:0] _RAND_936;
  reg [31:0] _RAND_937;
  reg [31:0] _RAND_938;
  reg [31:0] _RAND_939;
  reg [63:0] _RAND_940;
  reg [31:0] _RAND_941;
  reg [31:0] _RAND_942;
  reg [31:0] _RAND_943;
  reg [31:0] _RAND_944;
  reg [31:0] _RAND_945;
  reg [31:0] _RAND_946;
  reg [31:0] _RAND_947;
  reg [31:0] _RAND_948;
  reg [31:0] _RAND_949;
  reg [31:0] _RAND_950;
  reg [31:0] _RAND_951;
  reg [31:0] _RAND_952;
  reg [31:0] _RAND_953;
  reg [31:0] _RAND_954;
  reg [31:0] _RAND_955;
  reg [31:0] _RAND_956;
  reg [31:0] _RAND_957;
  reg [31:0] _RAND_958;
  reg [31:0] _RAND_959;
  reg [31:0] _RAND_960;
  reg [31:0] _RAND_961;
  reg [31:0] _RAND_962;
  reg [31:0] _RAND_963;
  reg [31:0] _RAND_964;
  reg [31:0] _RAND_965;
  reg [31:0] _RAND_966;
  reg [31:0] _RAND_967;
  reg [31:0] _RAND_968;
  reg [31:0] _RAND_969;
  reg [31:0] _RAND_970;
  reg [31:0] _RAND_971;
  reg [31:0] _RAND_972;
  reg [31:0] _RAND_973;
  reg [31:0] _RAND_974;
  reg [31:0] _RAND_975;
  reg [31:0] _RAND_976;
  reg [31:0] _RAND_977;
  reg [31:0] _RAND_978;
  reg [31:0] _RAND_979;
  reg [31:0] _RAND_980;
  reg [31:0] _RAND_981;
  reg [31:0] _RAND_982;
  reg [31:0] _RAND_983;
  reg [31:0] _RAND_984;
  reg [31:0] _RAND_985;
  reg [31:0] _RAND_986;
  reg [31:0] _RAND_987;
  reg [31:0] _RAND_988;
  reg [31:0] _RAND_989;
  reg [31:0] _RAND_990;
  reg [31:0] _RAND_991;
  reg [31:0] _RAND_992;
  reg [31:0] _RAND_993;
  reg [31:0] _RAND_994;
  reg [31:0] _RAND_995;
  reg [31:0] _RAND_996;
  reg [31:0] _RAND_997;
  reg [31:0] _RAND_998;
  reg [31:0] _RAND_999;
  reg [31:0] _RAND_1000;
  reg [31:0] _RAND_1001;
  reg [31:0] _RAND_1002;
  reg [31:0] _RAND_1003;
  reg [31:0] _RAND_1004;
  reg [31:0] _RAND_1005;
  reg [31:0] _RAND_1006;
  reg [31:0] _RAND_1007;
  reg [31:0] _RAND_1008;
  reg [31:0] _RAND_1009;
  reg [31:0] _RAND_1010;
  reg [31:0] _RAND_1011;
  reg [31:0] _RAND_1012;
  reg [31:0] _RAND_1013;
  reg [31:0] _RAND_1014;
  reg [31:0] _RAND_1015;
  reg [63:0] _RAND_1016;
  reg [31:0] _RAND_1017;
  reg [31:0] _RAND_1018;
  reg [31:0] _RAND_1019;
  reg [31:0] _RAND_1020;
  reg [31:0] _RAND_1021;
  reg [31:0] _RAND_1022;
  reg [31:0] _RAND_1023;
  reg [31:0] _RAND_1024;
  reg [31:0] _RAND_1025;
  reg [31:0] _RAND_1026;
  reg [31:0] _RAND_1027;
  reg [31:0] _RAND_1028;
  reg [31:0] _RAND_1029;
  reg [31:0] _RAND_1030;
  reg [31:0] _RAND_1031;
  reg [31:0] _RAND_1032;
  reg [31:0] _RAND_1033;
  reg [31:0] _RAND_1034;
  reg [31:0] _RAND_1035;
  reg [31:0] _RAND_1036;
  reg [31:0] _RAND_1037;
  reg [31:0] _RAND_1038;
  reg [31:0] _RAND_1039;
  reg [31:0] _RAND_1040;
  reg [31:0] _RAND_1041;
  reg [31:0] _RAND_1042;
  reg [31:0] _RAND_1043;
  reg [31:0] _RAND_1044;
  reg [31:0] _RAND_1045;
  reg [31:0] _RAND_1046;
  reg [31:0] _RAND_1047;
  reg [31:0] _RAND_1048;
  reg [31:0] _RAND_1049;
  reg [31:0] _RAND_1050;
  reg [31:0] _RAND_1051;
  reg [31:0] _RAND_1052;
  reg [31:0] _RAND_1053;
  reg [31:0] _RAND_1054;
  reg [31:0] _RAND_1055;
  reg [31:0] _RAND_1056;
  reg [31:0] _RAND_1057;
  reg [31:0] _RAND_1058;
  reg [31:0] _RAND_1059;
  reg [31:0] _RAND_1060;
  reg [31:0] _RAND_1061;
  reg [31:0] _RAND_1062;
  reg [31:0] _RAND_1063;
  reg [31:0] _RAND_1064;
  reg [31:0] _RAND_1065;
  reg [31:0] _RAND_1066;
  reg [31:0] _RAND_1067;
  reg [31:0] _RAND_1068;
  reg [31:0] _RAND_1069;
  reg [31:0] _RAND_1070;
  reg [31:0] _RAND_1071;
  reg [31:0] _RAND_1072;
  reg [31:0] _RAND_1073;
  reg [31:0] _RAND_1074;
  reg [31:0] _RAND_1075;
  reg [31:0] _RAND_1076;
  reg [31:0] _RAND_1077;
  reg [31:0] _RAND_1078;
  reg [31:0] _RAND_1079;
  reg [31:0] _RAND_1080;
  reg [31:0] _RAND_1081;
  reg [31:0] _RAND_1082;
  reg [31:0] _RAND_1083;
  reg [31:0] _RAND_1084;
  reg [31:0] _RAND_1085;
  reg [31:0] _RAND_1086;
  reg [31:0] _RAND_1087;
  reg [31:0] _RAND_1088;
  reg [31:0] _RAND_1089;
  reg [31:0] _RAND_1090;
  reg [31:0] _RAND_1091;
  reg [63:0] _RAND_1092;
  reg [31:0] _RAND_1093;
  reg [31:0] _RAND_1094;
  reg [31:0] _RAND_1095;
  reg [31:0] _RAND_1096;
  reg [31:0] _RAND_1097;
  reg [31:0] _RAND_1098;
  reg [31:0] _RAND_1099;
  reg [31:0] _RAND_1100;
  reg [31:0] _RAND_1101;
  reg [31:0] _RAND_1102;
  reg [31:0] _RAND_1103;
  reg [31:0] _RAND_1104;
  reg [31:0] _RAND_1105;
  reg [31:0] _RAND_1106;
  reg [31:0] _RAND_1107;
  reg [31:0] _RAND_1108;
  reg [31:0] _RAND_1109;
  reg [31:0] _RAND_1110;
  reg [31:0] _RAND_1111;
  reg [31:0] _RAND_1112;
  reg [31:0] _RAND_1113;
  reg [31:0] _RAND_1114;
  reg [31:0] _RAND_1115;
  reg [31:0] _RAND_1116;
  reg [31:0] _RAND_1117;
  reg [31:0] _RAND_1118;
  reg [31:0] _RAND_1119;
  reg [31:0] _RAND_1120;
  reg [31:0] _RAND_1121;
  reg [31:0] _RAND_1122;
  reg [31:0] _RAND_1123;
  reg [31:0] _RAND_1124;
  reg [31:0] _RAND_1125;
  reg [31:0] _RAND_1126;
  reg [31:0] _RAND_1127;
  reg [31:0] _RAND_1128;
  reg [31:0] _RAND_1129;
  reg [31:0] _RAND_1130;
  reg [31:0] _RAND_1131;
  reg [31:0] _RAND_1132;
  reg [31:0] _RAND_1133;
  reg [31:0] _RAND_1134;
  reg [31:0] _RAND_1135;
  reg [31:0] _RAND_1136;
  reg [31:0] _RAND_1137;
  reg [31:0] _RAND_1138;
  reg [31:0] _RAND_1139;
  reg [31:0] _RAND_1140;
  reg [31:0] _RAND_1141;
  reg [31:0] _RAND_1142;
  reg [31:0] _RAND_1143;
  reg [31:0] _RAND_1144;
  reg [31:0] _RAND_1145;
  reg [31:0] _RAND_1146;
  reg [31:0] _RAND_1147;
  reg [31:0] _RAND_1148;
  reg [31:0] _RAND_1149;
  reg [31:0] _RAND_1150;
  reg [31:0] _RAND_1151;
  reg [31:0] _RAND_1152;
  reg [31:0] _RAND_1153;
  reg [31:0] _RAND_1154;
  reg [31:0] _RAND_1155;
  reg [31:0] _RAND_1156;
  reg [31:0] _RAND_1157;
  reg [31:0] _RAND_1158;
  reg [31:0] _RAND_1159;
  reg [31:0] _RAND_1160;
  reg [31:0] _RAND_1161;
  reg [31:0] _RAND_1162;
  reg [31:0] _RAND_1163;
  reg [31:0] _RAND_1164;
  reg [31:0] _RAND_1165;
  reg [31:0] _RAND_1166;
  reg [31:0] _RAND_1167;
  reg [63:0] _RAND_1168;
  reg [31:0] _RAND_1169;
  reg [31:0] _RAND_1170;
  reg [31:0] _RAND_1171;
  reg [31:0] _RAND_1172;
  reg [31:0] _RAND_1173;
  reg [31:0] _RAND_1174;
  reg [31:0] _RAND_1175;
  reg [31:0] _RAND_1176;
  reg [31:0] _RAND_1177;
  reg [31:0] _RAND_1178;
  reg [31:0] _RAND_1179;
  reg [31:0] _RAND_1180;
  reg [31:0] _RAND_1181;
  reg [31:0] _RAND_1182;
  reg [31:0] _RAND_1183;
  reg [31:0] _RAND_1184;
  reg [31:0] _RAND_1185;
  reg [31:0] _RAND_1186;
  reg [31:0] _RAND_1187;
  reg [31:0] _RAND_1188;
  reg [31:0] _RAND_1189;
  reg [31:0] _RAND_1190;
  reg [31:0] _RAND_1191;
  reg [31:0] _RAND_1192;
  reg [31:0] _RAND_1193;
  reg [31:0] _RAND_1194;
  reg [31:0] _RAND_1195;
  reg [31:0] _RAND_1196;
  reg [31:0] _RAND_1197;
  reg [31:0] _RAND_1198;
  reg [31:0] _RAND_1199;
  reg [31:0] _RAND_1200;
  reg [31:0] _RAND_1201;
  reg [31:0] _RAND_1202;
  reg [31:0] _RAND_1203;
  reg [31:0] _RAND_1204;
  reg [31:0] _RAND_1205;
  reg [31:0] _RAND_1206;
  reg [31:0] _RAND_1207;
  reg [31:0] _RAND_1208;
  reg [31:0] _RAND_1209;
  reg [31:0] _RAND_1210;
  reg [31:0] _RAND_1211;
  reg [31:0] _RAND_1212;
  reg [31:0] _RAND_1213;
  reg [31:0] _RAND_1214;
  reg [31:0] _RAND_1215;
  reg [31:0] _RAND_1216;
  reg [31:0] _RAND_1217;
  reg [31:0] _RAND_1218;
  reg [31:0] _RAND_1219;
  reg [31:0] _RAND_1220;
  reg [31:0] _RAND_1221;
  reg [31:0] _RAND_1222;
  reg [31:0] _RAND_1223;
  reg [31:0] _RAND_1224;
  reg [31:0] _RAND_1225;
  reg [31:0] _RAND_1226;
  reg [31:0] _RAND_1227;
  reg [31:0] _RAND_1228;
  reg [31:0] _RAND_1229;
  reg [31:0] _RAND_1230;
  reg [31:0] _RAND_1231;
  reg [31:0] _RAND_1232;
  reg [31:0] _RAND_1233;
  reg [31:0] _RAND_1234;
  reg [31:0] _RAND_1235;
  reg [31:0] _RAND_1236;
  reg [31:0] _RAND_1237;
  reg [31:0] _RAND_1238;
  reg [31:0] _RAND_1239;
  reg [31:0] _RAND_1240;
  reg [31:0] _RAND_1241;
  reg [31:0] _RAND_1242;
  reg [31:0] _RAND_1243;
  reg [63:0] _RAND_1244;
  reg [31:0] _RAND_1245;
  reg [31:0] _RAND_1246;
  reg [31:0] _RAND_1247;
  reg [31:0] _RAND_1248;
  reg [31:0] _RAND_1249;
  reg [31:0] _RAND_1250;
  reg [31:0] _RAND_1251;
  reg [31:0] _RAND_1252;
  reg [31:0] _RAND_1253;
  reg [31:0] _RAND_1254;
  reg [31:0] _RAND_1255;
  reg [31:0] _RAND_1256;
  reg [31:0] _RAND_1257;
  reg [31:0] _RAND_1258;
  reg [31:0] _RAND_1259;
  reg [31:0] _RAND_1260;
  reg [31:0] _RAND_1261;
  reg [31:0] _RAND_1262;
  reg [31:0] _RAND_1263;
  reg [31:0] _RAND_1264;
  reg [31:0] _RAND_1265;
  reg [31:0] _RAND_1266;
  reg [31:0] _RAND_1267;
  reg [31:0] _RAND_1268;
  reg [31:0] _RAND_1269;
  reg [31:0] _RAND_1270;
  reg [31:0] _RAND_1271;
  reg [31:0] _RAND_1272;
  reg [31:0] _RAND_1273;
  reg [31:0] _RAND_1274;
  reg [31:0] _RAND_1275;
  reg [31:0] _RAND_1276;
  reg [31:0] _RAND_1277;
  reg [31:0] _RAND_1278;
  reg [31:0] _RAND_1279;
  reg [31:0] _RAND_1280;
  reg [31:0] _RAND_1281;
  reg [31:0] _RAND_1282;
  reg [31:0] _RAND_1283;
  reg [31:0] _RAND_1284;
  reg [31:0] _RAND_1285;
  reg [31:0] _RAND_1286;
  reg [31:0] _RAND_1287;
  reg [31:0] _RAND_1288;
  reg [31:0] _RAND_1289;
  reg [31:0] _RAND_1290;
  reg [31:0] _RAND_1291;
  reg [31:0] _RAND_1292;
  reg [31:0] _RAND_1293;
  reg [31:0] _RAND_1294;
  reg [31:0] _RAND_1295;
  reg [31:0] _RAND_1296;
  reg [31:0] _RAND_1297;
  reg [31:0] _RAND_1298;
  reg [31:0] _RAND_1299;
  reg [31:0] _RAND_1300;
  reg [31:0] _RAND_1301;
  reg [31:0] _RAND_1302;
  reg [31:0] _RAND_1303;
  reg [31:0] _RAND_1304;
  reg [31:0] _RAND_1305;
  reg [31:0] _RAND_1306;
  reg [31:0] _RAND_1307;
  reg [31:0] _RAND_1308;
  reg [31:0] _RAND_1309;
  reg [31:0] _RAND_1310;
  reg [31:0] _RAND_1311;
  reg [31:0] _RAND_1312;
  reg [31:0] _RAND_1313;
  reg [31:0] _RAND_1314;
  reg [31:0] _RAND_1315;
  reg [31:0] _RAND_1316;
  reg [31:0] _RAND_1317;
  reg [31:0] _RAND_1318;
  reg [31:0] _RAND_1319;
  reg [63:0] _RAND_1320;
  reg [31:0] _RAND_1321;
  reg [31:0] _RAND_1322;
  reg [31:0] _RAND_1323;
  reg [31:0] _RAND_1324;
  reg [31:0] _RAND_1325;
  reg [31:0] _RAND_1326;
  reg [31:0] _RAND_1327;
  reg [31:0] _RAND_1328;
  reg [31:0] _RAND_1329;
  reg [31:0] _RAND_1330;
  reg [31:0] _RAND_1331;
  reg [31:0] _RAND_1332;
  reg [31:0] _RAND_1333;
  reg [31:0] _RAND_1334;
  reg [31:0] _RAND_1335;
  reg [31:0] _RAND_1336;
  reg [31:0] _RAND_1337;
  reg [31:0] _RAND_1338;
  reg [31:0] _RAND_1339;
  reg [31:0] _RAND_1340;
  reg [31:0] _RAND_1341;
  reg [31:0] _RAND_1342;
  reg [31:0] _RAND_1343;
  reg [31:0] _RAND_1344;
  reg [31:0] _RAND_1345;
  reg [31:0] _RAND_1346;
  reg [31:0] _RAND_1347;
  reg [31:0] _RAND_1348;
  reg [31:0] _RAND_1349;
  reg [31:0] _RAND_1350;
  reg [31:0] _RAND_1351;
  reg [31:0] _RAND_1352;
  reg [31:0] _RAND_1353;
  reg [31:0] _RAND_1354;
  reg [31:0] _RAND_1355;
  reg [31:0] _RAND_1356;
  reg [31:0] _RAND_1357;
  reg [31:0] _RAND_1358;
  reg [31:0] _RAND_1359;
  reg [31:0] _RAND_1360;
  reg [31:0] _RAND_1361;
  reg [31:0] _RAND_1362;
  reg [31:0] _RAND_1363;
  reg [31:0] _RAND_1364;
  reg [31:0] _RAND_1365;
  reg [31:0] _RAND_1366;
  reg [31:0] _RAND_1367;
  reg [31:0] _RAND_1368;
  reg [31:0] _RAND_1369;
  reg [31:0] _RAND_1370;
  reg [31:0] _RAND_1371;
  reg [31:0] _RAND_1372;
  reg [31:0] _RAND_1373;
  reg [31:0] _RAND_1374;
  reg [31:0] _RAND_1375;
  reg [31:0] _RAND_1376;
  reg [31:0] _RAND_1377;
  reg [31:0] _RAND_1378;
  reg [31:0] _RAND_1379;
  reg [31:0] _RAND_1380;
  reg [31:0] _RAND_1381;
  reg [31:0] _RAND_1382;
  reg [31:0] _RAND_1383;
  reg [31:0] _RAND_1384;
  reg [31:0] _RAND_1385;
  reg [31:0] _RAND_1386;
  reg [31:0] _RAND_1387;
  reg [31:0] _RAND_1388;
  reg [31:0] _RAND_1389;
  reg [31:0] _RAND_1390;
  reg [31:0] _RAND_1391;
  reg [31:0] _RAND_1392;
  reg [31:0] _RAND_1393;
  reg [31:0] _RAND_1394;
  reg [31:0] _RAND_1395;
  reg [63:0] _RAND_1396;
  reg [31:0] _RAND_1397;
  reg [31:0] _RAND_1398;
  reg [31:0] _RAND_1399;
  reg [31:0] _RAND_1400;
  reg [31:0] _RAND_1401;
  reg [31:0] _RAND_1402;
  reg [31:0] _RAND_1403;
  reg [31:0] _RAND_1404;
  reg [31:0] _RAND_1405;
  reg [31:0] _RAND_1406;
  reg [31:0] _RAND_1407;
  reg [31:0] _RAND_1408;
  reg [31:0] _RAND_1409;
  reg [31:0] _RAND_1410;
  reg [31:0] _RAND_1411;
  reg [31:0] _RAND_1412;
  reg [31:0] _RAND_1413;
  reg [31:0] _RAND_1414;
  reg [31:0] _RAND_1415;
  reg [31:0] _RAND_1416;
  reg [31:0] _RAND_1417;
  reg [31:0] _RAND_1418;
  reg [31:0] _RAND_1419;
  reg [31:0] _RAND_1420;
  reg [31:0] _RAND_1421;
  reg [31:0] _RAND_1422;
  reg [31:0] _RAND_1423;
  reg [31:0] _RAND_1424;
  reg [31:0] _RAND_1425;
  reg [31:0] _RAND_1426;
  reg [31:0] _RAND_1427;
  reg [31:0] _RAND_1428;
  reg [31:0] _RAND_1429;
  reg [31:0] _RAND_1430;
  reg [31:0] _RAND_1431;
  reg [31:0] _RAND_1432;
  reg [31:0] _RAND_1433;
  reg [31:0] _RAND_1434;
  reg [31:0] _RAND_1435;
  reg [31:0] _RAND_1436;
  reg [31:0] _RAND_1437;
  reg [31:0] _RAND_1438;
  reg [31:0] _RAND_1439;
  reg [31:0] _RAND_1440;
  reg [31:0] _RAND_1441;
  reg [31:0] _RAND_1442;
  reg [31:0] _RAND_1443;
  reg [31:0] _RAND_1444;
  reg [31:0] _RAND_1445;
  reg [31:0] _RAND_1446;
  reg [31:0] _RAND_1447;
  reg [31:0] _RAND_1448;
  reg [31:0] _RAND_1449;
  reg [31:0] _RAND_1450;
  reg [31:0] _RAND_1451;
  reg [31:0] _RAND_1452;
  reg [31:0] _RAND_1453;
  reg [31:0] _RAND_1454;
  reg [31:0] _RAND_1455;
  reg [31:0] _RAND_1456;
  reg [31:0] _RAND_1457;
  reg [31:0] _RAND_1458;
  reg [31:0] _RAND_1459;
  reg [31:0] _RAND_1460;
  reg [31:0] _RAND_1461;
  reg [31:0] _RAND_1462;
  reg [31:0] _RAND_1463;
  reg [31:0] _RAND_1464;
  reg [31:0] _RAND_1465;
  reg [31:0] _RAND_1466;
  reg [31:0] _RAND_1467;
  reg [31:0] _RAND_1468;
  reg [31:0] _RAND_1469;
  reg [31:0] _RAND_1470;
  reg [31:0] _RAND_1471;
  reg [63:0] _RAND_1472;
  reg [31:0] _RAND_1473;
  reg [31:0] _RAND_1474;
  reg [31:0] _RAND_1475;
  reg [31:0] _RAND_1476;
  reg [31:0] _RAND_1477;
  reg [31:0] _RAND_1478;
  reg [31:0] _RAND_1479;
  reg [31:0] _RAND_1480;
  reg [31:0] _RAND_1481;
  reg [31:0] _RAND_1482;
  reg [31:0] _RAND_1483;
  reg [31:0] _RAND_1484;
  reg [31:0] _RAND_1485;
  reg [31:0] _RAND_1486;
  reg [31:0] _RAND_1487;
  reg [31:0] _RAND_1488;
  reg [31:0] _RAND_1489;
  reg [31:0] _RAND_1490;
  reg [31:0] _RAND_1491;
  reg [31:0] _RAND_1492;
  reg [31:0] _RAND_1493;
  reg [31:0] _RAND_1494;
  reg [31:0] _RAND_1495;
  reg [31:0] _RAND_1496;
  reg [31:0] _RAND_1497;
  reg [31:0] _RAND_1498;
  reg [31:0] _RAND_1499;
  reg [31:0] _RAND_1500;
  reg [31:0] _RAND_1501;
  reg [31:0] _RAND_1502;
  reg [31:0] _RAND_1503;
  reg [31:0] _RAND_1504;
  reg [31:0] _RAND_1505;
  reg [31:0] _RAND_1506;
  reg [31:0] _RAND_1507;
  reg [31:0] _RAND_1508;
  reg [31:0] _RAND_1509;
  reg [31:0] _RAND_1510;
  reg [31:0] _RAND_1511;
  reg [31:0] _RAND_1512;
  reg [31:0] _RAND_1513;
  reg [31:0] _RAND_1514;
  reg [31:0] _RAND_1515;
  reg [31:0] _RAND_1516;
  reg [31:0] _RAND_1517;
  reg [31:0] _RAND_1518;
  reg [31:0] _RAND_1519;
  reg [31:0] _RAND_1520;
  reg [31:0] _RAND_1521;
  reg [31:0] _RAND_1522;
  reg [31:0] _RAND_1523;
  reg [31:0] _RAND_1524;
  reg [31:0] _RAND_1525;
  reg [31:0] _RAND_1526;
  reg [31:0] _RAND_1527;
  reg [31:0] _RAND_1528;
  reg [31:0] _RAND_1529;
  reg [31:0] _RAND_1530;
  reg [31:0] _RAND_1531;
  reg [31:0] _RAND_1532;
  reg [31:0] _RAND_1533;
  reg [31:0] _RAND_1534;
  reg [31:0] _RAND_1535;
  reg [31:0] _RAND_1536;
  reg [31:0] _RAND_1537;
  reg [31:0] _RAND_1538;
  reg [31:0] _RAND_1539;
  reg [31:0] _RAND_1540;
  reg [31:0] _RAND_1541;
  reg [31:0] _RAND_1542;
  reg [31:0] _RAND_1543;
  reg [31:0] _RAND_1544;
  reg [31:0] _RAND_1545;
  reg [31:0] _RAND_1546;
`endif // RANDOMIZE_REG_INIT
  wire  l2_clock; // @[PageTableCache.scala 155:18]
  wire  l2_io_rreq_valid; // @[PageTableCache.scala 155:18]
  wire [1:0] l2_io_rreq_bits_setIdx; // @[PageTableCache.scala 155:18]
  wire [12:0] l2_io_rresp_data_0_entries_tag; // @[PageTableCache.scala 155:18]
  wire [15:0] l2_io_rresp_data_0_entries_asid; // @[PageTableCache.scala 155:18]
  wire [23:0] l2_io_rresp_data_0_entries_ppns_0; // @[PageTableCache.scala 155:18]
  wire [23:0] l2_io_rresp_data_0_entries_ppns_1; // @[PageTableCache.scala 155:18]
  wire [23:0] l2_io_rresp_data_0_entries_ppns_2; // @[PageTableCache.scala 155:18]
  wire [23:0] l2_io_rresp_data_0_entries_ppns_3; // @[PageTableCache.scala 155:18]
  wire [23:0] l2_io_rresp_data_0_entries_ppns_4; // @[PageTableCache.scala 155:18]
  wire [23:0] l2_io_rresp_data_0_entries_ppns_5; // @[PageTableCache.scala 155:18]
  wire [23:0] l2_io_rresp_data_0_entries_ppns_6; // @[PageTableCache.scala 155:18]
  wire [23:0] l2_io_rresp_data_0_entries_ppns_7; // @[PageTableCache.scala 155:18]
  wire  l2_io_rresp_data_0_entries_vs_0; // @[PageTableCache.scala 155:18]
  wire  l2_io_rresp_data_0_entries_vs_1; // @[PageTableCache.scala 155:18]
  wire  l2_io_rresp_data_0_entries_vs_2; // @[PageTableCache.scala 155:18]
  wire  l2_io_rresp_data_0_entries_vs_3; // @[PageTableCache.scala 155:18]
  wire  l2_io_rresp_data_0_entries_vs_4; // @[PageTableCache.scala 155:18]
  wire  l2_io_rresp_data_0_entries_vs_5; // @[PageTableCache.scala 155:18]
  wire  l2_io_rresp_data_0_entries_vs_6; // @[PageTableCache.scala 155:18]
  wire  l2_io_rresp_data_0_entries_vs_7; // @[PageTableCache.scala 155:18]
  wire  l2_io_rresp_data_0_entries_prefetch; // @[PageTableCache.scala 155:18]
  wire [30:0] l2_io_rresp_data_0_ecc; // @[PageTableCache.scala 155:18]
  wire [12:0] l2_io_rresp_data_1_entries_tag; // @[PageTableCache.scala 155:18]
  wire [15:0] l2_io_rresp_data_1_entries_asid; // @[PageTableCache.scala 155:18]
  wire [23:0] l2_io_rresp_data_1_entries_ppns_0; // @[PageTableCache.scala 155:18]
  wire [23:0] l2_io_rresp_data_1_entries_ppns_1; // @[PageTableCache.scala 155:18]
  wire [23:0] l2_io_rresp_data_1_entries_ppns_2; // @[PageTableCache.scala 155:18]
  wire [23:0] l2_io_rresp_data_1_entries_ppns_3; // @[PageTableCache.scala 155:18]
  wire [23:0] l2_io_rresp_data_1_entries_ppns_4; // @[PageTableCache.scala 155:18]
  wire [23:0] l2_io_rresp_data_1_entries_ppns_5; // @[PageTableCache.scala 155:18]
  wire [23:0] l2_io_rresp_data_1_entries_ppns_6; // @[PageTableCache.scala 155:18]
  wire [23:0] l2_io_rresp_data_1_entries_ppns_7; // @[PageTableCache.scala 155:18]
  wire  l2_io_rresp_data_1_entries_vs_0; // @[PageTableCache.scala 155:18]
  wire  l2_io_rresp_data_1_entries_vs_1; // @[PageTableCache.scala 155:18]
  wire  l2_io_rresp_data_1_entries_vs_2; // @[PageTableCache.scala 155:18]
  wire  l2_io_rresp_data_1_entries_vs_3; // @[PageTableCache.scala 155:18]
  wire  l2_io_rresp_data_1_entries_vs_4; // @[PageTableCache.scala 155:18]
  wire  l2_io_rresp_data_1_entries_vs_5; // @[PageTableCache.scala 155:18]
  wire  l2_io_rresp_data_1_entries_vs_6; // @[PageTableCache.scala 155:18]
  wire  l2_io_rresp_data_1_entries_vs_7; // @[PageTableCache.scala 155:18]
  wire  l2_io_rresp_data_1_entries_prefetch; // @[PageTableCache.scala 155:18]
  wire [30:0] l2_io_rresp_data_1_ecc; // @[PageTableCache.scala 155:18]
  wire [12:0] l2_io_rresp_data_2_entries_tag; // @[PageTableCache.scala 155:18]
  wire [15:0] l2_io_rresp_data_2_entries_asid; // @[PageTableCache.scala 155:18]
  wire [23:0] l2_io_rresp_data_2_entries_ppns_0; // @[PageTableCache.scala 155:18]
  wire [23:0] l2_io_rresp_data_2_entries_ppns_1; // @[PageTableCache.scala 155:18]
  wire [23:0] l2_io_rresp_data_2_entries_ppns_2; // @[PageTableCache.scala 155:18]
  wire [23:0] l2_io_rresp_data_2_entries_ppns_3; // @[PageTableCache.scala 155:18]
  wire [23:0] l2_io_rresp_data_2_entries_ppns_4; // @[PageTableCache.scala 155:18]
  wire [23:0] l2_io_rresp_data_2_entries_ppns_5; // @[PageTableCache.scala 155:18]
  wire [23:0] l2_io_rresp_data_2_entries_ppns_6; // @[PageTableCache.scala 155:18]
  wire [23:0] l2_io_rresp_data_2_entries_ppns_7; // @[PageTableCache.scala 155:18]
  wire  l2_io_rresp_data_2_entries_vs_0; // @[PageTableCache.scala 155:18]
  wire  l2_io_rresp_data_2_entries_vs_1; // @[PageTableCache.scala 155:18]
  wire  l2_io_rresp_data_2_entries_vs_2; // @[PageTableCache.scala 155:18]
  wire  l2_io_rresp_data_2_entries_vs_3; // @[PageTableCache.scala 155:18]
  wire  l2_io_rresp_data_2_entries_vs_4; // @[PageTableCache.scala 155:18]
  wire  l2_io_rresp_data_2_entries_vs_5; // @[PageTableCache.scala 155:18]
  wire  l2_io_rresp_data_2_entries_vs_6; // @[PageTableCache.scala 155:18]
  wire  l2_io_rresp_data_2_entries_vs_7; // @[PageTableCache.scala 155:18]
  wire  l2_io_rresp_data_2_entries_prefetch; // @[PageTableCache.scala 155:18]
  wire [30:0] l2_io_rresp_data_2_ecc; // @[PageTableCache.scala 155:18]
  wire [12:0] l2_io_rresp_data_3_entries_tag; // @[PageTableCache.scala 155:18]
  wire [15:0] l2_io_rresp_data_3_entries_asid; // @[PageTableCache.scala 155:18]
  wire [23:0] l2_io_rresp_data_3_entries_ppns_0; // @[PageTableCache.scala 155:18]
  wire [23:0] l2_io_rresp_data_3_entries_ppns_1; // @[PageTableCache.scala 155:18]
  wire [23:0] l2_io_rresp_data_3_entries_ppns_2; // @[PageTableCache.scala 155:18]
  wire [23:0] l2_io_rresp_data_3_entries_ppns_3; // @[PageTableCache.scala 155:18]
  wire [23:0] l2_io_rresp_data_3_entries_ppns_4; // @[PageTableCache.scala 155:18]
  wire [23:0] l2_io_rresp_data_3_entries_ppns_5; // @[PageTableCache.scala 155:18]
  wire [23:0] l2_io_rresp_data_3_entries_ppns_6; // @[PageTableCache.scala 155:18]
  wire [23:0] l2_io_rresp_data_3_entries_ppns_7; // @[PageTableCache.scala 155:18]
  wire  l2_io_rresp_data_3_entries_vs_0; // @[PageTableCache.scala 155:18]
  wire  l2_io_rresp_data_3_entries_vs_1; // @[PageTableCache.scala 155:18]
  wire  l2_io_rresp_data_3_entries_vs_2; // @[PageTableCache.scala 155:18]
  wire  l2_io_rresp_data_3_entries_vs_3; // @[PageTableCache.scala 155:18]
  wire  l2_io_rresp_data_3_entries_vs_4; // @[PageTableCache.scala 155:18]
  wire  l2_io_rresp_data_3_entries_vs_5; // @[PageTableCache.scala 155:18]
  wire  l2_io_rresp_data_3_entries_vs_6; // @[PageTableCache.scala 155:18]
  wire  l2_io_rresp_data_3_entries_vs_7; // @[PageTableCache.scala 155:18]
  wire  l2_io_rresp_data_3_entries_prefetch; // @[PageTableCache.scala 155:18]
  wire [30:0] l2_io_rresp_data_3_ecc; // @[PageTableCache.scala 155:18]
  wire  l2_io_wreq_valid; // @[PageTableCache.scala 155:18]
  wire [1:0] l2_io_wreq_bits_setIdx; // @[PageTableCache.scala 155:18]
  wire [12:0] l2_io_wreq_bits_data_0_entries_tag; // @[PageTableCache.scala 155:18]
  wire [15:0] l2_io_wreq_bits_data_0_entries_asid; // @[PageTableCache.scala 155:18]
  wire [23:0] l2_io_wreq_bits_data_0_entries_ppns_0; // @[PageTableCache.scala 155:18]
  wire [23:0] l2_io_wreq_bits_data_0_entries_ppns_1; // @[PageTableCache.scala 155:18]
  wire [23:0] l2_io_wreq_bits_data_0_entries_ppns_2; // @[PageTableCache.scala 155:18]
  wire [23:0] l2_io_wreq_bits_data_0_entries_ppns_3; // @[PageTableCache.scala 155:18]
  wire [23:0] l2_io_wreq_bits_data_0_entries_ppns_4; // @[PageTableCache.scala 155:18]
  wire [23:0] l2_io_wreq_bits_data_0_entries_ppns_5; // @[PageTableCache.scala 155:18]
  wire [23:0] l2_io_wreq_bits_data_0_entries_ppns_6; // @[PageTableCache.scala 155:18]
  wire [23:0] l2_io_wreq_bits_data_0_entries_ppns_7; // @[PageTableCache.scala 155:18]
  wire  l2_io_wreq_bits_data_0_entries_vs_0; // @[PageTableCache.scala 155:18]
  wire  l2_io_wreq_bits_data_0_entries_vs_1; // @[PageTableCache.scala 155:18]
  wire  l2_io_wreq_bits_data_0_entries_vs_2; // @[PageTableCache.scala 155:18]
  wire  l2_io_wreq_bits_data_0_entries_vs_3; // @[PageTableCache.scala 155:18]
  wire  l2_io_wreq_bits_data_0_entries_vs_4; // @[PageTableCache.scala 155:18]
  wire  l2_io_wreq_bits_data_0_entries_vs_5; // @[PageTableCache.scala 155:18]
  wire  l2_io_wreq_bits_data_0_entries_vs_6; // @[PageTableCache.scala 155:18]
  wire  l2_io_wreq_bits_data_0_entries_vs_7; // @[PageTableCache.scala 155:18]
  wire  l2_io_wreq_bits_data_0_entries_prefetch; // @[PageTableCache.scala 155:18]
  wire [30:0] l2_io_wreq_bits_data_0_ecc; // @[PageTableCache.scala 155:18]
  wire [12:0] l2_io_wreq_bits_data_1_entries_tag; // @[PageTableCache.scala 155:18]
  wire [15:0] l2_io_wreq_bits_data_1_entries_asid; // @[PageTableCache.scala 155:18]
  wire [23:0] l2_io_wreq_bits_data_1_entries_ppns_0; // @[PageTableCache.scala 155:18]
  wire [23:0] l2_io_wreq_bits_data_1_entries_ppns_1; // @[PageTableCache.scala 155:18]
  wire [23:0] l2_io_wreq_bits_data_1_entries_ppns_2; // @[PageTableCache.scala 155:18]
  wire [23:0] l2_io_wreq_bits_data_1_entries_ppns_3; // @[PageTableCache.scala 155:18]
  wire [23:0] l2_io_wreq_bits_data_1_entries_ppns_4; // @[PageTableCache.scala 155:18]
  wire [23:0] l2_io_wreq_bits_data_1_entries_ppns_5; // @[PageTableCache.scala 155:18]
  wire [23:0] l2_io_wreq_bits_data_1_entries_ppns_6; // @[PageTableCache.scala 155:18]
  wire [23:0] l2_io_wreq_bits_data_1_entries_ppns_7; // @[PageTableCache.scala 155:18]
  wire  l2_io_wreq_bits_data_1_entries_vs_0; // @[PageTableCache.scala 155:18]
  wire  l2_io_wreq_bits_data_1_entries_vs_1; // @[PageTableCache.scala 155:18]
  wire  l2_io_wreq_bits_data_1_entries_vs_2; // @[PageTableCache.scala 155:18]
  wire  l2_io_wreq_bits_data_1_entries_vs_3; // @[PageTableCache.scala 155:18]
  wire  l2_io_wreq_bits_data_1_entries_vs_4; // @[PageTableCache.scala 155:18]
  wire  l2_io_wreq_bits_data_1_entries_vs_5; // @[PageTableCache.scala 155:18]
  wire  l2_io_wreq_bits_data_1_entries_vs_6; // @[PageTableCache.scala 155:18]
  wire  l2_io_wreq_bits_data_1_entries_vs_7; // @[PageTableCache.scala 155:18]
  wire  l2_io_wreq_bits_data_1_entries_prefetch; // @[PageTableCache.scala 155:18]
  wire [30:0] l2_io_wreq_bits_data_1_ecc; // @[PageTableCache.scala 155:18]
  wire [12:0] l2_io_wreq_bits_data_2_entries_tag; // @[PageTableCache.scala 155:18]
  wire [15:0] l2_io_wreq_bits_data_2_entries_asid; // @[PageTableCache.scala 155:18]
  wire [23:0] l2_io_wreq_bits_data_2_entries_ppns_0; // @[PageTableCache.scala 155:18]
  wire [23:0] l2_io_wreq_bits_data_2_entries_ppns_1; // @[PageTableCache.scala 155:18]
  wire [23:0] l2_io_wreq_bits_data_2_entries_ppns_2; // @[PageTableCache.scala 155:18]
  wire [23:0] l2_io_wreq_bits_data_2_entries_ppns_3; // @[PageTableCache.scala 155:18]
  wire [23:0] l2_io_wreq_bits_data_2_entries_ppns_4; // @[PageTableCache.scala 155:18]
  wire [23:0] l2_io_wreq_bits_data_2_entries_ppns_5; // @[PageTableCache.scala 155:18]
  wire [23:0] l2_io_wreq_bits_data_2_entries_ppns_6; // @[PageTableCache.scala 155:18]
  wire [23:0] l2_io_wreq_bits_data_2_entries_ppns_7; // @[PageTableCache.scala 155:18]
  wire  l2_io_wreq_bits_data_2_entries_vs_0; // @[PageTableCache.scala 155:18]
  wire  l2_io_wreq_bits_data_2_entries_vs_1; // @[PageTableCache.scala 155:18]
  wire  l2_io_wreq_bits_data_2_entries_vs_2; // @[PageTableCache.scala 155:18]
  wire  l2_io_wreq_bits_data_2_entries_vs_3; // @[PageTableCache.scala 155:18]
  wire  l2_io_wreq_bits_data_2_entries_vs_4; // @[PageTableCache.scala 155:18]
  wire  l2_io_wreq_bits_data_2_entries_vs_5; // @[PageTableCache.scala 155:18]
  wire  l2_io_wreq_bits_data_2_entries_vs_6; // @[PageTableCache.scala 155:18]
  wire  l2_io_wreq_bits_data_2_entries_vs_7; // @[PageTableCache.scala 155:18]
  wire  l2_io_wreq_bits_data_2_entries_prefetch; // @[PageTableCache.scala 155:18]
  wire [30:0] l2_io_wreq_bits_data_2_ecc; // @[PageTableCache.scala 155:18]
  wire [12:0] l2_io_wreq_bits_data_3_entries_tag; // @[PageTableCache.scala 155:18]
  wire [15:0] l2_io_wreq_bits_data_3_entries_asid; // @[PageTableCache.scala 155:18]
  wire [23:0] l2_io_wreq_bits_data_3_entries_ppns_0; // @[PageTableCache.scala 155:18]
  wire [23:0] l2_io_wreq_bits_data_3_entries_ppns_1; // @[PageTableCache.scala 155:18]
  wire [23:0] l2_io_wreq_bits_data_3_entries_ppns_2; // @[PageTableCache.scala 155:18]
  wire [23:0] l2_io_wreq_bits_data_3_entries_ppns_3; // @[PageTableCache.scala 155:18]
  wire [23:0] l2_io_wreq_bits_data_3_entries_ppns_4; // @[PageTableCache.scala 155:18]
  wire [23:0] l2_io_wreq_bits_data_3_entries_ppns_5; // @[PageTableCache.scala 155:18]
  wire [23:0] l2_io_wreq_bits_data_3_entries_ppns_6; // @[PageTableCache.scala 155:18]
  wire [23:0] l2_io_wreq_bits_data_3_entries_ppns_7; // @[PageTableCache.scala 155:18]
  wire  l2_io_wreq_bits_data_3_entries_vs_0; // @[PageTableCache.scala 155:18]
  wire  l2_io_wreq_bits_data_3_entries_vs_1; // @[PageTableCache.scala 155:18]
  wire  l2_io_wreq_bits_data_3_entries_vs_2; // @[PageTableCache.scala 155:18]
  wire  l2_io_wreq_bits_data_3_entries_vs_3; // @[PageTableCache.scala 155:18]
  wire  l2_io_wreq_bits_data_3_entries_vs_4; // @[PageTableCache.scala 155:18]
  wire  l2_io_wreq_bits_data_3_entries_vs_5; // @[PageTableCache.scala 155:18]
  wire  l2_io_wreq_bits_data_3_entries_vs_6; // @[PageTableCache.scala 155:18]
  wire  l2_io_wreq_bits_data_3_entries_vs_7; // @[PageTableCache.scala 155:18]
  wire  l2_io_wreq_bits_data_3_entries_prefetch; // @[PageTableCache.scala 155:18]
  wire [30:0] l2_io_wreq_bits_data_3_ecc; // @[PageTableCache.scala 155:18]
  wire [3:0] l2_io_wreq_bits_waymask; // @[PageTableCache.scala 155:18]
  wire  l3_clock; // @[PageTableCache.scala 179:18]
  wire  l3_io_rreq_valid; // @[PageTableCache.scala 179:18]
  wire [1:0] l3_io_rreq_bits_setIdx; // @[PageTableCache.scala 179:18]
  wire [21:0] l3_io_rresp_data_0_entries_tag; // @[PageTableCache.scala 179:18]
  wire [15:0] l3_io_rresp_data_0_entries_asid; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_rresp_data_0_entries_ppns_0; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_rresp_data_0_entries_ppns_1; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_rresp_data_0_entries_ppns_2; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_rresp_data_0_entries_ppns_3; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_rresp_data_0_entries_ppns_4; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_rresp_data_0_entries_ppns_5; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_rresp_data_0_entries_ppns_6; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_rresp_data_0_entries_ppns_7; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_0_entries_vs_0; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_0_entries_vs_1; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_0_entries_vs_2; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_0_entries_vs_3; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_0_entries_vs_4; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_0_entries_vs_5; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_0_entries_vs_6; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_0_entries_vs_7; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_0_entries_perms_0_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_0_entries_perms_0_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_0_entries_perms_0_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_0_entries_perms_0_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_0_entries_perms_0_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_0_entries_perms_0_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_0_entries_perms_0_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_0_entries_perms_1_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_0_entries_perms_1_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_0_entries_perms_1_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_0_entries_perms_1_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_0_entries_perms_1_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_0_entries_perms_1_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_0_entries_perms_1_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_0_entries_perms_2_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_0_entries_perms_2_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_0_entries_perms_2_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_0_entries_perms_2_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_0_entries_perms_2_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_0_entries_perms_2_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_0_entries_perms_2_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_0_entries_perms_3_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_0_entries_perms_3_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_0_entries_perms_3_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_0_entries_perms_3_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_0_entries_perms_3_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_0_entries_perms_3_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_0_entries_perms_3_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_0_entries_perms_4_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_0_entries_perms_4_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_0_entries_perms_4_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_0_entries_perms_4_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_0_entries_perms_4_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_0_entries_perms_4_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_0_entries_perms_4_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_0_entries_perms_5_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_0_entries_perms_5_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_0_entries_perms_5_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_0_entries_perms_5_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_0_entries_perms_5_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_0_entries_perms_5_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_0_entries_perms_5_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_0_entries_perms_6_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_0_entries_perms_6_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_0_entries_perms_6_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_0_entries_perms_6_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_0_entries_perms_6_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_0_entries_perms_6_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_0_entries_perms_6_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_0_entries_perms_7_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_0_entries_perms_7_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_0_entries_perms_7_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_0_entries_perms_7_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_0_entries_perms_7_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_0_entries_perms_7_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_0_entries_perms_7_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_0_entries_prefetch; // @[PageTableCache.scala 179:18]
  wire [38:0] l3_io_rresp_data_0_ecc; // @[PageTableCache.scala 179:18]
  wire [21:0] l3_io_rresp_data_1_entries_tag; // @[PageTableCache.scala 179:18]
  wire [15:0] l3_io_rresp_data_1_entries_asid; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_rresp_data_1_entries_ppns_0; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_rresp_data_1_entries_ppns_1; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_rresp_data_1_entries_ppns_2; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_rresp_data_1_entries_ppns_3; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_rresp_data_1_entries_ppns_4; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_rresp_data_1_entries_ppns_5; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_rresp_data_1_entries_ppns_6; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_rresp_data_1_entries_ppns_7; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_1_entries_vs_0; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_1_entries_vs_1; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_1_entries_vs_2; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_1_entries_vs_3; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_1_entries_vs_4; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_1_entries_vs_5; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_1_entries_vs_6; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_1_entries_vs_7; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_1_entries_perms_0_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_1_entries_perms_0_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_1_entries_perms_0_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_1_entries_perms_0_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_1_entries_perms_0_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_1_entries_perms_0_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_1_entries_perms_0_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_1_entries_perms_1_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_1_entries_perms_1_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_1_entries_perms_1_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_1_entries_perms_1_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_1_entries_perms_1_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_1_entries_perms_1_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_1_entries_perms_1_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_1_entries_perms_2_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_1_entries_perms_2_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_1_entries_perms_2_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_1_entries_perms_2_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_1_entries_perms_2_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_1_entries_perms_2_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_1_entries_perms_2_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_1_entries_perms_3_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_1_entries_perms_3_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_1_entries_perms_3_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_1_entries_perms_3_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_1_entries_perms_3_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_1_entries_perms_3_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_1_entries_perms_3_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_1_entries_perms_4_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_1_entries_perms_4_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_1_entries_perms_4_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_1_entries_perms_4_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_1_entries_perms_4_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_1_entries_perms_4_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_1_entries_perms_4_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_1_entries_perms_5_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_1_entries_perms_5_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_1_entries_perms_5_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_1_entries_perms_5_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_1_entries_perms_5_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_1_entries_perms_5_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_1_entries_perms_5_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_1_entries_perms_6_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_1_entries_perms_6_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_1_entries_perms_6_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_1_entries_perms_6_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_1_entries_perms_6_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_1_entries_perms_6_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_1_entries_perms_6_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_1_entries_perms_7_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_1_entries_perms_7_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_1_entries_perms_7_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_1_entries_perms_7_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_1_entries_perms_7_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_1_entries_perms_7_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_1_entries_perms_7_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_1_entries_prefetch; // @[PageTableCache.scala 179:18]
  wire [38:0] l3_io_rresp_data_1_ecc; // @[PageTableCache.scala 179:18]
  wire [21:0] l3_io_rresp_data_2_entries_tag; // @[PageTableCache.scala 179:18]
  wire [15:0] l3_io_rresp_data_2_entries_asid; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_rresp_data_2_entries_ppns_0; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_rresp_data_2_entries_ppns_1; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_rresp_data_2_entries_ppns_2; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_rresp_data_2_entries_ppns_3; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_rresp_data_2_entries_ppns_4; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_rresp_data_2_entries_ppns_5; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_rresp_data_2_entries_ppns_6; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_rresp_data_2_entries_ppns_7; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_2_entries_vs_0; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_2_entries_vs_1; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_2_entries_vs_2; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_2_entries_vs_3; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_2_entries_vs_4; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_2_entries_vs_5; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_2_entries_vs_6; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_2_entries_vs_7; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_2_entries_perms_0_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_2_entries_perms_0_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_2_entries_perms_0_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_2_entries_perms_0_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_2_entries_perms_0_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_2_entries_perms_0_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_2_entries_perms_0_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_2_entries_perms_1_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_2_entries_perms_1_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_2_entries_perms_1_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_2_entries_perms_1_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_2_entries_perms_1_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_2_entries_perms_1_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_2_entries_perms_1_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_2_entries_perms_2_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_2_entries_perms_2_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_2_entries_perms_2_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_2_entries_perms_2_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_2_entries_perms_2_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_2_entries_perms_2_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_2_entries_perms_2_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_2_entries_perms_3_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_2_entries_perms_3_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_2_entries_perms_3_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_2_entries_perms_3_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_2_entries_perms_3_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_2_entries_perms_3_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_2_entries_perms_3_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_2_entries_perms_4_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_2_entries_perms_4_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_2_entries_perms_4_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_2_entries_perms_4_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_2_entries_perms_4_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_2_entries_perms_4_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_2_entries_perms_4_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_2_entries_perms_5_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_2_entries_perms_5_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_2_entries_perms_5_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_2_entries_perms_5_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_2_entries_perms_5_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_2_entries_perms_5_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_2_entries_perms_5_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_2_entries_perms_6_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_2_entries_perms_6_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_2_entries_perms_6_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_2_entries_perms_6_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_2_entries_perms_6_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_2_entries_perms_6_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_2_entries_perms_6_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_2_entries_perms_7_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_2_entries_perms_7_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_2_entries_perms_7_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_2_entries_perms_7_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_2_entries_perms_7_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_2_entries_perms_7_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_2_entries_perms_7_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_2_entries_prefetch; // @[PageTableCache.scala 179:18]
  wire [38:0] l3_io_rresp_data_2_ecc; // @[PageTableCache.scala 179:18]
  wire [21:0] l3_io_rresp_data_3_entries_tag; // @[PageTableCache.scala 179:18]
  wire [15:0] l3_io_rresp_data_3_entries_asid; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_rresp_data_3_entries_ppns_0; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_rresp_data_3_entries_ppns_1; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_rresp_data_3_entries_ppns_2; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_rresp_data_3_entries_ppns_3; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_rresp_data_3_entries_ppns_4; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_rresp_data_3_entries_ppns_5; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_rresp_data_3_entries_ppns_6; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_rresp_data_3_entries_ppns_7; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_3_entries_vs_0; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_3_entries_vs_1; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_3_entries_vs_2; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_3_entries_vs_3; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_3_entries_vs_4; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_3_entries_vs_5; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_3_entries_vs_6; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_3_entries_vs_7; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_3_entries_perms_0_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_3_entries_perms_0_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_3_entries_perms_0_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_3_entries_perms_0_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_3_entries_perms_0_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_3_entries_perms_0_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_3_entries_perms_0_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_3_entries_perms_1_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_3_entries_perms_1_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_3_entries_perms_1_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_3_entries_perms_1_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_3_entries_perms_1_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_3_entries_perms_1_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_3_entries_perms_1_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_3_entries_perms_2_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_3_entries_perms_2_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_3_entries_perms_2_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_3_entries_perms_2_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_3_entries_perms_2_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_3_entries_perms_2_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_3_entries_perms_2_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_3_entries_perms_3_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_3_entries_perms_3_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_3_entries_perms_3_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_3_entries_perms_3_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_3_entries_perms_3_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_3_entries_perms_3_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_3_entries_perms_3_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_3_entries_perms_4_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_3_entries_perms_4_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_3_entries_perms_4_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_3_entries_perms_4_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_3_entries_perms_4_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_3_entries_perms_4_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_3_entries_perms_4_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_3_entries_perms_5_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_3_entries_perms_5_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_3_entries_perms_5_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_3_entries_perms_5_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_3_entries_perms_5_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_3_entries_perms_5_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_3_entries_perms_5_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_3_entries_perms_6_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_3_entries_perms_6_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_3_entries_perms_6_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_3_entries_perms_6_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_3_entries_perms_6_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_3_entries_perms_6_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_3_entries_perms_6_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_3_entries_perms_7_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_3_entries_perms_7_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_3_entries_perms_7_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_3_entries_perms_7_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_3_entries_perms_7_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_3_entries_perms_7_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_3_entries_perms_7_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_3_entries_prefetch; // @[PageTableCache.scala 179:18]
  wire [38:0] l3_io_rresp_data_3_ecc; // @[PageTableCache.scala 179:18]
  wire [21:0] l3_io_rresp_data_4_entries_tag; // @[PageTableCache.scala 179:18]
  wire [15:0] l3_io_rresp_data_4_entries_asid; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_rresp_data_4_entries_ppns_0; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_rresp_data_4_entries_ppns_1; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_rresp_data_4_entries_ppns_2; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_rresp_data_4_entries_ppns_3; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_rresp_data_4_entries_ppns_4; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_rresp_data_4_entries_ppns_5; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_rresp_data_4_entries_ppns_6; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_rresp_data_4_entries_ppns_7; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_4_entries_vs_0; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_4_entries_vs_1; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_4_entries_vs_2; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_4_entries_vs_3; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_4_entries_vs_4; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_4_entries_vs_5; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_4_entries_vs_6; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_4_entries_vs_7; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_4_entries_perms_0_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_4_entries_perms_0_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_4_entries_perms_0_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_4_entries_perms_0_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_4_entries_perms_0_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_4_entries_perms_0_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_4_entries_perms_0_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_4_entries_perms_1_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_4_entries_perms_1_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_4_entries_perms_1_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_4_entries_perms_1_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_4_entries_perms_1_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_4_entries_perms_1_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_4_entries_perms_1_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_4_entries_perms_2_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_4_entries_perms_2_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_4_entries_perms_2_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_4_entries_perms_2_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_4_entries_perms_2_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_4_entries_perms_2_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_4_entries_perms_2_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_4_entries_perms_3_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_4_entries_perms_3_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_4_entries_perms_3_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_4_entries_perms_3_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_4_entries_perms_3_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_4_entries_perms_3_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_4_entries_perms_3_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_4_entries_perms_4_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_4_entries_perms_4_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_4_entries_perms_4_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_4_entries_perms_4_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_4_entries_perms_4_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_4_entries_perms_4_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_4_entries_perms_4_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_4_entries_perms_5_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_4_entries_perms_5_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_4_entries_perms_5_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_4_entries_perms_5_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_4_entries_perms_5_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_4_entries_perms_5_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_4_entries_perms_5_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_4_entries_perms_6_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_4_entries_perms_6_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_4_entries_perms_6_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_4_entries_perms_6_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_4_entries_perms_6_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_4_entries_perms_6_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_4_entries_perms_6_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_4_entries_perms_7_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_4_entries_perms_7_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_4_entries_perms_7_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_4_entries_perms_7_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_4_entries_perms_7_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_4_entries_perms_7_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_4_entries_perms_7_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_4_entries_prefetch; // @[PageTableCache.scala 179:18]
  wire [38:0] l3_io_rresp_data_4_ecc; // @[PageTableCache.scala 179:18]
  wire [21:0] l3_io_rresp_data_5_entries_tag; // @[PageTableCache.scala 179:18]
  wire [15:0] l3_io_rresp_data_5_entries_asid; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_rresp_data_5_entries_ppns_0; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_rresp_data_5_entries_ppns_1; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_rresp_data_5_entries_ppns_2; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_rresp_data_5_entries_ppns_3; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_rresp_data_5_entries_ppns_4; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_rresp_data_5_entries_ppns_5; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_rresp_data_5_entries_ppns_6; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_rresp_data_5_entries_ppns_7; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_5_entries_vs_0; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_5_entries_vs_1; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_5_entries_vs_2; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_5_entries_vs_3; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_5_entries_vs_4; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_5_entries_vs_5; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_5_entries_vs_6; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_5_entries_vs_7; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_5_entries_perms_0_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_5_entries_perms_0_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_5_entries_perms_0_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_5_entries_perms_0_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_5_entries_perms_0_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_5_entries_perms_0_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_5_entries_perms_0_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_5_entries_perms_1_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_5_entries_perms_1_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_5_entries_perms_1_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_5_entries_perms_1_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_5_entries_perms_1_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_5_entries_perms_1_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_5_entries_perms_1_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_5_entries_perms_2_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_5_entries_perms_2_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_5_entries_perms_2_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_5_entries_perms_2_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_5_entries_perms_2_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_5_entries_perms_2_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_5_entries_perms_2_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_5_entries_perms_3_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_5_entries_perms_3_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_5_entries_perms_3_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_5_entries_perms_3_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_5_entries_perms_3_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_5_entries_perms_3_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_5_entries_perms_3_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_5_entries_perms_4_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_5_entries_perms_4_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_5_entries_perms_4_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_5_entries_perms_4_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_5_entries_perms_4_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_5_entries_perms_4_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_5_entries_perms_4_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_5_entries_perms_5_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_5_entries_perms_5_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_5_entries_perms_5_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_5_entries_perms_5_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_5_entries_perms_5_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_5_entries_perms_5_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_5_entries_perms_5_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_5_entries_perms_6_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_5_entries_perms_6_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_5_entries_perms_6_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_5_entries_perms_6_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_5_entries_perms_6_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_5_entries_perms_6_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_5_entries_perms_6_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_5_entries_perms_7_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_5_entries_perms_7_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_5_entries_perms_7_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_5_entries_perms_7_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_5_entries_perms_7_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_5_entries_perms_7_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_5_entries_perms_7_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_5_entries_prefetch; // @[PageTableCache.scala 179:18]
  wire [38:0] l3_io_rresp_data_5_ecc; // @[PageTableCache.scala 179:18]
  wire [21:0] l3_io_rresp_data_6_entries_tag; // @[PageTableCache.scala 179:18]
  wire [15:0] l3_io_rresp_data_6_entries_asid; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_rresp_data_6_entries_ppns_0; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_rresp_data_6_entries_ppns_1; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_rresp_data_6_entries_ppns_2; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_rresp_data_6_entries_ppns_3; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_rresp_data_6_entries_ppns_4; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_rresp_data_6_entries_ppns_5; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_rresp_data_6_entries_ppns_6; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_rresp_data_6_entries_ppns_7; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_6_entries_vs_0; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_6_entries_vs_1; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_6_entries_vs_2; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_6_entries_vs_3; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_6_entries_vs_4; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_6_entries_vs_5; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_6_entries_vs_6; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_6_entries_vs_7; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_6_entries_perms_0_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_6_entries_perms_0_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_6_entries_perms_0_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_6_entries_perms_0_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_6_entries_perms_0_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_6_entries_perms_0_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_6_entries_perms_0_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_6_entries_perms_1_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_6_entries_perms_1_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_6_entries_perms_1_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_6_entries_perms_1_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_6_entries_perms_1_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_6_entries_perms_1_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_6_entries_perms_1_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_6_entries_perms_2_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_6_entries_perms_2_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_6_entries_perms_2_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_6_entries_perms_2_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_6_entries_perms_2_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_6_entries_perms_2_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_6_entries_perms_2_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_6_entries_perms_3_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_6_entries_perms_3_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_6_entries_perms_3_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_6_entries_perms_3_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_6_entries_perms_3_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_6_entries_perms_3_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_6_entries_perms_3_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_6_entries_perms_4_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_6_entries_perms_4_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_6_entries_perms_4_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_6_entries_perms_4_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_6_entries_perms_4_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_6_entries_perms_4_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_6_entries_perms_4_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_6_entries_perms_5_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_6_entries_perms_5_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_6_entries_perms_5_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_6_entries_perms_5_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_6_entries_perms_5_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_6_entries_perms_5_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_6_entries_perms_5_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_6_entries_perms_6_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_6_entries_perms_6_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_6_entries_perms_6_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_6_entries_perms_6_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_6_entries_perms_6_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_6_entries_perms_6_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_6_entries_perms_6_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_6_entries_perms_7_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_6_entries_perms_7_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_6_entries_perms_7_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_6_entries_perms_7_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_6_entries_perms_7_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_6_entries_perms_7_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_6_entries_perms_7_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_6_entries_prefetch; // @[PageTableCache.scala 179:18]
  wire [38:0] l3_io_rresp_data_6_ecc; // @[PageTableCache.scala 179:18]
  wire [21:0] l3_io_rresp_data_7_entries_tag; // @[PageTableCache.scala 179:18]
  wire [15:0] l3_io_rresp_data_7_entries_asid; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_rresp_data_7_entries_ppns_0; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_rresp_data_7_entries_ppns_1; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_rresp_data_7_entries_ppns_2; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_rresp_data_7_entries_ppns_3; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_rresp_data_7_entries_ppns_4; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_rresp_data_7_entries_ppns_5; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_rresp_data_7_entries_ppns_6; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_rresp_data_7_entries_ppns_7; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_7_entries_vs_0; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_7_entries_vs_1; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_7_entries_vs_2; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_7_entries_vs_3; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_7_entries_vs_4; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_7_entries_vs_5; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_7_entries_vs_6; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_7_entries_vs_7; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_7_entries_perms_0_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_7_entries_perms_0_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_7_entries_perms_0_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_7_entries_perms_0_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_7_entries_perms_0_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_7_entries_perms_0_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_7_entries_perms_0_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_7_entries_perms_1_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_7_entries_perms_1_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_7_entries_perms_1_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_7_entries_perms_1_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_7_entries_perms_1_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_7_entries_perms_1_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_7_entries_perms_1_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_7_entries_perms_2_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_7_entries_perms_2_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_7_entries_perms_2_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_7_entries_perms_2_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_7_entries_perms_2_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_7_entries_perms_2_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_7_entries_perms_2_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_7_entries_perms_3_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_7_entries_perms_3_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_7_entries_perms_3_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_7_entries_perms_3_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_7_entries_perms_3_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_7_entries_perms_3_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_7_entries_perms_3_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_7_entries_perms_4_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_7_entries_perms_4_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_7_entries_perms_4_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_7_entries_perms_4_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_7_entries_perms_4_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_7_entries_perms_4_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_7_entries_perms_4_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_7_entries_perms_5_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_7_entries_perms_5_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_7_entries_perms_5_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_7_entries_perms_5_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_7_entries_perms_5_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_7_entries_perms_5_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_7_entries_perms_5_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_7_entries_perms_6_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_7_entries_perms_6_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_7_entries_perms_6_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_7_entries_perms_6_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_7_entries_perms_6_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_7_entries_perms_6_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_7_entries_perms_6_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_7_entries_perms_7_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_7_entries_perms_7_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_7_entries_perms_7_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_7_entries_perms_7_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_7_entries_perms_7_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_7_entries_perms_7_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_7_entries_perms_7_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_rresp_data_7_entries_prefetch; // @[PageTableCache.scala 179:18]
  wire [38:0] l3_io_rresp_data_7_ecc; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_valid; // @[PageTableCache.scala 179:18]
  wire [1:0] l3_io_wreq_bits_setIdx; // @[PageTableCache.scala 179:18]
  wire [21:0] l3_io_wreq_bits_data_0_entries_tag; // @[PageTableCache.scala 179:18]
  wire [15:0] l3_io_wreq_bits_data_0_entries_asid; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_wreq_bits_data_0_entries_ppns_0; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_wreq_bits_data_0_entries_ppns_1; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_wreq_bits_data_0_entries_ppns_2; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_wreq_bits_data_0_entries_ppns_3; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_wreq_bits_data_0_entries_ppns_4; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_wreq_bits_data_0_entries_ppns_5; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_wreq_bits_data_0_entries_ppns_6; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_wreq_bits_data_0_entries_ppns_7; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_0_entries_vs_0; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_0_entries_vs_1; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_0_entries_vs_2; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_0_entries_vs_3; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_0_entries_vs_4; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_0_entries_vs_5; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_0_entries_vs_6; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_0_entries_vs_7; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_0_entries_perms_0_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_0_entries_perms_0_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_0_entries_perms_0_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_0_entries_perms_0_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_0_entries_perms_0_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_0_entries_perms_0_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_0_entries_perms_0_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_0_entries_perms_1_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_0_entries_perms_1_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_0_entries_perms_1_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_0_entries_perms_1_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_0_entries_perms_1_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_0_entries_perms_1_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_0_entries_perms_1_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_0_entries_perms_2_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_0_entries_perms_2_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_0_entries_perms_2_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_0_entries_perms_2_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_0_entries_perms_2_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_0_entries_perms_2_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_0_entries_perms_2_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_0_entries_perms_3_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_0_entries_perms_3_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_0_entries_perms_3_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_0_entries_perms_3_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_0_entries_perms_3_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_0_entries_perms_3_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_0_entries_perms_3_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_0_entries_perms_4_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_0_entries_perms_4_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_0_entries_perms_4_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_0_entries_perms_4_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_0_entries_perms_4_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_0_entries_perms_4_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_0_entries_perms_4_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_0_entries_perms_5_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_0_entries_perms_5_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_0_entries_perms_5_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_0_entries_perms_5_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_0_entries_perms_5_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_0_entries_perms_5_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_0_entries_perms_5_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_0_entries_perms_6_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_0_entries_perms_6_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_0_entries_perms_6_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_0_entries_perms_6_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_0_entries_perms_6_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_0_entries_perms_6_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_0_entries_perms_6_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_0_entries_perms_7_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_0_entries_perms_7_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_0_entries_perms_7_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_0_entries_perms_7_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_0_entries_perms_7_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_0_entries_perms_7_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_0_entries_perms_7_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_0_entries_prefetch; // @[PageTableCache.scala 179:18]
  wire [38:0] l3_io_wreq_bits_data_0_ecc; // @[PageTableCache.scala 179:18]
  wire [21:0] l3_io_wreq_bits_data_1_entries_tag; // @[PageTableCache.scala 179:18]
  wire [15:0] l3_io_wreq_bits_data_1_entries_asid; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_wreq_bits_data_1_entries_ppns_0; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_wreq_bits_data_1_entries_ppns_1; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_wreq_bits_data_1_entries_ppns_2; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_wreq_bits_data_1_entries_ppns_3; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_wreq_bits_data_1_entries_ppns_4; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_wreq_bits_data_1_entries_ppns_5; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_wreq_bits_data_1_entries_ppns_6; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_wreq_bits_data_1_entries_ppns_7; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_1_entries_vs_0; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_1_entries_vs_1; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_1_entries_vs_2; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_1_entries_vs_3; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_1_entries_vs_4; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_1_entries_vs_5; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_1_entries_vs_6; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_1_entries_vs_7; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_1_entries_perms_0_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_1_entries_perms_0_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_1_entries_perms_0_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_1_entries_perms_0_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_1_entries_perms_0_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_1_entries_perms_0_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_1_entries_perms_0_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_1_entries_perms_1_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_1_entries_perms_1_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_1_entries_perms_1_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_1_entries_perms_1_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_1_entries_perms_1_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_1_entries_perms_1_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_1_entries_perms_1_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_1_entries_perms_2_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_1_entries_perms_2_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_1_entries_perms_2_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_1_entries_perms_2_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_1_entries_perms_2_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_1_entries_perms_2_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_1_entries_perms_2_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_1_entries_perms_3_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_1_entries_perms_3_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_1_entries_perms_3_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_1_entries_perms_3_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_1_entries_perms_3_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_1_entries_perms_3_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_1_entries_perms_3_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_1_entries_perms_4_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_1_entries_perms_4_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_1_entries_perms_4_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_1_entries_perms_4_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_1_entries_perms_4_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_1_entries_perms_4_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_1_entries_perms_4_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_1_entries_perms_5_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_1_entries_perms_5_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_1_entries_perms_5_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_1_entries_perms_5_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_1_entries_perms_5_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_1_entries_perms_5_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_1_entries_perms_5_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_1_entries_perms_6_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_1_entries_perms_6_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_1_entries_perms_6_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_1_entries_perms_6_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_1_entries_perms_6_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_1_entries_perms_6_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_1_entries_perms_6_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_1_entries_perms_7_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_1_entries_perms_7_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_1_entries_perms_7_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_1_entries_perms_7_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_1_entries_perms_7_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_1_entries_perms_7_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_1_entries_perms_7_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_1_entries_prefetch; // @[PageTableCache.scala 179:18]
  wire [38:0] l3_io_wreq_bits_data_1_ecc; // @[PageTableCache.scala 179:18]
  wire [21:0] l3_io_wreq_bits_data_2_entries_tag; // @[PageTableCache.scala 179:18]
  wire [15:0] l3_io_wreq_bits_data_2_entries_asid; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_wreq_bits_data_2_entries_ppns_0; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_wreq_bits_data_2_entries_ppns_1; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_wreq_bits_data_2_entries_ppns_2; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_wreq_bits_data_2_entries_ppns_3; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_wreq_bits_data_2_entries_ppns_4; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_wreq_bits_data_2_entries_ppns_5; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_wreq_bits_data_2_entries_ppns_6; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_wreq_bits_data_2_entries_ppns_7; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_2_entries_vs_0; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_2_entries_vs_1; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_2_entries_vs_2; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_2_entries_vs_3; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_2_entries_vs_4; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_2_entries_vs_5; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_2_entries_vs_6; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_2_entries_vs_7; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_2_entries_perms_0_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_2_entries_perms_0_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_2_entries_perms_0_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_2_entries_perms_0_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_2_entries_perms_0_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_2_entries_perms_0_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_2_entries_perms_0_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_2_entries_perms_1_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_2_entries_perms_1_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_2_entries_perms_1_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_2_entries_perms_1_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_2_entries_perms_1_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_2_entries_perms_1_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_2_entries_perms_1_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_2_entries_perms_2_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_2_entries_perms_2_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_2_entries_perms_2_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_2_entries_perms_2_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_2_entries_perms_2_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_2_entries_perms_2_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_2_entries_perms_2_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_2_entries_perms_3_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_2_entries_perms_3_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_2_entries_perms_3_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_2_entries_perms_3_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_2_entries_perms_3_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_2_entries_perms_3_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_2_entries_perms_3_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_2_entries_perms_4_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_2_entries_perms_4_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_2_entries_perms_4_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_2_entries_perms_4_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_2_entries_perms_4_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_2_entries_perms_4_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_2_entries_perms_4_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_2_entries_perms_5_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_2_entries_perms_5_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_2_entries_perms_5_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_2_entries_perms_5_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_2_entries_perms_5_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_2_entries_perms_5_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_2_entries_perms_5_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_2_entries_perms_6_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_2_entries_perms_6_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_2_entries_perms_6_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_2_entries_perms_6_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_2_entries_perms_6_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_2_entries_perms_6_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_2_entries_perms_6_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_2_entries_perms_7_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_2_entries_perms_7_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_2_entries_perms_7_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_2_entries_perms_7_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_2_entries_perms_7_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_2_entries_perms_7_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_2_entries_perms_7_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_2_entries_prefetch; // @[PageTableCache.scala 179:18]
  wire [38:0] l3_io_wreq_bits_data_2_ecc; // @[PageTableCache.scala 179:18]
  wire [21:0] l3_io_wreq_bits_data_3_entries_tag; // @[PageTableCache.scala 179:18]
  wire [15:0] l3_io_wreq_bits_data_3_entries_asid; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_wreq_bits_data_3_entries_ppns_0; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_wreq_bits_data_3_entries_ppns_1; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_wreq_bits_data_3_entries_ppns_2; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_wreq_bits_data_3_entries_ppns_3; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_wreq_bits_data_3_entries_ppns_4; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_wreq_bits_data_3_entries_ppns_5; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_wreq_bits_data_3_entries_ppns_6; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_wreq_bits_data_3_entries_ppns_7; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_3_entries_vs_0; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_3_entries_vs_1; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_3_entries_vs_2; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_3_entries_vs_3; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_3_entries_vs_4; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_3_entries_vs_5; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_3_entries_vs_6; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_3_entries_vs_7; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_3_entries_perms_0_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_3_entries_perms_0_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_3_entries_perms_0_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_3_entries_perms_0_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_3_entries_perms_0_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_3_entries_perms_0_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_3_entries_perms_0_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_3_entries_perms_1_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_3_entries_perms_1_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_3_entries_perms_1_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_3_entries_perms_1_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_3_entries_perms_1_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_3_entries_perms_1_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_3_entries_perms_1_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_3_entries_perms_2_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_3_entries_perms_2_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_3_entries_perms_2_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_3_entries_perms_2_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_3_entries_perms_2_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_3_entries_perms_2_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_3_entries_perms_2_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_3_entries_perms_3_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_3_entries_perms_3_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_3_entries_perms_3_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_3_entries_perms_3_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_3_entries_perms_3_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_3_entries_perms_3_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_3_entries_perms_3_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_3_entries_perms_4_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_3_entries_perms_4_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_3_entries_perms_4_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_3_entries_perms_4_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_3_entries_perms_4_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_3_entries_perms_4_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_3_entries_perms_4_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_3_entries_perms_5_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_3_entries_perms_5_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_3_entries_perms_5_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_3_entries_perms_5_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_3_entries_perms_5_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_3_entries_perms_5_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_3_entries_perms_5_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_3_entries_perms_6_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_3_entries_perms_6_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_3_entries_perms_6_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_3_entries_perms_6_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_3_entries_perms_6_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_3_entries_perms_6_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_3_entries_perms_6_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_3_entries_perms_7_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_3_entries_perms_7_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_3_entries_perms_7_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_3_entries_perms_7_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_3_entries_perms_7_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_3_entries_perms_7_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_3_entries_perms_7_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_3_entries_prefetch; // @[PageTableCache.scala 179:18]
  wire [38:0] l3_io_wreq_bits_data_3_ecc; // @[PageTableCache.scala 179:18]
  wire [21:0] l3_io_wreq_bits_data_4_entries_tag; // @[PageTableCache.scala 179:18]
  wire [15:0] l3_io_wreq_bits_data_4_entries_asid; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_wreq_bits_data_4_entries_ppns_0; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_wreq_bits_data_4_entries_ppns_1; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_wreq_bits_data_4_entries_ppns_2; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_wreq_bits_data_4_entries_ppns_3; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_wreq_bits_data_4_entries_ppns_4; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_wreq_bits_data_4_entries_ppns_5; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_wreq_bits_data_4_entries_ppns_6; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_wreq_bits_data_4_entries_ppns_7; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_4_entries_vs_0; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_4_entries_vs_1; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_4_entries_vs_2; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_4_entries_vs_3; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_4_entries_vs_4; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_4_entries_vs_5; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_4_entries_vs_6; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_4_entries_vs_7; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_4_entries_perms_0_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_4_entries_perms_0_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_4_entries_perms_0_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_4_entries_perms_0_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_4_entries_perms_0_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_4_entries_perms_0_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_4_entries_perms_0_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_4_entries_perms_1_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_4_entries_perms_1_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_4_entries_perms_1_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_4_entries_perms_1_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_4_entries_perms_1_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_4_entries_perms_1_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_4_entries_perms_1_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_4_entries_perms_2_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_4_entries_perms_2_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_4_entries_perms_2_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_4_entries_perms_2_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_4_entries_perms_2_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_4_entries_perms_2_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_4_entries_perms_2_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_4_entries_perms_3_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_4_entries_perms_3_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_4_entries_perms_3_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_4_entries_perms_3_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_4_entries_perms_3_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_4_entries_perms_3_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_4_entries_perms_3_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_4_entries_perms_4_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_4_entries_perms_4_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_4_entries_perms_4_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_4_entries_perms_4_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_4_entries_perms_4_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_4_entries_perms_4_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_4_entries_perms_4_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_4_entries_perms_5_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_4_entries_perms_5_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_4_entries_perms_5_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_4_entries_perms_5_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_4_entries_perms_5_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_4_entries_perms_5_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_4_entries_perms_5_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_4_entries_perms_6_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_4_entries_perms_6_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_4_entries_perms_6_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_4_entries_perms_6_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_4_entries_perms_6_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_4_entries_perms_6_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_4_entries_perms_6_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_4_entries_perms_7_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_4_entries_perms_7_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_4_entries_perms_7_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_4_entries_perms_7_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_4_entries_perms_7_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_4_entries_perms_7_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_4_entries_perms_7_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_4_entries_prefetch; // @[PageTableCache.scala 179:18]
  wire [38:0] l3_io_wreq_bits_data_4_ecc; // @[PageTableCache.scala 179:18]
  wire [21:0] l3_io_wreq_bits_data_5_entries_tag; // @[PageTableCache.scala 179:18]
  wire [15:0] l3_io_wreq_bits_data_5_entries_asid; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_wreq_bits_data_5_entries_ppns_0; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_wreq_bits_data_5_entries_ppns_1; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_wreq_bits_data_5_entries_ppns_2; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_wreq_bits_data_5_entries_ppns_3; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_wreq_bits_data_5_entries_ppns_4; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_wreq_bits_data_5_entries_ppns_5; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_wreq_bits_data_5_entries_ppns_6; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_wreq_bits_data_5_entries_ppns_7; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_5_entries_vs_0; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_5_entries_vs_1; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_5_entries_vs_2; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_5_entries_vs_3; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_5_entries_vs_4; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_5_entries_vs_5; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_5_entries_vs_6; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_5_entries_vs_7; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_5_entries_perms_0_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_5_entries_perms_0_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_5_entries_perms_0_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_5_entries_perms_0_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_5_entries_perms_0_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_5_entries_perms_0_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_5_entries_perms_0_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_5_entries_perms_1_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_5_entries_perms_1_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_5_entries_perms_1_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_5_entries_perms_1_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_5_entries_perms_1_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_5_entries_perms_1_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_5_entries_perms_1_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_5_entries_perms_2_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_5_entries_perms_2_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_5_entries_perms_2_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_5_entries_perms_2_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_5_entries_perms_2_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_5_entries_perms_2_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_5_entries_perms_2_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_5_entries_perms_3_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_5_entries_perms_3_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_5_entries_perms_3_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_5_entries_perms_3_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_5_entries_perms_3_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_5_entries_perms_3_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_5_entries_perms_3_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_5_entries_perms_4_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_5_entries_perms_4_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_5_entries_perms_4_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_5_entries_perms_4_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_5_entries_perms_4_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_5_entries_perms_4_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_5_entries_perms_4_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_5_entries_perms_5_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_5_entries_perms_5_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_5_entries_perms_5_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_5_entries_perms_5_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_5_entries_perms_5_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_5_entries_perms_5_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_5_entries_perms_5_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_5_entries_perms_6_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_5_entries_perms_6_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_5_entries_perms_6_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_5_entries_perms_6_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_5_entries_perms_6_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_5_entries_perms_6_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_5_entries_perms_6_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_5_entries_perms_7_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_5_entries_perms_7_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_5_entries_perms_7_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_5_entries_perms_7_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_5_entries_perms_7_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_5_entries_perms_7_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_5_entries_perms_7_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_5_entries_prefetch; // @[PageTableCache.scala 179:18]
  wire [38:0] l3_io_wreq_bits_data_5_ecc; // @[PageTableCache.scala 179:18]
  wire [21:0] l3_io_wreq_bits_data_6_entries_tag; // @[PageTableCache.scala 179:18]
  wire [15:0] l3_io_wreq_bits_data_6_entries_asid; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_wreq_bits_data_6_entries_ppns_0; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_wreq_bits_data_6_entries_ppns_1; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_wreq_bits_data_6_entries_ppns_2; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_wreq_bits_data_6_entries_ppns_3; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_wreq_bits_data_6_entries_ppns_4; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_wreq_bits_data_6_entries_ppns_5; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_wreq_bits_data_6_entries_ppns_6; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_wreq_bits_data_6_entries_ppns_7; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_6_entries_vs_0; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_6_entries_vs_1; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_6_entries_vs_2; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_6_entries_vs_3; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_6_entries_vs_4; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_6_entries_vs_5; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_6_entries_vs_6; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_6_entries_vs_7; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_6_entries_perms_0_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_6_entries_perms_0_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_6_entries_perms_0_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_6_entries_perms_0_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_6_entries_perms_0_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_6_entries_perms_0_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_6_entries_perms_0_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_6_entries_perms_1_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_6_entries_perms_1_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_6_entries_perms_1_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_6_entries_perms_1_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_6_entries_perms_1_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_6_entries_perms_1_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_6_entries_perms_1_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_6_entries_perms_2_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_6_entries_perms_2_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_6_entries_perms_2_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_6_entries_perms_2_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_6_entries_perms_2_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_6_entries_perms_2_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_6_entries_perms_2_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_6_entries_perms_3_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_6_entries_perms_3_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_6_entries_perms_3_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_6_entries_perms_3_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_6_entries_perms_3_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_6_entries_perms_3_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_6_entries_perms_3_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_6_entries_perms_4_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_6_entries_perms_4_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_6_entries_perms_4_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_6_entries_perms_4_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_6_entries_perms_4_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_6_entries_perms_4_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_6_entries_perms_4_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_6_entries_perms_5_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_6_entries_perms_5_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_6_entries_perms_5_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_6_entries_perms_5_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_6_entries_perms_5_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_6_entries_perms_5_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_6_entries_perms_5_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_6_entries_perms_6_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_6_entries_perms_6_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_6_entries_perms_6_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_6_entries_perms_6_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_6_entries_perms_6_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_6_entries_perms_6_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_6_entries_perms_6_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_6_entries_perms_7_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_6_entries_perms_7_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_6_entries_perms_7_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_6_entries_perms_7_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_6_entries_perms_7_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_6_entries_perms_7_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_6_entries_perms_7_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_6_entries_prefetch; // @[PageTableCache.scala 179:18]
  wire [38:0] l3_io_wreq_bits_data_6_ecc; // @[PageTableCache.scala 179:18]
  wire [21:0] l3_io_wreq_bits_data_7_entries_tag; // @[PageTableCache.scala 179:18]
  wire [15:0] l3_io_wreq_bits_data_7_entries_asid; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_wreq_bits_data_7_entries_ppns_0; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_wreq_bits_data_7_entries_ppns_1; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_wreq_bits_data_7_entries_ppns_2; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_wreq_bits_data_7_entries_ppns_3; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_wreq_bits_data_7_entries_ppns_4; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_wreq_bits_data_7_entries_ppns_5; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_wreq_bits_data_7_entries_ppns_6; // @[PageTableCache.scala 179:18]
  wire [23:0] l3_io_wreq_bits_data_7_entries_ppns_7; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_7_entries_vs_0; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_7_entries_vs_1; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_7_entries_vs_2; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_7_entries_vs_3; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_7_entries_vs_4; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_7_entries_vs_5; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_7_entries_vs_6; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_7_entries_vs_7; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_7_entries_perms_0_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_7_entries_perms_0_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_7_entries_perms_0_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_7_entries_perms_0_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_7_entries_perms_0_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_7_entries_perms_0_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_7_entries_perms_0_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_7_entries_perms_1_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_7_entries_perms_1_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_7_entries_perms_1_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_7_entries_perms_1_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_7_entries_perms_1_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_7_entries_perms_1_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_7_entries_perms_1_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_7_entries_perms_2_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_7_entries_perms_2_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_7_entries_perms_2_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_7_entries_perms_2_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_7_entries_perms_2_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_7_entries_perms_2_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_7_entries_perms_2_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_7_entries_perms_3_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_7_entries_perms_3_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_7_entries_perms_3_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_7_entries_perms_3_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_7_entries_perms_3_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_7_entries_perms_3_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_7_entries_perms_3_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_7_entries_perms_4_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_7_entries_perms_4_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_7_entries_perms_4_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_7_entries_perms_4_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_7_entries_perms_4_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_7_entries_perms_4_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_7_entries_perms_4_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_7_entries_perms_5_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_7_entries_perms_5_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_7_entries_perms_5_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_7_entries_perms_5_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_7_entries_perms_5_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_7_entries_perms_5_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_7_entries_perms_5_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_7_entries_perms_6_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_7_entries_perms_6_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_7_entries_perms_6_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_7_entries_perms_6_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_7_entries_perms_6_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_7_entries_perms_6_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_7_entries_perms_6_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_7_entries_perms_7_d; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_7_entries_perms_7_a; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_7_entries_perms_7_g; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_7_entries_perms_7_u; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_7_entries_perms_7_x; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_7_entries_perms_7_w; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_7_entries_perms_7_r; // @[PageTableCache.scala 179:18]
  wire  l3_io_wreq_bits_data_7_entries_prefetch; // @[PageTableCache.scala 179:18]
  wire [38:0] l3_io_wreq_bits_data_7_ecc; // @[PageTableCache.scala 179:18]
  wire [7:0] l3_io_wreq_bits_waymask; // @[PageTableCache.scala 179:18]
  wire  refill_prefetch_dup_0 = io_refill_bits_req_info_dup_0_source == 2'h2; // @[MMUConst.scala 254:13]
  wire  refill_prefetch_dup_1 = io_refill_bits_req_info_dup_1_source == 2'h2; // @[MMUConst.scala 254:13]
  wire  refill_prefetch_dup_2 = io_refill_bits_req_info_dup_2_source == 2'h2; // @[MMUConst.scala 254:13]
  wire  flush = io_sfence_dup_0_valid | io_csr_dup_0_satp_changed; // @[PageTableCache.scala 122:66]
  wire  flush_dup_1 = io_sfence_dup_1_valid | io_csr_dup_1_satp_changed; // @[PageTableCache.scala 122:66]
  wire  flush_dup_2 = io_sfence_dup_2_valid | io_csr_dup_2_satp_changed; // @[PageTableCache.scala 122:66]
  reg  valid; // @[PipelineConnect.scala 108:24]
  reg  valid_1; // @[PipelineConnect.scala 108:24]
  reg  valid_2; // @[PipelineConnect.scala 108:24]
  wire  stageResp_ready = ~valid_2 | io_resp_ready; // @[PageTableCache.scala 146:39]
  wire  stageCheck_0_ready = ~valid_1 | stageResp_ready; // @[PageTableCache.scala 653:27]
  wire  stageDelay_0_ready = ~valid | stageCheck_0_ready; // @[PageTableCache.scala 653:27]
  wire  _stageReq_ready_T = ~io_refill_valid; // @[PipelineConnect.scala 114:34]
  wire  stageReq_ready = stageDelay_0_ready & ~io_refill_valid; // @[PipelineConnect.scala 114:31]
  wire  _stageDelay_valid_1cycle_T = stageReq_ready & io_req_valid; // @[Decoupled.scala 50:35]
  reg  stageDelay_valid_1cycle; // @[Hold.scala 54:24]
  wire  _GEN_0 = stageDelay_valid_1cycle ? 1'h0 : stageDelay_valid_1cycle; // @[Hold.scala 55:18 54:24 55:26]
  wire  _GEN_1 = _stageDelay_valid_1cycle_T | _GEN_0; // @[Hold.scala 56:{17,25}]
  wire  _stageCheck_valid_1cycle_T = stageCheck_0_ready & valid; // @[Decoupled.scala 50:35]
  reg  stageCheck_valid_1cycle; // @[Hold.scala 54:24]
  wire  _GEN_3 = stageCheck_valid_1cycle ? 1'h0 : stageCheck_valid_1cycle; // @[Hold.scala 55:18 54:24 55:26]
  wire  _GEN_4 = _stageCheck_valid_1cycle_T | _GEN_3; // @[Hold.scala 56:{17,25}]
  wire  _stageResp_valid_1cycle_dup_0_T = stageResp_ready & valid_1; // @[Decoupled.scala 50:35]
  reg  stageResp_valid_1cycle_dup_0_valid; // @[Hold.scala 54:24]
  wire  _GEN_6 = stageResp_valid_1cycle_dup_0_valid ? 1'h0 : stageResp_valid_1cycle_dup_0_valid; // @[Hold.scala 55:18 54:24 55:26]
  wire  _GEN_7 = _stageResp_valid_1cycle_dup_0_T | _GEN_6; // @[Hold.scala 56:{17,25}]
  reg  stageResp_valid_1cycle_dup_1_valid; // @[Hold.scala 54:24]
  wire  _GEN_9 = stageResp_valid_1cycle_dup_1_valid ? 1'h0 : stageResp_valid_1cycle_dup_1_valid; // @[Hold.scala 55:18 54:24 55:26]
  wire  _GEN_10 = _stageResp_valid_1cycle_dup_0_T | _GEN_9; // @[Hold.scala 56:{17,25}]
  wire  leftFire = io_req_valid & stageDelay_0_ready & _stageReq_ready_T; // @[PipelineConnect.scala 109:46]
  wire  _GEN_12 = stageCheck_0_ready ? 1'h0 : valid; // @[PipelineConnect.scala 108:24 110:{25,33}]
  wire  _GEN_13 = leftFire | _GEN_12; // @[PipelineConnect.scala 111:{21,29}]
  reg [26:0] data_req_info_vpn; // @[Reg.scala 16:16]
  reg [1:0] data_req_info_source; // @[Reg.scala 16:16]
  reg  data_isFirst; // @[Reg.scala 16:16]
  reg  bypassed_reg; // @[PageTableCache.scala 657:29]
  wire  _bypassed_wire_T_4 = io_refill_bits_req_info_dup_0_vpn[26:21] == data_req_info_vpn[26:21]; // @[PageTableCache.scala 221:44]
  wire  _bypassed_wire_T_5 = io_refill_valid & 2'h0 == io_refill_bits_level_dup_0 & _bypassed_wire_T_4; // @[PageTableCache.scala 225:66]
  wire  bypassed_wire = _bypassed_wire_T_5 & io_refill_valid; // @[PageTableCache.scala 658:66]
  wire  stageDelay_1_bits_bypassed_0 = bypassed_wire | bypassed_reg & ~stageDelay_valid_1cycle; // @[PageTableCache.scala 662:38]
  reg  bypassed_reg_1; // @[PageTableCache.scala 657:29]
  wire  _bypassed_wire_T_10 = io_refill_bits_req_info_dup_0_vpn[26:12] == data_req_info_vpn[26:12]; // @[PageTableCache.scala 221:44]
  wire  _bypassed_wire_T_11 = io_refill_valid & 2'h1 == io_refill_bits_level_dup_0 & _bypassed_wire_T_10; // @[PageTableCache.scala 225:66]
  wire  bypassed_wire_1 = _bypassed_wire_T_11 & io_refill_valid; // @[PageTableCache.scala 658:66]
  wire  stageDelay_1_bits_bypassed_1 = bypassed_wire_1 | bypassed_reg_1 & ~stageDelay_valid_1cycle; // @[PageTableCache.scala 662:38]
  reg  bypassed_reg_2; // @[PageTableCache.scala 657:29]
  wire  _bypassed_wire_T_16 = io_refill_bits_req_info_dup_0_vpn[26:3] == data_req_info_vpn[26:3]; // @[PageTableCache.scala 221:44]
  wire  _bypassed_wire_T_17 = io_refill_valid & 2'h2 == io_refill_bits_level_dup_0 & _bypassed_wire_T_16; // @[PageTableCache.scala 225:66]
  wire  bypassed_wire_2 = _bypassed_wire_T_17 & io_refill_valid; // @[PageTableCache.scala 658:66]
  wire  stageDelay_1_bits_bypassed_2 = bypassed_wire_2 | bypassed_reg_2 & ~stageDelay_valid_1cycle; // @[PageTableCache.scala 662:38]
  wire  leftFire_1 = valid & stageCheck_0_ready; // @[PipelineConnect.scala 109:31]
  wire  _GEN_27 = stageResp_ready ? 1'h0 : valid_1; // @[PipelineConnect.scala 108:24 110:{25,33}]
  wire  _GEN_28 = leftFire_1 | _GEN_27; // @[PipelineConnect.scala 111:{21,29}]
  reg [26:0] data_1_req_info_vpn; // @[Reg.scala 16:16]
  reg [1:0] data_1_req_info_source; // @[Reg.scala 16:16]
  reg  data_1_isFirst; // @[Reg.scala 16:16]
  reg  data_1_bypassed_0; // @[Reg.scala 16:16]
  reg  data_1_bypassed_1; // @[Reg.scala 16:16]
  reg  data_1_bypassed_2; // @[Reg.scala 16:16]
  reg  bypassed_reg_3; // @[PageTableCache.scala 657:29]
  wire  _bypassed_wire_T_22 = io_refill_bits_req_info_dup_0_vpn[26:21] == data_1_req_info_vpn[26:21]; // @[PageTableCache.scala 221:44]
  wire  _bypassed_wire_T_23 = io_refill_valid & 2'h0 == io_refill_bits_level_dup_0 & _bypassed_wire_T_22; // @[PageTableCache.scala 225:66]
  wire  bypassed_wire_3 = _bypassed_wire_T_23 & io_refill_valid; // @[PageTableCache.scala 658:66]
  wire  stageCheck_1_bits_bypassed_0 = data_1_bypassed_0 | (bypassed_wire_3 | bypassed_reg_3 & ~stageCheck_valid_1cycle)
    ; // @[PageTableCache.scala 662:20]
  reg  bypassed_reg_4; // @[PageTableCache.scala 657:29]
  wire  _bypassed_wire_T_28 = io_refill_bits_req_info_dup_0_vpn[26:12] == data_1_req_info_vpn[26:12]; // @[PageTableCache.scala 221:44]
  wire  _bypassed_wire_T_29 = io_refill_valid & 2'h1 == io_refill_bits_level_dup_0 & _bypassed_wire_T_28; // @[PageTableCache.scala 225:66]
  wire  bypassed_wire_4 = _bypassed_wire_T_29 & io_refill_valid; // @[PageTableCache.scala 658:66]
  wire  stageCheck_1_bits_bypassed_1 = data_1_bypassed_1 | (bypassed_wire_4 | bypassed_reg_4 & ~stageCheck_valid_1cycle)
    ; // @[PageTableCache.scala 662:20]
  reg  bypassed_reg_5; // @[PageTableCache.scala 657:29]
  wire  _bypassed_wire_T_34 = io_refill_bits_req_info_dup_0_vpn[26:3] == data_1_req_info_vpn[26:3]; // @[PageTableCache.scala 221:44]
  wire  _bypassed_wire_T_35 = io_refill_valid & 2'h2 == io_refill_bits_level_dup_0 & _bypassed_wire_T_34; // @[PageTableCache.scala 225:66]
  wire  bypassed_wire_5 = _bypassed_wire_T_35 & io_refill_valid; // @[PageTableCache.scala 658:66]
  wire  stageCheck_1_bits_bypassed_2 = data_1_bypassed_2 | (bypassed_wire_5 | bypassed_reg_5 & ~stageCheck_valid_1cycle)
    ; // @[PageTableCache.scala 662:20]
  wire  leftFire_2 = valid_1 & stageResp_ready; // @[PipelineConnect.scala 109:31]
  wire  _GEN_42 = io_resp_ready ? 1'h0 : valid_2; // @[PipelineConnect.scala 108:24 110:{25,33}]
  wire  _GEN_43 = leftFire_2 | _GEN_42; // @[PipelineConnect.scala 111:{21,29}]
  reg [26:0] data_2_req_info_vpn; // @[Reg.scala 16:16]
  reg [1:0] data_2_req_info_source; // @[Reg.scala 16:16]
  reg  data_2_isFirst; // @[Reg.scala 16:16]
  reg  data_2_bypassed_0; // @[Reg.scala 16:16]
  reg  data_2_bypassed_1; // @[Reg.scala 16:16]
  reg  data_2_bypassed_2; // @[Reg.scala 16:16]
  reg [8:0] l1_0_tag; // @[PageTableCache.scala 149:15]
  reg [15:0] l1_0_asid; // @[PageTableCache.scala 149:15]
  reg [23:0] l1_0_ppn; // @[PageTableCache.scala 149:15]
  reg [8:0] l1_1_tag; // @[PageTableCache.scala 149:15]
  reg [15:0] l1_1_asid; // @[PageTableCache.scala 149:15]
  reg [23:0] l1_1_ppn; // @[PageTableCache.scala 149:15]
  reg [8:0] l1_2_tag; // @[PageTableCache.scala 149:15]
  reg [15:0] l1_2_asid; // @[PageTableCache.scala 149:15]
  reg [23:0] l1_2_ppn; // @[PageTableCache.scala 149:15]
  reg [8:0] l1_3_tag; // @[PageTableCache.scala 149:15]
  reg [15:0] l1_3_asid; // @[PageTableCache.scala 149:15]
  reg [23:0] l1_3_ppn; // @[PageTableCache.scala 149:15]
  reg [3:0] l1v; // @[PageTableCache.scala 150:20]
  reg [3:0] l1g; // @[PageTableCache.scala 151:16]
  reg [15:0] l2v; // @[PageTableCache.scala 161:20]
  reg [15:0] l2g; // @[PageTableCache.scala 162:16]
  reg [31:0] l3v; // @[PageTableCache.scala 185:20]
  reg [31:0] l3g; // @[PageTableCache.scala 186:16]
  reg [17:0] sp_0_tag; // @[PageTableCache.scala 203:15]
  reg [15:0] sp_0_asid; // @[PageTableCache.scala 203:15]
  reg [23:0] sp_0_ppn; // @[PageTableCache.scala 203:15]
  reg  sp_0_perm_d; // @[PageTableCache.scala 203:15]
  reg  sp_0_perm_a; // @[PageTableCache.scala 203:15]
  reg  sp_0_perm_g; // @[PageTableCache.scala 203:15]
  reg  sp_0_perm_u; // @[PageTableCache.scala 203:15]
  reg  sp_0_perm_x; // @[PageTableCache.scala 203:15]
  reg  sp_0_perm_w; // @[PageTableCache.scala 203:15]
  reg  sp_0_perm_r; // @[PageTableCache.scala 203:15]
  reg [1:0] sp_0_level; // @[PageTableCache.scala 203:15]
  reg  sp_0_prefetch; // @[PageTableCache.scala 203:15]
  reg  sp_0_v; // @[PageTableCache.scala 203:15]
  reg [17:0] sp_1_tag; // @[PageTableCache.scala 203:15]
  reg [15:0] sp_1_asid; // @[PageTableCache.scala 203:15]
  reg [23:0] sp_1_ppn; // @[PageTableCache.scala 203:15]
  reg  sp_1_perm_d; // @[PageTableCache.scala 203:15]
  reg  sp_1_perm_a; // @[PageTableCache.scala 203:15]
  reg  sp_1_perm_g; // @[PageTableCache.scala 203:15]
  reg  sp_1_perm_u; // @[PageTableCache.scala 203:15]
  reg  sp_1_perm_x; // @[PageTableCache.scala 203:15]
  reg  sp_1_perm_w; // @[PageTableCache.scala 203:15]
  reg  sp_1_perm_r; // @[PageTableCache.scala 203:15]
  reg [1:0] sp_1_level; // @[PageTableCache.scala 203:15]
  reg  sp_1_prefetch; // @[PageTableCache.scala 203:15]
  reg  sp_1_v; // @[PageTableCache.scala 203:15]
  reg [1:0] spv; // @[PageTableCache.scala 204:20]
  reg [1:0] spg; // @[PageTableCache.scala 205:16]
  reg [2:0] state_reg; // @[Replacement.scala 168:70]
  wire  asid_hit = l1_0_asid == io_csr_dup_0_satp_asid; // @[MMUBundle.scala 578:59]
  wire  _T_2 = asid_hit & l1_0_tag == io_req_bits_req_info_vpn[26:18]; // @[MMUBundle.scala 592:16]
  wire  l1_hitVecT_0 = _T_2 & l1v[0]; // @[PageTableCache.scala 231:115]
  wire  asid_hit_1 = l1_1_asid == io_csr_dup_0_satp_asid; // @[MMUBundle.scala 578:59]
  wire  _T_7 = asid_hit_1 & l1_1_tag == io_req_bits_req_info_vpn[26:18]; // @[MMUBundle.scala 592:16]
  wire  l1_hitVecT_1 = _T_7 & l1v[1]; // @[PageTableCache.scala 231:115]
  wire  asid_hit_2 = l1_2_asid == io_csr_dup_0_satp_asid; // @[MMUBundle.scala 578:59]
  wire  _T_12 = asid_hit_2 & l1_2_tag == io_req_bits_req_info_vpn[26:18]; // @[MMUBundle.scala 592:16]
  wire  l1_hitVecT_2 = _T_12 & l1v[2]; // @[PageTableCache.scala 231:115]
  wire  asid_hit_3 = l1_3_asid == io_csr_dup_0_satp_asid; // @[MMUBundle.scala 578:59]
  wire  _T_17 = asid_hit_3 & l1_3_tag == io_req_bits_req_info_vpn[26:18]; // @[MMUBundle.scala 592:16]
  wire  l1_hitVecT_3 = _T_17 & l1v[3]; // @[PageTableCache.scala 231:115]
  reg  r; // @[Reg.scala 16:16]
  reg  r_1; // @[Reg.scala 16:16]
  reg  r_2; // @[Reg.scala 16:16]
  reg  r_3; // @[Reg.scala 16:16]
  wire  _T_28 = r | r_1 | (r_2 | r_3); // @[ParallelMux.scala 90:65]
  reg [23:0] r_4; // @[Reg.scala 16:16]
  reg  r_6; // @[Reg.scala 16:16]
  wire  _GEN_57 = stageDelay_valid_1cycle ? _T_28 : r_6; // @[Reg.scala 16:16 17:{18,22}]
  wire [3:0] _T_43 = {r_3,r_2,r_1,r}; // @[Cat.scala 31:58]
  wire [1:0] hi_1 = _T_43[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] lo_1 = _T_43[1:0]; // @[OneHot.scala 31:18]
  wire  _T_44 = |hi_1; // @[OneHot.scala 32:14]
  wire [1:0] _T_45 = hi_1 | lo_1; // @[OneHot.scala 32:28]
  wire [1:0] state_reg_touch_way_sized = {_T_44,_T_45[1]}; // @[Cat.scala 31:58]
  wire  state_reg_set_left_older = ~state_reg_touch_way_sized[1]; // @[Replacement.scala 196:33]
  wire  state_reg_left_subtree_state = state_reg[1]; // @[package.scala 154:13]
  wire  state_reg_right_subtree_state = state_reg[0]; // @[Replacement.scala 198:38]
  wire  _state_reg_T_2 = ~state_reg_touch_way_sized[0]; // @[Replacement.scala 218:7]
  wire  _state_reg_T_3 = state_reg_set_left_older ? state_reg_left_subtree_state : _state_reg_T_2; // @[Replacement.scala 203:16]
  wire  _state_reg_T_7 = state_reg_set_left_older ? _state_reg_T_2 : state_reg_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_reg_T_8 = {state_reg_set_left_older,_state_reg_T_3,_state_reg_T_7}; // @[Cat.scala 31:58]
  reg  l1Hit; // @[Reg.scala 16:16]
  reg [23:0] l1HitPPN; // @[Reg.scala 16:16]
  reg [2:0] state_vec__0; // @[Replacement.scala 305:17]
  reg [2:0] state_vec__1; // @[Replacement.scala 305:17]
  reg [2:0] state_vec__2; // @[Replacement.scala 305:17]
  reg [2:0] state_vec__3; // @[Replacement.scala 305:17]
  wire [1:0] l2_ridx = io_req_bits_req_info_vpn[13:12]; // @[MMUConst.scala 210:21]
  wire [3:0] l2vVec_0 = l2v[3:0]; // @[PageTableCache.scala 168:30]
  wire [3:0] l2vVec_1 = l2v[7:4]; // @[PageTableCache.scala 168:30]
  wire [3:0] l2vVec_2 = l2v[11:8]; // @[PageTableCache.scala 168:30]
  wire [3:0] l2vVec_3 = l2v[15:12]; // @[PageTableCache.scala 168:30]
  reg [12:0] r_7_0_entries_tag; // @[Reg.scala 16:16]
  reg [15:0] r_7_0_entries_asid; // @[Reg.scala 16:16]
  reg [23:0] r_7_0_entries_ppns_0; // @[Reg.scala 16:16]
  reg [23:0] r_7_0_entries_ppns_1; // @[Reg.scala 16:16]
  reg [23:0] r_7_0_entries_ppns_2; // @[Reg.scala 16:16]
  reg [23:0] r_7_0_entries_ppns_3; // @[Reg.scala 16:16]
  reg [23:0] r_7_0_entries_ppns_4; // @[Reg.scala 16:16]
  reg [23:0] r_7_0_entries_ppns_5; // @[Reg.scala 16:16]
  reg [23:0] r_7_0_entries_ppns_6; // @[Reg.scala 16:16]
  reg [23:0] r_7_0_entries_ppns_7; // @[Reg.scala 16:16]
  reg  r_7_0_entries_vs_0; // @[Reg.scala 16:16]
  reg  r_7_0_entries_vs_1; // @[Reg.scala 16:16]
  reg  r_7_0_entries_vs_2; // @[Reg.scala 16:16]
  reg  r_7_0_entries_vs_3; // @[Reg.scala 16:16]
  reg  r_7_0_entries_vs_4; // @[Reg.scala 16:16]
  reg  r_7_0_entries_vs_5; // @[Reg.scala 16:16]
  reg  r_7_0_entries_vs_6; // @[Reg.scala 16:16]
  reg  r_7_0_entries_vs_7; // @[Reg.scala 16:16]
  reg  r_7_0_entries_prefetch; // @[Reg.scala 16:16]
  reg [30:0] r_7_0_ecc; // @[Reg.scala 16:16]
  reg [12:0] r_7_1_entries_tag; // @[Reg.scala 16:16]
  reg [15:0] r_7_1_entries_asid; // @[Reg.scala 16:16]
  reg [23:0] r_7_1_entries_ppns_0; // @[Reg.scala 16:16]
  reg [23:0] r_7_1_entries_ppns_1; // @[Reg.scala 16:16]
  reg [23:0] r_7_1_entries_ppns_2; // @[Reg.scala 16:16]
  reg [23:0] r_7_1_entries_ppns_3; // @[Reg.scala 16:16]
  reg [23:0] r_7_1_entries_ppns_4; // @[Reg.scala 16:16]
  reg [23:0] r_7_1_entries_ppns_5; // @[Reg.scala 16:16]
  reg [23:0] r_7_1_entries_ppns_6; // @[Reg.scala 16:16]
  reg [23:0] r_7_1_entries_ppns_7; // @[Reg.scala 16:16]
  reg  r_7_1_entries_vs_0; // @[Reg.scala 16:16]
  reg  r_7_1_entries_vs_1; // @[Reg.scala 16:16]
  reg  r_7_1_entries_vs_2; // @[Reg.scala 16:16]
  reg  r_7_1_entries_vs_3; // @[Reg.scala 16:16]
  reg  r_7_1_entries_vs_4; // @[Reg.scala 16:16]
  reg  r_7_1_entries_vs_5; // @[Reg.scala 16:16]
  reg  r_7_1_entries_vs_6; // @[Reg.scala 16:16]
  reg  r_7_1_entries_vs_7; // @[Reg.scala 16:16]
  reg  r_7_1_entries_prefetch; // @[Reg.scala 16:16]
  reg [30:0] r_7_1_ecc; // @[Reg.scala 16:16]
  reg [12:0] r_7_2_entries_tag; // @[Reg.scala 16:16]
  reg [15:0] r_7_2_entries_asid; // @[Reg.scala 16:16]
  reg [23:0] r_7_2_entries_ppns_0; // @[Reg.scala 16:16]
  reg [23:0] r_7_2_entries_ppns_1; // @[Reg.scala 16:16]
  reg [23:0] r_7_2_entries_ppns_2; // @[Reg.scala 16:16]
  reg [23:0] r_7_2_entries_ppns_3; // @[Reg.scala 16:16]
  reg [23:0] r_7_2_entries_ppns_4; // @[Reg.scala 16:16]
  reg [23:0] r_7_2_entries_ppns_5; // @[Reg.scala 16:16]
  reg [23:0] r_7_2_entries_ppns_6; // @[Reg.scala 16:16]
  reg [23:0] r_7_2_entries_ppns_7; // @[Reg.scala 16:16]
  reg  r_7_2_entries_vs_0; // @[Reg.scala 16:16]
  reg  r_7_2_entries_vs_1; // @[Reg.scala 16:16]
  reg  r_7_2_entries_vs_2; // @[Reg.scala 16:16]
  reg  r_7_2_entries_vs_3; // @[Reg.scala 16:16]
  reg  r_7_2_entries_vs_4; // @[Reg.scala 16:16]
  reg  r_7_2_entries_vs_5; // @[Reg.scala 16:16]
  reg  r_7_2_entries_vs_6; // @[Reg.scala 16:16]
  reg  r_7_2_entries_vs_7; // @[Reg.scala 16:16]
  reg  r_7_2_entries_prefetch; // @[Reg.scala 16:16]
  reg [30:0] r_7_2_ecc; // @[Reg.scala 16:16]
  reg [12:0] r_7_3_entries_tag; // @[Reg.scala 16:16]
  reg [15:0] r_7_3_entries_asid; // @[Reg.scala 16:16]
  reg [23:0] r_7_3_entries_ppns_0; // @[Reg.scala 16:16]
  reg [23:0] r_7_3_entries_ppns_1; // @[Reg.scala 16:16]
  reg [23:0] r_7_3_entries_ppns_2; // @[Reg.scala 16:16]
  reg [23:0] r_7_3_entries_ppns_3; // @[Reg.scala 16:16]
  reg [23:0] r_7_3_entries_ppns_4; // @[Reg.scala 16:16]
  reg [23:0] r_7_3_entries_ppns_5; // @[Reg.scala 16:16]
  reg [23:0] r_7_3_entries_ppns_6; // @[Reg.scala 16:16]
  reg [23:0] r_7_3_entries_ppns_7; // @[Reg.scala 16:16]
  reg  r_7_3_entries_vs_0; // @[Reg.scala 16:16]
  reg  r_7_3_entries_vs_1; // @[Reg.scala 16:16]
  reg  r_7_3_entries_vs_2; // @[Reg.scala 16:16]
  reg  r_7_3_entries_vs_3; // @[Reg.scala 16:16]
  reg  r_7_3_entries_vs_4; // @[Reg.scala 16:16]
  reg  r_7_3_entries_vs_5; // @[Reg.scala 16:16]
  reg  r_7_3_entries_vs_6; // @[Reg.scala 16:16]
  reg  r_7_3_entries_vs_7; // @[Reg.scala 16:16]
  reg  r_7_3_entries_prefetch; // @[Reg.scala 16:16]
  reg [30:0] r_7_3_ecc; // @[Reg.scala 16:16]
  wire [12:0] _GEN_62 = stageDelay_valid_1cycle ? l2_io_rresp_data_0_entries_tag : r_7_0_entries_tag; // @[Reg.scala 16:16 17:{18,22}]
  wire [15:0] _GEN_63 = stageDelay_valid_1cycle ? l2_io_rresp_data_0_entries_asid : r_7_0_entries_asid; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_72 = stageDelay_valid_1cycle ? l2_io_rresp_data_0_entries_vs_0 : r_7_0_entries_vs_0; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_73 = stageDelay_valid_1cycle ? l2_io_rresp_data_0_entries_vs_1 : r_7_0_entries_vs_1; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_74 = stageDelay_valid_1cycle ? l2_io_rresp_data_0_entries_vs_2 : r_7_0_entries_vs_2; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_75 = stageDelay_valid_1cycle ? l2_io_rresp_data_0_entries_vs_3 : r_7_0_entries_vs_3; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_76 = stageDelay_valid_1cycle ? l2_io_rresp_data_0_entries_vs_4 : r_7_0_entries_vs_4; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_77 = stageDelay_valid_1cycle ? l2_io_rresp_data_0_entries_vs_5 : r_7_0_entries_vs_5; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_78 = stageDelay_valid_1cycle ? l2_io_rresp_data_0_entries_vs_6 : r_7_0_entries_vs_6; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_79 = stageDelay_valid_1cycle ? l2_io_rresp_data_0_entries_vs_7 : r_7_0_entries_vs_7; // @[Reg.scala 16:16 17:{18,22}]
  wire [12:0] _GEN_82 = stageDelay_valid_1cycle ? l2_io_rresp_data_1_entries_tag : r_7_1_entries_tag; // @[Reg.scala 16:16 17:{18,22}]
  wire [15:0] _GEN_83 = stageDelay_valid_1cycle ? l2_io_rresp_data_1_entries_asid : r_7_1_entries_asid; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_92 = stageDelay_valid_1cycle ? l2_io_rresp_data_1_entries_vs_0 : r_7_1_entries_vs_0; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_93 = stageDelay_valid_1cycle ? l2_io_rresp_data_1_entries_vs_1 : r_7_1_entries_vs_1; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_94 = stageDelay_valid_1cycle ? l2_io_rresp_data_1_entries_vs_2 : r_7_1_entries_vs_2; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_95 = stageDelay_valid_1cycle ? l2_io_rresp_data_1_entries_vs_3 : r_7_1_entries_vs_3; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_96 = stageDelay_valid_1cycle ? l2_io_rresp_data_1_entries_vs_4 : r_7_1_entries_vs_4; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_97 = stageDelay_valid_1cycle ? l2_io_rresp_data_1_entries_vs_5 : r_7_1_entries_vs_5; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_98 = stageDelay_valid_1cycle ? l2_io_rresp_data_1_entries_vs_6 : r_7_1_entries_vs_6; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_99 = stageDelay_valid_1cycle ? l2_io_rresp_data_1_entries_vs_7 : r_7_1_entries_vs_7; // @[Reg.scala 16:16 17:{18,22}]
  wire [12:0] _GEN_102 = stageDelay_valid_1cycle ? l2_io_rresp_data_2_entries_tag : r_7_2_entries_tag; // @[Reg.scala 16:16 17:{18,22}]
  wire [15:0] _GEN_103 = stageDelay_valid_1cycle ? l2_io_rresp_data_2_entries_asid : r_7_2_entries_asid; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_112 = stageDelay_valid_1cycle ? l2_io_rresp_data_2_entries_vs_0 : r_7_2_entries_vs_0; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_113 = stageDelay_valid_1cycle ? l2_io_rresp_data_2_entries_vs_1 : r_7_2_entries_vs_1; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_114 = stageDelay_valid_1cycle ? l2_io_rresp_data_2_entries_vs_2 : r_7_2_entries_vs_2; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_115 = stageDelay_valid_1cycle ? l2_io_rresp_data_2_entries_vs_3 : r_7_2_entries_vs_3; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_116 = stageDelay_valid_1cycle ? l2_io_rresp_data_2_entries_vs_4 : r_7_2_entries_vs_4; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_117 = stageDelay_valid_1cycle ? l2_io_rresp_data_2_entries_vs_5 : r_7_2_entries_vs_5; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_118 = stageDelay_valid_1cycle ? l2_io_rresp_data_2_entries_vs_6 : r_7_2_entries_vs_6; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_119 = stageDelay_valid_1cycle ? l2_io_rresp_data_2_entries_vs_7 : r_7_2_entries_vs_7; // @[Reg.scala 16:16 17:{18,22}]
  wire [12:0] _GEN_122 = stageDelay_valid_1cycle ? l2_io_rresp_data_3_entries_tag : r_7_3_entries_tag; // @[Reg.scala 16:16 17:{18,22}]
  wire [15:0] _GEN_123 = stageDelay_valid_1cycle ? l2_io_rresp_data_3_entries_asid : r_7_3_entries_asid; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_132 = stageDelay_valid_1cycle ? l2_io_rresp_data_3_entries_vs_0 : r_7_3_entries_vs_0; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_133 = stageDelay_valid_1cycle ? l2_io_rresp_data_3_entries_vs_1 : r_7_3_entries_vs_1; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_134 = stageDelay_valid_1cycle ? l2_io_rresp_data_3_entries_vs_2 : r_7_3_entries_vs_2; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_135 = stageDelay_valid_1cycle ? l2_io_rresp_data_3_entries_vs_3 : r_7_3_entries_vs_3; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_136 = stageDelay_valid_1cycle ? l2_io_rresp_data_3_entries_vs_4 : r_7_3_entries_vs_4; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_137 = stageDelay_valid_1cycle ? l2_io_rresp_data_3_entries_vs_5 : r_7_3_entries_vs_5; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_138 = stageDelay_valid_1cycle ? l2_io_rresp_data_3_entries_vs_6 : r_7_3_entries_vs_6; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_139 = stageDelay_valid_1cycle ? l2_io_rresp_data_3_entries_vs_7 : r_7_3_entries_vs_7; // @[Reg.scala 16:16 17:{18,22}]
  reg [3:0] r_8; // @[Reg.scala 16:16]
  wire  asid_hit_8 = _GEN_63 == io_csr_dup_1_satp_asid; // @[MMUBundle.scala 654:59]
  wire  _GEN_148 = 3'h1 == data_req_info_vpn[11:9] ? _GEN_73 : _GEN_72; // @[MMUBundle.scala 655:{38,38}]
  wire  _GEN_149 = 3'h2 == data_req_info_vpn[11:9] ? _GEN_74 : _GEN_148; // @[MMUBundle.scala 655:{38,38}]
  wire  _GEN_150 = 3'h3 == data_req_info_vpn[11:9] ? _GEN_75 : _GEN_149; // @[MMUBundle.scala 655:{38,38}]
  wire  _GEN_151 = 3'h4 == data_req_info_vpn[11:9] ? _GEN_76 : _GEN_150; // @[MMUBundle.scala 655:{38,38}]
  wire  _GEN_152 = 3'h5 == data_req_info_vpn[11:9] ? _GEN_77 : _GEN_151; // @[MMUBundle.scala 655:{38,38}]
  wire  _GEN_153 = 3'h6 == data_req_info_vpn[11:9] ? _GEN_78 : _GEN_152; // @[MMUBundle.scala 655:{38,38}]
  wire  _GEN_154 = 3'h7 == data_req_info_vpn[11:9] ? _GEN_79 : _GEN_153; // @[MMUBundle.scala 655:{38,38}]
  wire  _T_83 = asid_hit_8 & _GEN_62 == data_req_info_vpn[26:14] & _GEN_154; // @[MMUBundle.scala 655:38]
  wire  _T_84 = _T_83 & r_8[0]; // @[PageTableCache.scala 270:63]
  wire  asid_hit_9 = _GEN_83 == io_csr_dup_1_satp_asid; // @[MMUBundle.scala 654:59]
  wire  _GEN_156 = 3'h1 == data_req_info_vpn[11:9] ? _GEN_93 : _GEN_92; // @[MMUBundle.scala 655:{38,38}]
  wire  _GEN_157 = 3'h2 == data_req_info_vpn[11:9] ? _GEN_94 : _GEN_156; // @[MMUBundle.scala 655:{38,38}]
  wire  _GEN_158 = 3'h3 == data_req_info_vpn[11:9] ? _GEN_95 : _GEN_157; // @[MMUBundle.scala 655:{38,38}]
  wire  _GEN_159 = 3'h4 == data_req_info_vpn[11:9] ? _GEN_96 : _GEN_158; // @[MMUBundle.scala 655:{38,38}]
  wire  _GEN_160 = 3'h5 == data_req_info_vpn[11:9] ? _GEN_97 : _GEN_159; // @[MMUBundle.scala 655:{38,38}]
  wire  _GEN_161 = 3'h6 == data_req_info_vpn[11:9] ? _GEN_98 : _GEN_160; // @[MMUBundle.scala 655:{38,38}]
  wire  _GEN_162 = 3'h7 == data_req_info_vpn[11:9] ? _GEN_99 : _GEN_161; // @[MMUBundle.scala 655:{38,38}]
  wire  _T_90 = asid_hit_9 & _GEN_82 == data_req_info_vpn[26:14] & _GEN_162; // @[MMUBundle.scala 655:38]
  wire  _T_91 = _T_90 & r_8[1]; // @[PageTableCache.scala 270:63]
  wire  asid_hit_10 = _GEN_103 == io_csr_dup_1_satp_asid; // @[MMUBundle.scala 654:59]
  wire  _GEN_164 = 3'h1 == data_req_info_vpn[11:9] ? _GEN_113 : _GEN_112; // @[MMUBundle.scala 655:{38,38}]
  wire  _GEN_165 = 3'h2 == data_req_info_vpn[11:9] ? _GEN_114 : _GEN_164; // @[MMUBundle.scala 655:{38,38}]
  wire  _GEN_166 = 3'h3 == data_req_info_vpn[11:9] ? _GEN_115 : _GEN_165; // @[MMUBundle.scala 655:{38,38}]
  wire  _GEN_167 = 3'h4 == data_req_info_vpn[11:9] ? _GEN_116 : _GEN_166; // @[MMUBundle.scala 655:{38,38}]
  wire  _GEN_168 = 3'h5 == data_req_info_vpn[11:9] ? _GEN_117 : _GEN_167; // @[MMUBundle.scala 655:{38,38}]
  wire  _GEN_169 = 3'h6 == data_req_info_vpn[11:9] ? _GEN_118 : _GEN_168; // @[MMUBundle.scala 655:{38,38}]
  wire  _GEN_170 = 3'h7 == data_req_info_vpn[11:9] ? _GEN_119 : _GEN_169; // @[MMUBundle.scala 655:{38,38}]
  wire  _T_97 = asid_hit_10 & _GEN_102 == data_req_info_vpn[26:14] & _GEN_170; // @[MMUBundle.scala 655:38]
  wire  _T_98 = _T_97 & r_8[2]; // @[PageTableCache.scala 270:63]
  wire  asid_hit_11 = _GEN_123 == io_csr_dup_1_satp_asid; // @[MMUBundle.scala 654:59]
  wire  _GEN_172 = 3'h1 == data_req_info_vpn[11:9] ? _GEN_133 : _GEN_132; // @[MMUBundle.scala 655:{38,38}]
  wire  _GEN_173 = 3'h2 == data_req_info_vpn[11:9] ? _GEN_134 : _GEN_172; // @[MMUBundle.scala 655:{38,38}]
  wire  _GEN_174 = 3'h3 == data_req_info_vpn[11:9] ? _GEN_135 : _GEN_173; // @[MMUBundle.scala 655:{38,38}]
  wire  _GEN_175 = 3'h4 == data_req_info_vpn[11:9] ? _GEN_136 : _GEN_174; // @[MMUBundle.scala 655:{38,38}]
  wire  _GEN_176 = 3'h5 == data_req_info_vpn[11:9] ? _GEN_137 : _GEN_175; // @[MMUBundle.scala 655:{38,38}]
  wire  _GEN_177 = 3'h6 == data_req_info_vpn[11:9] ? _GEN_138 : _GEN_176; // @[MMUBundle.scala 655:{38,38}]
  wire  _GEN_178 = 3'h7 == data_req_info_vpn[11:9] ? _GEN_139 : _GEN_177; // @[MMUBundle.scala 655:{38,38}]
  wire  _T_104 = asid_hit_11 & _GEN_122 == data_req_info_vpn[26:14] & _GEN_178; // @[MMUBundle.scala 655:38]
  wire  _T_105 = _T_104 & r_8[3]; // @[PageTableCache.scala 270:63]
  reg [12:0] l2_ramDatas_0_entries_tag; // @[Reg.scala 16:16]
  reg [15:0] l2_ramDatas_0_entries_asid; // @[Reg.scala 16:16]
  reg [23:0] l2_ramDatas_0_entries_ppns_0; // @[Reg.scala 16:16]
  reg [23:0] l2_ramDatas_0_entries_ppns_1; // @[Reg.scala 16:16]
  reg [23:0] l2_ramDatas_0_entries_ppns_2; // @[Reg.scala 16:16]
  reg [23:0] l2_ramDatas_0_entries_ppns_3; // @[Reg.scala 16:16]
  reg [23:0] l2_ramDatas_0_entries_ppns_4; // @[Reg.scala 16:16]
  reg [23:0] l2_ramDatas_0_entries_ppns_5; // @[Reg.scala 16:16]
  reg [23:0] l2_ramDatas_0_entries_ppns_6; // @[Reg.scala 16:16]
  reg [23:0] l2_ramDatas_0_entries_ppns_7; // @[Reg.scala 16:16]
  reg  l2_ramDatas_0_entries_vs_0; // @[Reg.scala 16:16]
  reg  l2_ramDatas_0_entries_vs_1; // @[Reg.scala 16:16]
  reg  l2_ramDatas_0_entries_vs_2; // @[Reg.scala 16:16]
  reg  l2_ramDatas_0_entries_vs_3; // @[Reg.scala 16:16]
  reg  l2_ramDatas_0_entries_vs_4; // @[Reg.scala 16:16]
  reg  l2_ramDatas_0_entries_vs_5; // @[Reg.scala 16:16]
  reg  l2_ramDatas_0_entries_vs_6; // @[Reg.scala 16:16]
  reg  l2_ramDatas_0_entries_vs_7; // @[Reg.scala 16:16]
  reg  l2_ramDatas_0_entries_prefetch; // @[Reg.scala 16:16]
  reg [30:0] l2_ramDatas_0_ecc; // @[Reg.scala 16:16]
  reg [12:0] l2_ramDatas_1_entries_tag; // @[Reg.scala 16:16]
  reg [15:0] l2_ramDatas_1_entries_asid; // @[Reg.scala 16:16]
  reg [23:0] l2_ramDatas_1_entries_ppns_0; // @[Reg.scala 16:16]
  reg [23:0] l2_ramDatas_1_entries_ppns_1; // @[Reg.scala 16:16]
  reg [23:0] l2_ramDatas_1_entries_ppns_2; // @[Reg.scala 16:16]
  reg [23:0] l2_ramDatas_1_entries_ppns_3; // @[Reg.scala 16:16]
  reg [23:0] l2_ramDatas_1_entries_ppns_4; // @[Reg.scala 16:16]
  reg [23:0] l2_ramDatas_1_entries_ppns_5; // @[Reg.scala 16:16]
  reg [23:0] l2_ramDatas_1_entries_ppns_6; // @[Reg.scala 16:16]
  reg [23:0] l2_ramDatas_1_entries_ppns_7; // @[Reg.scala 16:16]
  reg  l2_ramDatas_1_entries_vs_0; // @[Reg.scala 16:16]
  reg  l2_ramDatas_1_entries_vs_1; // @[Reg.scala 16:16]
  reg  l2_ramDatas_1_entries_vs_2; // @[Reg.scala 16:16]
  reg  l2_ramDatas_1_entries_vs_3; // @[Reg.scala 16:16]
  reg  l2_ramDatas_1_entries_vs_4; // @[Reg.scala 16:16]
  reg  l2_ramDatas_1_entries_vs_5; // @[Reg.scala 16:16]
  reg  l2_ramDatas_1_entries_vs_6; // @[Reg.scala 16:16]
  reg  l2_ramDatas_1_entries_vs_7; // @[Reg.scala 16:16]
  reg  l2_ramDatas_1_entries_prefetch; // @[Reg.scala 16:16]
  reg [30:0] l2_ramDatas_1_ecc; // @[Reg.scala 16:16]
  reg [12:0] l2_ramDatas_2_entries_tag; // @[Reg.scala 16:16]
  reg [15:0] l2_ramDatas_2_entries_asid; // @[Reg.scala 16:16]
  reg [23:0] l2_ramDatas_2_entries_ppns_0; // @[Reg.scala 16:16]
  reg [23:0] l2_ramDatas_2_entries_ppns_1; // @[Reg.scala 16:16]
  reg [23:0] l2_ramDatas_2_entries_ppns_2; // @[Reg.scala 16:16]
  reg [23:0] l2_ramDatas_2_entries_ppns_3; // @[Reg.scala 16:16]
  reg [23:0] l2_ramDatas_2_entries_ppns_4; // @[Reg.scala 16:16]
  reg [23:0] l2_ramDatas_2_entries_ppns_5; // @[Reg.scala 16:16]
  reg [23:0] l2_ramDatas_2_entries_ppns_6; // @[Reg.scala 16:16]
  reg [23:0] l2_ramDatas_2_entries_ppns_7; // @[Reg.scala 16:16]
  reg  l2_ramDatas_2_entries_vs_0; // @[Reg.scala 16:16]
  reg  l2_ramDatas_2_entries_vs_1; // @[Reg.scala 16:16]
  reg  l2_ramDatas_2_entries_vs_2; // @[Reg.scala 16:16]
  reg  l2_ramDatas_2_entries_vs_3; // @[Reg.scala 16:16]
  reg  l2_ramDatas_2_entries_vs_4; // @[Reg.scala 16:16]
  reg  l2_ramDatas_2_entries_vs_5; // @[Reg.scala 16:16]
  reg  l2_ramDatas_2_entries_vs_6; // @[Reg.scala 16:16]
  reg  l2_ramDatas_2_entries_vs_7; // @[Reg.scala 16:16]
  reg  l2_ramDatas_2_entries_prefetch; // @[Reg.scala 16:16]
  reg [30:0] l2_ramDatas_2_ecc; // @[Reg.scala 16:16]
  reg [12:0] l2_ramDatas_3_entries_tag; // @[Reg.scala 16:16]
  reg [15:0] l2_ramDatas_3_entries_asid; // @[Reg.scala 16:16]
  reg [23:0] l2_ramDatas_3_entries_ppns_0; // @[Reg.scala 16:16]
  reg [23:0] l2_ramDatas_3_entries_ppns_1; // @[Reg.scala 16:16]
  reg [23:0] l2_ramDatas_3_entries_ppns_2; // @[Reg.scala 16:16]
  reg [23:0] l2_ramDatas_3_entries_ppns_3; // @[Reg.scala 16:16]
  reg [23:0] l2_ramDatas_3_entries_ppns_4; // @[Reg.scala 16:16]
  reg [23:0] l2_ramDatas_3_entries_ppns_5; // @[Reg.scala 16:16]
  reg [23:0] l2_ramDatas_3_entries_ppns_6; // @[Reg.scala 16:16]
  reg [23:0] l2_ramDatas_3_entries_ppns_7; // @[Reg.scala 16:16]
  reg  l2_ramDatas_3_entries_vs_0; // @[Reg.scala 16:16]
  reg  l2_ramDatas_3_entries_vs_1; // @[Reg.scala 16:16]
  reg  l2_ramDatas_3_entries_vs_2; // @[Reg.scala 16:16]
  reg  l2_ramDatas_3_entries_vs_3; // @[Reg.scala 16:16]
  reg  l2_ramDatas_3_entries_vs_4; // @[Reg.scala 16:16]
  reg  l2_ramDatas_3_entries_vs_5; // @[Reg.scala 16:16]
  reg  l2_ramDatas_3_entries_vs_6; // @[Reg.scala 16:16]
  reg  l2_ramDatas_3_entries_vs_7; // @[Reg.scala 16:16]
  reg  l2_ramDatas_3_entries_prefetch; // @[Reg.scala 16:16]
  reg [30:0] l2_ramDatas_3_ecc; // @[Reg.scala 16:16]
  reg  l2_hitVec_0; // @[Reg.scala 16:16]
  reg  l2_hitVec_1; // @[Reg.scala 16:16]
  reg  l2_hitVec_2; // @[Reg.scala 16:16]
  reg  l2_hitVec_3; // @[Reg.scala 16:16]
  wire  _T_113 = l2_hitVec_0 | l2_hitVec_1; // @[ParallelMux.scala 90:65]
  wire [12:0] _T_114_entries_tag = l2_hitVec_0 ? l2_ramDatas_0_entries_tag : l2_ramDatas_1_entries_tag; // @[ParallelMux.scala 90:77]
  wire [15:0] _T_114_entries_asid = l2_hitVec_0 ? l2_ramDatas_0_entries_asid : l2_ramDatas_1_entries_asid; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_114_entries_ppns_0 = l2_hitVec_0 ? l2_ramDatas_0_entries_ppns_0 : l2_ramDatas_1_entries_ppns_0; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_114_entries_ppns_1 = l2_hitVec_0 ? l2_ramDatas_0_entries_ppns_1 : l2_ramDatas_1_entries_ppns_1; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_114_entries_ppns_2 = l2_hitVec_0 ? l2_ramDatas_0_entries_ppns_2 : l2_ramDatas_1_entries_ppns_2; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_114_entries_ppns_3 = l2_hitVec_0 ? l2_ramDatas_0_entries_ppns_3 : l2_ramDatas_1_entries_ppns_3; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_114_entries_ppns_4 = l2_hitVec_0 ? l2_ramDatas_0_entries_ppns_4 : l2_ramDatas_1_entries_ppns_4; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_114_entries_ppns_5 = l2_hitVec_0 ? l2_ramDatas_0_entries_ppns_5 : l2_ramDatas_1_entries_ppns_5; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_114_entries_ppns_6 = l2_hitVec_0 ? l2_ramDatas_0_entries_ppns_6 : l2_ramDatas_1_entries_ppns_6; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_114_entries_ppns_7 = l2_hitVec_0 ? l2_ramDatas_0_entries_ppns_7 : l2_ramDatas_1_entries_ppns_7; // @[ParallelMux.scala 90:77]
  wire  _T_114_entries_vs_0 = l2_hitVec_0 ? l2_ramDatas_0_entries_vs_0 : l2_ramDatas_1_entries_vs_0; // @[ParallelMux.scala 90:77]
  wire  _T_114_entries_vs_1 = l2_hitVec_0 ? l2_ramDatas_0_entries_vs_1 : l2_ramDatas_1_entries_vs_1; // @[ParallelMux.scala 90:77]
  wire  _T_114_entries_vs_2 = l2_hitVec_0 ? l2_ramDatas_0_entries_vs_2 : l2_ramDatas_1_entries_vs_2; // @[ParallelMux.scala 90:77]
  wire  _T_114_entries_vs_3 = l2_hitVec_0 ? l2_ramDatas_0_entries_vs_3 : l2_ramDatas_1_entries_vs_3; // @[ParallelMux.scala 90:77]
  wire  _T_114_entries_vs_4 = l2_hitVec_0 ? l2_ramDatas_0_entries_vs_4 : l2_ramDatas_1_entries_vs_4; // @[ParallelMux.scala 90:77]
  wire  _T_114_entries_vs_5 = l2_hitVec_0 ? l2_ramDatas_0_entries_vs_5 : l2_ramDatas_1_entries_vs_5; // @[ParallelMux.scala 90:77]
  wire  _T_114_entries_vs_6 = l2_hitVec_0 ? l2_ramDatas_0_entries_vs_6 : l2_ramDatas_1_entries_vs_6; // @[ParallelMux.scala 90:77]
  wire  _T_114_entries_vs_7 = l2_hitVec_0 ? l2_ramDatas_0_entries_vs_7 : l2_ramDatas_1_entries_vs_7; // @[ParallelMux.scala 90:77]
  wire  _T_114_entries_prefetch = l2_hitVec_0 ? l2_ramDatas_0_entries_prefetch : l2_ramDatas_1_entries_prefetch; // @[ParallelMux.scala 90:77]
  wire [30:0] _T_114_ecc = l2_hitVec_0 ? l2_ramDatas_0_ecc : l2_ramDatas_1_ecc; // @[ParallelMux.scala 90:77]
  wire  _T_115 = l2_hitVec_2 | l2_hitVec_3; // @[ParallelMux.scala 90:65]
  wire [12:0] _T_116_entries_tag = l2_hitVec_2 ? l2_ramDatas_2_entries_tag : l2_ramDatas_3_entries_tag; // @[ParallelMux.scala 90:77]
  wire [15:0] _T_116_entries_asid = l2_hitVec_2 ? l2_ramDatas_2_entries_asid : l2_ramDatas_3_entries_asid; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_116_entries_ppns_0 = l2_hitVec_2 ? l2_ramDatas_2_entries_ppns_0 : l2_ramDatas_3_entries_ppns_0; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_116_entries_ppns_1 = l2_hitVec_2 ? l2_ramDatas_2_entries_ppns_1 : l2_ramDatas_3_entries_ppns_1; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_116_entries_ppns_2 = l2_hitVec_2 ? l2_ramDatas_2_entries_ppns_2 : l2_ramDatas_3_entries_ppns_2; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_116_entries_ppns_3 = l2_hitVec_2 ? l2_ramDatas_2_entries_ppns_3 : l2_ramDatas_3_entries_ppns_3; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_116_entries_ppns_4 = l2_hitVec_2 ? l2_ramDatas_2_entries_ppns_4 : l2_ramDatas_3_entries_ppns_4; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_116_entries_ppns_5 = l2_hitVec_2 ? l2_ramDatas_2_entries_ppns_5 : l2_ramDatas_3_entries_ppns_5; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_116_entries_ppns_6 = l2_hitVec_2 ? l2_ramDatas_2_entries_ppns_6 : l2_ramDatas_3_entries_ppns_6; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_116_entries_ppns_7 = l2_hitVec_2 ? l2_ramDatas_2_entries_ppns_7 : l2_ramDatas_3_entries_ppns_7; // @[ParallelMux.scala 90:77]
  wire  _T_116_entries_vs_0 = l2_hitVec_2 ? l2_ramDatas_2_entries_vs_0 : l2_ramDatas_3_entries_vs_0; // @[ParallelMux.scala 90:77]
  wire  _T_116_entries_vs_1 = l2_hitVec_2 ? l2_ramDatas_2_entries_vs_1 : l2_ramDatas_3_entries_vs_1; // @[ParallelMux.scala 90:77]
  wire  _T_116_entries_vs_2 = l2_hitVec_2 ? l2_ramDatas_2_entries_vs_2 : l2_ramDatas_3_entries_vs_2; // @[ParallelMux.scala 90:77]
  wire  _T_116_entries_vs_3 = l2_hitVec_2 ? l2_ramDatas_2_entries_vs_3 : l2_ramDatas_3_entries_vs_3; // @[ParallelMux.scala 90:77]
  wire  _T_116_entries_vs_4 = l2_hitVec_2 ? l2_ramDatas_2_entries_vs_4 : l2_ramDatas_3_entries_vs_4; // @[ParallelMux.scala 90:77]
  wire  _T_116_entries_vs_5 = l2_hitVec_2 ? l2_ramDatas_2_entries_vs_5 : l2_ramDatas_3_entries_vs_5; // @[ParallelMux.scala 90:77]
  wire  _T_116_entries_vs_6 = l2_hitVec_2 ? l2_ramDatas_2_entries_vs_6 : l2_ramDatas_3_entries_vs_6; // @[ParallelMux.scala 90:77]
  wire  _T_116_entries_vs_7 = l2_hitVec_2 ? l2_ramDatas_2_entries_vs_7 : l2_ramDatas_3_entries_vs_7; // @[ParallelMux.scala 90:77]
  wire  _T_116_entries_prefetch = l2_hitVec_2 ? l2_ramDatas_2_entries_prefetch : l2_ramDatas_3_entries_prefetch; // @[ParallelMux.scala 90:77]
  wire [30:0] _T_116_ecc = l2_hitVec_2 ? l2_ramDatas_2_ecc : l2_ramDatas_3_ecc; // @[ParallelMux.scala 90:77]
  wire  _T_117 = l2_hitVec_0 | l2_hitVec_1 | (l2_hitVec_2 | l2_hitVec_3); // @[ParallelMux.scala 90:65]
  wire [12:0] _T_118_entries_tag = l2_hitVec_0 | l2_hitVec_1 ? _T_114_entries_tag : _T_116_entries_tag; // @[ParallelMux.scala 90:77]
  wire [15:0] _T_118_entries_asid = l2_hitVec_0 | l2_hitVec_1 ? _T_114_entries_asid : _T_116_entries_asid; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_118_entries_ppns_0 = l2_hitVec_0 | l2_hitVec_1 ? _T_114_entries_ppns_0 : _T_116_entries_ppns_0; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_118_entries_ppns_1 = l2_hitVec_0 | l2_hitVec_1 ? _T_114_entries_ppns_1 : _T_116_entries_ppns_1; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_118_entries_ppns_2 = l2_hitVec_0 | l2_hitVec_1 ? _T_114_entries_ppns_2 : _T_116_entries_ppns_2; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_118_entries_ppns_3 = l2_hitVec_0 | l2_hitVec_1 ? _T_114_entries_ppns_3 : _T_116_entries_ppns_3; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_118_entries_ppns_4 = l2_hitVec_0 | l2_hitVec_1 ? _T_114_entries_ppns_4 : _T_116_entries_ppns_4; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_118_entries_ppns_5 = l2_hitVec_0 | l2_hitVec_1 ? _T_114_entries_ppns_5 : _T_116_entries_ppns_5; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_118_entries_ppns_6 = l2_hitVec_0 | l2_hitVec_1 ? _T_114_entries_ppns_6 : _T_116_entries_ppns_6; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_118_entries_ppns_7 = l2_hitVec_0 | l2_hitVec_1 ? _T_114_entries_ppns_7 : _T_116_entries_ppns_7; // @[ParallelMux.scala 90:77]
  wire  _T_118_entries_vs_0 = l2_hitVec_0 | l2_hitVec_1 ? _T_114_entries_vs_0 : _T_116_entries_vs_0; // @[ParallelMux.scala 90:77]
  wire  _T_118_entries_vs_1 = l2_hitVec_0 | l2_hitVec_1 ? _T_114_entries_vs_1 : _T_116_entries_vs_1; // @[ParallelMux.scala 90:77]
  wire  _T_118_entries_vs_2 = l2_hitVec_0 | l2_hitVec_1 ? _T_114_entries_vs_2 : _T_116_entries_vs_2; // @[ParallelMux.scala 90:77]
  wire  _T_118_entries_vs_3 = l2_hitVec_0 | l2_hitVec_1 ? _T_114_entries_vs_3 : _T_116_entries_vs_3; // @[ParallelMux.scala 90:77]
  wire  _T_118_entries_vs_4 = l2_hitVec_0 | l2_hitVec_1 ? _T_114_entries_vs_4 : _T_116_entries_vs_4; // @[ParallelMux.scala 90:77]
  wire  _T_118_entries_vs_5 = l2_hitVec_0 | l2_hitVec_1 ? _T_114_entries_vs_5 : _T_116_entries_vs_5; // @[ParallelMux.scala 90:77]
  wire  _T_118_entries_vs_6 = l2_hitVec_0 | l2_hitVec_1 ? _T_114_entries_vs_6 : _T_116_entries_vs_6; // @[ParallelMux.scala 90:77]
  wire  _T_118_entries_vs_7 = l2_hitVec_0 | l2_hitVec_1 ? _T_114_entries_vs_7 : _T_116_entries_vs_7; // @[ParallelMux.scala 90:77]
  wire  check_res_l2_pre = l2_hitVec_0 | l2_hitVec_1 ? _T_114_entries_prefetch : _T_116_entries_prefetch; // @[ParallelMux.scala 90:77]
  wire [30:0] _T_118_ecc = l2_hitVec_0 | l2_hitVec_1 ? _T_114_ecc : _T_116_ecc; // @[ParallelMux.scala 90:77]
  wire [1:0] _T_123 = l2_hitVec_0 ? 2'h0 : 2'h1; // @[ParallelMux.scala 90:77]
  wire [1:0] _T_125 = l2_hitVec_2 ? 2'h2 : 2'h3; // @[ParallelMux.scala 90:77]
  wire [1:0] l2_hitWay = l2_hitVec_0 | l2_hitVec_1 ? _T_123 : _T_125; // @[ParallelMux.scala 90:77]
  wire [220:0] data_hi = {_T_118_entries_tag,_T_118_entries_asid,_T_118_entries_ppns_7,_T_118_entries_ppns_6,
    _T_118_entries_ppns_5,_T_118_entries_ppns_4,_T_118_entries_ppns_3,_T_118_entries_ppns_2,_T_118_entries_ppns_1,
    _T_118_entries_ppns_0}; // @[MMUBundle.scala 717:30]
  wire [229:0] data_3 = {data_hi,_T_118_entries_vs_7,_T_118_entries_vs_6,_T_118_entries_vs_5,_T_118_entries_vs_4,
    _T_118_entries_vs_3,_T_118_entries_vs_2,_T_118_entries_vs_1,_T_118_entries_vs_0,check_res_l2_pre}; // @[MMUBundle.scala 717:30]
  wire [71:0] _res_0_T_2 = {_T_118_ecc[7:0],data_3[63:0]}; // @[Cat.scala 31:58]
  wire [70:0] _res_0_syndromeUInt_T = 71'h1ab55555556aaad5b & _res_0_T_2[70:0]; // @[ECC.scala 156:66]
  wire [70:0] _res_0_syndromeUInt_T_2 = 71'h2cd9999999b33366d & _res_0_T_2[70:0]; // @[ECC.scala 156:66]
  wire [70:0] _res_0_syndromeUInt_T_4 = 71'h4f1e1e1e1e3c3c78e & _res_0_T_2[70:0]; // @[ECC.scala 156:66]
  wire [70:0] _res_0_syndromeUInt_T_6 = 71'h801fe01fe03fc07f0 & _res_0_T_2[70:0]; // @[ECC.scala 156:66]
  wire [70:0] _res_0_syndromeUInt_T_8 = 71'h1001fffe0003fff800 & _res_0_T_2[70:0]; // @[ECC.scala 156:66]
  wire [70:0] _res_0_syndromeUInt_T_10 = 71'h2001fffffffc000000 & _res_0_T_2[70:0]; // @[ECC.scala 156:66]
  wire [70:0] _res_0_syndromeUInt_T_12 = 71'h40fe00000000000000 & _res_0_T_2[70:0]; // @[ECC.scala 156:66]
  wire [6:0] res_0_syndromeUInt = {^_res_0_syndromeUInt_T_12,^_res_0_syndromeUInt_T_10,^_res_0_syndromeUInt_T_8,^
    _res_0_syndromeUInt_T_6,^_res_0_syndromeUInt_T_4,^_res_0_syndromeUInt_T_2,^_res_0_syndromeUInt_T}; // @[ECC.scala 156:78]
  wire  res_0_correctable = |res_0_syndromeUInt; // @[ECC.scala 163:36]
  wire  res_0_uncorrectable_1 = ^_res_0_T_2; // @[ECC.scala 87:27]
  wire  res_0_uncorrectable_2 = ~res_0_uncorrectable_1 & res_0_correctable; // @[ECC.scala 195:47]
  wire  res__0 = res_0_uncorrectable_1 | res_0_uncorrectable_2; // @[ECC.scala 31:27]
  wire [71:0] _res_1_T_2 = {_T_118_ecc[15:8],data_3[127:64]}; // @[Cat.scala 31:58]
  wire [70:0] _res_1_syndromeUInt_T = 71'h1ab55555556aaad5b & _res_1_T_2[70:0]; // @[ECC.scala 156:66]
  wire [70:0] _res_1_syndromeUInt_T_2 = 71'h2cd9999999b33366d & _res_1_T_2[70:0]; // @[ECC.scala 156:66]
  wire [70:0] _res_1_syndromeUInt_T_4 = 71'h4f1e1e1e1e3c3c78e & _res_1_T_2[70:0]; // @[ECC.scala 156:66]
  wire [70:0] _res_1_syndromeUInt_T_6 = 71'h801fe01fe03fc07f0 & _res_1_T_2[70:0]; // @[ECC.scala 156:66]
  wire [70:0] _res_1_syndromeUInt_T_8 = 71'h1001fffe0003fff800 & _res_1_T_2[70:0]; // @[ECC.scala 156:66]
  wire [70:0] _res_1_syndromeUInt_T_10 = 71'h2001fffffffc000000 & _res_1_T_2[70:0]; // @[ECC.scala 156:66]
  wire [70:0] _res_1_syndromeUInt_T_12 = 71'h40fe00000000000000 & _res_1_T_2[70:0]; // @[ECC.scala 156:66]
  wire [6:0] res_1_syndromeUInt = {^_res_1_syndromeUInt_T_12,^_res_1_syndromeUInt_T_10,^_res_1_syndromeUInt_T_8,^
    _res_1_syndromeUInt_T_6,^_res_1_syndromeUInt_T_4,^_res_1_syndromeUInt_T_2,^_res_1_syndromeUInt_T}; // @[ECC.scala 156:78]
  wire  res_1_correctable = |res_1_syndromeUInt; // @[ECC.scala 163:36]
  wire  res_1_uncorrectable_1 = ^_res_1_T_2; // @[ECC.scala 87:27]
  wire  res_1_uncorrectable_2 = ~res_1_uncorrectable_1 & res_1_correctable; // @[ECC.scala 195:47]
  wire  res__1 = res_1_uncorrectable_1 | res_1_uncorrectable_2; // @[ECC.scala 31:27]
  wire [71:0] _res_2_T_2 = {_T_118_ecc[23:16],data_3[191:128]}; // @[Cat.scala 31:58]
  wire [70:0] _res_2_syndromeUInt_T = 71'h1ab55555556aaad5b & _res_2_T_2[70:0]; // @[ECC.scala 156:66]
  wire [70:0] _res_2_syndromeUInt_T_2 = 71'h2cd9999999b33366d & _res_2_T_2[70:0]; // @[ECC.scala 156:66]
  wire [70:0] _res_2_syndromeUInt_T_4 = 71'h4f1e1e1e1e3c3c78e & _res_2_T_2[70:0]; // @[ECC.scala 156:66]
  wire [70:0] _res_2_syndromeUInt_T_6 = 71'h801fe01fe03fc07f0 & _res_2_T_2[70:0]; // @[ECC.scala 156:66]
  wire [70:0] _res_2_syndromeUInt_T_8 = 71'h1001fffe0003fff800 & _res_2_T_2[70:0]; // @[ECC.scala 156:66]
  wire [70:0] _res_2_syndromeUInt_T_10 = 71'h2001fffffffc000000 & _res_2_T_2[70:0]; // @[ECC.scala 156:66]
  wire [70:0] _res_2_syndromeUInt_T_12 = 71'h40fe00000000000000 & _res_2_T_2[70:0]; // @[ECC.scala 156:66]
  wire [6:0] res_2_syndromeUInt = {^_res_2_syndromeUInt_T_12,^_res_2_syndromeUInt_T_10,^_res_2_syndromeUInt_T_8,^
    _res_2_syndromeUInt_T_6,^_res_2_syndromeUInt_T_4,^_res_2_syndromeUInt_T_2,^_res_2_syndromeUInt_T}; // @[ECC.scala 156:78]
  wire  res_2_correctable = |res_2_syndromeUInt; // @[ECC.scala 163:36]
  wire  res_2_uncorrectable_1 = ^_res_2_T_2; // @[ECC.scala 87:27]
  wire  res_2_uncorrectable_2 = ~res_2_uncorrectable_1 & res_2_correctable; // @[ECC.scala 195:47]
  wire  res__2 = res_2_uncorrectable_1 | res_2_uncorrectable_2; // @[ECC.scala 31:27]
  wire [44:0] _res_3_T_2 = {_T_118_ecc[30:24],data_3[229:192]}; // @[Cat.scala 31:58]
  wire [43:0] _res_3_syndromeUInt_T = 44'h5556aaad5b & _res_3_T_2[43:0]; // @[ECC.scala 156:66]
  wire [43:0] _res_3_syndromeUInt_T_2 = 44'h999b33366d & _res_3_T_2[43:0]; // @[ECC.scala 156:66]
  wire [43:0] _res_3_syndromeUInt_T_4 = 44'h121e3c3c78e & _res_3_T_2[43:0]; // @[ECC.scala 156:66]
  wire [43:0] _res_3_syndromeUInt_T_6 = 44'h23e03fc07f0 & _res_3_T_2[43:0]; // @[ECC.scala 156:66]
  wire [43:0] _res_3_syndromeUInt_T_8 = 44'h40003fff800 & _res_3_T_2[43:0]; // @[ECC.scala 156:66]
  wire [43:0] _res_3_syndromeUInt_T_10 = 44'h83ffc000000 & _res_3_T_2[43:0]; // @[ECC.scala 156:66]
  wire [5:0] res_3_syndromeUInt = {^_res_3_syndromeUInt_T_10,^_res_3_syndromeUInt_T_8,^_res_3_syndromeUInt_T_6,^
    _res_3_syndromeUInt_T_4,^_res_3_syndromeUInt_T_2,^_res_3_syndromeUInt_T}; // @[ECC.scala 156:78]
  wire  res_3_correctable = |res_3_syndromeUInt; // @[ECC.scala 163:36]
  wire  res_3_uncorrectable_1 = ^_res_3_T_2; // @[ECC.scala 87:27]
  wire  res_3_uncorrectable_2 = ~res_3_uncorrectable_1 & res_3_correctable; // @[ECC.scala 195:47]
  wire  res__3 = res_3_uncorrectable_1 | res_3_uncorrectable_2; // @[ECC.scala 31:27]
  wire [3:0] _T_127 = {res__0,res__1,res__2,res__3}; // @[Cat.scala 31:58]
  wire  l2eccError = |_T_127; // @[MMUBundle.scala 727:14]
  wire  state_vec_set_left_older = ~l2_hitWay[1]; // @[Replacement.scala 196:33]
  wire [2:0] _GEN_265 = 2'h1 == data_1_req_info_vpn[13:12] ? state_vec__1 : state_vec__0; // @[package.scala 154:{13,13}]
  wire [2:0] _GEN_266 = 2'h2 == data_1_req_info_vpn[13:12] ? state_vec__2 : _GEN_265; // @[package.scala 154:{13,13}]
  wire [2:0] _GEN_267 = 2'h3 == data_1_req_info_vpn[13:12] ? state_vec__3 : _GEN_266; // @[package.scala 154:{13,13}]
  wire  state_vec_left_subtree_state = _GEN_267[1]; // @[package.scala 154:13]
  wire  state_vec_right_subtree_state = _GEN_267[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_T_2 = ~l2_hitWay[0]; // @[Replacement.scala 218:7]
  wire  _state_vec_T_3 = state_vec_set_left_older ? state_vec_left_subtree_state : _state_vec_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_T_7 = state_vec_set_left_older ? _state_vec_T_2 : state_vec_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_T_8 = {state_vec_set_left_older,_state_vec_T_3,_state_vec_T_7}; // @[Cat.scala 31:58]
  wire [2:0] _GEN_268 = 2'h0 == data_1_req_info_vpn[13:12] ? _state_vec_T_8 : state_vec__0; // @[Replacement.scala 305:17 308:{20,20}]
  wire [2:0] _GEN_269 = 2'h1 == data_1_req_info_vpn[13:12] ? _state_vec_T_8 : state_vec__1; // @[Replacement.scala 305:17 308:{20,20}]
  wire [2:0] _GEN_270 = 2'h2 == data_1_req_info_vpn[13:12] ? _state_vec_T_8 : state_vec__2; // @[Replacement.scala 305:17 308:{20,20}]
  wire [2:0] _GEN_271 = 2'h3 == data_1_req_info_vpn[13:12] ? _state_vec_T_8 : state_vec__3; // @[Replacement.scala 305:17 308:{20,20}]
  wire [2:0] _GEN_272 = _T_117 & stageCheck_valid_1cycle ? _GEN_268 : state_vec__0; // @[PageTableCache.scala 290:43 Replacement.scala 305:17]
  wire [2:0] _GEN_273 = _T_117 & stageCheck_valid_1cycle ? _GEN_269 : state_vec__1; // @[PageTableCache.scala 290:43 Replacement.scala 305:17]
  wire [2:0] _GEN_274 = _T_117 & stageCheck_valid_1cycle ? _GEN_270 : state_vec__2; // @[PageTableCache.scala 290:43 Replacement.scala 305:17]
  wire [2:0] _GEN_275 = _T_117 & stageCheck_valid_1cycle ? _GEN_271 : state_vec__3; // @[PageTableCache.scala 290:43 Replacement.scala 305:17]
  reg [6:0] state_vec_1_0; // @[Replacement.scala 305:17]
  reg [6:0] state_vec_1_1; // @[Replacement.scala 305:17]
  reg [6:0] state_vec_1_2; // @[Replacement.scala 305:17]
  reg [6:0] state_vec_1_3; // @[Replacement.scala 305:17]
  wire [1:0] l3_ridx = io_req_bits_req_info_vpn[4:3]; // @[MMUConst.scala 226:21]
  wire [7:0] l3vVec_0 = l3v[7:0]; // @[PageTableCache.scala 192:30]
  wire [7:0] l3vVec_1 = l3v[15:8]; // @[PageTableCache.scala 192:30]
  wire [7:0] l3vVec_2 = l3v[23:16]; // @[PageTableCache.scala 192:30]
  wire [7:0] l3vVec_3 = l3v[31:24]; // @[PageTableCache.scala 192:30]
  reg [21:0] r_10_0_entries_tag; // @[Reg.scala 16:16]
  reg [15:0] r_10_0_entries_asid; // @[Reg.scala 16:16]
  reg [23:0] r_10_0_entries_ppns_0; // @[Reg.scala 16:16]
  reg [23:0] r_10_0_entries_ppns_1; // @[Reg.scala 16:16]
  reg [23:0] r_10_0_entries_ppns_2; // @[Reg.scala 16:16]
  reg [23:0] r_10_0_entries_ppns_3; // @[Reg.scala 16:16]
  reg [23:0] r_10_0_entries_ppns_4; // @[Reg.scala 16:16]
  reg [23:0] r_10_0_entries_ppns_5; // @[Reg.scala 16:16]
  reg [23:0] r_10_0_entries_ppns_6; // @[Reg.scala 16:16]
  reg [23:0] r_10_0_entries_ppns_7; // @[Reg.scala 16:16]
  reg  r_10_0_entries_vs_0; // @[Reg.scala 16:16]
  reg  r_10_0_entries_vs_1; // @[Reg.scala 16:16]
  reg  r_10_0_entries_vs_2; // @[Reg.scala 16:16]
  reg  r_10_0_entries_vs_3; // @[Reg.scala 16:16]
  reg  r_10_0_entries_vs_4; // @[Reg.scala 16:16]
  reg  r_10_0_entries_vs_5; // @[Reg.scala 16:16]
  reg  r_10_0_entries_vs_6; // @[Reg.scala 16:16]
  reg  r_10_0_entries_vs_7; // @[Reg.scala 16:16]
  reg  r_10_0_entries_perms_0_d; // @[Reg.scala 16:16]
  reg  r_10_0_entries_perms_0_a; // @[Reg.scala 16:16]
  reg  r_10_0_entries_perms_0_g; // @[Reg.scala 16:16]
  reg  r_10_0_entries_perms_0_u; // @[Reg.scala 16:16]
  reg  r_10_0_entries_perms_0_x; // @[Reg.scala 16:16]
  reg  r_10_0_entries_perms_0_w; // @[Reg.scala 16:16]
  reg  r_10_0_entries_perms_0_r; // @[Reg.scala 16:16]
  reg  r_10_0_entries_perms_1_d; // @[Reg.scala 16:16]
  reg  r_10_0_entries_perms_1_a; // @[Reg.scala 16:16]
  reg  r_10_0_entries_perms_1_g; // @[Reg.scala 16:16]
  reg  r_10_0_entries_perms_1_u; // @[Reg.scala 16:16]
  reg  r_10_0_entries_perms_1_x; // @[Reg.scala 16:16]
  reg  r_10_0_entries_perms_1_w; // @[Reg.scala 16:16]
  reg  r_10_0_entries_perms_1_r; // @[Reg.scala 16:16]
  reg  r_10_0_entries_perms_2_d; // @[Reg.scala 16:16]
  reg  r_10_0_entries_perms_2_a; // @[Reg.scala 16:16]
  reg  r_10_0_entries_perms_2_g; // @[Reg.scala 16:16]
  reg  r_10_0_entries_perms_2_u; // @[Reg.scala 16:16]
  reg  r_10_0_entries_perms_2_x; // @[Reg.scala 16:16]
  reg  r_10_0_entries_perms_2_w; // @[Reg.scala 16:16]
  reg  r_10_0_entries_perms_2_r; // @[Reg.scala 16:16]
  reg  r_10_0_entries_perms_3_d; // @[Reg.scala 16:16]
  reg  r_10_0_entries_perms_3_a; // @[Reg.scala 16:16]
  reg  r_10_0_entries_perms_3_g; // @[Reg.scala 16:16]
  reg  r_10_0_entries_perms_3_u; // @[Reg.scala 16:16]
  reg  r_10_0_entries_perms_3_x; // @[Reg.scala 16:16]
  reg  r_10_0_entries_perms_3_w; // @[Reg.scala 16:16]
  reg  r_10_0_entries_perms_3_r; // @[Reg.scala 16:16]
  reg  r_10_0_entries_perms_4_d; // @[Reg.scala 16:16]
  reg  r_10_0_entries_perms_4_a; // @[Reg.scala 16:16]
  reg  r_10_0_entries_perms_4_g; // @[Reg.scala 16:16]
  reg  r_10_0_entries_perms_4_u; // @[Reg.scala 16:16]
  reg  r_10_0_entries_perms_4_x; // @[Reg.scala 16:16]
  reg  r_10_0_entries_perms_4_w; // @[Reg.scala 16:16]
  reg  r_10_0_entries_perms_4_r; // @[Reg.scala 16:16]
  reg  r_10_0_entries_perms_5_d; // @[Reg.scala 16:16]
  reg  r_10_0_entries_perms_5_a; // @[Reg.scala 16:16]
  reg  r_10_0_entries_perms_5_g; // @[Reg.scala 16:16]
  reg  r_10_0_entries_perms_5_u; // @[Reg.scala 16:16]
  reg  r_10_0_entries_perms_5_x; // @[Reg.scala 16:16]
  reg  r_10_0_entries_perms_5_w; // @[Reg.scala 16:16]
  reg  r_10_0_entries_perms_5_r; // @[Reg.scala 16:16]
  reg  r_10_0_entries_perms_6_d; // @[Reg.scala 16:16]
  reg  r_10_0_entries_perms_6_a; // @[Reg.scala 16:16]
  reg  r_10_0_entries_perms_6_g; // @[Reg.scala 16:16]
  reg  r_10_0_entries_perms_6_u; // @[Reg.scala 16:16]
  reg  r_10_0_entries_perms_6_x; // @[Reg.scala 16:16]
  reg  r_10_0_entries_perms_6_w; // @[Reg.scala 16:16]
  reg  r_10_0_entries_perms_6_r; // @[Reg.scala 16:16]
  reg  r_10_0_entries_perms_7_d; // @[Reg.scala 16:16]
  reg  r_10_0_entries_perms_7_a; // @[Reg.scala 16:16]
  reg  r_10_0_entries_perms_7_g; // @[Reg.scala 16:16]
  reg  r_10_0_entries_perms_7_u; // @[Reg.scala 16:16]
  reg  r_10_0_entries_perms_7_x; // @[Reg.scala 16:16]
  reg  r_10_0_entries_perms_7_w; // @[Reg.scala 16:16]
  reg  r_10_0_entries_perms_7_r; // @[Reg.scala 16:16]
  reg  r_10_0_entries_prefetch; // @[Reg.scala 16:16]
  reg [38:0] r_10_0_ecc; // @[Reg.scala 16:16]
  reg [21:0] r_10_1_entries_tag; // @[Reg.scala 16:16]
  reg [15:0] r_10_1_entries_asid; // @[Reg.scala 16:16]
  reg [23:0] r_10_1_entries_ppns_0; // @[Reg.scala 16:16]
  reg [23:0] r_10_1_entries_ppns_1; // @[Reg.scala 16:16]
  reg [23:0] r_10_1_entries_ppns_2; // @[Reg.scala 16:16]
  reg [23:0] r_10_1_entries_ppns_3; // @[Reg.scala 16:16]
  reg [23:0] r_10_1_entries_ppns_4; // @[Reg.scala 16:16]
  reg [23:0] r_10_1_entries_ppns_5; // @[Reg.scala 16:16]
  reg [23:0] r_10_1_entries_ppns_6; // @[Reg.scala 16:16]
  reg [23:0] r_10_1_entries_ppns_7; // @[Reg.scala 16:16]
  reg  r_10_1_entries_vs_0; // @[Reg.scala 16:16]
  reg  r_10_1_entries_vs_1; // @[Reg.scala 16:16]
  reg  r_10_1_entries_vs_2; // @[Reg.scala 16:16]
  reg  r_10_1_entries_vs_3; // @[Reg.scala 16:16]
  reg  r_10_1_entries_vs_4; // @[Reg.scala 16:16]
  reg  r_10_1_entries_vs_5; // @[Reg.scala 16:16]
  reg  r_10_1_entries_vs_6; // @[Reg.scala 16:16]
  reg  r_10_1_entries_vs_7; // @[Reg.scala 16:16]
  reg  r_10_1_entries_perms_0_d; // @[Reg.scala 16:16]
  reg  r_10_1_entries_perms_0_a; // @[Reg.scala 16:16]
  reg  r_10_1_entries_perms_0_g; // @[Reg.scala 16:16]
  reg  r_10_1_entries_perms_0_u; // @[Reg.scala 16:16]
  reg  r_10_1_entries_perms_0_x; // @[Reg.scala 16:16]
  reg  r_10_1_entries_perms_0_w; // @[Reg.scala 16:16]
  reg  r_10_1_entries_perms_0_r; // @[Reg.scala 16:16]
  reg  r_10_1_entries_perms_1_d; // @[Reg.scala 16:16]
  reg  r_10_1_entries_perms_1_a; // @[Reg.scala 16:16]
  reg  r_10_1_entries_perms_1_g; // @[Reg.scala 16:16]
  reg  r_10_1_entries_perms_1_u; // @[Reg.scala 16:16]
  reg  r_10_1_entries_perms_1_x; // @[Reg.scala 16:16]
  reg  r_10_1_entries_perms_1_w; // @[Reg.scala 16:16]
  reg  r_10_1_entries_perms_1_r; // @[Reg.scala 16:16]
  reg  r_10_1_entries_perms_2_d; // @[Reg.scala 16:16]
  reg  r_10_1_entries_perms_2_a; // @[Reg.scala 16:16]
  reg  r_10_1_entries_perms_2_g; // @[Reg.scala 16:16]
  reg  r_10_1_entries_perms_2_u; // @[Reg.scala 16:16]
  reg  r_10_1_entries_perms_2_x; // @[Reg.scala 16:16]
  reg  r_10_1_entries_perms_2_w; // @[Reg.scala 16:16]
  reg  r_10_1_entries_perms_2_r; // @[Reg.scala 16:16]
  reg  r_10_1_entries_perms_3_d; // @[Reg.scala 16:16]
  reg  r_10_1_entries_perms_3_a; // @[Reg.scala 16:16]
  reg  r_10_1_entries_perms_3_g; // @[Reg.scala 16:16]
  reg  r_10_1_entries_perms_3_u; // @[Reg.scala 16:16]
  reg  r_10_1_entries_perms_3_x; // @[Reg.scala 16:16]
  reg  r_10_1_entries_perms_3_w; // @[Reg.scala 16:16]
  reg  r_10_1_entries_perms_3_r; // @[Reg.scala 16:16]
  reg  r_10_1_entries_perms_4_d; // @[Reg.scala 16:16]
  reg  r_10_1_entries_perms_4_a; // @[Reg.scala 16:16]
  reg  r_10_1_entries_perms_4_g; // @[Reg.scala 16:16]
  reg  r_10_1_entries_perms_4_u; // @[Reg.scala 16:16]
  reg  r_10_1_entries_perms_4_x; // @[Reg.scala 16:16]
  reg  r_10_1_entries_perms_4_w; // @[Reg.scala 16:16]
  reg  r_10_1_entries_perms_4_r; // @[Reg.scala 16:16]
  reg  r_10_1_entries_perms_5_d; // @[Reg.scala 16:16]
  reg  r_10_1_entries_perms_5_a; // @[Reg.scala 16:16]
  reg  r_10_1_entries_perms_5_g; // @[Reg.scala 16:16]
  reg  r_10_1_entries_perms_5_u; // @[Reg.scala 16:16]
  reg  r_10_1_entries_perms_5_x; // @[Reg.scala 16:16]
  reg  r_10_1_entries_perms_5_w; // @[Reg.scala 16:16]
  reg  r_10_1_entries_perms_5_r; // @[Reg.scala 16:16]
  reg  r_10_1_entries_perms_6_d; // @[Reg.scala 16:16]
  reg  r_10_1_entries_perms_6_a; // @[Reg.scala 16:16]
  reg  r_10_1_entries_perms_6_g; // @[Reg.scala 16:16]
  reg  r_10_1_entries_perms_6_u; // @[Reg.scala 16:16]
  reg  r_10_1_entries_perms_6_x; // @[Reg.scala 16:16]
  reg  r_10_1_entries_perms_6_w; // @[Reg.scala 16:16]
  reg  r_10_1_entries_perms_6_r; // @[Reg.scala 16:16]
  reg  r_10_1_entries_perms_7_d; // @[Reg.scala 16:16]
  reg  r_10_1_entries_perms_7_a; // @[Reg.scala 16:16]
  reg  r_10_1_entries_perms_7_g; // @[Reg.scala 16:16]
  reg  r_10_1_entries_perms_7_u; // @[Reg.scala 16:16]
  reg  r_10_1_entries_perms_7_x; // @[Reg.scala 16:16]
  reg  r_10_1_entries_perms_7_w; // @[Reg.scala 16:16]
  reg  r_10_1_entries_perms_7_r; // @[Reg.scala 16:16]
  reg  r_10_1_entries_prefetch; // @[Reg.scala 16:16]
  reg [38:0] r_10_1_ecc; // @[Reg.scala 16:16]
  reg [21:0] r_10_2_entries_tag; // @[Reg.scala 16:16]
  reg [15:0] r_10_2_entries_asid; // @[Reg.scala 16:16]
  reg [23:0] r_10_2_entries_ppns_0; // @[Reg.scala 16:16]
  reg [23:0] r_10_2_entries_ppns_1; // @[Reg.scala 16:16]
  reg [23:0] r_10_2_entries_ppns_2; // @[Reg.scala 16:16]
  reg [23:0] r_10_2_entries_ppns_3; // @[Reg.scala 16:16]
  reg [23:0] r_10_2_entries_ppns_4; // @[Reg.scala 16:16]
  reg [23:0] r_10_2_entries_ppns_5; // @[Reg.scala 16:16]
  reg [23:0] r_10_2_entries_ppns_6; // @[Reg.scala 16:16]
  reg [23:0] r_10_2_entries_ppns_7; // @[Reg.scala 16:16]
  reg  r_10_2_entries_vs_0; // @[Reg.scala 16:16]
  reg  r_10_2_entries_vs_1; // @[Reg.scala 16:16]
  reg  r_10_2_entries_vs_2; // @[Reg.scala 16:16]
  reg  r_10_2_entries_vs_3; // @[Reg.scala 16:16]
  reg  r_10_2_entries_vs_4; // @[Reg.scala 16:16]
  reg  r_10_2_entries_vs_5; // @[Reg.scala 16:16]
  reg  r_10_2_entries_vs_6; // @[Reg.scala 16:16]
  reg  r_10_2_entries_vs_7; // @[Reg.scala 16:16]
  reg  r_10_2_entries_perms_0_d; // @[Reg.scala 16:16]
  reg  r_10_2_entries_perms_0_a; // @[Reg.scala 16:16]
  reg  r_10_2_entries_perms_0_g; // @[Reg.scala 16:16]
  reg  r_10_2_entries_perms_0_u; // @[Reg.scala 16:16]
  reg  r_10_2_entries_perms_0_x; // @[Reg.scala 16:16]
  reg  r_10_2_entries_perms_0_w; // @[Reg.scala 16:16]
  reg  r_10_2_entries_perms_0_r; // @[Reg.scala 16:16]
  reg  r_10_2_entries_perms_1_d; // @[Reg.scala 16:16]
  reg  r_10_2_entries_perms_1_a; // @[Reg.scala 16:16]
  reg  r_10_2_entries_perms_1_g; // @[Reg.scala 16:16]
  reg  r_10_2_entries_perms_1_u; // @[Reg.scala 16:16]
  reg  r_10_2_entries_perms_1_x; // @[Reg.scala 16:16]
  reg  r_10_2_entries_perms_1_w; // @[Reg.scala 16:16]
  reg  r_10_2_entries_perms_1_r; // @[Reg.scala 16:16]
  reg  r_10_2_entries_perms_2_d; // @[Reg.scala 16:16]
  reg  r_10_2_entries_perms_2_a; // @[Reg.scala 16:16]
  reg  r_10_2_entries_perms_2_g; // @[Reg.scala 16:16]
  reg  r_10_2_entries_perms_2_u; // @[Reg.scala 16:16]
  reg  r_10_2_entries_perms_2_x; // @[Reg.scala 16:16]
  reg  r_10_2_entries_perms_2_w; // @[Reg.scala 16:16]
  reg  r_10_2_entries_perms_2_r; // @[Reg.scala 16:16]
  reg  r_10_2_entries_perms_3_d; // @[Reg.scala 16:16]
  reg  r_10_2_entries_perms_3_a; // @[Reg.scala 16:16]
  reg  r_10_2_entries_perms_3_g; // @[Reg.scala 16:16]
  reg  r_10_2_entries_perms_3_u; // @[Reg.scala 16:16]
  reg  r_10_2_entries_perms_3_x; // @[Reg.scala 16:16]
  reg  r_10_2_entries_perms_3_w; // @[Reg.scala 16:16]
  reg  r_10_2_entries_perms_3_r; // @[Reg.scala 16:16]
  reg  r_10_2_entries_perms_4_d; // @[Reg.scala 16:16]
  reg  r_10_2_entries_perms_4_a; // @[Reg.scala 16:16]
  reg  r_10_2_entries_perms_4_g; // @[Reg.scala 16:16]
  reg  r_10_2_entries_perms_4_u; // @[Reg.scala 16:16]
  reg  r_10_2_entries_perms_4_x; // @[Reg.scala 16:16]
  reg  r_10_2_entries_perms_4_w; // @[Reg.scala 16:16]
  reg  r_10_2_entries_perms_4_r; // @[Reg.scala 16:16]
  reg  r_10_2_entries_perms_5_d; // @[Reg.scala 16:16]
  reg  r_10_2_entries_perms_5_a; // @[Reg.scala 16:16]
  reg  r_10_2_entries_perms_5_g; // @[Reg.scala 16:16]
  reg  r_10_2_entries_perms_5_u; // @[Reg.scala 16:16]
  reg  r_10_2_entries_perms_5_x; // @[Reg.scala 16:16]
  reg  r_10_2_entries_perms_5_w; // @[Reg.scala 16:16]
  reg  r_10_2_entries_perms_5_r; // @[Reg.scala 16:16]
  reg  r_10_2_entries_perms_6_d; // @[Reg.scala 16:16]
  reg  r_10_2_entries_perms_6_a; // @[Reg.scala 16:16]
  reg  r_10_2_entries_perms_6_g; // @[Reg.scala 16:16]
  reg  r_10_2_entries_perms_6_u; // @[Reg.scala 16:16]
  reg  r_10_2_entries_perms_6_x; // @[Reg.scala 16:16]
  reg  r_10_2_entries_perms_6_w; // @[Reg.scala 16:16]
  reg  r_10_2_entries_perms_6_r; // @[Reg.scala 16:16]
  reg  r_10_2_entries_perms_7_d; // @[Reg.scala 16:16]
  reg  r_10_2_entries_perms_7_a; // @[Reg.scala 16:16]
  reg  r_10_2_entries_perms_7_g; // @[Reg.scala 16:16]
  reg  r_10_2_entries_perms_7_u; // @[Reg.scala 16:16]
  reg  r_10_2_entries_perms_7_x; // @[Reg.scala 16:16]
  reg  r_10_2_entries_perms_7_w; // @[Reg.scala 16:16]
  reg  r_10_2_entries_perms_7_r; // @[Reg.scala 16:16]
  reg  r_10_2_entries_prefetch; // @[Reg.scala 16:16]
  reg [38:0] r_10_2_ecc; // @[Reg.scala 16:16]
  reg [21:0] r_10_3_entries_tag; // @[Reg.scala 16:16]
  reg [15:0] r_10_3_entries_asid; // @[Reg.scala 16:16]
  reg [23:0] r_10_3_entries_ppns_0; // @[Reg.scala 16:16]
  reg [23:0] r_10_3_entries_ppns_1; // @[Reg.scala 16:16]
  reg [23:0] r_10_3_entries_ppns_2; // @[Reg.scala 16:16]
  reg [23:0] r_10_3_entries_ppns_3; // @[Reg.scala 16:16]
  reg [23:0] r_10_3_entries_ppns_4; // @[Reg.scala 16:16]
  reg [23:0] r_10_3_entries_ppns_5; // @[Reg.scala 16:16]
  reg [23:0] r_10_3_entries_ppns_6; // @[Reg.scala 16:16]
  reg [23:0] r_10_3_entries_ppns_7; // @[Reg.scala 16:16]
  reg  r_10_3_entries_vs_0; // @[Reg.scala 16:16]
  reg  r_10_3_entries_vs_1; // @[Reg.scala 16:16]
  reg  r_10_3_entries_vs_2; // @[Reg.scala 16:16]
  reg  r_10_3_entries_vs_3; // @[Reg.scala 16:16]
  reg  r_10_3_entries_vs_4; // @[Reg.scala 16:16]
  reg  r_10_3_entries_vs_5; // @[Reg.scala 16:16]
  reg  r_10_3_entries_vs_6; // @[Reg.scala 16:16]
  reg  r_10_3_entries_vs_7; // @[Reg.scala 16:16]
  reg  r_10_3_entries_perms_0_d; // @[Reg.scala 16:16]
  reg  r_10_3_entries_perms_0_a; // @[Reg.scala 16:16]
  reg  r_10_3_entries_perms_0_g; // @[Reg.scala 16:16]
  reg  r_10_3_entries_perms_0_u; // @[Reg.scala 16:16]
  reg  r_10_3_entries_perms_0_x; // @[Reg.scala 16:16]
  reg  r_10_3_entries_perms_0_w; // @[Reg.scala 16:16]
  reg  r_10_3_entries_perms_0_r; // @[Reg.scala 16:16]
  reg  r_10_3_entries_perms_1_d; // @[Reg.scala 16:16]
  reg  r_10_3_entries_perms_1_a; // @[Reg.scala 16:16]
  reg  r_10_3_entries_perms_1_g; // @[Reg.scala 16:16]
  reg  r_10_3_entries_perms_1_u; // @[Reg.scala 16:16]
  reg  r_10_3_entries_perms_1_x; // @[Reg.scala 16:16]
  reg  r_10_3_entries_perms_1_w; // @[Reg.scala 16:16]
  reg  r_10_3_entries_perms_1_r; // @[Reg.scala 16:16]
  reg  r_10_3_entries_perms_2_d; // @[Reg.scala 16:16]
  reg  r_10_3_entries_perms_2_a; // @[Reg.scala 16:16]
  reg  r_10_3_entries_perms_2_g; // @[Reg.scala 16:16]
  reg  r_10_3_entries_perms_2_u; // @[Reg.scala 16:16]
  reg  r_10_3_entries_perms_2_x; // @[Reg.scala 16:16]
  reg  r_10_3_entries_perms_2_w; // @[Reg.scala 16:16]
  reg  r_10_3_entries_perms_2_r; // @[Reg.scala 16:16]
  reg  r_10_3_entries_perms_3_d; // @[Reg.scala 16:16]
  reg  r_10_3_entries_perms_3_a; // @[Reg.scala 16:16]
  reg  r_10_3_entries_perms_3_g; // @[Reg.scala 16:16]
  reg  r_10_3_entries_perms_3_u; // @[Reg.scala 16:16]
  reg  r_10_3_entries_perms_3_x; // @[Reg.scala 16:16]
  reg  r_10_3_entries_perms_3_w; // @[Reg.scala 16:16]
  reg  r_10_3_entries_perms_3_r; // @[Reg.scala 16:16]
  reg  r_10_3_entries_perms_4_d; // @[Reg.scala 16:16]
  reg  r_10_3_entries_perms_4_a; // @[Reg.scala 16:16]
  reg  r_10_3_entries_perms_4_g; // @[Reg.scala 16:16]
  reg  r_10_3_entries_perms_4_u; // @[Reg.scala 16:16]
  reg  r_10_3_entries_perms_4_x; // @[Reg.scala 16:16]
  reg  r_10_3_entries_perms_4_w; // @[Reg.scala 16:16]
  reg  r_10_3_entries_perms_4_r; // @[Reg.scala 16:16]
  reg  r_10_3_entries_perms_5_d; // @[Reg.scala 16:16]
  reg  r_10_3_entries_perms_5_a; // @[Reg.scala 16:16]
  reg  r_10_3_entries_perms_5_g; // @[Reg.scala 16:16]
  reg  r_10_3_entries_perms_5_u; // @[Reg.scala 16:16]
  reg  r_10_3_entries_perms_5_x; // @[Reg.scala 16:16]
  reg  r_10_3_entries_perms_5_w; // @[Reg.scala 16:16]
  reg  r_10_3_entries_perms_5_r; // @[Reg.scala 16:16]
  reg  r_10_3_entries_perms_6_d; // @[Reg.scala 16:16]
  reg  r_10_3_entries_perms_6_a; // @[Reg.scala 16:16]
  reg  r_10_3_entries_perms_6_g; // @[Reg.scala 16:16]
  reg  r_10_3_entries_perms_6_u; // @[Reg.scala 16:16]
  reg  r_10_3_entries_perms_6_x; // @[Reg.scala 16:16]
  reg  r_10_3_entries_perms_6_w; // @[Reg.scala 16:16]
  reg  r_10_3_entries_perms_6_r; // @[Reg.scala 16:16]
  reg  r_10_3_entries_perms_7_d; // @[Reg.scala 16:16]
  reg  r_10_3_entries_perms_7_a; // @[Reg.scala 16:16]
  reg  r_10_3_entries_perms_7_g; // @[Reg.scala 16:16]
  reg  r_10_3_entries_perms_7_u; // @[Reg.scala 16:16]
  reg  r_10_3_entries_perms_7_x; // @[Reg.scala 16:16]
  reg  r_10_3_entries_perms_7_w; // @[Reg.scala 16:16]
  reg  r_10_3_entries_perms_7_r; // @[Reg.scala 16:16]
  reg  r_10_3_entries_prefetch; // @[Reg.scala 16:16]
  reg [38:0] r_10_3_ecc; // @[Reg.scala 16:16]
  reg [21:0] r_10_4_entries_tag; // @[Reg.scala 16:16]
  reg [15:0] r_10_4_entries_asid; // @[Reg.scala 16:16]
  reg [23:0] r_10_4_entries_ppns_0; // @[Reg.scala 16:16]
  reg [23:0] r_10_4_entries_ppns_1; // @[Reg.scala 16:16]
  reg [23:0] r_10_4_entries_ppns_2; // @[Reg.scala 16:16]
  reg [23:0] r_10_4_entries_ppns_3; // @[Reg.scala 16:16]
  reg [23:0] r_10_4_entries_ppns_4; // @[Reg.scala 16:16]
  reg [23:0] r_10_4_entries_ppns_5; // @[Reg.scala 16:16]
  reg [23:0] r_10_4_entries_ppns_6; // @[Reg.scala 16:16]
  reg [23:0] r_10_4_entries_ppns_7; // @[Reg.scala 16:16]
  reg  r_10_4_entries_vs_0; // @[Reg.scala 16:16]
  reg  r_10_4_entries_vs_1; // @[Reg.scala 16:16]
  reg  r_10_4_entries_vs_2; // @[Reg.scala 16:16]
  reg  r_10_4_entries_vs_3; // @[Reg.scala 16:16]
  reg  r_10_4_entries_vs_4; // @[Reg.scala 16:16]
  reg  r_10_4_entries_vs_5; // @[Reg.scala 16:16]
  reg  r_10_4_entries_vs_6; // @[Reg.scala 16:16]
  reg  r_10_4_entries_vs_7; // @[Reg.scala 16:16]
  reg  r_10_4_entries_perms_0_d; // @[Reg.scala 16:16]
  reg  r_10_4_entries_perms_0_a; // @[Reg.scala 16:16]
  reg  r_10_4_entries_perms_0_g; // @[Reg.scala 16:16]
  reg  r_10_4_entries_perms_0_u; // @[Reg.scala 16:16]
  reg  r_10_4_entries_perms_0_x; // @[Reg.scala 16:16]
  reg  r_10_4_entries_perms_0_w; // @[Reg.scala 16:16]
  reg  r_10_4_entries_perms_0_r; // @[Reg.scala 16:16]
  reg  r_10_4_entries_perms_1_d; // @[Reg.scala 16:16]
  reg  r_10_4_entries_perms_1_a; // @[Reg.scala 16:16]
  reg  r_10_4_entries_perms_1_g; // @[Reg.scala 16:16]
  reg  r_10_4_entries_perms_1_u; // @[Reg.scala 16:16]
  reg  r_10_4_entries_perms_1_x; // @[Reg.scala 16:16]
  reg  r_10_4_entries_perms_1_w; // @[Reg.scala 16:16]
  reg  r_10_4_entries_perms_1_r; // @[Reg.scala 16:16]
  reg  r_10_4_entries_perms_2_d; // @[Reg.scala 16:16]
  reg  r_10_4_entries_perms_2_a; // @[Reg.scala 16:16]
  reg  r_10_4_entries_perms_2_g; // @[Reg.scala 16:16]
  reg  r_10_4_entries_perms_2_u; // @[Reg.scala 16:16]
  reg  r_10_4_entries_perms_2_x; // @[Reg.scala 16:16]
  reg  r_10_4_entries_perms_2_w; // @[Reg.scala 16:16]
  reg  r_10_4_entries_perms_2_r; // @[Reg.scala 16:16]
  reg  r_10_4_entries_perms_3_d; // @[Reg.scala 16:16]
  reg  r_10_4_entries_perms_3_a; // @[Reg.scala 16:16]
  reg  r_10_4_entries_perms_3_g; // @[Reg.scala 16:16]
  reg  r_10_4_entries_perms_3_u; // @[Reg.scala 16:16]
  reg  r_10_4_entries_perms_3_x; // @[Reg.scala 16:16]
  reg  r_10_4_entries_perms_3_w; // @[Reg.scala 16:16]
  reg  r_10_4_entries_perms_3_r; // @[Reg.scala 16:16]
  reg  r_10_4_entries_perms_4_d; // @[Reg.scala 16:16]
  reg  r_10_4_entries_perms_4_a; // @[Reg.scala 16:16]
  reg  r_10_4_entries_perms_4_g; // @[Reg.scala 16:16]
  reg  r_10_4_entries_perms_4_u; // @[Reg.scala 16:16]
  reg  r_10_4_entries_perms_4_x; // @[Reg.scala 16:16]
  reg  r_10_4_entries_perms_4_w; // @[Reg.scala 16:16]
  reg  r_10_4_entries_perms_4_r; // @[Reg.scala 16:16]
  reg  r_10_4_entries_perms_5_d; // @[Reg.scala 16:16]
  reg  r_10_4_entries_perms_5_a; // @[Reg.scala 16:16]
  reg  r_10_4_entries_perms_5_g; // @[Reg.scala 16:16]
  reg  r_10_4_entries_perms_5_u; // @[Reg.scala 16:16]
  reg  r_10_4_entries_perms_5_x; // @[Reg.scala 16:16]
  reg  r_10_4_entries_perms_5_w; // @[Reg.scala 16:16]
  reg  r_10_4_entries_perms_5_r; // @[Reg.scala 16:16]
  reg  r_10_4_entries_perms_6_d; // @[Reg.scala 16:16]
  reg  r_10_4_entries_perms_6_a; // @[Reg.scala 16:16]
  reg  r_10_4_entries_perms_6_g; // @[Reg.scala 16:16]
  reg  r_10_4_entries_perms_6_u; // @[Reg.scala 16:16]
  reg  r_10_4_entries_perms_6_x; // @[Reg.scala 16:16]
  reg  r_10_4_entries_perms_6_w; // @[Reg.scala 16:16]
  reg  r_10_4_entries_perms_6_r; // @[Reg.scala 16:16]
  reg  r_10_4_entries_perms_7_d; // @[Reg.scala 16:16]
  reg  r_10_4_entries_perms_7_a; // @[Reg.scala 16:16]
  reg  r_10_4_entries_perms_7_g; // @[Reg.scala 16:16]
  reg  r_10_4_entries_perms_7_u; // @[Reg.scala 16:16]
  reg  r_10_4_entries_perms_7_x; // @[Reg.scala 16:16]
  reg  r_10_4_entries_perms_7_w; // @[Reg.scala 16:16]
  reg  r_10_4_entries_perms_7_r; // @[Reg.scala 16:16]
  reg  r_10_4_entries_prefetch; // @[Reg.scala 16:16]
  reg [38:0] r_10_4_ecc; // @[Reg.scala 16:16]
  reg [21:0] r_10_5_entries_tag; // @[Reg.scala 16:16]
  reg [15:0] r_10_5_entries_asid; // @[Reg.scala 16:16]
  reg [23:0] r_10_5_entries_ppns_0; // @[Reg.scala 16:16]
  reg [23:0] r_10_5_entries_ppns_1; // @[Reg.scala 16:16]
  reg [23:0] r_10_5_entries_ppns_2; // @[Reg.scala 16:16]
  reg [23:0] r_10_5_entries_ppns_3; // @[Reg.scala 16:16]
  reg [23:0] r_10_5_entries_ppns_4; // @[Reg.scala 16:16]
  reg [23:0] r_10_5_entries_ppns_5; // @[Reg.scala 16:16]
  reg [23:0] r_10_5_entries_ppns_6; // @[Reg.scala 16:16]
  reg [23:0] r_10_5_entries_ppns_7; // @[Reg.scala 16:16]
  reg  r_10_5_entries_vs_0; // @[Reg.scala 16:16]
  reg  r_10_5_entries_vs_1; // @[Reg.scala 16:16]
  reg  r_10_5_entries_vs_2; // @[Reg.scala 16:16]
  reg  r_10_5_entries_vs_3; // @[Reg.scala 16:16]
  reg  r_10_5_entries_vs_4; // @[Reg.scala 16:16]
  reg  r_10_5_entries_vs_5; // @[Reg.scala 16:16]
  reg  r_10_5_entries_vs_6; // @[Reg.scala 16:16]
  reg  r_10_5_entries_vs_7; // @[Reg.scala 16:16]
  reg  r_10_5_entries_perms_0_d; // @[Reg.scala 16:16]
  reg  r_10_5_entries_perms_0_a; // @[Reg.scala 16:16]
  reg  r_10_5_entries_perms_0_g; // @[Reg.scala 16:16]
  reg  r_10_5_entries_perms_0_u; // @[Reg.scala 16:16]
  reg  r_10_5_entries_perms_0_x; // @[Reg.scala 16:16]
  reg  r_10_5_entries_perms_0_w; // @[Reg.scala 16:16]
  reg  r_10_5_entries_perms_0_r; // @[Reg.scala 16:16]
  reg  r_10_5_entries_perms_1_d; // @[Reg.scala 16:16]
  reg  r_10_5_entries_perms_1_a; // @[Reg.scala 16:16]
  reg  r_10_5_entries_perms_1_g; // @[Reg.scala 16:16]
  reg  r_10_5_entries_perms_1_u; // @[Reg.scala 16:16]
  reg  r_10_5_entries_perms_1_x; // @[Reg.scala 16:16]
  reg  r_10_5_entries_perms_1_w; // @[Reg.scala 16:16]
  reg  r_10_5_entries_perms_1_r; // @[Reg.scala 16:16]
  reg  r_10_5_entries_perms_2_d; // @[Reg.scala 16:16]
  reg  r_10_5_entries_perms_2_a; // @[Reg.scala 16:16]
  reg  r_10_5_entries_perms_2_g; // @[Reg.scala 16:16]
  reg  r_10_5_entries_perms_2_u; // @[Reg.scala 16:16]
  reg  r_10_5_entries_perms_2_x; // @[Reg.scala 16:16]
  reg  r_10_5_entries_perms_2_w; // @[Reg.scala 16:16]
  reg  r_10_5_entries_perms_2_r; // @[Reg.scala 16:16]
  reg  r_10_5_entries_perms_3_d; // @[Reg.scala 16:16]
  reg  r_10_5_entries_perms_3_a; // @[Reg.scala 16:16]
  reg  r_10_5_entries_perms_3_g; // @[Reg.scala 16:16]
  reg  r_10_5_entries_perms_3_u; // @[Reg.scala 16:16]
  reg  r_10_5_entries_perms_3_x; // @[Reg.scala 16:16]
  reg  r_10_5_entries_perms_3_w; // @[Reg.scala 16:16]
  reg  r_10_5_entries_perms_3_r; // @[Reg.scala 16:16]
  reg  r_10_5_entries_perms_4_d; // @[Reg.scala 16:16]
  reg  r_10_5_entries_perms_4_a; // @[Reg.scala 16:16]
  reg  r_10_5_entries_perms_4_g; // @[Reg.scala 16:16]
  reg  r_10_5_entries_perms_4_u; // @[Reg.scala 16:16]
  reg  r_10_5_entries_perms_4_x; // @[Reg.scala 16:16]
  reg  r_10_5_entries_perms_4_w; // @[Reg.scala 16:16]
  reg  r_10_5_entries_perms_4_r; // @[Reg.scala 16:16]
  reg  r_10_5_entries_perms_5_d; // @[Reg.scala 16:16]
  reg  r_10_5_entries_perms_5_a; // @[Reg.scala 16:16]
  reg  r_10_5_entries_perms_5_g; // @[Reg.scala 16:16]
  reg  r_10_5_entries_perms_5_u; // @[Reg.scala 16:16]
  reg  r_10_5_entries_perms_5_x; // @[Reg.scala 16:16]
  reg  r_10_5_entries_perms_5_w; // @[Reg.scala 16:16]
  reg  r_10_5_entries_perms_5_r; // @[Reg.scala 16:16]
  reg  r_10_5_entries_perms_6_d; // @[Reg.scala 16:16]
  reg  r_10_5_entries_perms_6_a; // @[Reg.scala 16:16]
  reg  r_10_5_entries_perms_6_g; // @[Reg.scala 16:16]
  reg  r_10_5_entries_perms_6_u; // @[Reg.scala 16:16]
  reg  r_10_5_entries_perms_6_x; // @[Reg.scala 16:16]
  reg  r_10_5_entries_perms_6_w; // @[Reg.scala 16:16]
  reg  r_10_5_entries_perms_6_r; // @[Reg.scala 16:16]
  reg  r_10_5_entries_perms_7_d; // @[Reg.scala 16:16]
  reg  r_10_5_entries_perms_7_a; // @[Reg.scala 16:16]
  reg  r_10_5_entries_perms_7_g; // @[Reg.scala 16:16]
  reg  r_10_5_entries_perms_7_u; // @[Reg.scala 16:16]
  reg  r_10_5_entries_perms_7_x; // @[Reg.scala 16:16]
  reg  r_10_5_entries_perms_7_w; // @[Reg.scala 16:16]
  reg  r_10_5_entries_perms_7_r; // @[Reg.scala 16:16]
  reg  r_10_5_entries_prefetch; // @[Reg.scala 16:16]
  reg [38:0] r_10_5_ecc; // @[Reg.scala 16:16]
  reg [21:0] r_10_6_entries_tag; // @[Reg.scala 16:16]
  reg [15:0] r_10_6_entries_asid; // @[Reg.scala 16:16]
  reg [23:0] r_10_6_entries_ppns_0; // @[Reg.scala 16:16]
  reg [23:0] r_10_6_entries_ppns_1; // @[Reg.scala 16:16]
  reg [23:0] r_10_6_entries_ppns_2; // @[Reg.scala 16:16]
  reg [23:0] r_10_6_entries_ppns_3; // @[Reg.scala 16:16]
  reg [23:0] r_10_6_entries_ppns_4; // @[Reg.scala 16:16]
  reg [23:0] r_10_6_entries_ppns_5; // @[Reg.scala 16:16]
  reg [23:0] r_10_6_entries_ppns_6; // @[Reg.scala 16:16]
  reg [23:0] r_10_6_entries_ppns_7; // @[Reg.scala 16:16]
  reg  r_10_6_entries_vs_0; // @[Reg.scala 16:16]
  reg  r_10_6_entries_vs_1; // @[Reg.scala 16:16]
  reg  r_10_6_entries_vs_2; // @[Reg.scala 16:16]
  reg  r_10_6_entries_vs_3; // @[Reg.scala 16:16]
  reg  r_10_6_entries_vs_4; // @[Reg.scala 16:16]
  reg  r_10_6_entries_vs_5; // @[Reg.scala 16:16]
  reg  r_10_6_entries_vs_6; // @[Reg.scala 16:16]
  reg  r_10_6_entries_vs_7; // @[Reg.scala 16:16]
  reg  r_10_6_entries_perms_0_d; // @[Reg.scala 16:16]
  reg  r_10_6_entries_perms_0_a; // @[Reg.scala 16:16]
  reg  r_10_6_entries_perms_0_g; // @[Reg.scala 16:16]
  reg  r_10_6_entries_perms_0_u; // @[Reg.scala 16:16]
  reg  r_10_6_entries_perms_0_x; // @[Reg.scala 16:16]
  reg  r_10_6_entries_perms_0_w; // @[Reg.scala 16:16]
  reg  r_10_6_entries_perms_0_r; // @[Reg.scala 16:16]
  reg  r_10_6_entries_perms_1_d; // @[Reg.scala 16:16]
  reg  r_10_6_entries_perms_1_a; // @[Reg.scala 16:16]
  reg  r_10_6_entries_perms_1_g; // @[Reg.scala 16:16]
  reg  r_10_6_entries_perms_1_u; // @[Reg.scala 16:16]
  reg  r_10_6_entries_perms_1_x; // @[Reg.scala 16:16]
  reg  r_10_6_entries_perms_1_w; // @[Reg.scala 16:16]
  reg  r_10_6_entries_perms_1_r; // @[Reg.scala 16:16]
  reg  r_10_6_entries_perms_2_d; // @[Reg.scala 16:16]
  reg  r_10_6_entries_perms_2_a; // @[Reg.scala 16:16]
  reg  r_10_6_entries_perms_2_g; // @[Reg.scala 16:16]
  reg  r_10_6_entries_perms_2_u; // @[Reg.scala 16:16]
  reg  r_10_6_entries_perms_2_x; // @[Reg.scala 16:16]
  reg  r_10_6_entries_perms_2_w; // @[Reg.scala 16:16]
  reg  r_10_6_entries_perms_2_r; // @[Reg.scala 16:16]
  reg  r_10_6_entries_perms_3_d; // @[Reg.scala 16:16]
  reg  r_10_6_entries_perms_3_a; // @[Reg.scala 16:16]
  reg  r_10_6_entries_perms_3_g; // @[Reg.scala 16:16]
  reg  r_10_6_entries_perms_3_u; // @[Reg.scala 16:16]
  reg  r_10_6_entries_perms_3_x; // @[Reg.scala 16:16]
  reg  r_10_6_entries_perms_3_w; // @[Reg.scala 16:16]
  reg  r_10_6_entries_perms_3_r; // @[Reg.scala 16:16]
  reg  r_10_6_entries_perms_4_d; // @[Reg.scala 16:16]
  reg  r_10_6_entries_perms_4_a; // @[Reg.scala 16:16]
  reg  r_10_6_entries_perms_4_g; // @[Reg.scala 16:16]
  reg  r_10_6_entries_perms_4_u; // @[Reg.scala 16:16]
  reg  r_10_6_entries_perms_4_x; // @[Reg.scala 16:16]
  reg  r_10_6_entries_perms_4_w; // @[Reg.scala 16:16]
  reg  r_10_6_entries_perms_4_r; // @[Reg.scala 16:16]
  reg  r_10_6_entries_perms_5_d; // @[Reg.scala 16:16]
  reg  r_10_6_entries_perms_5_a; // @[Reg.scala 16:16]
  reg  r_10_6_entries_perms_5_g; // @[Reg.scala 16:16]
  reg  r_10_6_entries_perms_5_u; // @[Reg.scala 16:16]
  reg  r_10_6_entries_perms_5_x; // @[Reg.scala 16:16]
  reg  r_10_6_entries_perms_5_w; // @[Reg.scala 16:16]
  reg  r_10_6_entries_perms_5_r; // @[Reg.scala 16:16]
  reg  r_10_6_entries_perms_6_d; // @[Reg.scala 16:16]
  reg  r_10_6_entries_perms_6_a; // @[Reg.scala 16:16]
  reg  r_10_6_entries_perms_6_g; // @[Reg.scala 16:16]
  reg  r_10_6_entries_perms_6_u; // @[Reg.scala 16:16]
  reg  r_10_6_entries_perms_6_x; // @[Reg.scala 16:16]
  reg  r_10_6_entries_perms_6_w; // @[Reg.scala 16:16]
  reg  r_10_6_entries_perms_6_r; // @[Reg.scala 16:16]
  reg  r_10_6_entries_perms_7_d; // @[Reg.scala 16:16]
  reg  r_10_6_entries_perms_7_a; // @[Reg.scala 16:16]
  reg  r_10_6_entries_perms_7_g; // @[Reg.scala 16:16]
  reg  r_10_6_entries_perms_7_u; // @[Reg.scala 16:16]
  reg  r_10_6_entries_perms_7_x; // @[Reg.scala 16:16]
  reg  r_10_6_entries_perms_7_w; // @[Reg.scala 16:16]
  reg  r_10_6_entries_perms_7_r; // @[Reg.scala 16:16]
  reg  r_10_6_entries_prefetch; // @[Reg.scala 16:16]
  reg [38:0] r_10_6_ecc; // @[Reg.scala 16:16]
  reg [21:0] r_10_7_entries_tag; // @[Reg.scala 16:16]
  reg [15:0] r_10_7_entries_asid; // @[Reg.scala 16:16]
  reg [23:0] r_10_7_entries_ppns_0; // @[Reg.scala 16:16]
  reg [23:0] r_10_7_entries_ppns_1; // @[Reg.scala 16:16]
  reg [23:0] r_10_7_entries_ppns_2; // @[Reg.scala 16:16]
  reg [23:0] r_10_7_entries_ppns_3; // @[Reg.scala 16:16]
  reg [23:0] r_10_7_entries_ppns_4; // @[Reg.scala 16:16]
  reg [23:0] r_10_7_entries_ppns_5; // @[Reg.scala 16:16]
  reg [23:0] r_10_7_entries_ppns_6; // @[Reg.scala 16:16]
  reg [23:0] r_10_7_entries_ppns_7; // @[Reg.scala 16:16]
  reg  r_10_7_entries_vs_0; // @[Reg.scala 16:16]
  reg  r_10_7_entries_vs_1; // @[Reg.scala 16:16]
  reg  r_10_7_entries_vs_2; // @[Reg.scala 16:16]
  reg  r_10_7_entries_vs_3; // @[Reg.scala 16:16]
  reg  r_10_7_entries_vs_4; // @[Reg.scala 16:16]
  reg  r_10_7_entries_vs_5; // @[Reg.scala 16:16]
  reg  r_10_7_entries_vs_6; // @[Reg.scala 16:16]
  reg  r_10_7_entries_vs_7; // @[Reg.scala 16:16]
  reg  r_10_7_entries_perms_0_d; // @[Reg.scala 16:16]
  reg  r_10_7_entries_perms_0_a; // @[Reg.scala 16:16]
  reg  r_10_7_entries_perms_0_g; // @[Reg.scala 16:16]
  reg  r_10_7_entries_perms_0_u; // @[Reg.scala 16:16]
  reg  r_10_7_entries_perms_0_x; // @[Reg.scala 16:16]
  reg  r_10_7_entries_perms_0_w; // @[Reg.scala 16:16]
  reg  r_10_7_entries_perms_0_r; // @[Reg.scala 16:16]
  reg  r_10_7_entries_perms_1_d; // @[Reg.scala 16:16]
  reg  r_10_7_entries_perms_1_a; // @[Reg.scala 16:16]
  reg  r_10_7_entries_perms_1_g; // @[Reg.scala 16:16]
  reg  r_10_7_entries_perms_1_u; // @[Reg.scala 16:16]
  reg  r_10_7_entries_perms_1_x; // @[Reg.scala 16:16]
  reg  r_10_7_entries_perms_1_w; // @[Reg.scala 16:16]
  reg  r_10_7_entries_perms_1_r; // @[Reg.scala 16:16]
  reg  r_10_7_entries_perms_2_d; // @[Reg.scala 16:16]
  reg  r_10_7_entries_perms_2_a; // @[Reg.scala 16:16]
  reg  r_10_7_entries_perms_2_g; // @[Reg.scala 16:16]
  reg  r_10_7_entries_perms_2_u; // @[Reg.scala 16:16]
  reg  r_10_7_entries_perms_2_x; // @[Reg.scala 16:16]
  reg  r_10_7_entries_perms_2_w; // @[Reg.scala 16:16]
  reg  r_10_7_entries_perms_2_r; // @[Reg.scala 16:16]
  reg  r_10_7_entries_perms_3_d; // @[Reg.scala 16:16]
  reg  r_10_7_entries_perms_3_a; // @[Reg.scala 16:16]
  reg  r_10_7_entries_perms_3_g; // @[Reg.scala 16:16]
  reg  r_10_7_entries_perms_3_u; // @[Reg.scala 16:16]
  reg  r_10_7_entries_perms_3_x; // @[Reg.scala 16:16]
  reg  r_10_7_entries_perms_3_w; // @[Reg.scala 16:16]
  reg  r_10_7_entries_perms_3_r; // @[Reg.scala 16:16]
  reg  r_10_7_entries_perms_4_d; // @[Reg.scala 16:16]
  reg  r_10_7_entries_perms_4_a; // @[Reg.scala 16:16]
  reg  r_10_7_entries_perms_4_g; // @[Reg.scala 16:16]
  reg  r_10_7_entries_perms_4_u; // @[Reg.scala 16:16]
  reg  r_10_7_entries_perms_4_x; // @[Reg.scala 16:16]
  reg  r_10_7_entries_perms_4_w; // @[Reg.scala 16:16]
  reg  r_10_7_entries_perms_4_r; // @[Reg.scala 16:16]
  reg  r_10_7_entries_perms_5_d; // @[Reg.scala 16:16]
  reg  r_10_7_entries_perms_5_a; // @[Reg.scala 16:16]
  reg  r_10_7_entries_perms_5_g; // @[Reg.scala 16:16]
  reg  r_10_7_entries_perms_5_u; // @[Reg.scala 16:16]
  reg  r_10_7_entries_perms_5_x; // @[Reg.scala 16:16]
  reg  r_10_7_entries_perms_5_w; // @[Reg.scala 16:16]
  reg  r_10_7_entries_perms_5_r; // @[Reg.scala 16:16]
  reg  r_10_7_entries_perms_6_d; // @[Reg.scala 16:16]
  reg  r_10_7_entries_perms_6_a; // @[Reg.scala 16:16]
  reg  r_10_7_entries_perms_6_g; // @[Reg.scala 16:16]
  reg  r_10_7_entries_perms_6_u; // @[Reg.scala 16:16]
  reg  r_10_7_entries_perms_6_x; // @[Reg.scala 16:16]
  reg  r_10_7_entries_perms_6_w; // @[Reg.scala 16:16]
  reg  r_10_7_entries_perms_6_r; // @[Reg.scala 16:16]
  reg  r_10_7_entries_perms_7_d; // @[Reg.scala 16:16]
  reg  r_10_7_entries_perms_7_a; // @[Reg.scala 16:16]
  reg  r_10_7_entries_perms_7_g; // @[Reg.scala 16:16]
  reg  r_10_7_entries_perms_7_u; // @[Reg.scala 16:16]
  reg  r_10_7_entries_perms_7_x; // @[Reg.scala 16:16]
  reg  r_10_7_entries_perms_7_w; // @[Reg.scala 16:16]
  reg  r_10_7_entries_perms_7_r; // @[Reg.scala 16:16]
  reg  r_10_7_entries_prefetch; // @[Reg.scala 16:16]
  reg [38:0] r_10_7_ecc; // @[Reg.scala 16:16]
  wire [21:0] _GEN_276 = stageDelay_valid_1cycle ? l3_io_rresp_data_0_entries_tag : r_10_0_entries_tag; // @[Reg.scala 16:16 17:{18,22}]
  wire [15:0] _GEN_277 = stageDelay_valid_1cycle ? l3_io_rresp_data_0_entries_asid : r_10_0_entries_asid; // @[Reg.scala 16:16 17:{18,22}]
  wire [21:0] _GEN_352 = stageDelay_valid_1cycle ? l3_io_rresp_data_1_entries_tag : r_10_1_entries_tag; // @[Reg.scala 16:16 17:{18,22}]
  wire [15:0] _GEN_353 = stageDelay_valid_1cycle ? l3_io_rresp_data_1_entries_asid : r_10_1_entries_asid; // @[Reg.scala 16:16 17:{18,22}]
  wire [21:0] _GEN_428 = stageDelay_valid_1cycle ? l3_io_rresp_data_2_entries_tag : r_10_2_entries_tag; // @[Reg.scala 16:16 17:{18,22}]
  wire [15:0] _GEN_429 = stageDelay_valid_1cycle ? l3_io_rresp_data_2_entries_asid : r_10_2_entries_asid; // @[Reg.scala 16:16 17:{18,22}]
  wire [21:0] _GEN_504 = stageDelay_valid_1cycle ? l3_io_rresp_data_3_entries_tag : r_10_3_entries_tag; // @[Reg.scala 16:16 17:{18,22}]
  wire [15:0] _GEN_505 = stageDelay_valid_1cycle ? l3_io_rresp_data_3_entries_asid : r_10_3_entries_asid; // @[Reg.scala 16:16 17:{18,22}]
  wire [21:0] _GEN_580 = stageDelay_valid_1cycle ? l3_io_rresp_data_4_entries_tag : r_10_4_entries_tag; // @[Reg.scala 16:16 17:{18,22}]
  wire [15:0] _GEN_581 = stageDelay_valid_1cycle ? l3_io_rresp_data_4_entries_asid : r_10_4_entries_asid; // @[Reg.scala 16:16 17:{18,22}]
  wire [21:0] _GEN_656 = stageDelay_valid_1cycle ? l3_io_rresp_data_5_entries_tag : r_10_5_entries_tag; // @[Reg.scala 16:16 17:{18,22}]
  wire [15:0] _GEN_657 = stageDelay_valid_1cycle ? l3_io_rresp_data_5_entries_asid : r_10_5_entries_asid; // @[Reg.scala 16:16 17:{18,22}]
  wire [21:0] _GEN_732 = stageDelay_valid_1cycle ? l3_io_rresp_data_6_entries_tag : r_10_6_entries_tag; // @[Reg.scala 16:16 17:{18,22}]
  wire [15:0] _GEN_733 = stageDelay_valid_1cycle ? l3_io_rresp_data_6_entries_asid : r_10_6_entries_asid; // @[Reg.scala 16:16 17:{18,22}]
  wire [21:0] _GEN_808 = stageDelay_valid_1cycle ? l3_io_rresp_data_7_entries_tag : r_10_7_entries_tag; // @[Reg.scala 16:16 17:{18,22}]
  wire [15:0] _GEN_809 = stageDelay_valid_1cycle ? l3_io_rresp_data_7_entries_asid : r_10_7_entries_asid; // @[Reg.scala 16:16 17:{18,22}]
  reg [7:0] r_11; // @[Reg.scala 16:16]
  wire  asid_hit_12 = _GEN_277 == io_csr_dup_2_satp_asid; // @[MMUBundle.scala 654:59]
  wire  _T_156 = asid_hit_12 & _GEN_276 == data_req_info_vpn[26:5]; // @[MMUBundle.scala 655:14]
  wire  _T_158 = _T_156 & r_11[0]; // @[PageTableCache.scala 315:63]
  wire  asid_hit_13 = _GEN_353 == io_csr_dup_2_satp_asid; // @[MMUBundle.scala 654:59]
  wire  _T_161 = asid_hit_13 & _GEN_352 == data_req_info_vpn[26:5]; // @[MMUBundle.scala 655:14]
  wire  _T_163 = _T_161 & r_11[1]; // @[PageTableCache.scala 315:63]
  wire  asid_hit_14 = _GEN_429 == io_csr_dup_2_satp_asid; // @[MMUBundle.scala 654:59]
  wire  _T_166 = asid_hit_14 & _GEN_428 == data_req_info_vpn[26:5]; // @[MMUBundle.scala 655:14]
  wire  _T_168 = _T_166 & r_11[2]; // @[PageTableCache.scala 315:63]
  wire  asid_hit_15 = _GEN_505 == io_csr_dup_2_satp_asid; // @[MMUBundle.scala 654:59]
  wire  _T_171 = asid_hit_15 & _GEN_504 == data_req_info_vpn[26:5]; // @[MMUBundle.scala 655:14]
  wire  _T_173 = _T_171 & r_11[3]; // @[PageTableCache.scala 315:63]
  wire  asid_hit_16 = _GEN_581 == io_csr_dup_2_satp_asid; // @[MMUBundle.scala 654:59]
  wire  _T_176 = asid_hit_16 & _GEN_580 == data_req_info_vpn[26:5]; // @[MMUBundle.scala 655:14]
  wire  _T_178 = _T_176 & r_11[4]; // @[PageTableCache.scala 315:63]
  wire  asid_hit_17 = _GEN_657 == io_csr_dup_2_satp_asid; // @[MMUBundle.scala 654:59]
  wire  _T_181 = asid_hit_17 & _GEN_656 == data_req_info_vpn[26:5]; // @[MMUBundle.scala 655:14]
  wire  _T_183 = _T_181 & r_11[5]; // @[PageTableCache.scala 315:63]
  wire  asid_hit_18 = _GEN_733 == io_csr_dup_2_satp_asid; // @[MMUBundle.scala 654:59]
  wire  _T_186 = asid_hit_18 & _GEN_732 == data_req_info_vpn[26:5]; // @[MMUBundle.scala 655:14]
  wire  _T_188 = _T_186 & r_11[6]; // @[PageTableCache.scala 315:63]
  wire  asid_hit_19 = _GEN_809 == io_csr_dup_2_satp_asid; // @[MMUBundle.scala 654:59]
  wire  _T_191 = asid_hit_19 & _GEN_808 == data_req_info_vpn[26:5]; // @[MMUBundle.scala 655:14]
  wire  _T_193 = _T_191 & r_11[7]; // @[PageTableCache.scala 315:63]
  reg [21:0] l3_ramDatas_0_entries_tag; // @[Reg.scala 16:16]
  reg [15:0] l3_ramDatas_0_entries_asid; // @[Reg.scala 16:16]
  reg [23:0] l3_ramDatas_0_entries_ppns_0; // @[Reg.scala 16:16]
  reg [23:0] l3_ramDatas_0_entries_ppns_1; // @[Reg.scala 16:16]
  reg [23:0] l3_ramDatas_0_entries_ppns_2; // @[Reg.scala 16:16]
  reg [23:0] l3_ramDatas_0_entries_ppns_3; // @[Reg.scala 16:16]
  reg [23:0] l3_ramDatas_0_entries_ppns_4; // @[Reg.scala 16:16]
  reg [23:0] l3_ramDatas_0_entries_ppns_5; // @[Reg.scala 16:16]
  reg [23:0] l3_ramDatas_0_entries_ppns_6; // @[Reg.scala 16:16]
  reg [23:0] l3_ramDatas_0_entries_ppns_7; // @[Reg.scala 16:16]
  reg  l3_ramDatas_0_entries_vs_0; // @[Reg.scala 16:16]
  reg  l3_ramDatas_0_entries_vs_1; // @[Reg.scala 16:16]
  reg  l3_ramDatas_0_entries_vs_2; // @[Reg.scala 16:16]
  reg  l3_ramDatas_0_entries_vs_3; // @[Reg.scala 16:16]
  reg  l3_ramDatas_0_entries_vs_4; // @[Reg.scala 16:16]
  reg  l3_ramDatas_0_entries_vs_5; // @[Reg.scala 16:16]
  reg  l3_ramDatas_0_entries_vs_6; // @[Reg.scala 16:16]
  reg  l3_ramDatas_0_entries_vs_7; // @[Reg.scala 16:16]
  reg  l3_ramDatas_0_entries_perms_0_d; // @[Reg.scala 16:16]
  reg  l3_ramDatas_0_entries_perms_0_a; // @[Reg.scala 16:16]
  reg  l3_ramDatas_0_entries_perms_0_g; // @[Reg.scala 16:16]
  reg  l3_ramDatas_0_entries_perms_0_u; // @[Reg.scala 16:16]
  reg  l3_ramDatas_0_entries_perms_0_x; // @[Reg.scala 16:16]
  reg  l3_ramDatas_0_entries_perms_0_w; // @[Reg.scala 16:16]
  reg  l3_ramDatas_0_entries_perms_0_r; // @[Reg.scala 16:16]
  reg  l3_ramDatas_0_entries_perms_1_d; // @[Reg.scala 16:16]
  reg  l3_ramDatas_0_entries_perms_1_a; // @[Reg.scala 16:16]
  reg  l3_ramDatas_0_entries_perms_1_g; // @[Reg.scala 16:16]
  reg  l3_ramDatas_0_entries_perms_1_u; // @[Reg.scala 16:16]
  reg  l3_ramDatas_0_entries_perms_1_x; // @[Reg.scala 16:16]
  reg  l3_ramDatas_0_entries_perms_1_w; // @[Reg.scala 16:16]
  reg  l3_ramDatas_0_entries_perms_1_r; // @[Reg.scala 16:16]
  reg  l3_ramDatas_0_entries_perms_2_d; // @[Reg.scala 16:16]
  reg  l3_ramDatas_0_entries_perms_2_a; // @[Reg.scala 16:16]
  reg  l3_ramDatas_0_entries_perms_2_g; // @[Reg.scala 16:16]
  reg  l3_ramDatas_0_entries_perms_2_u; // @[Reg.scala 16:16]
  reg  l3_ramDatas_0_entries_perms_2_x; // @[Reg.scala 16:16]
  reg  l3_ramDatas_0_entries_perms_2_w; // @[Reg.scala 16:16]
  reg  l3_ramDatas_0_entries_perms_2_r; // @[Reg.scala 16:16]
  reg  l3_ramDatas_0_entries_perms_3_d; // @[Reg.scala 16:16]
  reg  l3_ramDatas_0_entries_perms_3_a; // @[Reg.scala 16:16]
  reg  l3_ramDatas_0_entries_perms_3_g; // @[Reg.scala 16:16]
  reg  l3_ramDatas_0_entries_perms_3_u; // @[Reg.scala 16:16]
  reg  l3_ramDatas_0_entries_perms_3_x; // @[Reg.scala 16:16]
  reg  l3_ramDatas_0_entries_perms_3_w; // @[Reg.scala 16:16]
  reg  l3_ramDatas_0_entries_perms_3_r; // @[Reg.scala 16:16]
  reg  l3_ramDatas_0_entries_perms_4_d; // @[Reg.scala 16:16]
  reg  l3_ramDatas_0_entries_perms_4_a; // @[Reg.scala 16:16]
  reg  l3_ramDatas_0_entries_perms_4_g; // @[Reg.scala 16:16]
  reg  l3_ramDatas_0_entries_perms_4_u; // @[Reg.scala 16:16]
  reg  l3_ramDatas_0_entries_perms_4_x; // @[Reg.scala 16:16]
  reg  l3_ramDatas_0_entries_perms_4_w; // @[Reg.scala 16:16]
  reg  l3_ramDatas_0_entries_perms_4_r; // @[Reg.scala 16:16]
  reg  l3_ramDatas_0_entries_perms_5_d; // @[Reg.scala 16:16]
  reg  l3_ramDatas_0_entries_perms_5_a; // @[Reg.scala 16:16]
  reg  l3_ramDatas_0_entries_perms_5_g; // @[Reg.scala 16:16]
  reg  l3_ramDatas_0_entries_perms_5_u; // @[Reg.scala 16:16]
  reg  l3_ramDatas_0_entries_perms_5_x; // @[Reg.scala 16:16]
  reg  l3_ramDatas_0_entries_perms_5_w; // @[Reg.scala 16:16]
  reg  l3_ramDatas_0_entries_perms_5_r; // @[Reg.scala 16:16]
  reg  l3_ramDatas_0_entries_perms_6_d; // @[Reg.scala 16:16]
  reg  l3_ramDatas_0_entries_perms_6_a; // @[Reg.scala 16:16]
  reg  l3_ramDatas_0_entries_perms_6_g; // @[Reg.scala 16:16]
  reg  l3_ramDatas_0_entries_perms_6_u; // @[Reg.scala 16:16]
  reg  l3_ramDatas_0_entries_perms_6_x; // @[Reg.scala 16:16]
  reg  l3_ramDatas_0_entries_perms_6_w; // @[Reg.scala 16:16]
  reg  l3_ramDatas_0_entries_perms_6_r; // @[Reg.scala 16:16]
  reg  l3_ramDatas_0_entries_perms_7_d; // @[Reg.scala 16:16]
  reg  l3_ramDatas_0_entries_perms_7_a; // @[Reg.scala 16:16]
  reg  l3_ramDatas_0_entries_perms_7_g; // @[Reg.scala 16:16]
  reg  l3_ramDatas_0_entries_perms_7_u; // @[Reg.scala 16:16]
  reg  l3_ramDatas_0_entries_perms_7_x; // @[Reg.scala 16:16]
  reg  l3_ramDatas_0_entries_perms_7_w; // @[Reg.scala 16:16]
  reg  l3_ramDatas_0_entries_perms_7_r; // @[Reg.scala 16:16]
  reg  l3_ramDatas_0_entries_prefetch; // @[Reg.scala 16:16]
  reg [38:0] l3_ramDatas_0_ecc; // @[Reg.scala 16:16]
  reg [21:0] l3_ramDatas_1_entries_tag; // @[Reg.scala 16:16]
  reg [15:0] l3_ramDatas_1_entries_asid; // @[Reg.scala 16:16]
  reg [23:0] l3_ramDatas_1_entries_ppns_0; // @[Reg.scala 16:16]
  reg [23:0] l3_ramDatas_1_entries_ppns_1; // @[Reg.scala 16:16]
  reg [23:0] l3_ramDatas_1_entries_ppns_2; // @[Reg.scala 16:16]
  reg [23:0] l3_ramDatas_1_entries_ppns_3; // @[Reg.scala 16:16]
  reg [23:0] l3_ramDatas_1_entries_ppns_4; // @[Reg.scala 16:16]
  reg [23:0] l3_ramDatas_1_entries_ppns_5; // @[Reg.scala 16:16]
  reg [23:0] l3_ramDatas_1_entries_ppns_6; // @[Reg.scala 16:16]
  reg [23:0] l3_ramDatas_1_entries_ppns_7; // @[Reg.scala 16:16]
  reg  l3_ramDatas_1_entries_vs_0; // @[Reg.scala 16:16]
  reg  l3_ramDatas_1_entries_vs_1; // @[Reg.scala 16:16]
  reg  l3_ramDatas_1_entries_vs_2; // @[Reg.scala 16:16]
  reg  l3_ramDatas_1_entries_vs_3; // @[Reg.scala 16:16]
  reg  l3_ramDatas_1_entries_vs_4; // @[Reg.scala 16:16]
  reg  l3_ramDatas_1_entries_vs_5; // @[Reg.scala 16:16]
  reg  l3_ramDatas_1_entries_vs_6; // @[Reg.scala 16:16]
  reg  l3_ramDatas_1_entries_vs_7; // @[Reg.scala 16:16]
  reg  l3_ramDatas_1_entries_perms_0_d; // @[Reg.scala 16:16]
  reg  l3_ramDatas_1_entries_perms_0_a; // @[Reg.scala 16:16]
  reg  l3_ramDatas_1_entries_perms_0_g; // @[Reg.scala 16:16]
  reg  l3_ramDatas_1_entries_perms_0_u; // @[Reg.scala 16:16]
  reg  l3_ramDatas_1_entries_perms_0_x; // @[Reg.scala 16:16]
  reg  l3_ramDatas_1_entries_perms_0_w; // @[Reg.scala 16:16]
  reg  l3_ramDatas_1_entries_perms_0_r; // @[Reg.scala 16:16]
  reg  l3_ramDatas_1_entries_perms_1_d; // @[Reg.scala 16:16]
  reg  l3_ramDatas_1_entries_perms_1_a; // @[Reg.scala 16:16]
  reg  l3_ramDatas_1_entries_perms_1_g; // @[Reg.scala 16:16]
  reg  l3_ramDatas_1_entries_perms_1_u; // @[Reg.scala 16:16]
  reg  l3_ramDatas_1_entries_perms_1_x; // @[Reg.scala 16:16]
  reg  l3_ramDatas_1_entries_perms_1_w; // @[Reg.scala 16:16]
  reg  l3_ramDatas_1_entries_perms_1_r; // @[Reg.scala 16:16]
  reg  l3_ramDatas_1_entries_perms_2_d; // @[Reg.scala 16:16]
  reg  l3_ramDatas_1_entries_perms_2_a; // @[Reg.scala 16:16]
  reg  l3_ramDatas_1_entries_perms_2_g; // @[Reg.scala 16:16]
  reg  l3_ramDatas_1_entries_perms_2_u; // @[Reg.scala 16:16]
  reg  l3_ramDatas_1_entries_perms_2_x; // @[Reg.scala 16:16]
  reg  l3_ramDatas_1_entries_perms_2_w; // @[Reg.scala 16:16]
  reg  l3_ramDatas_1_entries_perms_2_r; // @[Reg.scala 16:16]
  reg  l3_ramDatas_1_entries_perms_3_d; // @[Reg.scala 16:16]
  reg  l3_ramDatas_1_entries_perms_3_a; // @[Reg.scala 16:16]
  reg  l3_ramDatas_1_entries_perms_3_g; // @[Reg.scala 16:16]
  reg  l3_ramDatas_1_entries_perms_3_u; // @[Reg.scala 16:16]
  reg  l3_ramDatas_1_entries_perms_3_x; // @[Reg.scala 16:16]
  reg  l3_ramDatas_1_entries_perms_3_w; // @[Reg.scala 16:16]
  reg  l3_ramDatas_1_entries_perms_3_r; // @[Reg.scala 16:16]
  reg  l3_ramDatas_1_entries_perms_4_d; // @[Reg.scala 16:16]
  reg  l3_ramDatas_1_entries_perms_4_a; // @[Reg.scala 16:16]
  reg  l3_ramDatas_1_entries_perms_4_g; // @[Reg.scala 16:16]
  reg  l3_ramDatas_1_entries_perms_4_u; // @[Reg.scala 16:16]
  reg  l3_ramDatas_1_entries_perms_4_x; // @[Reg.scala 16:16]
  reg  l3_ramDatas_1_entries_perms_4_w; // @[Reg.scala 16:16]
  reg  l3_ramDatas_1_entries_perms_4_r; // @[Reg.scala 16:16]
  reg  l3_ramDatas_1_entries_perms_5_d; // @[Reg.scala 16:16]
  reg  l3_ramDatas_1_entries_perms_5_a; // @[Reg.scala 16:16]
  reg  l3_ramDatas_1_entries_perms_5_g; // @[Reg.scala 16:16]
  reg  l3_ramDatas_1_entries_perms_5_u; // @[Reg.scala 16:16]
  reg  l3_ramDatas_1_entries_perms_5_x; // @[Reg.scala 16:16]
  reg  l3_ramDatas_1_entries_perms_5_w; // @[Reg.scala 16:16]
  reg  l3_ramDatas_1_entries_perms_5_r; // @[Reg.scala 16:16]
  reg  l3_ramDatas_1_entries_perms_6_d; // @[Reg.scala 16:16]
  reg  l3_ramDatas_1_entries_perms_6_a; // @[Reg.scala 16:16]
  reg  l3_ramDatas_1_entries_perms_6_g; // @[Reg.scala 16:16]
  reg  l3_ramDatas_1_entries_perms_6_u; // @[Reg.scala 16:16]
  reg  l3_ramDatas_1_entries_perms_6_x; // @[Reg.scala 16:16]
  reg  l3_ramDatas_1_entries_perms_6_w; // @[Reg.scala 16:16]
  reg  l3_ramDatas_1_entries_perms_6_r; // @[Reg.scala 16:16]
  reg  l3_ramDatas_1_entries_perms_7_d; // @[Reg.scala 16:16]
  reg  l3_ramDatas_1_entries_perms_7_a; // @[Reg.scala 16:16]
  reg  l3_ramDatas_1_entries_perms_7_g; // @[Reg.scala 16:16]
  reg  l3_ramDatas_1_entries_perms_7_u; // @[Reg.scala 16:16]
  reg  l3_ramDatas_1_entries_perms_7_x; // @[Reg.scala 16:16]
  reg  l3_ramDatas_1_entries_perms_7_w; // @[Reg.scala 16:16]
  reg  l3_ramDatas_1_entries_perms_7_r; // @[Reg.scala 16:16]
  reg  l3_ramDatas_1_entries_prefetch; // @[Reg.scala 16:16]
  reg [38:0] l3_ramDatas_1_ecc; // @[Reg.scala 16:16]
  reg [21:0] l3_ramDatas_2_entries_tag; // @[Reg.scala 16:16]
  reg [15:0] l3_ramDatas_2_entries_asid; // @[Reg.scala 16:16]
  reg [23:0] l3_ramDatas_2_entries_ppns_0; // @[Reg.scala 16:16]
  reg [23:0] l3_ramDatas_2_entries_ppns_1; // @[Reg.scala 16:16]
  reg [23:0] l3_ramDatas_2_entries_ppns_2; // @[Reg.scala 16:16]
  reg [23:0] l3_ramDatas_2_entries_ppns_3; // @[Reg.scala 16:16]
  reg [23:0] l3_ramDatas_2_entries_ppns_4; // @[Reg.scala 16:16]
  reg [23:0] l3_ramDatas_2_entries_ppns_5; // @[Reg.scala 16:16]
  reg [23:0] l3_ramDatas_2_entries_ppns_6; // @[Reg.scala 16:16]
  reg [23:0] l3_ramDatas_2_entries_ppns_7; // @[Reg.scala 16:16]
  reg  l3_ramDatas_2_entries_vs_0; // @[Reg.scala 16:16]
  reg  l3_ramDatas_2_entries_vs_1; // @[Reg.scala 16:16]
  reg  l3_ramDatas_2_entries_vs_2; // @[Reg.scala 16:16]
  reg  l3_ramDatas_2_entries_vs_3; // @[Reg.scala 16:16]
  reg  l3_ramDatas_2_entries_vs_4; // @[Reg.scala 16:16]
  reg  l3_ramDatas_2_entries_vs_5; // @[Reg.scala 16:16]
  reg  l3_ramDatas_2_entries_vs_6; // @[Reg.scala 16:16]
  reg  l3_ramDatas_2_entries_vs_7; // @[Reg.scala 16:16]
  reg  l3_ramDatas_2_entries_perms_0_d; // @[Reg.scala 16:16]
  reg  l3_ramDatas_2_entries_perms_0_a; // @[Reg.scala 16:16]
  reg  l3_ramDatas_2_entries_perms_0_g; // @[Reg.scala 16:16]
  reg  l3_ramDatas_2_entries_perms_0_u; // @[Reg.scala 16:16]
  reg  l3_ramDatas_2_entries_perms_0_x; // @[Reg.scala 16:16]
  reg  l3_ramDatas_2_entries_perms_0_w; // @[Reg.scala 16:16]
  reg  l3_ramDatas_2_entries_perms_0_r; // @[Reg.scala 16:16]
  reg  l3_ramDatas_2_entries_perms_1_d; // @[Reg.scala 16:16]
  reg  l3_ramDatas_2_entries_perms_1_a; // @[Reg.scala 16:16]
  reg  l3_ramDatas_2_entries_perms_1_g; // @[Reg.scala 16:16]
  reg  l3_ramDatas_2_entries_perms_1_u; // @[Reg.scala 16:16]
  reg  l3_ramDatas_2_entries_perms_1_x; // @[Reg.scala 16:16]
  reg  l3_ramDatas_2_entries_perms_1_w; // @[Reg.scala 16:16]
  reg  l3_ramDatas_2_entries_perms_1_r; // @[Reg.scala 16:16]
  reg  l3_ramDatas_2_entries_perms_2_d; // @[Reg.scala 16:16]
  reg  l3_ramDatas_2_entries_perms_2_a; // @[Reg.scala 16:16]
  reg  l3_ramDatas_2_entries_perms_2_g; // @[Reg.scala 16:16]
  reg  l3_ramDatas_2_entries_perms_2_u; // @[Reg.scala 16:16]
  reg  l3_ramDatas_2_entries_perms_2_x; // @[Reg.scala 16:16]
  reg  l3_ramDatas_2_entries_perms_2_w; // @[Reg.scala 16:16]
  reg  l3_ramDatas_2_entries_perms_2_r; // @[Reg.scala 16:16]
  reg  l3_ramDatas_2_entries_perms_3_d; // @[Reg.scala 16:16]
  reg  l3_ramDatas_2_entries_perms_3_a; // @[Reg.scala 16:16]
  reg  l3_ramDatas_2_entries_perms_3_g; // @[Reg.scala 16:16]
  reg  l3_ramDatas_2_entries_perms_3_u; // @[Reg.scala 16:16]
  reg  l3_ramDatas_2_entries_perms_3_x; // @[Reg.scala 16:16]
  reg  l3_ramDatas_2_entries_perms_3_w; // @[Reg.scala 16:16]
  reg  l3_ramDatas_2_entries_perms_3_r; // @[Reg.scala 16:16]
  reg  l3_ramDatas_2_entries_perms_4_d; // @[Reg.scala 16:16]
  reg  l3_ramDatas_2_entries_perms_4_a; // @[Reg.scala 16:16]
  reg  l3_ramDatas_2_entries_perms_4_g; // @[Reg.scala 16:16]
  reg  l3_ramDatas_2_entries_perms_4_u; // @[Reg.scala 16:16]
  reg  l3_ramDatas_2_entries_perms_4_x; // @[Reg.scala 16:16]
  reg  l3_ramDatas_2_entries_perms_4_w; // @[Reg.scala 16:16]
  reg  l3_ramDatas_2_entries_perms_4_r; // @[Reg.scala 16:16]
  reg  l3_ramDatas_2_entries_perms_5_d; // @[Reg.scala 16:16]
  reg  l3_ramDatas_2_entries_perms_5_a; // @[Reg.scala 16:16]
  reg  l3_ramDatas_2_entries_perms_5_g; // @[Reg.scala 16:16]
  reg  l3_ramDatas_2_entries_perms_5_u; // @[Reg.scala 16:16]
  reg  l3_ramDatas_2_entries_perms_5_x; // @[Reg.scala 16:16]
  reg  l3_ramDatas_2_entries_perms_5_w; // @[Reg.scala 16:16]
  reg  l3_ramDatas_2_entries_perms_5_r; // @[Reg.scala 16:16]
  reg  l3_ramDatas_2_entries_perms_6_d; // @[Reg.scala 16:16]
  reg  l3_ramDatas_2_entries_perms_6_a; // @[Reg.scala 16:16]
  reg  l3_ramDatas_2_entries_perms_6_g; // @[Reg.scala 16:16]
  reg  l3_ramDatas_2_entries_perms_6_u; // @[Reg.scala 16:16]
  reg  l3_ramDatas_2_entries_perms_6_x; // @[Reg.scala 16:16]
  reg  l3_ramDatas_2_entries_perms_6_w; // @[Reg.scala 16:16]
  reg  l3_ramDatas_2_entries_perms_6_r; // @[Reg.scala 16:16]
  reg  l3_ramDatas_2_entries_perms_7_d; // @[Reg.scala 16:16]
  reg  l3_ramDatas_2_entries_perms_7_a; // @[Reg.scala 16:16]
  reg  l3_ramDatas_2_entries_perms_7_g; // @[Reg.scala 16:16]
  reg  l3_ramDatas_2_entries_perms_7_u; // @[Reg.scala 16:16]
  reg  l3_ramDatas_2_entries_perms_7_x; // @[Reg.scala 16:16]
  reg  l3_ramDatas_2_entries_perms_7_w; // @[Reg.scala 16:16]
  reg  l3_ramDatas_2_entries_perms_7_r; // @[Reg.scala 16:16]
  reg  l3_ramDatas_2_entries_prefetch; // @[Reg.scala 16:16]
  reg [38:0] l3_ramDatas_2_ecc; // @[Reg.scala 16:16]
  reg [21:0] l3_ramDatas_3_entries_tag; // @[Reg.scala 16:16]
  reg [15:0] l3_ramDatas_3_entries_asid; // @[Reg.scala 16:16]
  reg [23:0] l3_ramDatas_3_entries_ppns_0; // @[Reg.scala 16:16]
  reg [23:0] l3_ramDatas_3_entries_ppns_1; // @[Reg.scala 16:16]
  reg [23:0] l3_ramDatas_3_entries_ppns_2; // @[Reg.scala 16:16]
  reg [23:0] l3_ramDatas_3_entries_ppns_3; // @[Reg.scala 16:16]
  reg [23:0] l3_ramDatas_3_entries_ppns_4; // @[Reg.scala 16:16]
  reg [23:0] l3_ramDatas_3_entries_ppns_5; // @[Reg.scala 16:16]
  reg [23:0] l3_ramDatas_3_entries_ppns_6; // @[Reg.scala 16:16]
  reg [23:0] l3_ramDatas_3_entries_ppns_7; // @[Reg.scala 16:16]
  reg  l3_ramDatas_3_entries_vs_0; // @[Reg.scala 16:16]
  reg  l3_ramDatas_3_entries_vs_1; // @[Reg.scala 16:16]
  reg  l3_ramDatas_3_entries_vs_2; // @[Reg.scala 16:16]
  reg  l3_ramDatas_3_entries_vs_3; // @[Reg.scala 16:16]
  reg  l3_ramDatas_3_entries_vs_4; // @[Reg.scala 16:16]
  reg  l3_ramDatas_3_entries_vs_5; // @[Reg.scala 16:16]
  reg  l3_ramDatas_3_entries_vs_6; // @[Reg.scala 16:16]
  reg  l3_ramDatas_3_entries_vs_7; // @[Reg.scala 16:16]
  reg  l3_ramDatas_3_entries_perms_0_d; // @[Reg.scala 16:16]
  reg  l3_ramDatas_3_entries_perms_0_a; // @[Reg.scala 16:16]
  reg  l3_ramDatas_3_entries_perms_0_g; // @[Reg.scala 16:16]
  reg  l3_ramDatas_3_entries_perms_0_u; // @[Reg.scala 16:16]
  reg  l3_ramDatas_3_entries_perms_0_x; // @[Reg.scala 16:16]
  reg  l3_ramDatas_3_entries_perms_0_w; // @[Reg.scala 16:16]
  reg  l3_ramDatas_3_entries_perms_0_r; // @[Reg.scala 16:16]
  reg  l3_ramDatas_3_entries_perms_1_d; // @[Reg.scala 16:16]
  reg  l3_ramDatas_3_entries_perms_1_a; // @[Reg.scala 16:16]
  reg  l3_ramDatas_3_entries_perms_1_g; // @[Reg.scala 16:16]
  reg  l3_ramDatas_3_entries_perms_1_u; // @[Reg.scala 16:16]
  reg  l3_ramDatas_3_entries_perms_1_x; // @[Reg.scala 16:16]
  reg  l3_ramDatas_3_entries_perms_1_w; // @[Reg.scala 16:16]
  reg  l3_ramDatas_3_entries_perms_1_r; // @[Reg.scala 16:16]
  reg  l3_ramDatas_3_entries_perms_2_d; // @[Reg.scala 16:16]
  reg  l3_ramDatas_3_entries_perms_2_a; // @[Reg.scala 16:16]
  reg  l3_ramDatas_3_entries_perms_2_g; // @[Reg.scala 16:16]
  reg  l3_ramDatas_3_entries_perms_2_u; // @[Reg.scala 16:16]
  reg  l3_ramDatas_3_entries_perms_2_x; // @[Reg.scala 16:16]
  reg  l3_ramDatas_3_entries_perms_2_w; // @[Reg.scala 16:16]
  reg  l3_ramDatas_3_entries_perms_2_r; // @[Reg.scala 16:16]
  reg  l3_ramDatas_3_entries_perms_3_d; // @[Reg.scala 16:16]
  reg  l3_ramDatas_3_entries_perms_3_a; // @[Reg.scala 16:16]
  reg  l3_ramDatas_3_entries_perms_3_g; // @[Reg.scala 16:16]
  reg  l3_ramDatas_3_entries_perms_3_u; // @[Reg.scala 16:16]
  reg  l3_ramDatas_3_entries_perms_3_x; // @[Reg.scala 16:16]
  reg  l3_ramDatas_3_entries_perms_3_w; // @[Reg.scala 16:16]
  reg  l3_ramDatas_3_entries_perms_3_r; // @[Reg.scala 16:16]
  reg  l3_ramDatas_3_entries_perms_4_d; // @[Reg.scala 16:16]
  reg  l3_ramDatas_3_entries_perms_4_a; // @[Reg.scala 16:16]
  reg  l3_ramDatas_3_entries_perms_4_g; // @[Reg.scala 16:16]
  reg  l3_ramDatas_3_entries_perms_4_u; // @[Reg.scala 16:16]
  reg  l3_ramDatas_3_entries_perms_4_x; // @[Reg.scala 16:16]
  reg  l3_ramDatas_3_entries_perms_4_w; // @[Reg.scala 16:16]
  reg  l3_ramDatas_3_entries_perms_4_r; // @[Reg.scala 16:16]
  reg  l3_ramDatas_3_entries_perms_5_d; // @[Reg.scala 16:16]
  reg  l3_ramDatas_3_entries_perms_5_a; // @[Reg.scala 16:16]
  reg  l3_ramDatas_3_entries_perms_5_g; // @[Reg.scala 16:16]
  reg  l3_ramDatas_3_entries_perms_5_u; // @[Reg.scala 16:16]
  reg  l3_ramDatas_3_entries_perms_5_x; // @[Reg.scala 16:16]
  reg  l3_ramDatas_3_entries_perms_5_w; // @[Reg.scala 16:16]
  reg  l3_ramDatas_3_entries_perms_5_r; // @[Reg.scala 16:16]
  reg  l3_ramDatas_3_entries_perms_6_d; // @[Reg.scala 16:16]
  reg  l3_ramDatas_3_entries_perms_6_a; // @[Reg.scala 16:16]
  reg  l3_ramDatas_3_entries_perms_6_g; // @[Reg.scala 16:16]
  reg  l3_ramDatas_3_entries_perms_6_u; // @[Reg.scala 16:16]
  reg  l3_ramDatas_3_entries_perms_6_x; // @[Reg.scala 16:16]
  reg  l3_ramDatas_3_entries_perms_6_w; // @[Reg.scala 16:16]
  reg  l3_ramDatas_3_entries_perms_6_r; // @[Reg.scala 16:16]
  reg  l3_ramDatas_3_entries_perms_7_d; // @[Reg.scala 16:16]
  reg  l3_ramDatas_3_entries_perms_7_a; // @[Reg.scala 16:16]
  reg  l3_ramDatas_3_entries_perms_7_g; // @[Reg.scala 16:16]
  reg  l3_ramDatas_3_entries_perms_7_u; // @[Reg.scala 16:16]
  reg  l3_ramDatas_3_entries_perms_7_x; // @[Reg.scala 16:16]
  reg  l3_ramDatas_3_entries_perms_7_w; // @[Reg.scala 16:16]
  reg  l3_ramDatas_3_entries_perms_7_r; // @[Reg.scala 16:16]
  reg  l3_ramDatas_3_entries_prefetch; // @[Reg.scala 16:16]
  reg [38:0] l3_ramDatas_3_ecc; // @[Reg.scala 16:16]
  reg [21:0] l3_ramDatas_4_entries_tag; // @[Reg.scala 16:16]
  reg [15:0] l3_ramDatas_4_entries_asid; // @[Reg.scala 16:16]
  reg [23:0] l3_ramDatas_4_entries_ppns_0; // @[Reg.scala 16:16]
  reg [23:0] l3_ramDatas_4_entries_ppns_1; // @[Reg.scala 16:16]
  reg [23:0] l3_ramDatas_4_entries_ppns_2; // @[Reg.scala 16:16]
  reg [23:0] l3_ramDatas_4_entries_ppns_3; // @[Reg.scala 16:16]
  reg [23:0] l3_ramDatas_4_entries_ppns_4; // @[Reg.scala 16:16]
  reg [23:0] l3_ramDatas_4_entries_ppns_5; // @[Reg.scala 16:16]
  reg [23:0] l3_ramDatas_4_entries_ppns_6; // @[Reg.scala 16:16]
  reg [23:0] l3_ramDatas_4_entries_ppns_7; // @[Reg.scala 16:16]
  reg  l3_ramDatas_4_entries_vs_0; // @[Reg.scala 16:16]
  reg  l3_ramDatas_4_entries_vs_1; // @[Reg.scala 16:16]
  reg  l3_ramDatas_4_entries_vs_2; // @[Reg.scala 16:16]
  reg  l3_ramDatas_4_entries_vs_3; // @[Reg.scala 16:16]
  reg  l3_ramDatas_4_entries_vs_4; // @[Reg.scala 16:16]
  reg  l3_ramDatas_4_entries_vs_5; // @[Reg.scala 16:16]
  reg  l3_ramDatas_4_entries_vs_6; // @[Reg.scala 16:16]
  reg  l3_ramDatas_4_entries_vs_7; // @[Reg.scala 16:16]
  reg  l3_ramDatas_4_entries_perms_0_d; // @[Reg.scala 16:16]
  reg  l3_ramDatas_4_entries_perms_0_a; // @[Reg.scala 16:16]
  reg  l3_ramDatas_4_entries_perms_0_g; // @[Reg.scala 16:16]
  reg  l3_ramDatas_4_entries_perms_0_u; // @[Reg.scala 16:16]
  reg  l3_ramDatas_4_entries_perms_0_x; // @[Reg.scala 16:16]
  reg  l3_ramDatas_4_entries_perms_0_w; // @[Reg.scala 16:16]
  reg  l3_ramDatas_4_entries_perms_0_r; // @[Reg.scala 16:16]
  reg  l3_ramDatas_4_entries_perms_1_d; // @[Reg.scala 16:16]
  reg  l3_ramDatas_4_entries_perms_1_a; // @[Reg.scala 16:16]
  reg  l3_ramDatas_4_entries_perms_1_g; // @[Reg.scala 16:16]
  reg  l3_ramDatas_4_entries_perms_1_u; // @[Reg.scala 16:16]
  reg  l3_ramDatas_4_entries_perms_1_x; // @[Reg.scala 16:16]
  reg  l3_ramDatas_4_entries_perms_1_w; // @[Reg.scala 16:16]
  reg  l3_ramDatas_4_entries_perms_1_r; // @[Reg.scala 16:16]
  reg  l3_ramDatas_4_entries_perms_2_d; // @[Reg.scala 16:16]
  reg  l3_ramDatas_4_entries_perms_2_a; // @[Reg.scala 16:16]
  reg  l3_ramDatas_4_entries_perms_2_g; // @[Reg.scala 16:16]
  reg  l3_ramDatas_4_entries_perms_2_u; // @[Reg.scala 16:16]
  reg  l3_ramDatas_4_entries_perms_2_x; // @[Reg.scala 16:16]
  reg  l3_ramDatas_4_entries_perms_2_w; // @[Reg.scala 16:16]
  reg  l3_ramDatas_4_entries_perms_2_r; // @[Reg.scala 16:16]
  reg  l3_ramDatas_4_entries_perms_3_d; // @[Reg.scala 16:16]
  reg  l3_ramDatas_4_entries_perms_3_a; // @[Reg.scala 16:16]
  reg  l3_ramDatas_4_entries_perms_3_g; // @[Reg.scala 16:16]
  reg  l3_ramDatas_4_entries_perms_3_u; // @[Reg.scala 16:16]
  reg  l3_ramDatas_4_entries_perms_3_x; // @[Reg.scala 16:16]
  reg  l3_ramDatas_4_entries_perms_3_w; // @[Reg.scala 16:16]
  reg  l3_ramDatas_4_entries_perms_3_r; // @[Reg.scala 16:16]
  reg  l3_ramDatas_4_entries_perms_4_d; // @[Reg.scala 16:16]
  reg  l3_ramDatas_4_entries_perms_4_a; // @[Reg.scala 16:16]
  reg  l3_ramDatas_4_entries_perms_4_g; // @[Reg.scala 16:16]
  reg  l3_ramDatas_4_entries_perms_4_u; // @[Reg.scala 16:16]
  reg  l3_ramDatas_4_entries_perms_4_x; // @[Reg.scala 16:16]
  reg  l3_ramDatas_4_entries_perms_4_w; // @[Reg.scala 16:16]
  reg  l3_ramDatas_4_entries_perms_4_r; // @[Reg.scala 16:16]
  reg  l3_ramDatas_4_entries_perms_5_d; // @[Reg.scala 16:16]
  reg  l3_ramDatas_4_entries_perms_5_a; // @[Reg.scala 16:16]
  reg  l3_ramDatas_4_entries_perms_5_g; // @[Reg.scala 16:16]
  reg  l3_ramDatas_4_entries_perms_5_u; // @[Reg.scala 16:16]
  reg  l3_ramDatas_4_entries_perms_5_x; // @[Reg.scala 16:16]
  reg  l3_ramDatas_4_entries_perms_5_w; // @[Reg.scala 16:16]
  reg  l3_ramDatas_4_entries_perms_5_r; // @[Reg.scala 16:16]
  reg  l3_ramDatas_4_entries_perms_6_d; // @[Reg.scala 16:16]
  reg  l3_ramDatas_4_entries_perms_6_a; // @[Reg.scala 16:16]
  reg  l3_ramDatas_4_entries_perms_6_g; // @[Reg.scala 16:16]
  reg  l3_ramDatas_4_entries_perms_6_u; // @[Reg.scala 16:16]
  reg  l3_ramDatas_4_entries_perms_6_x; // @[Reg.scala 16:16]
  reg  l3_ramDatas_4_entries_perms_6_w; // @[Reg.scala 16:16]
  reg  l3_ramDatas_4_entries_perms_6_r; // @[Reg.scala 16:16]
  reg  l3_ramDatas_4_entries_perms_7_d; // @[Reg.scala 16:16]
  reg  l3_ramDatas_4_entries_perms_7_a; // @[Reg.scala 16:16]
  reg  l3_ramDatas_4_entries_perms_7_g; // @[Reg.scala 16:16]
  reg  l3_ramDatas_4_entries_perms_7_u; // @[Reg.scala 16:16]
  reg  l3_ramDatas_4_entries_perms_7_x; // @[Reg.scala 16:16]
  reg  l3_ramDatas_4_entries_perms_7_w; // @[Reg.scala 16:16]
  reg  l3_ramDatas_4_entries_perms_7_r; // @[Reg.scala 16:16]
  reg  l3_ramDatas_4_entries_prefetch; // @[Reg.scala 16:16]
  reg [38:0] l3_ramDatas_4_ecc; // @[Reg.scala 16:16]
  reg [21:0] l3_ramDatas_5_entries_tag; // @[Reg.scala 16:16]
  reg [15:0] l3_ramDatas_5_entries_asid; // @[Reg.scala 16:16]
  reg [23:0] l3_ramDatas_5_entries_ppns_0; // @[Reg.scala 16:16]
  reg [23:0] l3_ramDatas_5_entries_ppns_1; // @[Reg.scala 16:16]
  reg [23:0] l3_ramDatas_5_entries_ppns_2; // @[Reg.scala 16:16]
  reg [23:0] l3_ramDatas_5_entries_ppns_3; // @[Reg.scala 16:16]
  reg [23:0] l3_ramDatas_5_entries_ppns_4; // @[Reg.scala 16:16]
  reg [23:0] l3_ramDatas_5_entries_ppns_5; // @[Reg.scala 16:16]
  reg [23:0] l3_ramDatas_5_entries_ppns_6; // @[Reg.scala 16:16]
  reg [23:0] l3_ramDatas_5_entries_ppns_7; // @[Reg.scala 16:16]
  reg  l3_ramDatas_5_entries_vs_0; // @[Reg.scala 16:16]
  reg  l3_ramDatas_5_entries_vs_1; // @[Reg.scala 16:16]
  reg  l3_ramDatas_5_entries_vs_2; // @[Reg.scala 16:16]
  reg  l3_ramDatas_5_entries_vs_3; // @[Reg.scala 16:16]
  reg  l3_ramDatas_5_entries_vs_4; // @[Reg.scala 16:16]
  reg  l3_ramDatas_5_entries_vs_5; // @[Reg.scala 16:16]
  reg  l3_ramDatas_5_entries_vs_6; // @[Reg.scala 16:16]
  reg  l3_ramDatas_5_entries_vs_7; // @[Reg.scala 16:16]
  reg  l3_ramDatas_5_entries_perms_0_d; // @[Reg.scala 16:16]
  reg  l3_ramDatas_5_entries_perms_0_a; // @[Reg.scala 16:16]
  reg  l3_ramDatas_5_entries_perms_0_g; // @[Reg.scala 16:16]
  reg  l3_ramDatas_5_entries_perms_0_u; // @[Reg.scala 16:16]
  reg  l3_ramDatas_5_entries_perms_0_x; // @[Reg.scala 16:16]
  reg  l3_ramDatas_5_entries_perms_0_w; // @[Reg.scala 16:16]
  reg  l3_ramDatas_5_entries_perms_0_r; // @[Reg.scala 16:16]
  reg  l3_ramDatas_5_entries_perms_1_d; // @[Reg.scala 16:16]
  reg  l3_ramDatas_5_entries_perms_1_a; // @[Reg.scala 16:16]
  reg  l3_ramDatas_5_entries_perms_1_g; // @[Reg.scala 16:16]
  reg  l3_ramDatas_5_entries_perms_1_u; // @[Reg.scala 16:16]
  reg  l3_ramDatas_5_entries_perms_1_x; // @[Reg.scala 16:16]
  reg  l3_ramDatas_5_entries_perms_1_w; // @[Reg.scala 16:16]
  reg  l3_ramDatas_5_entries_perms_1_r; // @[Reg.scala 16:16]
  reg  l3_ramDatas_5_entries_perms_2_d; // @[Reg.scala 16:16]
  reg  l3_ramDatas_5_entries_perms_2_a; // @[Reg.scala 16:16]
  reg  l3_ramDatas_5_entries_perms_2_g; // @[Reg.scala 16:16]
  reg  l3_ramDatas_5_entries_perms_2_u; // @[Reg.scala 16:16]
  reg  l3_ramDatas_5_entries_perms_2_x; // @[Reg.scala 16:16]
  reg  l3_ramDatas_5_entries_perms_2_w; // @[Reg.scala 16:16]
  reg  l3_ramDatas_5_entries_perms_2_r; // @[Reg.scala 16:16]
  reg  l3_ramDatas_5_entries_perms_3_d; // @[Reg.scala 16:16]
  reg  l3_ramDatas_5_entries_perms_3_a; // @[Reg.scala 16:16]
  reg  l3_ramDatas_5_entries_perms_3_g; // @[Reg.scala 16:16]
  reg  l3_ramDatas_5_entries_perms_3_u; // @[Reg.scala 16:16]
  reg  l3_ramDatas_5_entries_perms_3_x; // @[Reg.scala 16:16]
  reg  l3_ramDatas_5_entries_perms_3_w; // @[Reg.scala 16:16]
  reg  l3_ramDatas_5_entries_perms_3_r; // @[Reg.scala 16:16]
  reg  l3_ramDatas_5_entries_perms_4_d; // @[Reg.scala 16:16]
  reg  l3_ramDatas_5_entries_perms_4_a; // @[Reg.scala 16:16]
  reg  l3_ramDatas_5_entries_perms_4_g; // @[Reg.scala 16:16]
  reg  l3_ramDatas_5_entries_perms_4_u; // @[Reg.scala 16:16]
  reg  l3_ramDatas_5_entries_perms_4_x; // @[Reg.scala 16:16]
  reg  l3_ramDatas_5_entries_perms_4_w; // @[Reg.scala 16:16]
  reg  l3_ramDatas_5_entries_perms_4_r; // @[Reg.scala 16:16]
  reg  l3_ramDatas_5_entries_perms_5_d; // @[Reg.scala 16:16]
  reg  l3_ramDatas_5_entries_perms_5_a; // @[Reg.scala 16:16]
  reg  l3_ramDatas_5_entries_perms_5_g; // @[Reg.scala 16:16]
  reg  l3_ramDatas_5_entries_perms_5_u; // @[Reg.scala 16:16]
  reg  l3_ramDatas_5_entries_perms_5_x; // @[Reg.scala 16:16]
  reg  l3_ramDatas_5_entries_perms_5_w; // @[Reg.scala 16:16]
  reg  l3_ramDatas_5_entries_perms_5_r; // @[Reg.scala 16:16]
  reg  l3_ramDatas_5_entries_perms_6_d; // @[Reg.scala 16:16]
  reg  l3_ramDatas_5_entries_perms_6_a; // @[Reg.scala 16:16]
  reg  l3_ramDatas_5_entries_perms_6_g; // @[Reg.scala 16:16]
  reg  l3_ramDatas_5_entries_perms_6_u; // @[Reg.scala 16:16]
  reg  l3_ramDatas_5_entries_perms_6_x; // @[Reg.scala 16:16]
  reg  l3_ramDatas_5_entries_perms_6_w; // @[Reg.scala 16:16]
  reg  l3_ramDatas_5_entries_perms_6_r; // @[Reg.scala 16:16]
  reg  l3_ramDatas_5_entries_perms_7_d; // @[Reg.scala 16:16]
  reg  l3_ramDatas_5_entries_perms_7_a; // @[Reg.scala 16:16]
  reg  l3_ramDatas_5_entries_perms_7_g; // @[Reg.scala 16:16]
  reg  l3_ramDatas_5_entries_perms_7_u; // @[Reg.scala 16:16]
  reg  l3_ramDatas_5_entries_perms_7_x; // @[Reg.scala 16:16]
  reg  l3_ramDatas_5_entries_perms_7_w; // @[Reg.scala 16:16]
  reg  l3_ramDatas_5_entries_perms_7_r; // @[Reg.scala 16:16]
  reg  l3_ramDatas_5_entries_prefetch; // @[Reg.scala 16:16]
  reg [38:0] l3_ramDatas_5_ecc; // @[Reg.scala 16:16]
  reg [21:0] l3_ramDatas_6_entries_tag; // @[Reg.scala 16:16]
  reg [15:0] l3_ramDatas_6_entries_asid; // @[Reg.scala 16:16]
  reg [23:0] l3_ramDatas_6_entries_ppns_0; // @[Reg.scala 16:16]
  reg [23:0] l3_ramDatas_6_entries_ppns_1; // @[Reg.scala 16:16]
  reg [23:0] l3_ramDatas_6_entries_ppns_2; // @[Reg.scala 16:16]
  reg [23:0] l3_ramDatas_6_entries_ppns_3; // @[Reg.scala 16:16]
  reg [23:0] l3_ramDatas_6_entries_ppns_4; // @[Reg.scala 16:16]
  reg [23:0] l3_ramDatas_6_entries_ppns_5; // @[Reg.scala 16:16]
  reg [23:0] l3_ramDatas_6_entries_ppns_6; // @[Reg.scala 16:16]
  reg [23:0] l3_ramDatas_6_entries_ppns_7; // @[Reg.scala 16:16]
  reg  l3_ramDatas_6_entries_vs_0; // @[Reg.scala 16:16]
  reg  l3_ramDatas_6_entries_vs_1; // @[Reg.scala 16:16]
  reg  l3_ramDatas_6_entries_vs_2; // @[Reg.scala 16:16]
  reg  l3_ramDatas_6_entries_vs_3; // @[Reg.scala 16:16]
  reg  l3_ramDatas_6_entries_vs_4; // @[Reg.scala 16:16]
  reg  l3_ramDatas_6_entries_vs_5; // @[Reg.scala 16:16]
  reg  l3_ramDatas_6_entries_vs_6; // @[Reg.scala 16:16]
  reg  l3_ramDatas_6_entries_vs_7; // @[Reg.scala 16:16]
  reg  l3_ramDatas_6_entries_perms_0_d; // @[Reg.scala 16:16]
  reg  l3_ramDatas_6_entries_perms_0_a; // @[Reg.scala 16:16]
  reg  l3_ramDatas_6_entries_perms_0_g; // @[Reg.scala 16:16]
  reg  l3_ramDatas_6_entries_perms_0_u; // @[Reg.scala 16:16]
  reg  l3_ramDatas_6_entries_perms_0_x; // @[Reg.scala 16:16]
  reg  l3_ramDatas_6_entries_perms_0_w; // @[Reg.scala 16:16]
  reg  l3_ramDatas_6_entries_perms_0_r; // @[Reg.scala 16:16]
  reg  l3_ramDatas_6_entries_perms_1_d; // @[Reg.scala 16:16]
  reg  l3_ramDatas_6_entries_perms_1_a; // @[Reg.scala 16:16]
  reg  l3_ramDatas_6_entries_perms_1_g; // @[Reg.scala 16:16]
  reg  l3_ramDatas_6_entries_perms_1_u; // @[Reg.scala 16:16]
  reg  l3_ramDatas_6_entries_perms_1_x; // @[Reg.scala 16:16]
  reg  l3_ramDatas_6_entries_perms_1_w; // @[Reg.scala 16:16]
  reg  l3_ramDatas_6_entries_perms_1_r; // @[Reg.scala 16:16]
  reg  l3_ramDatas_6_entries_perms_2_d; // @[Reg.scala 16:16]
  reg  l3_ramDatas_6_entries_perms_2_a; // @[Reg.scala 16:16]
  reg  l3_ramDatas_6_entries_perms_2_g; // @[Reg.scala 16:16]
  reg  l3_ramDatas_6_entries_perms_2_u; // @[Reg.scala 16:16]
  reg  l3_ramDatas_6_entries_perms_2_x; // @[Reg.scala 16:16]
  reg  l3_ramDatas_6_entries_perms_2_w; // @[Reg.scala 16:16]
  reg  l3_ramDatas_6_entries_perms_2_r; // @[Reg.scala 16:16]
  reg  l3_ramDatas_6_entries_perms_3_d; // @[Reg.scala 16:16]
  reg  l3_ramDatas_6_entries_perms_3_a; // @[Reg.scala 16:16]
  reg  l3_ramDatas_6_entries_perms_3_g; // @[Reg.scala 16:16]
  reg  l3_ramDatas_6_entries_perms_3_u; // @[Reg.scala 16:16]
  reg  l3_ramDatas_6_entries_perms_3_x; // @[Reg.scala 16:16]
  reg  l3_ramDatas_6_entries_perms_3_w; // @[Reg.scala 16:16]
  reg  l3_ramDatas_6_entries_perms_3_r; // @[Reg.scala 16:16]
  reg  l3_ramDatas_6_entries_perms_4_d; // @[Reg.scala 16:16]
  reg  l3_ramDatas_6_entries_perms_4_a; // @[Reg.scala 16:16]
  reg  l3_ramDatas_6_entries_perms_4_g; // @[Reg.scala 16:16]
  reg  l3_ramDatas_6_entries_perms_4_u; // @[Reg.scala 16:16]
  reg  l3_ramDatas_6_entries_perms_4_x; // @[Reg.scala 16:16]
  reg  l3_ramDatas_6_entries_perms_4_w; // @[Reg.scala 16:16]
  reg  l3_ramDatas_6_entries_perms_4_r; // @[Reg.scala 16:16]
  reg  l3_ramDatas_6_entries_perms_5_d; // @[Reg.scala 16:16]
  reg  l3_ramDatas_6_entries_perms_5_a; // @[Reg.scala 16:16]
  reg  l3_ramDatas_6_entries_perms_5_g; // @[Reg.scala 16:16]
  reg  l3_ramDatas_6_entries_perms_5_u; // @[Reg.scala 16:16]
  reg  l3_ramDatas_6_entries_perms_5_x; // @[Reg.scala 16:16]
  reg  l3_ramDatas_6_entries_perms_5_w; // @[Reg.scala 16:16]
  reg  l3_ramDatas_6_entries_perms_5_r; // @[Reg.scala 16:16]
  reg  l3_ramDatas_6_entries_perms_6_d; // @[Reg.scala 16:16]
  reg  l3_ramDatas_6_entries_perms_6_a; // @[Reg.scala 16:16]
  reg  l3_ramDatas_6_entries_perms_6_g; // @[Reg.scala 16:16]
  reg  l3_ramDatas_6_entries_perms_6_u; // @[Reg.scala 16:16]
  reg  l3_ramDatas_6_entries_perms_6_x; // @[Reg.scala 16:16]
  reg  l3_ramDatas_6_entries_perms_6_w; // @[Reg.scala 16:16]
  reg  l3_ramDatas_6_entries_perms_6_r; // @[Reg.scala 16:16]
  reg  l3_ramDatas_6_entries_perms_7_d; // @[Reg.scala 16:16]
  reg  l3_ramDatas_6_entries_perms_7_a; // @[Reg.scala 16:16]
  reg  l3_ramDatas_6_entries_perms_7_g; // @[Reg.scala 16:16]
  reg  l3_ramDatas_6_entries_perms_7_u; // @[Reg.scala 16:16]
  reg  l3_ramDatas_6_entries_perms_7_x; // @[Reg.scala 16:16]
  reg  l3_ramDatas_6_entries_perms_7_w; // @[Reg.scala 16:16]
  reg  l3_ramDatas_6_entries_perms_7_r; // @[Reg.scala 16:16]
  reg  l3_ramDatas_6_entries_prefetch; // @[Reg.scala 16:16]
  reg [38:0] l3_ramDatas_6_ecc; // @[Reg.scala 16:16]
  reg [21:0] l3_ramDatas_7_entries_tag; // @[Reg.scala 16:16]
  reg [15:0] l3_ramDatas_7_entries_asid; // @[Reg.scala 16:16]
  reg [23:0] l3_ramDatas_7_entries_ppns_0; // @[Reg.scala 16:16]
  reg [23:0] l3_ramDatas_7_entries_ppns_1; // @[Reg.scala 16:16]
  reg [23:0] l3_ramDatas_7_entries_ppns_2; // @[Reg.scala 16:16]
  reg [23:0] l3_ramDatas_7_entries_ppns_3; // @[Reg.scala 16:16]
  reg [23:0] l3_ramDatas_7_entries_ppns_4; // @[Reg.scala 16:16]
  reg [23:0] l3_ramDatas_7_entries_ppns_5; // @[Reg.scala 16:16]
  reg [23:0] l3_ramDatas_7_entries_ppns_6; // @[Reg.scala 16:16]
  reg [23:0] l3_ramDatas_7_entries_ppns_7; // @[Reg.scala 16:16]
  reg  l3_ramDatas_7_entries_vs_0; // @[Reg.scala 16:16]
  reg  l3_ramDatas_7_entries_vs_1; // @[Reg.scala 16:16]
  reg  l3_ramDatas_7_entries_vs_2; // @[Reg.scala 16:16]
  reg  l3_ramDatas_7_entries_vs_3; // @[Reg.scala 16:16]
  reg  l3_ramDatas_7_entries_vs_4; // @[Reg.scala 16:16]
  reg  l3_ramDatas_7_entries_vs_5; // @[Reg.scala 16:16]
  reg  l3_ramDatas_7_entries_vs_6; // @[Reg.scala 16:16]
  reg  l3_ramDatas_7_entries_vs_7; // @[Reg.scala 16:16]
  reg  l3_ramDatas_7_entries_perms_0_d; // @[Reg.scala 16:16]
  reg  l3_ramDatas_7_entries_perms_0_a; // @[Reg.scala 16:16]
  reg  l3_ramDatas_7_entries_perms_0_g; // @[Reg.scala 16:16]
  reg  l3_ramDatas_7_entries_perms_0_u; // @[Reg.scala 16:16]
  reg  l3_ramDatas_7_entries_perms_0_x; // @[Reg.scala 16:16]
  reg  l3_ramDatas_7_entries_perms_0_w; // @[Reg.scala 16:16]
  reg  l3_ramDatas_7_entries_perms_0_r; // @[Reg.scala 16:16]
  reg  l3_ramDatas_7_entries_perms_1_d; // @[Reg.scala 16:16]
  reg  l3_ramDatas_7_entries_perms_1_a; // @[Reg.scala 16:16]
  reg  l3_ramDatas_7_entries_perms_1_g; // @[Reg.scala 16:16]
  reg  l3_ramDatas_7_entries_perms_1_u; // @[Reg.scala 16:16]
  reg  l3_ramDatas_7_entries_perms_1_x; // @[Reg.scala 16:16]
  reg  l3_ramDatas_7_entries_perms_1_w; // @[Reg.scala 16:16]
  reg  l3_ramDatas_7_entries_perms_1_r; // @[Reg.scala 16:16]
  reg  l3_ramDatas_7_entries_perms_2_d; // @[Reg.scala 16:16]
  reg  l3_ramDatas_7_entries_perms_2_a; // @[Reg.scala 16:16]
  reg  l3_ramDatas_7_entries_perms_2_g; // @[Reg.scala 16:16]
  reg  l3_ramDatas_7_entries_perms_2_u; // @[Reg.scala 16:16]
  reg  l3_ramDatas_7_entries_perms_2_x; // @[Reg.scala 16:16]
  reg  l3_ramDatas_7_entries_perms_2_w; // @[Reg.scala 16:16]
  reg  l3_ramDatas_7_entries_perms_2_r; // @[Reg.scala 16:16]
  reg  l3_ramDatas_7_entries_perms_3_d; // @[Reg.scala 16:16]
  reg  l3_ramDatas_7_entries_perms_3_a; // @[Reg.scala 16:16]
  reg  l3_ramDatas_7_entries_perms_3_g; // @[Reg.scala 16:16]
  reg  l3_ramDatas_7_entries_perms_3_u; // @[Reg.scala 16:16]
  reg  l3_ramDatas_7_entries_perms_3_x; // @[Reg.scala 16:16]
  reg  l3_ramDatas_7_entries_perms_3_w; // @[Reg.scala 16:16]
  reg  l3_ramDatas_7_entries_perms_3_r; // @[Reg.scala 16:16]
  reg  l3_ramDatas_7_entries_perms_4_d; // @[Reg.scala 16:16]
  reg  l3_ramDatas_7_entries_perms_4_a; // @[Reg.scala 16:16]
  reg  l3_ramDatas_7_entries_perms_4_g; // @[Reg.scala 16:16]
  reg  l3_ramDatas_7_entries_perms_4_u; // @[Reg.scala 16:16]
  reg  l3_ramDatas_7_entries_perms_4_x; // @[Reg.scala 16:16]
  reg  l3_ramDatas_7_entries_perms_4_w; // @[Reg.scala 16:16]
  reg  l3_ramDatas_7_entries_perms_4_r; // @[Reg.scala 16:16]
  reg  l3_ramDatas_7_entries_perms_5_d; // @[Reg.scala 16:16]
  reg  l3_ramDatas_7_entries_perms_5_a; // @[Reg.scala 16:16]
  reg  l3_ramDatas_7_entries_perms_5_g; // @[Reg.scala 16:16]
  reg  l3_ramDatas_7_entries_perms_5_u; // @[Reg.scala 16:16]
  reg  l3_ramDatas_7_entries_perms_5_x; // @[Reg.scala 16:16]
  reg  l3_ramDatas_7_entries_perms_5_w; // @[Reg.scala 16:16]
  reg  l3_ramDatas_7_entries_perms_5_r; // @[Reg.scala 16:16]
  reg  l3_ramDatas_7_entries_perms_6_d; // @[Reg.scala 16:16]
  reg  l3_ramDatas_7_entries_perms_6_a; // @[Reg.scala 16:16]
  reg  l3_ramDatas_7_entries_perms_6_g; // @[Reg.scala 16:16]
  reg  l3_ramDatas_7_entries_perms_6_u; // @[Reg.scala 16:16]
  reg  l3_ramDatas_7_entries_perms_6_x; // @[Reg.scala 16:16]
  reg  l3_ramDatas_7_entries_perms_6_w; // @[Reg.scala 16:16]
  reg  l3_ramDatas_7_entries_perms_6_r; // @[Reg.scala 16:16]
  reg  l3_ramDatas_7_entries_perms_7_d; // @[Reg.scala 16:16]
  reg  l3_ramDatas_7_entries_perms_7_a; // @[Reg.scala 16:16]
  reg  l3_ramDatas_7_entries_perms_7_g; // @[Reg.scala 16:16]
  reg  l3_ramDatas_7_entries_perms_7_u; // @[Reg.scala 16:16]
  reg  l3_ramDatas_7_entries_perms_7_x; // @[Reg.scala 16:16]
  reg  l3_ramDatas_7_entries_perms_7_w; // @[Reg.scala 16:16]
  reg  l3_ramDatas_7_entries_perms_7_r; // @[Reg.scala 16:16]
  reg  l3_ramDatas_7_entries_prefetch; // @[Reg.scala 16:16]
  reg [38:0] l3_ramDatas_7_ecc; // @[Reg.scala 16:16]
  reg  l3_hitVec_0; // @[Reg.scala 16:16]
  reg  l3_hitVec_1; // @[Reg.scala 16:16]
  reg  l3_hitVec_2; // @[Reg.scala 16:16]
  reg  l3_hitVec_3; // @[Reg.scala 16:16]
  reg  l3_hitVec_4; // @[Reg.scala 16:16]
  reg  l3_hitVec_5; // @[Reg.scala 16:16]
  reg  l3_hitVec_6; // @[Reg.scala 16:16]
  reg  l3_hitVec_7; // @[Reg.scala 16:16]
  wire [21:0] _T_206_entries_tag = l3_hitVec_0 ? l3_ramDatas_0_entries_tag : l3_ramDatas_1_entries_tag; // @[ParallelMux.scala 90:77]
  wire [15:0] _T_206_entries_asid = l3_hitVec_0 ? l3_ramDatas_0_entries_asid : l3_ramDatas_1_entries_asid; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_206_entries_ppns_0 = l3_hitVec_0 ? l3_ramDatas_0_entries_ppns_0 : l3_ramDatas_1_entries_ppns_0; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_206_entries_ppns_1 = l3_hitVec_0 ? l3_ramDatas_0_entries_ppns_1 : l3_ramDatas_1_entries_ppns_1; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_206_entries_ppns_2 = l3_hitVec_0 ? l3_ramDatas_0_entries_ppns_2 : l3_ramDatas_1_entries_ppns_2; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_206_entries_ppns_3 = l3_hitVec_0 ? l3_ramDatas_0_entries_ppns_3 : l3_ramDatas_1_entries_ppns_3; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_206_entries_ppns_4 = l3_hitVec_0 ? l3_ramDatas_0_entries_ppns_4 : l3_ramDatas_1_entries_ppns_4; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_206_entries_ppns_5 = l3_hitVec_0 ? l3_ramDatas_0_entries_ppns_5 : l3_ramDatas_1_entries_ppns_5; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_206_entries_ppns_6 = l3_hitVec_0 ? l3_ramDatas_0_entries_ppns_6 : l3_ramDatas_1_entries_ppns_6; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_206_entries_ppns_7 = l3_hitVec_0 ? l3_ramDatas_0_entries_ppns_7 : l3_ramDatas_1_entries_ppns_7; // @[ParallelMux.scala 90:77]
  wire  _T_206_entries_vs_0 = l3_hitVec_0 ? l3_ramDatas_0_entries_vs_0 : l3_ramDatas_1_entries_vs_0; // @[ParallelMux.scala 90:77]
  wire  _T_206_entries_vs_1 = l3_hitVec_0 ? l3_ramDatas_0_entries_vs_1 : l3_ramDatas_1_entries_vs_1; // @[ParallelMux.scala 90:77]
  wire  _T_206_entries_vs_2 = l3_hitVec_0 ? l3_ramDatas_0_entries_vs_2 : l3_ramDatas_1_entries_vs_2; // @[ParallelMux.scala 90:77]
  wire  _T_206_entries_vs_3 = l3_hitVec_0 ? l3_ramDatas_0_entries_vs_3 : l3_ramDatas_1_entries_vs_3; // @[ParallelMux.scala 90:77]
  wire  _T_206_entries_vs_4 = l3_hitVec_0 ? l3_ramDatas_0_entries_vs_4 : l3_ramDatas_1_entries_vs_4; // @[ParallelMux.scala 90:77]
  wire  _T_206_entries_vs_5 = l3_hitVec_0 ? l3_ramDatas_0_entries_vs_5 : l3_ramDatas_1_entries_vs_5; // @[ParallelMux.scala 90:77]
  wire  _T_206_entries_vs_6 = l3_hitVec_0 ? l3_ramDatas_0_entries_vs_6 : l3_ramDatas_1_entries_vs_6; // @[ParallelMux.scala 90:77]
  wire  _T_206_entries_vs_7 = l3_hitVec_0 ? l3_ramDatas_0_entries_vs_7 : l3_ramDatas_1_entries_vs_7; // @[ParallelMux.scala 90:77]
  wire  _T_206_entries_perms_0_d = l3_hitVec_0 ? l3_ramDatas_0_entries_perms_0_d : l3_ramDatas_1_entries_perms_0_d; // @[ParallelMux.scala 90:77]
  wire  _T_206_entries_perms_0_a = l3_hitVec_0 ? l3_ramDatas_0_entries_perms_0_a : l3_ramDatas_1_entries_perms_0_a; // @[ParallelMux.scala 90:77]
  wire  _T_206_entries_perms_0_g = l3_hitVec_0 ? l3_ramDatas_0_entries_perms_0_g : l3_ramDatas_1_entries_perms_0_g; // @[ParallelMux.scala 90:77]
  wire  _T_206_entries_perms_0_u = l3_hitVec_0 ? l3_ramDatas_0_entries_perms_0_u : l3_ramDatas_1_entries_perms_0_u; // @[ParallelMux.scala 90:77]
  wire  _T_206_entries_perms_0_x = l3_hitVec_0 ? l3_ramDatas_0_entries_perms_0_x : l3_ramDatas_1_entries_perms_0_x; // @[ParallelMux.scala 90:77]
  wire  _T_206_entries_perms_0_w = l3_hitVec_0 ? l3_ramDatas_0_entries_perms_0_w : l3_ramDatas_1_entries_perms_0_w; // @[ParallelMux.scala 90:77]
  wire  _T_206_entries_perms_0_r = l3_hitVec_0 ? l3_ramDatas_0_entries_perms_0_r : l3_ramDatas_1_entries_perms_0_r; // @[ParallelMux.scala 90:77]
  wire  _T_206_entries_perms_1_d = l3_hitVec_0 ? l3_ramDatas_0_entries_perms_1_d : l3_ramDatas_1_entries_perms_1_d; // @[ParallelMux.scala 90:77]
  wire  _T_206_entries_perms_1_a = l3_hitVec_0 ? l3_ramDatas_0_entries_perms_1_a : l3_ramDatas_1_entries_perms_1_a; // @[ParallelMux.scala 90:77]
  wire  _T_206_entries_perms_1_g = l3_hitVec_0 ? l3_ramDatas_0_entries_perms_1_g : l3_ramDatas_1_entries_perms_1_g; // @[ParallelMux.scala 90:77]
  wire  _T_206_entries_perms_1_u = l3_hitVec_0 ? l3_ramDatas_0_entries_perms_1_u : l3_ramDatas_1_entries_perms_1_u; // @[ParallelMux.scala 90:77]
  wire  _T_206_entries_perms_1_x = l3_hitVec_0 ? l3_ramDatas_0_entries_perms_1_x : l3_ramDatas_1_entries_perms_1_x; // @[ParallelMux.scala 90:77]
  wire  _T_206_entries_perms_1_w = l3_hitVec_0 ? l3_ramDatas_0_entries_perms_1_w : l3_ramDatas_1_entries_perms_1_w; // @[ParallelMux.scala 90:77]
  wire  _T_206_entries_perms_1_r = l3_hitVec_0 ? l3_ramDatas_0_entries_perms_1_r : l3_ramDatas_1_entries_perms_1_r; // @[ParallelMux.scala 90:77]
  wire  _T_206_entries_perms_2_d = l3_hitVec_0 ? l3_ramDatas_0_entries_perms_2_d : l3_ramDatas_1_entries_perms_2_d; // @[ParallelMux.scala 90:77]
  wire  _T_206_entries_perms_2_a = l3_hitVec_0 ? l3_ramDatas_0_entries_perms_2_a : l3_ramDatas_1_entries_perms_2_a; // @[ParallelMux.scala 90:77]
  wire  _T_206_entries_perms_2_g = l3_hitVec_0 ? l3_ramDatas_0_entries_perms_2_g : l3_ramDatas_1_entries_perms_2_g; // @[ParallelMux.scala 90:77]
  wire  _T_206_entries_perms_2_u = l3_hitVec_0 ? l3_ramDatas_0_entries_perms_2_u : l3_ramDatas_1_entries_perms_2_u; // @[ParallelMux.scala 90:77]
  wire  _T_206_entries_perms_2_x = l3_hitVec_0 ? l3_ramDatas_0_entries_perms_2_x : l3_ramDatas_1_entries_perms_2_x; // @[ParallelMux.scala 90:77]
  wire  _T_206_entries_perms_2_w = l3_hitVec_0 ? l3_ramDatas_0_entries_perms_2_w : l3_ramDatas_1_entries_perms_2_w; // @[ParallelMux.scala 90:77]
  wire  _T_206_entries_perms_2_r = l3_hitVec_0 ? l3_ramDatas_0_entries_perms_2_r : l3_ramDatas_1_entries_perms_2_r; // @[ParallelMux.scala 90:77]
  wire  _T_206_entries_perms_3_d = l3_hitVec_0 ? l3_ramDatas_0_entries_perms_3_d : l3_ramDatas_1_entries_perms_3_d; // @[ParallelMux.scala 90:77]
  wire  _T_206_entries_perms_3_a = l3_hitVec_0 ? l3_ramDatas_0_entries_perms_3_a : l3_ramDatas_1_entries_perms_3_a; // @[ParallelMux.scala 90:77]
  wire  _T_206_entries_perms_3_g = l3_hitVec_0 ? l3_ramDatas_0_entries_perms_3_g : l3_ramDatas_1_entries_perms_3_g; // @[ParallelMux.scala 90:77]
  wire  _T_206_entries_perms_3_u = l3_hitVec_0 ? l3_ramDatas_0_entries_perms_3_u : l3_ramDatas_1_entries_perms_3_u; // @[ParallelMux.scala 90:77]
  wire  _T_206_entries_perms_3_x = l3_hitVec_0 ? l3_ramDatas_0_entries_perms_3_x : l3_ramDatas_1_entries_perms_3_x; // @[ParallelMux.scala 90:77]
  wire  _T_206_entries_perms_3_w = l3_hitVec_0 ? l3_ramDatas_0_entries_perms_3_w : l3_ramDatas_1_entries_perms_3_w; // @[ParallelMux.scala 90:77]
  wire  _T_206_entries_perms_3_r = l3_hitVec_0 ? l3_ramDatas_0_entries_perms_3_r : l3_ramDatas_1_entries_perms_3_r; // @[ParallelMux.scala 90:77]
  wire  _T_206_entries_perms_4_d = l3_hitVec_0 ? l3_ramDatas_0_entries_perms_4_d : l3_ramDatas_1_entries_perms_4_d; // @[ParallelMux.scala 90:77]
  wire  _T_206_entries_perms_4_a = l3_hitVec_0 ? l3_ramDatas_0_entries_perms_4_a : l3_ramDatas_1_entries_perms_4_a; // @[ParallelMux.scala 90:77]
  wire  _T_206_entries_perms_4_g = l3_hitVec_0 ? l3_ramDatas_0_entries_perms_4_g : l3_ramDatas_1_entries_perms_4_g; // @[ParallelMux.scala 90:77]
  wire  _T_206_entries_perms_4_u = l3_hitVec_0 ? l3_ramDatas_0_entries_perms_4_u : l3_ramDatas_1_entries_perms_4_u; // @[ParallelMux.scala 90:77]
  wire  _T_206_entries_perms_4_x = l3_hitVec_0 ? l3_ramDatas_0_entries_perms_4_x : l3_ramDatas_1_entries_perms_4_x; // @[ParallelMux.scala 90:77]
  wire  _T_206_entries_perms_4_w = l3_hitVec_0 ? l3_ramDatas_0_entries_perms_4_w : l3_ramDatas_1_entries_perms_4_w; // @[ParallelMux.scala 90:77]
  wire  _T_206_entries_perms_4_r = l3_hitVec_0 ? l3_ramDatas_0_entries_perms_4_r : l3_ramDatas_1_entries_perms_4_r; // @[ParallelMux.scala 90:77]
  wire  _T_206_entries_perms_5_d = l3_hitVec_0 ? l3_ramDatas_0_entries_perms_5_d : l3_ramDatas_1_entries_perms_5_d; // @[ParallelMux.scala 90:77]
  wire  _T_206_entries_perms_5_a = l3_hitVec_0 ? l3_ramDatas_0_entries_perms_5_a : l3_ramDatas_1_entries_perms_5_a; // @[ParallelMux.scala 90:77]
  wire  _T_206_entries_perms_5_g = l3_hitVec_0 ? l3_ramDatas_0_entries_perms_5_g : l3_ramDatas_1_entries_perms_5_g; // @[ParallelMux.scala 90:77]
  wire  _T_206_entries_perms_5_u = l3_hitVec_0 ? l3_ramDatas_0_entries_perms_5_u : l3_ramDatas_1_entries_perms_5_u; // @[ParallelMux.scala 90:77]
  wire  _T_206_entries_perms_5_x = l3_hitVec_0 ? l3_ramDatas_0_entries_perms_5_x : l3_ramDatas_1_entries_perms_5_x; // @[ParallelMux.scala 90:77]
  wire  _T_206_entries_perms_5_w = l3_hitVec_0 ? l3_ramDatas_0_entries_perms_5_w : l3_ramDatas_1_entries_perms_5_w; // @[ParallelMux.scala 90:77]
  wire  _T_206_entries_perms_5_r = l3_hitVec_0 ? l3_ramDatas_0_entries_perms_5_r : l3_ramDatas_1_entries_perms_5_r; // @[ParallelMux.scala 90:77]
  wire  _T_206_entries_perms_6_d = l3_hitVec_0 ? l3_ramDatas_0_entries_perms_6_d : l3_ramDatas_1_entries_perms_6_d; // @[ParallelMux.scala 90:77]
  wire  _T_206_entries_perms_6_a = l3_hitVec_0 ? l3_ramDatas_0_entries_perms_6_a : l3_ramDatas_1_entries_perms_6_a; // @[ParallelMux.scala 90:77]
  wire  _T_206_entries_perms_6_g = l3_hitVec_0 ? l3_ramDatas_0_entries_perms_6_g : l3_ramDatas_1_entries_perms_6_g; // @[ParallelMux.scala 90:77]
  wire  _T_206_entries_perms_6_u = l3_hitVec_0 ? l3_ramDatas_0_entries_perms_6_u : l3_ramDatas_1_entries_perms_6_u; // @[ParallelMux.scala 90:77]
  wire  _T_206_entries_perms_6_x = l3_hitVec_0 ? l3_ramDatas_0_entries_perms_6_x : l3_ramDatas_1_entries_perms_6_x; // @[ParallelMux.scala 90:77]
  wire  _T_206_entries_perms_6_w = l3_hitVec_0 ? l3_ramDatas_0_entries_perms_6_w : l3_ramDatas_1_entries_perms_6_w; // @[ParallelMux.scala 90:77]
  wire  _T_206_entries_perms_6_r = l3_hitVec_0 ? l3_ramDatas_0_entries_perms_6_r : l3_ramDatas_1_entries_perms_6_r; // @[ParallelMux.scala 90:77]
  wire  _T_206_entries_perms_7_d = l3_hitVec_0 ? l3_ramDatas_0_entries_perms_7_d : l3_ramDatas_1_entries_perms_7_d; // @[ParallelMux.scala 90:77]
  wire  _T_206_entries_perms_7_a = l3_hitVec_0 ? l3_ramDatas_0_entries_perms_7_a : l3_ramDatas_1_entries_perms_7_a; // @[ParallelMux.scala 90:77]
  wire  _T_206_entries_perms_7_g = l3_hitVec_0 ? l3_ramDatas_0_entries_perms_7_g : l3_ramDatas_1_entries_perms_7_g; // @[ParallelMux.scala 90:77]
  wire  _T_206_entries_perms_7_u = l3_hitVec_0 ? l3_ramDatas_0_entries_perms_7_u : l3_ramDatas_1_entries_perms_7_u; // @[ParallelMux.scala 90:77]
  wire  _T_206_entries_perms_7_x = l3_hitVec_0 ? l3_ramDatas_0_entries_perms_7_x : l3_ramDatas_1_entries_perms_7_x; // @[ParallelMux.scala 90:77]
  wire  _T_206_entries_perms_7_w = l3_hitVec_0 ? l3_ramDatas_0_entries_perms_7_w : l3_ramDatas_1_entries_perms_7_w; // @[ParallelMux.scala 90:77]
  wire  _T_206_entries_perms_7_r = l3_hitVec_0 ? l3_ramDatas_0_entries_perms_7_r : l3_ramDatas_1_entries_perms_7_r; // @[ParallelMux.scala 90:77]
  wire  _T_206_entries_prefetch = l3_hitVec_0 ? l3_ramDatas_0_entries_prefetch : l3_ramDatas_1_entries_prefetch; // @[ParallelMux.scala 90:77]
  wire [38:0] _T_206_ecc = l3_hitVec_0 ? l3_ramDatas_0_ecc : l3_ramDatas_1_ecc; // @[ParallelMux.scala 90:77]
  wire [21:0] _T_208_entries_tag = l3_hitVec_2 ? l3_ramDatas_2_entries_tag : l3_ramDatas_3_entries_tag; // @[ParallelMux.scala 90:77]
  wire [15:0] _T_208_entries_asid = l3_hitVec_2 ? l3_ramDatas_2_entries_asid : l3_ramDatas_3_entries_asid; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_208_entries_ppns_0 = l3_hitVec_2 ? l3_ramDatas_2_entries_ppns_0 : l3_ramDatas_3_entries_ppns_0; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_208_entries_ppns_1 = l3_hitVec_2 ? l3_ramDatas_2_entries_ppns_1 : l3_ramDatas_3_entries_ppns_1; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_208_entries_ppns_2 = l3_hitVec_2 ? l3_ramDatas_2_entries_ppns_2 : l3_ramDatas_3_entries_ppns_2; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_208_entries_ppns_3 = l3_hitVec_2 ? l3_ramDatas_2_entries_ppns_3 : l3_ramDatas_3_entries_ppns_3; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_208_entries_ppns_4 = l3_hitVec_2 ? l3_ramDatas_2_entries_ppns_4 : l3_ramDatas_3_entries_ppns_4; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_208_entries_ppns_5 = l3_hitVec_2 ? l3_ramDatas_2_entries_ppns_5 : l3_ramDatas_3_entries_ppns_5; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_208_entries_ppns_6 = l3_hitVec_2 ? l3_ramDatas_2_entries_ppns_6 : l3_ramDatas_3_entries_ppns_6; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_208_entries_ppns_7 = l3_hitVec_2 ? l3_ramDatas_2_entries_ppns_7 : l3_ramDatas_3_entries_ppns_7; // @[ParallelMux.scala 90:77]
  wire  _T_208_entries_vs_0 = l3_hitVec_2 ? l3_ramDatas_2_entries_vs_0 : l3_ramDatas_3_entries_vs_0; // @[ParallelMux.scala 90:77]
  wire  _T_208_entries_vs_1 = l3_hitVec_2 ? l3_ramDatas_2_entries_vs_1 : l3_ramDatas_3_entries_vs_1; // @[ParallelMux.scala 90:77]
  wire  _T_208_entries_vs_2 = l3_hitVec_2 ? l3_ramDatas_2_entries_vs_2 : l3_ramDatas_3_entries_vs_2; // @[ParallelMux.scala 90:77]
  wire  _T_208_entries_vs_3 = l3_hitVec_2 ? l3_ramDatas_2_entries_vs_3 : l3_ramDatas_3_entries_vs_3; // @[ParallelMux.scala 90:77]
  wire  _T_208_entries_vs_4 = l3_hitVec_2 ? l3_ramDatas_2_entries_vs_4 : l3_ramDatas_3_entries_vs_4; // @[ParallelMux.scala 90:77]
  wire  _T_208_entries_vs_5 = l3_hitVec_2 ? l3_ramDatas_2_entries_vs_5 : l3_ramDatas_3_entries_vs_5; // @[ParallelMux.scala 90:77]
  wire  _T_208_entries_vs_6 = l3_hitVec_2 ? l3_ramDatas_2_entries_vs_6 : l3_ramDatas_3_entries_vs_6; // @[ParallelMux.scala 90:77]
  wire  _T_208_entries_vs_7 = l3_hitVec_2 ? l3_ramDatas_2_entries_vs_7 : l3_ramDatas_3_entries_vs_7; // @[ParallelMux.scala 90:77]
  wire  _T_208_entries_perms_0_d = l3_hitVec_2 ? l3_ramDatas_2_entries_perms_0_d : l3_ramDatas_3_entries_perms_0_d; // @[ParallelMux.scala 90:77]
  wire  _T_208_entries_perms_0_a = l3_hitVec_2 ? l3_ramDatas_2_entries_perms_0_a : l3_ramDatas_3_entries_perms_0_a; // @[ParallelMux.scala 90:77]
  wire  _T_208_entries_perms_0_g = l3_hitVec_2 ? l3_ramDatas_2_entries_perms_0_g : l3_ramDatas_3_entries_perms_0_g; // @[ParallelMux.scala 90:77]
  wire  _T_208_entries_perms_0_u = l3_hitVec_2 ? l3_ramDatas_2_entries_perms_0_u : l3_ramDatas_3_entries_perms_0_u; // @[ParallelMux.scala 90:77]
  wire  _T_208_entries_perms_0_x = l3_hitVec_2 ? l3_ramDatas_2_entries_perms_0_x : l3_ramDatas_3_entries_perms_0_x; // @[ParallelMux.scala 90:77]
  wire  _T_208_entries_perms_0_w = l3_hitVec_2 ? l3_ramDatas_2_entries_perms_0_w : l3_ramDatas_3_entries_perms_0_w; // @[ParallelMux.scala 90:77]
  wire  _T_208_entries_perms_0_r = l3_hitVec_2 ? l3_ramDatas_2_entries_perms_0_r : l3_ramDatas_3_entries_perms_0_r; // @[ParallelMux.scala 90:77]
  wire  _T_208_entries_perms_1_d = l3_hitVec_2 ? l3_ramDatas_2_entries_perms_1_d : l3_ramDatas_3_entries_perms_1_d; // @[ParallelMux.scala 90:77]
  wire  _T_208_entries_perms_1_a = l3_hitVec_2 ? l3_ramDatas_2_entries_perms_1_a : l3_ramDatas_3_entries_perms_1_a; // @[ParallelMux.scala 90:77]
  wire  _T_208_entries_perms_1_g = l3_hitVec_2 ? l3_ramDatas_2_entries_perms_1_g : l3_ramDatas_3_entries_perms_1_g; // @[ParallelMux.scala 90:77]
  wire  _T_208_entries_perms_1_u = l3_hitVec_2 ? l3_ramDatas_2_entries_perms_1_u : l3_ramDatas_3_entries_perms_1_u; // @[ParallelMux.scala 90:77]
  wire  _T_208_entries_perms_1_x = l3_hitVec_2 ? l3_ramDatas_2_entries_perms_1_x : l3_ramDatas_3_entries_perms_1_x; // @[ParallelMux.scala 90:77]
  wire  _T_208_entries_perms_1_w = l3_hitVec_2 ? l3_ramDatas_2_entries_perms_1_w : l3_ramDatas_3_entries_perms_1_w; // @[ParallelMux.scala 90:77]
  wire  _T_208_entries_perms_1_r = l3_hitVec_2 ? l3_ramDatas_2_entries_perms_1_r : l3_ramDatas_3_entries_perms_1_r; // @[ParallelMux.scala 90:77]
  wire  _T_208_entries_perms_2_d = l3_hitVec_2 ? l3_ramDatas_2_entries_perms_2_d : l3_ramDatas_3_entries_perms_2_d; // @[ParallelMux.scala 90:77]
  wire  _T_208_entries_perms_2_a = l3_hitVec_2 ? l3_ramDatas_2_entries_perms_2_a : l3_ramDatas_3_entries_perms_2_a; // @[ParallelMux.scala 90:77]
  wire  _T_208_entries_perms_2_g = l3_hitVec_2 ? l3_ramDatas_2_entries_perms_2_g : l3_ramDatas_3_entries_perms_2_g; // @[ParallelMux.scala 90:77]
  wire  _T_208_entries_perms_2_u = l3_hitVec_2 ? l3_ramDatas_2_entries_perms_2_u : l3_ramDatas_3_entries_perms_2_u; // @[ParallelMux.scala 90:77]
  wire  _T_208_entries_perms_2_x = l3_hitVec_2 ? l3_ramDatas_2_entries_perms_2_x : l3_ramDatas_3_entries_perms_2_x; // @[ParallelMux.scala 90:77]
  wire  _T_208_entries_perms_2_w = l3_hitVec_2 ? l3_ramDatas_2_entries_perms_2_w : l3_ramDatas_3_entries_perms_2_w; // @[ParallelMux.scala 90:77]
  wire  _T_208_entries_perms_2_r = l3_hitVec_2 ? l3_ramDatas_2_entries_perms_2_r : l3_ramDatas_3_entries_perms_2_r; // @[ParallelMux.scala 90:77]
  wire  _T_208_entries_perms_3_d = l3_hitVec_2 ? l3_ramDatas_2_entries_perms_3_d : l3_ramDatas_3_entries_perms_3_d; // @[ParallelMux.scala 90:77]
  wire  _T_208_entries_perms_3_a = l3_hitVec_2 ? l3_ramDatas_2_entries_perms_3_a : l3_ramDatas_3_entries_perms_3_a; // @[ParallelMux.scala 90:77]
  wire  _T_208_entries_perms_3_g = l3_hitVec_2 ? l3_ramDatas_2_entries_perms_3_g : l3_ramDatas_3_entries_perms_3_g; // @[ParallelMux.scala 90:77]
  wire  _T_208_entries_perms_3_u = l3_hitVec_2 ? l3_ramDatas_2_entries_perms_3_u : l3_ramDatas_3_entries_perms_3_u; // @[ParallelMux.scala 90:77]
  wire  _T_208_entries_perms_3_x = l3_hitVec_2 ? l3_ramDatas_2_entries_perms_3_x : l3_ramDatas_3_entries_perms_3_x; // @[ParallelMux.scala 90:77]
  wire  _T_208_entries_perms_3_w = l3_hitVec_2 ? l3_ramDatas_2_entries_perms_3_w : l3_ramDatas_3_entries_perms_3_w; // @[ParallelMux.scala 90:77]
  wire  _T_208_entries_perms_3_r = l3_hitVec_2 ? l3_ramDatas_2_entries_perms_3_r : l3_ramDatas_3_entries_perms_3_r; // @[ParallelMux.scala 90:77]
  wire  _T_208_entries_perms_4_d = l3_hitVec_2 ? l3_ramDatas_2_entries_perms_4_d : l3_ramDatas_3_entries_perms_4_d; // @[ParallelMux.scala 90:77]
  wire  _T_208_entries_perms_4_a = l3_hitVec_2 ? l3_ramDatas_2_entries_perms_4_a : l3_ramDatas_3_entries_perms_4_a; // @[ParallelMux.scala 90:77]
  wire  _T_208_entries_perms_4_g = l3_hitVec_2 ? l3_ramDatas_2_entries_perms_4_g : l3_ramDatas_3_entries_perms_4_g; // @[ParallelMux.scala 90:77]
  wire  _T_208_entries_perms_4_u = l3_hitVec_2 ? l3_ramDatas_2_entries_perms_4_u : l3_ramDatas_3_entries_perms_4_u; // @[ParallelMux.scala 90:77]
  wire  _T_208_entries_perms_4_x = l3_hitVec_2 ? l3_ramDatas_2_entries_perms_4_x : l3_ramDatas_3_entries_perms_4_x; // @[ParallelMux.scala 90:77]
  wire  _T_208_entries_perms_4_w = l3_hitVec_2 ? l3_ramDatas_2_entries_perms_4_w : l3_ramDatas_3_entries_perms_4_w; // @[ParallelMux.scala 90:77]
  wire  _T_208_entries_perms_4_r = l3_hitVec_2 ? l3_ramDatas_2_entries_perms_4_r : l3_ramDatas_3_entries_perms_4_r; // @[ParallelMux.scala 90:77]
  wire  _T_208_entries_perms_5_d = l3_hitVec_2 ? l3_ramDatas_2_entries_perms_5_d : l3_ramDatas_3_entries_perms_5_d; // @[ParallelMux.scala 90:77]
  wire  _T_208_entries_perms_5_a = l3_hitVec_2 ? l3_ramDatas_2_entries_perms_5_a : l3_ramDatas_3_entries_perms_5_a; // @[ParallelMux.scala 90:77]
  wire  _T_208_entries_perms_5_g = l3_hitVec_2 ? l3_ramDatas_2_entries_perms_5_g : l3_ramDatas_3_entries_perms_5_g; // @[ParallelMux.scala 90:77]
  wire  _T_208_entries_perms_5_u = l3_hitVec_2 ? l3_ramDatas_2_entries_perms_5_u : l3_ramDatas_3_entries_perms_5_u; // @[ParallelMux.scala 90:77]
  wire  _T_208_entries_perms_5_x = l3_hitVec_2 ? l3_ramDatas_2_entries_perms_5_x : l3_ramDatas_3_entries_perms_5_x; // @[ParallelMux.scala 90:77]
  wire  _T_208_entries_perms_5_w = l3_hitVec_2 ? l3_ramDatas_2_entries_perms_5_w : l3_ramDatas_3_entries_perms_5_w; // @[ParallelMux.scala 90:77]
  wire  _T_208_entries_perms_5_r = l3_hitVec_2 ? l3_ramDatas_2_entries_perms_5_r : l3_ramDatas_3_entries_perms_5_r; // @[ParallelMux.scala 90:77]
  wire  _T_208_entries_perms_6_d = l3_hitVec_2 ? l3_ramDatas_2_entries_perms_6_d : l3_ramDatas_3_entries_perms_6_d; // @[ParallelMux.scala 90:77]
  wire  _T_208_entries_perms_6_a = l3_hitVec_2 ? l3_ramDatas_2_entries_perms_6_a : l3_ramDatas_3_entries_perms_6_a; // @[ParallelMux.scala 90:77]
  wire  _T_208_entries_perms_6_g = l3_hitVec_2 ? l3_ramDatas_2_entries_perms_6_g : l3_ramDatas_3_entries_perms_6_g; // @[ParallelMux.scala 90:77]
  wire  _T_208_entries_perms_6_u = l3_hitVec_2 ? l3_ramDatas_2_entries_perms_6_u : l3_ramDatas_3_entries_perms_6_u; // @[ParallelMux.scala 90:77]
  wire  _T_208_entries_perms_6_x = l3_hitVec_2 ? l3_ramDatas_2_entries_perms_6_x : l3_ramDatas_3_entries_perms_6_x; // @[ParallelMux.scala 90:77]
  wire  _T_208_entries_perms_6_w = l3_hitVec_2 ? l3_ramDatas_2_entries_perms_6_w : l3_ramDatas_3_entries_perms_6_w; // @[ParallelMux.scala 90:77]
  wire  _T_208_entries_perms_6_r = l3_hitVec_2 ? l3_ramDatas_2_entries_perms_6_r : l3_ramDatas_3_entries_perms_6_r; // @[ParallelMux.scala 90:77]
  wire  _T_208_entries_perms_7_d = l3_hitVec_2 ? l3_ramDatas_2_entries_perms_7_d : l3_ramDatas_3_entries_perms_7_d; // @[ParallelMux.scala 90:77]
  wire  _T_208_entries_perms_7_a = l3_hitVec_2 ? l3_ramDatas_2_entries_perms_7_a : l3_ramDatas_3_entries_perms_7_a; // @[ParallelMux.scala 90:77]
  wire  _T_208_entries_perms_7_g = l3_hitVec_2 ? l3_ramDatas_2_entries_perms_7_g : l3_ramDatas_3_entries_perms_7_g; // @[ParallelMux.scala 90:77]
  wire  _T_208_entries_perms_7_u = l3_hitVec_2 ? l3_ramDatas_2_entries_perms_7_u : l3_ramDatas_3_entries_perms_7_u; // @[ParallelMux.scala 90:77]
  wire  _T_208_entries_perms_7_x = l3_hitVec_2 ? l3_ramDatas_2_entries_perms_7_x : l3_ramDatas_3_entries_perms_7_x; // @[ParallelMux.scala 90:77]
  wire  _T_208_entries_perms_7_w = l3_hitVec_2 ? l3_ramDatas_2_entries_perms_7_w : l3_ramDatas_3_entries_perms_7_w; // @[ParallelMux.scala 90:77]
  wire  _T_208_entries_perms_7_r = l3_hitVec_2 ? l3_ramDatas_2_entries_perms_7_r : l3_ramDatas_3_entries_perms_7_r; // @[ParallelMux.scala 90:77]
  wire  _T_208_entries_prefetch = l3_hitVec_2 ? l3_ramDatas_2_entries_prefetch : l3_ramDatas_3_entries_prefetch; // @[ParallelMux.scala 90:77]
  wire [38:0] _T_208_ecc = l3_hitVec_2 ? l3_ramDatas_2_ecc : l3_ramDatas_3_ecc; // @[ParallelMux.scala 90:77]
  wire  _T_209 = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3); // @[ParallelMux.scala 90:65]
  wire [21:0] _T_210_entries_tag = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_tag : _T_208_entries_tag; // @[ParallelMux.scala 90:77]
  wire [15:0] _T_210_entries_asid = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_asid : _T_208_entries_asid; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_210_entries_ppns_0 = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_ppns_0 : _T_208_entries_ppns_0; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_210_entries_ppns_1 = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_ppns_1 : _T_208_entries_ppns_1; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_210_entries_ppns_2 = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_ppns_2 : _T_208_entries_ppns_2; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_210_entries_ppns_3 = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_ppns_3 : _T_208_entries_ppns_3; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_210_entries_ppns_4 = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_ppns_4 : _T_208_entries_ppns_4; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_210_entries_ppns_5 = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_ppns_5 : _T_208_entries_ppns_5; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_210_entries_ppns_6 = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_ppns_6 : _T_208_entries_ppns_6; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_210_entries_ppns_7 = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_ppns_7 : _T_208_entries_ppns_7; // @[ParallelMux.scala 90:77]
  wire  _T_210_entries_vs_0 = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_vs_0 : _T_208_entries_vs_0; // @[ParallelMux.scala 90:77]
  wire  _T_210_entries_vs_1 = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_vs_1 : _T_208_entries_vs_1; // @[ParallelMux.scala 90:77]
  wire  _T_210_entries_vs_2 = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_vs_2 : _T_208_entries_vs_2; // @[ParallelMux.scala 90:77]
  wire  _T_210_entries_vs_3 = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_vs_3 : _T_208_entries_vs_3; // @[ParallelMux.scala 90:77]
  wire  _T_210_entries_vs_4 = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_vs_4 : _T_208_entries_vs_4; // @[ParallelMux.scala 90:77]
  wire  _T_210_entries_vs_5 = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_vs_5 : _T_208_entries_vs_5; // @[ParallelMux.scala 90:77]
  wire  _T_210_entries_vs_6 = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_vs_6 : _T_208_entries_vs_6; // @[ParallelMux.scala 90:77]
  wire  _T_210_entries_vs_7 = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_vs_7 : _T_208_entries_vs_7; // @[ParallelMux.scala 90:77]
  wire  _T_210_entries_perms_0_d = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_perms_0_d : _T_208_entries_perms_0_d; // @[ParallelMux.scala 90:77]
  wire  _T_210_entries_perms_0_a = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_perms_0_a : _T_208_entries_perms_0_a; // @[ParallelMux.scala 90:77]
  wire  _T_210_entries_perms_0_g = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_perms_0_g : _T_208_entries_perms_0_g; // @[ParallelMux.scala 90:77]
  wire  _T_210_entries_perms_0_u = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_perms_0_u : _T_208_entries_perms_0_u; // @[ParallelMux.scala 90:77]
  wire  _T_210_entries_perms_0_x = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_perms_0_x : _T_208_entries_perms_0_x; // @[ParallelMux.scala 90:77]
  wire  _T_210_entries_perms_0_w = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_perms_0_w : _T_208_entries_perms_0_w; // @[ParallelMux.scala 90:77]
  wire  _T_210_entries_perms_0_r = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_perms_0_r : _T_208_entries_perms_0_r; // @[ParallelMux.scala 90:77]
  wire  _T_210_entries_perms_1_d = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_perms_1_d : _T_208_entries_perms_1_d; // @[ParallelMux.scala 90:77]
  wire  _T_210_entries_perms_1_a = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_perms_1_a : _T_208_entries_perms_1_a; // @[ParallelMux.scala 90:77]
  wire  _T_210_entries_perms_1_g = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_perms_1_g : _T_208_entries_perms_1_g; // @[ParallelMux.scala 90:77]
  wire  _T_210_entries_perms_1_u = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_perms_1_u : _T_208_entries_perms_1_u; // @[ParallelMux.scala 90:77]
  wire  _T_210_entries_perms_1_x = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_perms_1_x : _T_208_entries_perms_1_x; // @[ParallelMux.scala 90:77]
  wire  _T_210_entries_perms_1_w = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_perms_1_w : _T_208_entries_perms_1_w; // @[ParallelMux.scala 90:77]
  wire  _T_210_entries_perms_1_r = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_perms_1_r : _T_208_entries_perms_1_r; // @[ParallelMux.scala 90:77]
  wire  _T_210_entries_perms_2_d = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_perms_2_d : _T_208_entries_perms_2_d; // @[ParallelMux.scala 90:77]
  wire  _T_210_entries_perms_2_a = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_perms_2_a : _T_208_entries_perms_2_a; // @[ParallelMux.scala 90:77]
  wire  _T_210_entries_perms_2_g = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_perms_2_g : _T_208_entries_perms_2_g; // @[ParallelMux.scala 90:77]
  wire  _T_210_entries_perms_2_u = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_perms_2_u : _T_208_entries_perms_2_u; // @[ParallelMux.scala 90:77]
  wire  _T_210_entries_perms_2_x = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_perms_2_x : _T_208_entries_perms_2_x; // @[ParallelMux.scala 90:77]
  wire  _T_210_entries_perms_2_w = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_perms_2_w : _T_208_entries_perms_2_w; // @[ParallelMux.scala 90:77]
  wire  _T_210_entries_perms_2_r = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_perms_2_r : _T_208_entries_perms_2_r; // @[ParallelMux.scala 90:77]
  wire  _T_210_entries_perms_3_d = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_perms_3_d : _T_208_entries_perms_3_d; // @[ParallelMux.scala 90:77]
  wire  _T_210_entries_perms_3_a = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_perms_3_a : _T_208_entries_perms_3_a; // @[ParallelMux.scala 90:77]
  wire  _T_210_entries_perms_3_g = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_perms_3_g : _T_208_entries_perms_3_g; // @[ParallelMux.scala 90:77]
  wire  _T_210_entries_perms_3_u = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_perms_3_u : _T_208_entries_perms_3_u; // @[ParallelMux.scala 90:77]
  wire  _T_210_entries_perms_3_x = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_perms_3_x : _T_208_entries_perms_3_x; // @[ParallelMux.scala 90:77]
  wire  _T_210_entries_perms_3_w = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_perms_3_w : _T_208_entries_perms_3_w; // @[ParallelMux.scala 90:77]
  wire  _T_210_entries_perms_3_r = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_perms_3_r : _T_208_entries_perms_3_r; // @[ParallelMux.scala 90:77]
  wire  _T_210_entries_perms_4_d = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_perms_4_d : _T_208_entries_perms_4_d; // @[ParallelMux.scala 90:77]
  wire  _T_210_entries_perms_4_a = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_perms_4_a : _T_208_entries_perms_4_a; // @[ParallelMux.scala 90:77]
  wire  _T_210_entries_perms_4_g = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_perms_4_g : _T_208_entries_perms_4_g; // @[ParallelMux.scala 90:77]
  wire  _T_210_entries_perms_4_u = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_perms_4_u : _T_208_entries_perms_4_u; // @[ParallelMux.scala 90:77]
  wire  _T_210_entries_perms_4_x = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_perms_4_x : _T_208_entries_perms_4_x; // @[ParallelMux.scala 90:77]
  wire  _T_210_entries_perms_4_w = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_perms_4_w : _T_208_entries_perms_4_w; // @[ParallelMux.scala 90:77]
  wire  _T_210_entries_perms_4_r = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_perms_4_r : _T_208_entries_perms_4_r; // @[ParallelMux.scala 90:77]
  wire  _T_210_entries_perms_5_d = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_perms_5_d : _T_208_entries_perms_5_d; // @[ParallelMux.scala 90:77]
  wire  _T_210_entries_perms_5_a = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_perms_5_a : _T_208_entries_perms_5_a; // @[ParallelMux.scala 90:77]
  wire  _T_210_entries_perms_5_g = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_perms_5_g : _T_208_entries_perms_5_g; // @[ParallelMux.scala 90:77]
  wire  _T_210_entries_perms_5_u = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_perms_5_u : _T_208_entries_perms_5_u; // @[ParallelMux.scala 90:77]
  wire  _T_210_entries_perms_5_x = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_perms_5_x : _T_208_entries_perms_5_x; // @[ParallelMux.scala 90:77]
  wire  _T_210_entries_perms_5_w = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_perms_5_w : _T_208_entries_perms_5_w; // @[ParallelMux.scala 90:77]
  wire  _T_210_entries_perms_5_r = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_perms_5_r : _T_208_entries_perms_5_r; // @[ParallelMux.scala 90:77]
  wire  _T_210_entries_perms_6_d = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_perms_6_d : _T_208_entries_perms_6_d; // @[ParallelMux.scala 90:77]
  wire  _T_210_entries_perms_6_a = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_perms_6_a : _T_208_entries_perms_6_a; // @[ParallelMux.scala 90:77]
  wire  _T_210_entries_perms_6_g = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_perms_6_g : _T_208_entries_perms_6_g; // @[ParallelMux.scala 90:77]
  wire  _T_210_entries_perms_6_u = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_perms_6_u : _T_208_entries_perms_6_u; // @[ParallelMux.scala 90:77]
  wire  _T_210_entries_perms_6_x = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_perms_6_x : _T_208_entries_perms_6_x; // @[ParallelMux.scala 90:77]
  wire  _T_210_entries_perms_6_w = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_perms_6_w : _T_208_entries_perms_6_w; // @[ParallelMux.scala 90:77]
  wire  _T_210_entries_perms_6_r = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_perms_6_r : _T_208_entries_perms_6_r; // @[ParallelMux.scala 90:77]
  wire  _T_210_entries_perms_7_d = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_perms_7_d : _T_208_entries_perms_7_d; // @[ParallelMux.scala 90:77]
  wire  _T_210_entries_perms_7_a = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_perms_7_a : _T_208_entries_perms_7_a; // @[ParallelMux.scala 90:77]
  wire  _T_210_entries_perms_7_g = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_perms_7_g : _T_208_entries_perms_7_g; // @[ParallelMux.scala 90:77]
  wire  _T_210_entries_perms_7_u = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_perms_7_u : _T_208_entries_perms_7_u; // @[ParallelMux.scala 90:77]
  wire  _T_210_entries_perms_7_x = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_perms_7_x : _T_208_entries_perms_7_x; // @[ParallelMux.scala 90:77]
  wire  _T_210_entries_perms_7_w = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_perms_7_w : _T_208_entries_perms_7_w; // @[ParallelMux.scala 90:77]
  wire  _T_210_entries_perms_7_r = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_perms_7_r : _T_208_entries_perms_7_r; // @[ParallelMux.scala 90:77]
  wire  _T_210_entries_prefetch = l3_hitVec_0 | l3_hitVec_1 ? _T_206_entries_prefetch : _T_208_entries_prefetch; // @[ParallelMux.scala 90:77]
  wire [38:0] _T_210_ecc = l3_hitVec_0 | l3_hitVec_1 ? _T_206_ecc : _T_208_ecc; // @[ParallelMux.scala 90:77]
  wire [21:0] _T_212_entries_tag = l3_hitVec_4 ? l3_ramDatas_4_entries_tag : l3_ramDatas_5_entries_tag; // @[ParallelMux.scala 90:77]
  wire [15:0] _T_212_entries_asid = l3_hitVec_4 ? l3_ramDatas_4_entries_asid : l3_ramDatas_5_entries_asid; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_212_entries_ppns_0 = l3_hitVec_4 ? l3_ramDatas_4_entries_ppns_0 : l3_ramDatas_5_entries_ppns_0; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_212_entries_ppns_1 = l3_hitVec_4 ? l3_ramDatas_4_entries_ppns_1 : l3_ramDatas_5_entries_ppns_1; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_212_entries_ppns_2 = l3_hitVec_4 ? l3_ramDatas_4_entries_ppns_2 : l3_ramDatas_5_entries_ppns_2; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_212_entries_ppns_3 = l3_hitVec_4 ? l3_ramDatas_4_entries_ppns_3 : l3_ramDatas_5_entries_ppns_3; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_212_entries_ppns_4 = l3_hitVec_4 ? l3_ramDatas_4_entries_ppns_4 : l3_ramDatas_5_entries_ppns_4; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_212_entries_ppns_5 = l3_hitVec_4 ? l3_ramDatas_4_entries_ppns_5 : l3_ramDatas_5_entries_ppns_5; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_212_entries_ppns_6 = l3_hitVec_4 ? l3_ramDatas_4_entries_ppns_6 : l3_ramDatas_5_entries_ppns_6; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_212_entries_ppns_7 = l3_hitVec_4 ? l3_ramDatas_4_entries_ppns_7 : l3_ramDatas_5_entries_ppns_7; // @[ParallelMux.scala 90:77]
  wire  _T_212_entries_vs_0 = l3_hitVec_4 ? l3_ramDatas_4_entries_vs_0 : l3_ramDatas_5_entries_vs_0; // @[ParallelMux.scala 90:77]
  wire  _T_212_entries_vs_1 = l3_hitVec_4 ? l3_ramDatas_4_entries_vs_1 : l3_ramDatas_5_entries_vs_1; // @[ParallelMux.scala 90:77]
  wire  _T_212_entries_vs_2 = l3_hitVec_4 ? l3_ramDatas_4_entries_vs_2 : l3_ramDatas_5_entries_vs_2; // @[ParallelMux.scala 90:77]
  wire  _T_212_entries_vs_3 = l3_hitVec_4 ? l3_ramDatas_4_entries_vs_3 : l3_ramDatas_5_entries_vs_3; // @[ParallelMux.scala 90:77]
  wire  _T_212_entries_vs_4 = l3_hitVec_4 ? l3_ramDatas_4_entries_vs_4 : l3_ramDatas_5_entries_vs_4; // @[ParallelMux.scala 90:77]
  wire  _T_212_entries_vs_5 = l3_hitVec_4 ? l3_ramDatas_4_entries_vs_5 : l3_ramDatas_5_entries_vs_5; // @[ParallelMux.scala 90:77]
  wire  _T_212_entries_vs_6 = l3_hitVec_4 ? l3_ramDatas_4_entries_vs_6 : l3_ramDatas_5_entries_vs_6; // @[ParallelMux.scala 90:77]
  wire  _T_212_entries_vs_7 = l3_hitVec_4 ? l3_ramDatas_4_entries_vs_7 : l3_ramDatas_5_entries_vs_7; // @[ParallelMux.scala 90:77]
  wire  _T_212_entries_perms_0_d = l3_hitVec_4 ? l3_ramDatas_4_entries_perms_0_d : l3_ramDatas_5_entries_perms_0_d; // @[ParallelMux.scala 90:77]
  wire  _T_212_entries_perms_0_a = l3_hitVec_4 ? l3_ramDatas_4_entries_perms_0_a : l3_ramDatas_5_entries_perms_0_a; // @[ParallelMux.scala 90:77]
  wire  _T_212_entries_perms_0_g = l3_hitVec_4 ? l3_ramDatas_4_entries_perms_0_g : l3_ramDatas_5_entries_perms_0_g; // @[ParallelMux.scala 90:77]
  wire  _T_212_entries_perms_0_u = l3_hitVec_4 ? l3_ramDatas_4_entries_perms_0_u : l3_ramDatas_5_entries_perms_0_u; // @[ParallelMux.scala 90:77]
  wire  _T_212_entries_perms_0_x = l3_hitVec_4 ? l3_ramDatas_4_entries_perms_0_x : l3_ramDatas_5_entries_perms_0_x; // @[ParallelMux.scala 90:77]
  wire  _T_212_entries_perms_0_w = l3_hitVec_4 ? l3_ramDatas_4_entries_perms_0_w : l3_ramDatas_5_entries_perms_0_w; // @[ParallelMux.scala 90:77]
  wire  _T_212_entries_perms_0_r = l3_hitVec_4 ? l3_ramDatas_4_entries_perms_0_r : l3_ramDatas_5_entries_perms_0_r; // @[ParallelMux.scala 90:77]
  wire  _T_212_entries_perms_1_d = l3_hitVec_4 ? l3_ramDatas_4_entries_perms_1_d : l3_ramDatas_5_entries_perms_1_d; // @[ParallelMux.scala 90:77]
  wire  _T_212_entries_perms_1_a = l3_hitVec_4 ? l3_ramDatas_4_entries_perms_1_a : l3_ramDatas_5_entries_perms_1_a; // @[ParallelMux.scala 90:77]
  wire  _T_212_entries_perms_1_g = l3_hitVec_4 ? l3_ramDatas_4_entries_perms_1_g : l3_ramDatas_5_entries_perms_1_g; // @[ParallelMux.scala 90:77]
  wire  _T_212_entries_perms_1_u = l3_hitVec_4 ? l3_ramDatas_4_entries_perms_1_u : l3_ramDatas_5_entries_perms_1_u; // @[ParallelMux.scala 90:77]
  wire  _T_212_entries_perms_1_x = l3_hitVec_4 ? l3_ramDatas_4_entries_perms_1_x : l3_ramDatas_5_entries_perms_1_x; // @[ParallelMux.scala 90:77]
  wire  _T_212_entries_perms_1_w = l3_hitVec_4 ? l3_ramDatas_4_entries_perms_1_w : l3_ramDatas_5_entries_perms_1_w; // @[ParallelMux.scala 90:77]
  wire  _T_212_entries_perms_1_r = l3_hitVec_4 ? l3_ramDatas_4_entries_perms_1_r : l3_ramDatas_5_entries_perms_1_r; // @[ParallelMux.scala 90:77]
  wire  _T_212_entries_perms_2_d = l3_hitVec_4 ? l3_ramDatas_4_entries_perms_2_d : l3_ramDatas_5_entries_perms_2_d; // @[ParallelMux.scala 90:77]
  wire  _T_212_entries_perms_2_a = l3_hitVec_4 ? l3_ramDatas_4_entries_perms_2_a : l3_ramDatas_5_entries_perms_2_a; // @[ParallelMux.scala 90:77]
  wire  _T_212_entries_perms_2_g = l3_hitVec_4 ? l3_ramDatas_4_entries_perms_2_g : l3_ramDatas_5_entries_perms_2_g; // @[ParallelMux.scala 90:77]
  wire  _T_212_entries_perms_2_u = l3_hitVec_4 ? l3_ramDatas_4_entries_perms_2_u : l3_ramDatas_5_entries_perms_2_u; // @[ParallelMux.scala 90:77]
  wire  _T_212_entries_perms_2_x = l3_hitVec_4 ? l3_ramDatas_4_entries_perms_2_x : l3_ramDatas_5_entries_perms_2_x; // @[ParallelMux.scala 90:77]
  wire  _T_212_entries_perms_2_w = l3_hitVec_4 ? l3_ramDatas_4_entries_perms_2_w : l3_ramDatas_5_entries_perms_2_w; // @[ParallelMux.scala 90:77]
  wire  _T_212_entries_perms_2_r = l3_hitVec_4 ? l3_ramDatas_4_entries_perms_2_r : l3_ramDatas_5_entries_perms_2_r; // @[ParallelMux.scala 90:77]
  wire  _T_212_entries_perms_3_d = l3_hitVec_4 ? l3_ramDatas_4_entries_perms_3_d : l3_ramDatas_5_entries_perms_3_d; // @[ParallelMux.scala 90:77]
  wire  _T_212_entries_perms_3_a = l3_hitVec_4 ? l3_ramDatas_4_entries_perms_3_a : l3_ramDatas_5_entries_perms_3_a; // @[ParallelMux.scala 90:77]
  wire  _T_212_entries_perms_3_g = l3_hitVec_4 ? l3_ramDatas_4_entries_perms_3_g : l3_ramDatas_5_entries_perms_3_g; // @[ParallelMux.scala 90:77]
  wire  _T_212_entries_perms_3_u = l3_hitVec_4 ? l3_ramDatas_4_entries_perms_3_u : l3_ramDatas_5_entries_perms_3_u; // @[ParallelMux.scala 90:77]
  wire  _T_212_entries_perms_3_x = l3_hitVec_4 ? l3_ramDatas_4_entries_perms_3_x : l3_ramDatas_5_entries_perms_3_x; // @[ParallelMux.scala 90:77]
  wire  _T_212_entries_perms_3_w = l3_hitVec_4 ? l3_ramDatas_4_entries_perms_3_w : l3_ramDatas_5_entries_perms_3_w; // @[ParallelMux.scala 90:77]
  wire  _T_212_entries_perms_3_r = l3_hitVec_4 ? l3_ramDatas_4_entries_perms_3_r : l3_ramDatas_5_entries_perms_3_r; // @[ParallelMux.scala 90:77]
  wire  _T_212_entries_perms_4_d = l3_hitVec_4 ? l3_ramDatas_4_entries_perms_4_d : l3_ramDatas_5_entries_perms_4_d; // @[ParallelMux.scala 90:77]
  wire  _T_212_entries_perms_4_a = l3_hitVec_4 ? l3_ramDatas_4_entries_perms_4_a : l3_ramDatas_5_entries_perms_4_a; // @[ParallelMux.scala 90:77]
  wire  _T_212_entries_perms_4_g = l3_hitVec_4 ? l3_ramDatas_4_entries_perms_4_g : l3_ramDatas_5_entries_perms_4_g; // @[ParallelMux.scala 90:77]
  wire  _T_212_entries_perms_4_u = l3_hitVec_4 ? l3_ramDatas_4_entries_perms_4_u : l3_ramDatas_5_entries_perms_4_u; // @[ParallelMux.scala 90:77]
  wire  _T_212_entries_perms_4_x = l3_hitVec_4 ? l3_ramDatas_4_entries_perms_4_x : l3_ramDatas_5_entries_perms_4_x; // @[ParallelMux.scala 90:77]
  wire  _T_212_entries_perms_4_w = l3_hitVec_4 ? l3_ramDatas_4_entries_perms_4_w : l3_ramDatas_5_entries_perms_4_w; // @[ParallelMux.scala 90:77]
  wire  _T_212_entries_perms_4_r = l3_hitVec_4 ? l3_ramDatas_4_entries_perms_4_r : l3_ramDatas_5_entries_perms_4_r; // @[ParallelMux.scala 90:77]
  wire  _T_212_entries_perms_5_d = l3_hitVec_4 ? l3_ramDatas_4_entries_perms_5_d : l3_ramDatas_5_entries_perms_5_d; // @[ParallelMux.scala 90:77]
  wire  _T_212_entries_perms_5_a = l3_hitVec_4 ? l3_ramDatas_4_entries_perms_5_a : l3_ramDatas_5_entries_perms_5_a; // @[ParallelMux.scala 90:77]
  wire  _T_212_entries_perms_5_g = l3_hitVec_4 ? l3_ramDatas_4_entries_perms_5_g : l3_ramDatas_5_entries_perms_5_g; // @[ParallelMux.scala 90:77]
  wire  _T_212_entries_perms_5_u = l3_hitVec_4 ? l3_ramDatas_4_entries_perms_5_u : l3_ramDatas_5_entries_perms_5_u; // @[ParallelMux.scala 90:77]
  wire  _T_212_entries_perms_5_x = l3_hitVec_4 ? l3_ramDatas_4_entries_perms_5_x : l3_ramDatas_5_entries_perms_5_x; // @[ParallelMux.scala 90:77]
  wire  _T_212_entries_perms_5_w = l3_hitVec_4 ? l3_ramDatas_4_entries_perms_5_w : l3_ramDatas_5_entries_perms_5_w; // @[ParallelMux.scala 90:77]
  wire  _T_212_entries_perms_5_r = l3_hitVec_4 ? l3_ramDatas_4_entries_perms_5_r : l3_ramDatas_5_entries_perms_5_r; // @[ParallelMux.scala 90:77]
  wire  _T_212_entries_perms_6_d = l3_hitVec_4 ? l3_ramDatas_4_entries_perms_6_d : l3_ramDatas_5_entries_perms_6_d; // @[ParallelMux.scala 90:77]
  wire  _T_212_entries_perms_6_a = l3_hitVec_4 ? l3_ramDatas_4_entries_perms_6_a : l3_ramDatas_5_entries_perms_6_a; // @[ParallelMux.scala 90:77]
  wire  _T_212_entries_perms_6_g = l3_hitVec_4 ? l3_ramDatas_4_entries_perms_6_g : l3_ramDatas_5_entries_perms_6_g; // @[ParallelMux.scala 90:77]
  wire  _T_212_entries_perms_6_u = l3_hitVec_4 ? l3_ramDatas_4_entries_perms_6_u : l3_ramDatas_5_entries_perms_6_u; // @[ParallelMux.scala 90:77]
  wire  _T_212_entries_perms_6_x = l3_hitVec_4 ? l3_ramDatas_4_entries_perms_6_x : l3_ramDatas_5_entries_perms_6_x; // @[ParallelMux.scala 90:77]
  wire  _T_212_entries_perms_6_w = l3_hitVec_4 ? l3_ramDatas_4_entries_perms_6_w : l3_ramDatas_5_entries_perms_6_w; // @[ParallelMux.scala 90:77]
  wire  _T_212_entries_perms_6_r = l3_hitVec_4 ? l3_ramDatas_4_entries_perms_6_r : l3_ramDatas_5_entries_perms_6_r; // @[ParallelMux.scala 90:77]
  wire  _T_212_entries_perms_7_d = l3_hitVec_4 ? l3_ramDatas_4_entries_perms_7_d : l3_ramDatas_5_entries_perms_7_d; // @[ParallelMux.scala 90:77]
  wire  _T_212_entries_perms_7_a = l3_hitVec_4 ? l3_ramDatas_4_entries_perms_7_a : l3_ramDatas_5_entries_perms_7_a; // @[ParallelMux.scala 90:77]
  wire  _T_212_entries_perms_7_g = l3_hitVec_4 ? l3_ramDatas_4_entries_perms_7_g : l3_ramDatas_5_entries_perms_7_g; // @[ParallelMux.scala 90:77]
  wire  _T_212_entries_perms_7_u = l3_hitVec_4 ? l3_ramDatas_4_entries_perms_7_u : l3_ramDatas_5_entries_perms_7_u; // @[ParallelMux.scala 90:77]
  wire  _T_212_entries_perms_7_x = l3_hitVec_4 ? l3_ramDatas_4_entries_perms_7_x : l3_ramDatas_5_entries_perms_7_x; // @[ParallelMux.scala 90:77]
  wire  _T_212_entries_perms_7_w = l3_hitVec_4 ? l3_ramDatas_4_entries_perms_7_w : l3_ramDatas_5_entries_perms_7_w; // @[ParallelMux.scala 90:77]
  wire  _T_212_entries_perms_7_r = l3_hitVec_4 ? l3_ramDatas_4_entries_perms_7_r : l3_ramDatas_5_entries_perms_7_r; // @[ParallelMux.scala 90:77]
  wire  _T_212_entries_prefetch = l3_hitVec_4 ? l3_ramDatas_4_entries_prefetch : l3_ramDatas_5_entries_prefetch; // @[ParallelMux.scala 90:77]
  wire [38:0] _T_212_ecc = l3_hitVec_4 ? l3_ramDatas_4_ecc : l3_ramDatas_5_ecc; // @[ParallelMux.scala 90:77]
  wire [21:0] _T_214_entries_tag = l3_hitVec_6 ? l3_ramDatas_6_entries_tag : l3_ramDatas_7_entries_tag; // @[ParallelMux.scala 90:77]
  wire [15:0] _T_214_entries_asid = l3_hitVec_6 ? l3_ramDatas_6_entries_asid : l3_ramDatas_7_entries_asid; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_214_entries_ppns_0 = l3_hitVec_6 ? l3_ramDatas_6_entries_ppns_0 : l3_ramDatas_7_entries_ppns_0; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_214_entries_ppns_1 = l3_hitVec_6 ? l3_ramDatas_6_entries_ppns_1 : l3_ramDatas_7_entries_ppns_1; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_214_entries_ppns_2 = l3_hitVec_6 ? l3_ramDatas_6_entries_ppns_2 : l3_ramDatas_7_entries_ppns_2; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_214_entries_ppns_3 = l3_hitVec_6 ? l3_ramDatas_6_entries_ppns_3 : l3_ramDatas_7_entries_ppns_3; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_214_entries_ppns_4 = l3_hitVec_6 ? l3_ramDatas_6_entries_ppns_4 : l3_ramDatas_7_entries_ppns_4; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_214_entries_ppns_5 = l3_hitVec_6 ? l3_ramDatas_6_entries_ppns_5 : l3_ramDatas_7_entries_ppns_5; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_214_entries_ppns_6 = l3_hitVec_6 ? l3_ramDatas_6_entries_ppns_6 : l3_ramDatas_7_entries_ppns_6; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_214_entries_ppns_7 = l3_hitVec_6 ? l3_ramDatas_6_entries_ppns_7 : l3_ramDatas_7_entries_ppns_7; // @[ParallelMux.scala 90:77]
  wire  _T_214_entries_vs_0 = l3_hitVec_6 ? l3_ramDatas_6_entries_vs_0 : l3_ramDatas_7_entries_vs_0; // @[ParallelMux.scala 90:77]
  wire  _T_214_entries_vs_1 = l3_hitVec_6 ? l3_ramDatas_6_entries_vs_1 : l3_ramDatas_7_entries_vs_1; // @[ParallelMux.scala 90:77]
  wire  _T_214_entries_vs_2 = l3_hitVec_6 ? l3_ramDatas_6_entries_vs_2 : l3_ramDatas_7_entries_vs_2; // @[ParallelMux.scala 90:77]
  wire  _T_214_entries_vs_3 = l3_hitVec_6 ? l3_ramDatas_6_entries_vs_3 : l3_ramDatas_7_entries_vs_3; // @[ParallelMux.scala 90:77]
  wire  _T_214_entries_vs_4 = l3_hitVec_6 ? l3_ramDatas_6_entries_vs_4 : l3_ramDatas_7_entries_vs_4; // @[ParallelMux.scala 90:77]
  wire  _T_214_entries_vs_5 = l3_hitVec_6 ? l3_ramDatas_6_entries_vs_5 : l3_ramDatas_7_entries_vs_5; // @[ParallelMux.scala 90:77]
  wire  _T_214_entries_vs_6 = l3_hitVec_6 ? l3_ramDatas_6_entries_vs_6 : l3_ramDatas_7_entries_vs_6; // @[ParallelMux.scala 90:77]
  wire  _T_214_entries_vs_7 = l3_hitVec_6 ? l3_ramDatas_6_entries_vs_7 : l3_ramDatas_7_entries_vs_7; // @[ParallelMux.scala 90:77]
  wire  _T_214_entries_perms_0_d = l3_hitVec_6 ? l3_ramDatas_6_entries_perms_0_d : l3_ramDatas_7_entries_perms_0_d; // @[ParallelMux.scala 90:77]
  wire  _T_214_entries_perms_0_a = l3_hitVec_6 ? l3_ramDatas_6_entries_perms_0_a : l3_ramDatas_7_entries_perms_0_a; // @[ParallelMux.scala 90:77]
  wire  _T_214_entries_perms_0_g = l3_hitVec_6 ? l3_ramDatas_6_entries_perms_0_g : l3_ramDatas_7_entries_perms_0_g; // @[ParallelMux.scala 90:77]
  wire  _T_214_entries_perms_0_u = l3_hitVec_6 ? l3_ramDatas_6_entries_perms_0_u : l3_ramDatas_7_entries_perms_0_u; // @[ParallelMux.scala 90:77]
  wire  _T_214_entries_perms_0_x = l3_hitVec_6 ? l3_ramDatas_6_entries_perms_0_x : l3_ramDatas_7_entries_perms_0_x; // @[ParallelMux.scala 90:77]
  wire  _T_214_entries_perms_0_w = l3_hitVec_6 ? l3_ramDatas_6_entries_perms_0_w : l3_ramDatas_7_entries_perms_0_w; // @[ParallelMux.scala 90:77]
  wire  _T_214_entries_perms_0_r = l3_hitVec_6 ? l3_ramDatas_6_entries_perms_0_r : l3_ramDatas_7_entries_perms_0_r; // @[ParallelMux.scala 90:77]
  wire  _T_214_entries_perms_1_d = l3_hitVec_6 ? l3_ramDatas_6_entries_perms_1_d : l3_ramDatas_7_entries_perms_1_d; // @[ParallelMux.scala 90:77]
  wire  _T_214_entries_perms_1_a = l3_hitVec_6 ? l3_ramDatas_6_entries_perms_1_a : l3_ramDatas_7_entries_perms_1_a; // @[ParallelMux.scala 90:77]
  wire  _T_214_entries_perms_1_g = l3_hitVec_6 ? l3_ramDatas_6_entries_perms_1_g : l3_ramDatas_7_entries_perms_1_g; // @[ParallelMux.scala 90:77]
  wire  _T_214_entries_perms_1_u = l3_hitVec_6 ? l3_ramDatas_6_entries_perms_1_u : l3_ramDatas_7_entries_perms_1_u; // @[ParallelMux.scala 90:77]
  wire  _T_214_entries_perms_1_x = l3_hitVec_6 ? l3_ramDatas_6_entries_perms_1_x : l3_ramDatas_7_entries_perms_1_x; // @[ParallelMux.scala 90:77]
  wire  _T_214_entries_perms_1_w = l3_hitVec_6 ? l3_ramDatas_6_entries_perms_1_w : l3_ramDatas_7_entries_perms_1_w; // @[ParallelMux.scala 90:77]
  wire  _T_214_entries_perms_1_r = l3_hitVec_6 ? l3_ramDatas_6_entries_perms_1_r : l3_ramDatas_7_entries_perms_1_r; // @[ParallelMux.scala 90:77]
  wire  _T_214_entries_perms_2_d = l3_hitVec_6 ? l3_ramDatas_6_entries_perms_2_d : l3_ramDatas_7_entries_perms_2_d; // @[ParallelMux.scala 90:77]
  wire  _T_214_entries_perms_2_a = l3_hitVec_6 ? l3_ramDatas_6_entries_perms_2_a : l3_ramDatas_7_entries_perms_2_a; // @[ParallelMux.scala 90:77]
  wire  _T_214_entries_perms_2_g = l3_hitVec_6 ? l3_ramDatas_6_entries_perms_2_g : l3_ramDatas_7_entries_perms_2_g; // @[ParallelMux.scala 90:77]
  wire  _T_214_entries_perms_2_u = l3_hitVec_6 ? l3_ramDatas_6_entries_perms_2_u : l3_ramDatas_7_entries_perms_2_u; // @[ParallelMux.scala 90:77]
  wire  _T_214_entries_perms_2_x = l3_hitVec_6 ? l3_ramDatas_6_entries_perms_2_x : l3_ramDatas_7_entries_perms_2_x; // @[ParallelMux.scala 90:77]
  wire  _T_214_entries_perms_2_w = l3_hitVec_6 ? l3_ramDatas_6_entries_perms_2_w : l3_ramDatas_7_entries_perms_2_w; // @[ParallelMux.scala 90:77]
  wire  _T_214_entries_perms_2_r = l3_hitVec_6 ? l3_ramDatas_6_entries_perms_2_r : l3_ramDatas_7_entries_perms_2_r; // @[ParallelMux.scala 90:77]
  wire  _T_214_entries_perms_3_d = l3_hitVec_6 ? l3_ramDatas_6_entries_perms_3_d : l3_ramDatas_7_entries_perms_3_d; // @[ParallelMux.scala 90:77]
  wire  _T_214_entries_perms_3_a = l3_hitVec_6 ? l3_ramDatas_6_entries_perms_3_a : l3_ramDatas_7_entries_perms_3_a; // @[ParallelMux.scala 90:77]
  wire  _T_214_entries_perms_3_g = l3_hitVec_6 ? l3_ramDatas_6_entries_perms_3_g : l3_ramDatas_7_entries_perms_3_g; // @[ParallelMux.scala 90:77]
  wire  _T_214_entries_perms_3_u = l3_hitVec_6 ? l3_ramDatas_6_entries_perms_3_u : l3_ramDatas_7_entries_perms_3_u; // @[ParallelMux.scala 90:77]
  wire  _T_214_entries_perms_3_x = l3_hitVec_6 ? l3_ramDatas_6_entries_perms_3_x : l3_ramDatas_7_entries_perms_3_x; // @[ParallelMux.scala 90:77]
  wire  _T_214_entries_perms_3_w = l3_hitVec_6 ? l3_ramDatas_6_entries_perms_3_w : l3_ramDatas_7_entries_perms_3_w; // @[ParallelMux.scala 90:77]
  wire  _T_214_entries_perms_3_r = l3_hitVec_6 ? l3_ramDatas_6_entries_perms_3_r : l3_ramDatas_7_entries_perms_3_r; // @[ParallelMux.scala 90:77]
  wire  _T_214_entries_perms_4_d = l3_hitVec_6 ? l3_ramDatas_6_entries_perms_4_d : l3_ramDatas_7_entries_perms_4_d; // @[ParallelMux.scala 90:77]
  wire  _T_214_entries_perms_4_a = l3_hitVec_6 ? l3_ramDatas_6_entries_perms_4_a : l3_ramDatas_7_entries_perms_4_a; // @[ParallelMux.scala 90:77]
  wire  _T_214_entries_perms_4_g = l3_hitVec_6 ? l3_ramDatas_6_entries_perms_4_g : l3_ramDatas_7_entries_perms_4_g; // @[ParallelMux.scala 90:77]
  wire  _T_214_entries_perms_4_u = l3_hitVec_6 ? l3_ramDatas_6_entries_perms_4_u : l3_ramDatas_7_entries_perms_4_u; // @[ParallelMux.scala 90:77]
  wire  _T_214_entries_perms_4_x = l3_hitVec_6 ? l3_ramDatas_6_entries_perms_4_x : l3_ramDatas_7_entries_perms_4_x; // @[ParallelMux.scala 90:77]
  wire  _T_214_entries_perms_4_w = l3_hitVec_6 ? l3_ramDatas_6_entries_perms_4_w : l3_ramDatas_7_entries_perms_4_w; // @[ParallelMux.scala 90:77]
  wire  _T_214_entries_perms_4_r = l3_hitVec_6 ? l3_ramDatas_6_entries_perms_4_r : l3_ramDatas_7_entries_perms_4_r; // @[ParallelMux.scala 90:77]
  wire  _T_214_entries_perms_5_d = l3_hitVec_6 ? l3_ramDatas_6_entries_perms_5_d : l3_ramDatas_7_entries_perms_5_d; // @[ParallelMux.scala 90:77]
  wire  _T_214_entries_perms_5_a = l3_hitVec_6 ? l3_ramDatas_6_entries_perms_5_a : l3_ramDatas_7_entries_perms_5_a; // @[ParallelMux.scala 90:77]
  wire  _T_214_entries_perms_5_g = l3_hitVec_6 ? l3_ramDatas_6_entries_perms_5_g : l3_ramDatas_7_entries_perms_5_g; // @[ParallelMux.scala 90:77]
  wire  _T_214_entries_perms_5_u = l3_hitVec_6 ? l3_ramDatas_6_entries_perms_5_u : l3_ramDatas_7_entries_perms_5_u; // @[ParallelMux.scala 90:77]
  wire  _T_214_entries_perms_5_x = l3_hitVec_6 ? l3_ramDatas_6_entries_perms_5_x : l3_ramDatas_7_entries_perms_5_x; // @[ParallelMux.scala 90:77]
  wire  _T_214_entries_perms_5_w = l3_hitVec_6 ? l3_ramDatas_6_entries_perms_5_w : l3_ramDatas_7_entries_perms_5_w; // @[ParallelMux.scala 90:77]
  wire  _T_214_entries_perms_5_r = l3_hitVec_6 ? l3_ramDatas_6_entries_perms_5_r : l3_ramDatas_7_entries_perms_5_r; // @[ParallelMux.scala 90:77]
  wire  _T_214_entries_perms_6_d = l3_hitVec_6 ? l3_ramDatas_6_entries_perms_6_d : l3_ramDatas_7_entries_perms_6_d; // @[ParallelMux.scala 90:77]
  wire  _T_214_entries_perms_6_a = l3_hitVec_6 ? l3_ramDatas_6_entries_perms_6_a : l3_ramDatas_7_entries_perms_6_a; // @[ParallelMux.scala 90:77]
  wire  _T_214_entries_perms_6_g = l3_hitVec_6 ? l3_ramDatas_6_entries_perms_6_g : l3_ramDatas_7_entries_perms_6_g; // @[ParallelMux.scala 90:77]
  wire  _T_214_entries_perms_6_u = l3_hitVec_6 ? l3_ramDatas_6_entries_perms_6_u : l3_ramDatas_7_entries_perms_6_u; // @[ParallelMux.scala 90:77]
  wire  _T_214_entries_perms_6_x = l3_hitVec_6 ? l3_ramDatas_6_entries_perms_6_x : l3_ramDatas_7_entries_perms_6_x; // @[ParallelMux.scala 90:77]
  wire  _T_214_entries_perms_6_w = l3_hitVec_6 ? l3_ramDatas_6_entries_perms_6_w : l3_ramDatas_7_entries_perms_6_w; // @[ParallelMux.scala 90:77]
  wire  _T_214_entries_perms_6_r = l3_hitVec_6 ? l3_ramDatas_6_entries_perms_6_r : l3_ramDatas_7_entries_perms_6_r; // @[ParallelMux.scala 90:77]
  wire  _T_214_entries_perms_7_d = l3_hitVec_6 ? l3_ramDatas_6_entries_perms_7_d : l3_ramDatas_7_entries_perms_7_d; // @[ParallelMux.scala 90:77]
  wire  _T_214_entries_perms_7_a = l3_hitVec_6 ? l3_ramDatas_6_entries_perms_7_a : l3_ramDatas_7_entries_perms_7_a; // @[ParallelMux.scala 90:77]
  wire  _T_214_entries_perms_7_g = l3_hitVec_6 ? l3_ramDatas_6_entries_perms_7_g : l3_ramDatas_7_entries_perms_7_g; // @[ParallelMux.scala 90:77]
  wire  _T_214_entries_perms_7_u = l3_hitVec_6 ? l3_ramDatas_6_entries_perms_7_u : l3_ramDatas_7_entries_perms_7_u; // @[ParallelMux.scala 90:77]
  wire  _T_214_entries_perms_7_x = l3_hitVec_6 ? l3_ramDatas_6_entries_perms_7_x : l3_ramDatas_7_entries_perms_7_x; // @[ParallelMux.scala 90:77]
  wire  _T_214_entries_perms_7_w = l3_hitVec_6 ? l3_ramDatas_6_entries_perms_7_w : l3_ramDatas_7_entries_perms_7_w; // @[ParallelMux.scala 90:77]
  wire  _T_214_entries_perms_7_r = l3_hitVec_6 ? l3_ramDatas_6_entries_perms_7_r : l3_ramDatas_7_entries_perms_7_r; // @[ParallelMux.scala 90:77]
  wire  _T_214_entries_prefetch = l3_hitVec_6 ? l3_ramDatas_6_entries_prefetch : l3_ramDatas_7_entries_prefetch; // @[ParallelMux.scala 90:77]
  wire [38:0] _T_214_ecc = l3_hitVec_6 ? l3_ramDatas_6_ecc : l3_ramDatas_7_ecc; // @[ParallelMux.scala 90:77]
  wire  _T_215 = l3_hitVec_4 | l3_hitVec_5 | (l3_hitVec_6 | l3_hitVec_7); // @[ParallelMux.scala 90:65]
  wire [21:0] _T_216_entries_tag = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_tag : _T_214_entries_tag; // @[ParallelMux.scala 90:77]
  wire [15:0] _T_216_entries_asid = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_asid : _T_214_entries_asid; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_216_entries_ppns_0 = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_ppns_0 : _T_214_entries_ppns_0; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_216_entries_ppns_1 = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_ppns_1 : _T_214_entries_ppns_1; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_216_entries_ppns_2 = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_ppns_2 : _T_214_entries_ppns_2; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_216_entries_ppns_3 = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_ppns_3 : _T_214_entries_ppns_3; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_216_entries_ppns_4 = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_ppns_4 : _T_214_entries_ppns_4; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_216_entries_ppns_5 = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_ppns_5 : _T_214_entries_ppns_5; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_216_entries_ppns_6 = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_ppns_6 : _T_214_entries_ppns_6; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_216_entries_ppns_7 = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_ppns_7 : _T_214_entries_ppns_7; // @[ParallelMux.scala 90:77]
  wire  _T_216_entries_vs_0 = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_vs_0 : _T_214_entries_vs_0; // @[ParallelMux.scala 90:77]
  wire  _T_216_entries_vs_1 = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_vs_1 : _T_214_entries_vs_1; // @[ParallelMux.scala 90:77]
  wire  _T_216_entries_vs_2 = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_vs_2 : _T_214_entries_vs_2; // @[ParallelMux.scala 90:77]
  wire  _T_216_entries_vs_3 = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_vs_3 : _T_214_entries_vs_3; // @[ParallelMux.scala 90:77]
  wire  _T_216_entries_vs_4 = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_vs_4 : _T_214_entries_vs_4; // @[ParallelMux.scala 90:77]
  wire  _T_216_entries_vs_5 = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_vs_5 : _T_214_entries_vs_5; // @[ParallelMux.scala 90:77]
  wire  _T_216_entries_vs_6 = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_vs_6 : _T_214_entries_vs_6; // @[ParallelMux.scala 90:77]
  wire  _T_216_entries_vs_7 = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_vs_7 : _T_214_entries_vs_7; // @[ParallelMux.scala 90:77]
  wire  _T_216_entries_perms_0_d = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_perms_0_d : _T_214_entries_perms_0_d; // @[ParallelMux.scala 90:77]
  wire  _T_216_entries_perms_0_a = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_perms_0_a : _T_214_entries_perms_0_a; // @[ParallelMux.scala 90:77]
  wire  _T_216_entries_perms_0_g = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_perms_0_g : _T_214_entries_perms_0_g; // @[ParallelMux.scala 90:77]
  wire  _T_216_entries_perms_0_u = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_perms_0_u : _T_214_entries_perms_0_u; // @[ParallelMux.scala 90:77]
  wire  _T_216_entries_perms_0_x = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_perms_0_x : _T_214_entries_perms_0_x; // @[ParallelMux.scala 90:77]
  wire  _T_216_entries_perms_0_w = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_perms_0_w : _T_214_entries_perms_0_w; // @[ParallelMux.scala 90:77]
  wire  _T_216_entries_perms_0_r = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_perms_0_r : _T_214_entries_perms_0_r; // @[ParallelMux.scala 90:77]
  wire  _T_216_entries_perms_1_d = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_perms_1_d : _T_214_entries_perms_1_d; // @[ParallelMux.scala 90:77]
  wire  _T_216_entries_perms_1_a = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_perms_1_a : _T_214_entries_perms_1_a; // @[ParallelMux.scala 90:77]
  wire  _T_216_entries_perms_1_g = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_perms_1_g : _T_214_entries_perms_1_g; // @[ParallelMux.scala 90:77]
  wire  _T_216_entries_perms_1_u = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_perms_1_u : _T_214_entries_perms_1_u; // @[ParallelMux.scala 90:77]
  wire  _T_216_entries_perms_1_x = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_perms_1_x : _T_214_entries_perms_1_x; // @[ParallelMux.scala 90:77]
  wire  _T_216_entries_perms_1_w = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_perms_1_w : _T_214_entries_perms_1_w; // @[ParallelMux.scala 90:77]
  wire  _T_216_entries_perms_1_r = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_perms_1_r : _T_214_entries_perms_1_r; // @[ParallelMux.scala 90:77]
  wire  _T_216_entries_perms_2_d = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_perms_2_d : _T_214_entries_perms_2_d; // @[ParallelMux.scala 90:77]
  wire  _T_216_entries_perms_2_a = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_perms_2_a : _T_214_entries_perms_2_a; // @[ParallelMux.scala 90:77]
  wire  _T_216_entries_perms_2_g = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_perms_2_g : _T_214_entries_perms_2_g; // @[ParallelMux.scala 90:77]
  wire  _T_216_entries_perms_2_u = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_perms_2_u : _T_214_entries_perms_2_u; // @[ParallelMux.scala 90:77]
  wire  _T_216_entries_perms_2_x = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_perms_2_x : _T_214_entries_perms_2_x; // @[ParallelMux.scala 90:77]
  wire  _T_216_entries_perms_2_w = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_perms_2_w : _T_214_entries_perms_2_w; // @[ParallelMux.scala 90:77]
  wire  _T_216_entries_perms_2_r = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_perms_2_r : _T_214_entries_perms_2_r; // @[ParallelMux.scala 90:77]
  wire  _T_216_entries_perms_3_d = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_perms_3_d : _T_214_entries_perms_3_d; // @[ParallelMux.scala 90:77]
  wire  _T_216_entries_perms_3_a = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_perms_3_a : _T_214_entries_perms_3_a; // @[ParallelMux.scala 90:77]
  wire  _T_216_entries_perms_3_g = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_perms_3_g : _T_214_entries_perms_3_g; // @[ParallelMux.scala 90:77]
  wire  _T_216_entries_perms_3_u = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_perms_3_u : _T_214_entries_perms_3_u; // @[ParallelMux.scala 90:77]
  wire  _T_216_entries_perms_3_x = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_perms_3_x : _T_214_entries_perms_3_x; // @[ParallelMux.scala 90:77]
  wire  _T_216_entries_perms_3_w = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_perms_3_w : _T_214_entries_perms_3_w; // @[ParallelMux.scala 90:77]
  wire  _T_216_entries_perms_3_r = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_perms_3_r : _T_214_entries_perms_3_r; // @[ParallelMux.scala 90:77]
  wire  _T_216_entries_perms_4_d = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_perms_4_d : _T_214_entries_perms_4_d; // @[ParallelMux.scala 90:77]
  wire  _T_216_entries_perms_4_a = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_perms_4_a : _T_214_entries_perms_4_a; // @[ParallelMux.scala 90:77]
  wire  _T_216_entries_perms_4_g = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_perms_4_g : _T_214_entries_perms_4_g; // @[ParallelMux.scala 90:77]
  wire  _T_216_entries_perms_4_u = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_perms_4_u : _T_214_entries_perms_4_u; // @[ParallelMux.scala 90:77]
  wire  _T_216_entries_perms_4_x = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_perms_4_x : _T_214_entries_perms_4_x; // @[ParallelMux.scala 90:77]
  wire  _T_216_entries_perms_4_w = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_perms_4_w : _T_214_entries_perms_4_w; // @[ParallelMux.scala 90:77]
  wire  _T_216_entries_perms_4_r = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_perms_4_r : _T_214_entries_perms_4_r; // @[ParallelMux.scala 90:77]
  wire  _T_216_entries_perms_5_d = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_perms_5_d : _T_214_entries_perms_5_d; // @[ParallelMux.scala 90:77]
  wire  _T_216_entries_perms_5_a = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_perms_5_a : _T_214_entries_perms_5_a; // @[ParallelMux.scala 90:77]
  wire  _T_216_entries_perms_5_g = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_perms_5_g : _T_214_entries_perms_5_g; // @[ParallelMux.scala 90:77]
  wire  _T_216_entries_perms_5_u = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_perms_5_u : _T_214_entries_perms_5_u; // @[ParallelMux.scala 90:77]
  wire  _T_216_entries_perms_5_x = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_perms_5_x : _T_214_entries_perms_5_x; // @[ParallelMux.scala 90:77]
  wire  _T_216_entries_perms_5_w = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_perms_5_w : _T_214_entries_perms_5_w; // @[ParallelMux.scala 90:77]
  wire  _T_216_entries_perms_5_r = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_perms_5_r : _T_214_entries_perms_5_r; // @[ParallelMux.scala 90:77]
  wire  _T_216_entries_perms_6_d = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_perms_6_d : _T_214_entries_perms_6_d; // @[ParallelMux.scala 90:77]
  wire  _T_216_entries_perms_6_a = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_perms_6_a : _T_214_entries_perms_6_a; // @[ParallelMux.scala 90:77]
  wire  _T_216_entries_perms_6_g = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_perms_6_g : _T_214_entries_perms_6_g; // @[ParallelMux.scala 90:77]
  wire  _T_216_entries_perms_6_u = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_perms_6_u : _T_214_entries_perms_6_u; // @[ParallelMux.scala 90:77]
  wire  _T_216_entries_perms_6_x = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_perms_6_x : _T_214_entries_perms_6_x; // @[ParallelMux.scala 90:77]
  wire  _T_216_entries_perms_6_w = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_perms_6_w : _T_214_entries_perms_6_w; // @[ParallelMux.scala 90:77]
  wire  _T_216_entries_perms_6_r = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_perms_6_r : _T_214_entries_perms_6_r; // @[ParallelMux.scala 90:77]
  wire  _T_216_entries_perms_7_d = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_perms_7_d : _T_214_entries_perms_7_d; // @[ParallelMux.scala 90:77]
  wire  _T_216_entries_perms_7_a = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_perms_7_a : _T_214_entries_perms_7_a; // @[ParallelMux.scala 90:77]
  wire  _T_216_entries_perms_7_g = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_perms_7_g : _T_214_entries_perms_7_g; // @[ParallelMux.scala 90:77]
  wire  _T_216_entries_perms_7_u = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_perms_7_u : _T_214_entries_perms_7_u; // @[ParallelMux.scala 90:77]
  wire  _T_216_entries_perms_7_x = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_perms_7_x : _T_214_entries_perms_7_x; // @[ParallelMux.scala 90:77]
  wire  _T_216_entries_perms_7_w = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_perms_7_w : _T_214_entries_perms_7_w; // @[ParallelMux.scala 90:77]
  wire  _T_216_entries_perms_7_r = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_perms_7_r : _T_214_entries_perms_7_r; // @[ParallelMux.scala 90:77]
  wire  _T_216_entries_prefetch = l3_hitVec_4 | l3_hitVec_5 ? _T_212_entries_prefetch : _T_214_entries_prefetch; // @[ParallelMux.scala 90:77]
  wire [38:0] _T_216_ecc = l3_hitVec_4 | l3_hitVec_5 ? _T_212_ecc : _T_214_ecc; // @[ParallelMux.scala 90:77]
  wire  _T_217 = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) | (l3_hitVec_4 | l3_hitVec_5 | (l3_hitVec_6 |
    l3_hitVec_7)); // @[ParallelMux.scala 90:65]
  wire [21:0] _T_218_entries_tag = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_tag :
    _T_216_entries_tag; // @[ParallelMux.scala 90:77]
  wire [15:0] _T_218_entries_asid = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_asid :
    _T_216_entries_asid; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_218_entries_ppns_0 = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_ppns_0 :
    _T_216_entries_ppns_0; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_218_entries_ppns_1 = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_ppns_1 :
    _T_216_entries_ppns_1; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_218_entries_ppns_2 = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_ppns_2 :
    _T_216_entries_ppns_2; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_218_entries_ppns_3 = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_ppns_3 :
    _T_216_entries_ppns_3; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_218_entries_ppns_4 = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_ppns_4 :
    _T_216_entries_ppns_4; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_218_entries_ppns_5 = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_ppns_5 :
    _T_216_entries_ppns_5; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_218_entries_ppns_6 = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_ppns_6 :
    _T_216_entries_ppns_6; // @[ParallelMux.scala 90:77]
  wire [23:0] _T_218_entries_ppns_7 = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_ppns_7 :
    _T_216_entries_ppns_7; // @[ParallelMux.scala 90:77]
  wire  _T_218_entries_vs_0 = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_vs_0 :
    _T_216_entries_vs_0; // @[ParallelMux.scala 90:77]
  wire  _T_218_entries_vs_1 = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_vs_1 :
    _T_216_entries_vs_1; // @[ParallelMux.scala 90:77]
  wire  _T_218_entries_vs_2 = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_vs_2 :
    _T_216_entries_vs_2; // @[ParallelMux.scala 90:77]
  wire  _T_218_entries_vs_3 = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_vs_3 :
    _T_216_entries_vs_3; // @[ParallelMux.scala 90:77]
  wire  _T_218_entries_vs_4 = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_vs_4 :
    _T_216_entries_vs_4; // @[ParallelMux.scala 90:77]
  wire  _T_218_entries_vs_5 = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_vs_5 :
    _T_216_entries_vs_5; // @[ParallelMux.scala 90:77]
  wire  _T_218_entries_vs_6 = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_vs_6 :
    _T_216_entries_vs_6; // @[ParallelMux.scala 90:77]
  wire  _T_218_entries_vs_7 = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_vs_7 :
    _T_216_entries_vs_7; // @[ParallelMux.scala 90:77]
  wire  _T_218_entries_perms_0_d = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_perms_0_d :
    _T_216_entries_perms_0_d; // @[ParallelMux.scala 90:77]
  wire  _T_218_entries_perms_0_a = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_perms_0_a :
    _T_216_entries_perms_0_a; // @[ParallelMux.scala 90:77]
  wire  _T_218_entries_perms_0_g = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_perms_0_g :
    _T_216_entries_perms_0_g; // @[ParallelMux.scala 90:77]
  wire  _T_218_entries_perms_0_u = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_perms_0_u :
    _T_216_entries_perms_0_u; // @[ParallelMux.scala 90:77]
  wire  _T_218_entries_perms_0_x = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_perms_0_x :
    _T_216_entries_perms_0_x; // @[ParallelMux.scala 90:77]
  wire  _T_218_entries_perms_0_w = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_perms_0_w :
    _T_216_entries_perms_0_w; // @[ParallelMux.scala 90:77]
  wire  _T_218_entries_perms_0_r = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_perms_0_r :
    _T_216_entries_perms_0_r; // @[ParallelMux.scala 90:77]
  wire  _T_218_entries_perms_1_d = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_perms_1_d :
    _T_216_entries_perms_1_d; // @[ParallelMux.scala 90:77]
  wire  _T_218_entries_perms_1_a = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_perms_1_a :
    _T_216_entries_perms_1_a; // @[ParallelMux.scala 90:77]
  wire  _T_218_entries_perms_1_g = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_perms_1_g :
    _T_216_entries_perms_1_g; // @[ParallelMux.scala 90:77]
  wire  _T_218_entries_perms_1_u = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_perms_1_u :
    _T_216_entries_perms_1_u; // @[ParallelMux.scala 90:77]
  wire  _T_218_entries_perms_1_x = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_perms_1_x :
    _T_216_entries_perms_1_x; // @[ParallelMux.scala 90:77]
  wire  _T_218_entries_perms_1_w = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_perms_1_w :
    _T_216_entries_perms_1_w; // @[ParallelMux.scala 90:77]
  wire  _T_218_entries_perms_1_r = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_perms_1_r :
    _T_216_entries_perms_1_r; // @[ParallelMux.scala 90:77]
  wire  _T_218_entries_perms_2_d = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_perms_2_d :
    _T_216_entries_perms_2_d; // @[ParallelMux.scala 90:77]
  wire  _T_218_entries_perms_2_a = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_perms_2_a :
    _T_216_entries_perms_2_a; // @[ParallelMux.scala 90:77]
  wire  _T_218_entries_perms_2_g = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_perms_2_g :
    _T_216_entries_perms_2_g; // @[ParallelMux.scala 90:77]
  wire  _T_218_entries_perms_2_u = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_perms_2_u :
    _T_216_entries_perms_2_u; // @[ParallelMux.scala 90:77]
  wire  _T_218_entries_perms_2_x = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_perms_2_x :
    _T_216_entries_perms_2_x; // @[ParallelMux.scala 90:77]
  wire  _T_218_entries_perms_2_w = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_perms_2_w :
    _T_216_entries_perms_2_w; // @[ParallelMux.scala 90:77]
  wire  _T_218_entries_perms_2_r = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_perms_2_r :
    _T_216_entries_perms_2_r; // @[ParallelMux.scala 90:77]
  wire  _T_218_entries_perms_3_d = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_perms_3_d :
    _T_216_entries_perms_3_d; // @[ParallelMux.scala 90:77]
  wire  _T_218_entries_perms_3_a = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_perms_3_a :
    _T_216_entries_perms_3_a; // @[ParallelMux.scala 90:77]
  wire  _T_218_entries_perms_3_g = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_perms_3_g :
    _T_216_entries_perms_3_g; // @[ParallelMux.scala 90:77]
  wire  _T_218_entries_perms_3_u = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_perms_3_u :
    _T_216_entries_perms_3_u; // @[ParallelMux.scala 90:77]
  wire  _T_218_entries_perms_3_x = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_perms_3_x :
    _T_216_entries_perms_3_x; // @[ParallelMux.scala 90:77]
  wire  _T_218_entries_perms_3_w = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_perms_3_w :
    _T_216_entries_perms_3_w; // @[ParallelMux.scala 90:77]
  wire  _T_218_entries_perms_3_r = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_perms_3_r :
    _T_216_entries_perms_3_r; // @[ParallelMux.scala 90:77]
  wire  _T_218_entries_perms_4_d = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_perms_4_d :
    _T_216_entries_perms_4_d; // @[ParallelMux.scala 90:77]
  wire  _T_218_entries_perms_4_a = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_perms_4_a :
    _T_216_entries_perms_4_a; // @[ParallelMux.scala 90:77]
  wire  _T_218_entries_perms_4_g = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_perms_4_g :
    _T_216_entries_perms_4_g; // @[ParallelMux.scala 90:77]
  wire  _T_218_entries_perms_4_u = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_perms_4_u :
    _T_216_entries_perms_4_u; // @[ParallelMux.scala 90:77]
  wire  _T_218_entries_perms_4_x = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_perms_4_x :
    _T_216_entries_perms_4_x; // @[ParallelMux.scala 90:77]
  wire  _T_218_entries_perms_4_w = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_perms_4_w :
    _T_216_entries_perms_4_w; // @[ParallelMux.scala 90:77]
  wire  _T_218_entries_perms_4_r = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_perms_4_r :
    _T_216_entries_perms_4_r; // @[ParallelMux.scala 90:77]
  wire  _T_218_entries_perms_5_d = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_perms_5_d :
    _T_216_entries_perms_5_d; // @[ParallelMux.scala 90:77]
  wire  _T_218_entries_perms_5_a = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_perms_5_a :
    _T_216_entries_perms_5_a; // @[ParallelMux.scala 90:77]
  wire  _T_218_entries_perms_5_g = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_perms_5_g :
    _T_216_entries_perms_5_g; // @[ParallelMux.scala 90:77]
  wire  _T_218_entries_perms_5_u = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_perms_5_u :
    _T_216_entries_perms_5_u; // @[ParallelMux.scala 90:77]
  wire  _T_218_entries_perms_5_x = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_perms_5_x :
    _T_216_entries_perms_5_x; // @[ParallelMux.scala 90:77]
  wire  _T_218_entries_perms_5_w = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_perms_5_w :
    _T_216_entries_perms_5_w; // @[ParallelMux.scala 90:77]
  wire  _T_218_entries_perms_5_r = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_perms_5_r :
    _T_216_entries_perms_5_r; // @[ParallelMux.scala 90:77]
  wire  _T_218_entries_perms_6_d = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_perms_6_d :
    _T_216_entries_perms_6_d; // @[ParallelMux.scala 90:77]
  wire  _T_218_entries_perms_6_a = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_perms_6_a :
    _T_216_entries_perms_6_a; // @[ParallelMux.scala 90:77]
  wire  _T_218_entries_perms_6_g = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_perms_6_g :
    _T_216_entries_perms_6_g; // @[ParallelMux.scala 90:77]
  wire  _T_218_entries_perms_6_u = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_perms_6_u :
    _T_216_entries_perms_6_u; // @[ParallelMux.scala 90:77]
  wire  _T_218_entries_perms_6_x = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_perms_6_x :
    _T_216_entries_perms_6_x; // @[ParallelMux.scala 90:77]
  wire  _T_218_entries_perms_6_w = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_perms_6_w :
    _T_216_entries_perms_6_w; // @[ParallelMux.scala 90:77]
  wire  _T_218_entries_perms_6_r = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_perms_6_r :
    _T_216_entries_perms_6_r; // @[ParallelMux.scala 90:77]
  wire  _T_218_entries_perms_7_d = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_perms_7_d :
    _T_216_entries_perms_7_d; // @[ParallelMux.scala 90:77]
  wire  _T_218_entries_perms_7_a = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_perms_7_a :
    _T_216_entries_perms_7_a; // @[ParallelMux.scala 90:77]
  wire  _T_218_entries_perms_7_g = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_perms_7_g :
    _T_216_entries_perms_7_g; // @[ParallelMux.scala 90:77]
  wire  _T_218_entries_perms_7_u = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_perms_7_u :
    _T_216_entries_perms_7_u; // @[ParallelMux.scala 90:77]
  wire  _T_218_entries_perms_7_x = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_perms_7_x :
    _T_216_entries_perms_7_x; // @[ParallelMux.scala 90:77]
  wire  _T_218_entries_perms_7_w = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_perms_7_w :
    _T_216_entries_perms_7_w; // @[ParallelMux.scala 90:77]
  wire  _T_218_entries_perms_7_r = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_perms_7_r :
    _T_216_entries_perms_7_r; // @[ParallelMux.scala 90:77]
  wire  check_res_l3_pre = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_entries_prefetch :
    _T_216_entries_prefetch; // @[ParallelMux.scala 90:77]
  wire [38:0] _T_218_ecc = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_210_ecc : _T_216_ecc; // @[ParallelMux.scala 90:77]
  wire [2:0] _T_227 = l3_hitVec_0 ? 3'h0 : 3'h1; // @[ParallelMux.scala 90:77]
  wire [2:0] _T_229 = l3_hitVec_2 ? 3'h2 : 3'h3; // @[ParallelMux.scala 90:77]
  wire [2:0] _T_231 = l3_hitVec_0 | l3_hitVec_1 ? _T_227 : _T_229; // @[ParallelMux.scala 90:77]
  wire [2:0] _T_233 = l3_hitVec_4 ? 3'h4 : 3'h5; // @[ParallelMux.scala 90:77]
  wire [2:0] _T_235 = l3_hitVec_6 ? 3'h6 : 3'h7; // @[ParallelMux.scala 90:77]
  wire [2:0] _T_237 = l3_hitVec_4 | l3_hitVec_5 ? _T_233 : _T_235; // @[ParallelMux.scala 90:77]
  wire [2:0] l3_hitWay = l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3) ? _T_231 : _T_237; // @[ParallelMux.scala 90:77]
  wire [8:0] data_lo_lo_lo_1 = {_T_218_entries_perms_1_r,_T_218_entries_perms_0_d,_T_218_entries_perms_0_a,
    _T_218_entries_perms_0_g,_T_218_entries_perms_0_u,_T_218_entries_perms_0_x,_T_218_entries_perms_0_w,
    _T_218_entries_perms_0_r,check_res_l3_pre}; // @[MMUBundle.scala 717:30]
  wire [17:0] data_lo_lo_1 = {_T_218_entries_perms_2_x,_T_218_entries_perms_2_w,_T_218_entries_perms_2_r,
    _T_218_entries_perms_1_d,_T_218_entries_perms_1_a,_T_218_entries_perms_1_g,_T_218_entries_perms_1_u,
    _T_218_entries_perms_1_x,_T_218_entries_perms_1_w,data_lo_lo_lo_1}; // @[MMUBundle.scala 717:30]
  wire [9:0] data_lo_hi_hi_1 = {_T_218_entries_perms_5_r,_T_218_entries_perms_4_d,_T_218_entries_perms_4_a,
    _T_218_entries_perms_4_g,_T_218_entries_perms_4_u,_T_218_entries_perms_4_x,_T_218_entries_perms_4_w,
    _T_218_entries_perms_4_r,_T_218_entries_perms_3_d,_T_218_entries_perms_3_a}; // @[MMUBundle.scala 717:30]
  wire [18:0] data_lo_hi_1 = {data_lo_hi_hi_1,_T_218_entries_perms_3_g,_T_218_entries_perms_3_u,_T_218_entries_perms_3_x
    ,_T_218_entries_perms_3_w,_T_218_entries_perms_3_r,_T_218_entries_perms_2_d,_T_218_entries_perms_2_a,
    _T_218_entries_perms_2_g,_T_218_entries_perms_2_u}; // @[MMUBundle.scala 717:30]
  wire [9:0] data_hi_lo_hi_1 = {_T_218_entries_perms_7_a,_T_218_entries_perms_7_g,_T_218_entries_perms_7_u,
    _T_218_entries_perms_7_x,_T_218_entries_perms_7_w,_T_218_entries_perms_7_r,_T_218_entries_perms_6_d,
    _T_218_entries_perms_6_a,_T_218_entries_perms_6_g,_T_218_entries_perms_6_u}; // @[MMUBundle.scala 717:30]
  wire [18:0] data_hi_lo_1 = {data_hi_lo_hi_1,_T_218_entries_perms_6_x,_T_218_entries_perms_6_w,_T_218_entries_perms_6_r
    ,_T_218_entries_perms_5_d,_T_218_entries_perms_5_a,_T_218_entries_perms_5_g,_T_218_entries_perms_5_u,
    _T_218_entries_perms_5_x,_T_218_entries_perms_5_w}; // @[MMUBundle.scala 717:30]
  wire [229:0] data_hi_hi_hi_1 = {_T_218_entries_tag,_T_218_entries_asid,_T_218_entries_ppns_7,_T_218_entries_ppns_6,
    _T_218_entries_ppns_5,_T_218_entries_ppns_4,_T_218_entries_ppns_3,_T_218_entries_ppns_2,_T_218_entries_ppns_1,
    _T_218_entries_ppns_0}; // @[MMUBundle.scala 717:30]
  wire [238:0] data_hi_hi_1 = {data_hi_hi_hi_1,_T_218_entries_vs_7,_T_218_entries_vs_6,_T_218_entries_vs_5,
    _T_218_entries_vs_4,_T_218_entries_vs_3,_T_218_entries_vs_2,_T_218_entries_vs_1,_T_218_entries_vs_0,
    _T_218_entries_perms_7_d}; // @[MMUBundle.scala 717:30]
  wire [294:0] data_4 = {data_hi_hi_1,data_hi_lo_1,data_lo_hi_1,data_lo_lo_1}; // @[MMUBundle.scala 717:30]
  wire [71:0] _res_0_T_7 = {_T_218_ecc[7:0],data_4[63:0]}; // @[Cat.scala 31:58]
  wire [70:0] _res_0_syndromeUInt_T_14 = 71'h1ab55555556aaad5b & _res_0_T_7[70:0]; // @[ECC.scala 156:66]
  wire [70:0] _res_0_syndromeUInt_T_16 = 71'h2cd9999999b33366d & _res_0_T_7[70:0]; // @[ECC.scala 156:66]
  wire [70:0] _res_0_syndromeUInt_T_18 = 71'h4f1e1e1e1e3c3c78e & _res_0_T_7[70:0]; // @[ECC.scala 156:66]
  wire [70:0] _res_0_syndromeUInt_T_20 = 71'h801fe01fe03fc07f0 & _res_0_T_7[70:0]; // @[ECC.scala 156:66]
  wire [70:0] _res_0_syndromeUInt_T_22 = 71'h1001fffe0003fff800 & _res_0_T_7[70:0]; // @[ECC.scala 156:66]
  wire [70:0] _res_0_syndromeUInt_T_24 = 71'h2001fffffffc000000 & _res_0_T_7[70:0]; // @[ECC.scala 156:66]
  wire [70:0] _res_0_syndromeUInt_T_26 = 71'h40fe00000000000000 & _res_0_T_7[70:0]; // @[ECC.scala 156:66]
  wire [6:0] res_0_syndromeUInt_1 = {^_res_0_syndromeUInt_T_26,^_res_0_syndromeUInt_T_24,^_res_0_syndromeUInt_T_22,^
    _res_0_syndromeUInt_T_20,^_res_0_syndromeUInt_T_18,^_res_0_syndromeUInt_T_16,^_res_0_syndromeUInt_T_14}; // @[ECC.scala 156:78]
  wire  res_0_correctable_1 = |res_0_syndromeUInt_1; // @[ECC.scala 163:36]
  wire  res_0_uncorrectable_4 = ^_res_0_T_7; // @[ECC.scala 87:27]
  wire  res_0_uncorrectable_5 = ~res_0_uncorrectable_4 & res_0_correctable_1; // @[ECC.scala 195:47]
  wire  res_1_0 = res_0_uncorrectable_4 | res_0_uncorrectable_5; // @[ECC.scala 31:27]
  wire [71:0] _res_1_T_7 = {_T_218_ecc[15:8],data_4[127:64]}; // @[Cat.scala 31:58]
  wire [70:0] _res_1_syndromeUInt_T_14 = 71'h1ab55555556aaad5b & _res_1_T_7[70:0]; // @[ECC.scala 156:66]
  wire [70:0] _res_1_syndromeUInt_T_16 = 71'h2cd9999999b33366d & _res_1_T_7[70:0]; // @[ECC.scala 156:66]
  wire [70:0] _res_1_syndromeUInt_T_18 = 71'h4f1e1e1e1e3c3c78e & _res_1_T_7[70:0]; // @[ECC.scala 156:66]
  wire [70:0] _res_1_syndromeUInt_T_20 = 71'h801fe01fe03fc07f0 & _res_1_T_7[70:0]; // @[ECC.scala 156:66]
  wire [70:0] _res_1_syndromeUInt_T_22 = 71'h1001fffe0003fff800 & _res_1_T_7[70:0]; // @[ECC.scala 156:66]
  wire [70:0] _res_1_syndromeUInt_T_24 = 71'h2001fffffffc000000 & _res_1_T_7[70:0]; // @[ECC.scala 156:66]
  wire [70:0] _res_1_syndromeUInt_T_26 = 71'h40fe00000000000000 & _res_1_T_7[70:0]; // @[ECC.scala 156:66]
  wire [6:0] res_1_syndromeUInt_1 = {^_res_1_syndromeUInt_T_26,^_res_1_syndromeUInt_T_24,^_res_1_syndromeUInt_T_22,^
    _res_1_syndromeUInt_T_20,^_res_1_syndromeUInt_T_18,^_res_1_syndromeUInt_T_16,^_res_1_syndromeUInt_T_14}; // @[ECC.scala 156:78]
  wire  res_1_correctable_1 = |res_1_syndromeUInt_1; // @[ECC.scala 163:36]
  wire  res_1_uncorrectable_4 = ^_res_1_T_7; // @[ECC.scala 87:27]
  wire  res_1_uncorrectable_5 = ~res_1_uncorrectable_4 & res_1_correctable_1; // @[ECC.scala 195:47]
  wire  res_1_1 = res_1_uncorrectable_4 | res_1_uncorrectable_5; // @[ECC.scala 31:27]
  wire [71:0] _res_2_T_7 = {_T_218_ecc[23:16],data_4[191:128]}; // @[Cat.scala 31:58]
  wire [70:0] _res_2_syndromeUInt_T_14 = 71'h1ab55555556aaad5b & _res_2_T_7[70:0]; // @[ECC.scala 156:66]
  wire [70:0] _res_2_syndromeUInt_T_16 = 71'h2cd9999999b33366d & _res_2_T_7[70:0]; // @[ECC.scala 156:66]
  wire [70:0] _res_2_syndromeUInt_T_18 = 71'h4f1e1e1e1e3c3c78e & _res_2_T_7[70:0]; // @[ECC.scala 156:66]
  wire [70:0] _res_2_syndromeUInt_T_20 = 71'h801fe01fe03fc07f0 & _res_2_T_7[70:0]; // @[ECC.scala 156:66]
  wire [70:0] _res_2_syndromeUInt_T_22 = 71'h1001fffe0003fff800 & _res_2_T_7[70:0]; // @[ECC.scala 156:66]
  wire [70:0] _res_2_syndromeUInt_T_24 = 71'h2001fffffffc000000 & _res_2_T_7[70:0]; // @[ECC.scala 156:66]
  wire [70:0] _res_2_syndromeUInt_T_26 = 71'h40fe00000000000000 & _res_2_T_7[70:0]; // @[ECC.scala 156:66]
  wire [6:0] res_2_syndromeUInt_1 = {^_res_2_syndromeUInt_T_26,^_res_2_syndromeUInt_T_24,^_res_2_syndromeUInt_T_22,^
    _res_2_syndromeUInt_T_20,^_res_2_syndromeUInt_T_18,^_res_2_syndromeUInt_T_16,^_res_2_syndromeUInt_T_14}; // @[ECC.scala 156:78]
  wire  res_2_correctable_1 = |res_2_syndromeUInt_1; // @[ECC.scala 163:36]
  wire  res_2_uncorrectable_4 = ^_res_2_T_7; // @[ECC.scala 87:27]
  wire  res_2_uncorrectable_5 = ~res_2_uncorrectable_4 & res_2_correctable_1; // @[ECC.scala 195:47]
  wire  res_1_2 = res_2_uncorrectable_4 | res_2_uncorrectable_5; // @[ECC.scala 31:27]
  wire [71:0] _res_3_T_7 = {_T_218_ecc[31:24],data_4[255:192]}; // @[Cat.scala 31:58]
  wire [70:0] _res_3_syndromeUInt_T_12 = 71'h1ab55555556aaad5b & _res_3_T_7[70:0]; // @[ECC.scala 156:66]
  wire [70:0] _res_3_syndromeUInt_T_14 = 71'h2cd9999999b33366d & _res_3_T_7[70:0]; // @[ECC.scala 156:66]
  wire [70:0] _res_3_syndromeUInt_T_16 = 71'h4f1e1e1e1e3c3c78e & _res_3_T_7[70:0]; // @[ECC.scala 156:66]
  wire [70:0] _res_3_syndromeUInt_T_18 = 71'h801fe01fe03fc07f0 & _res_3_T_7[70:0]; // @[ECC.scala 156:66]
  wire [70:0] _res_3_syndromeUInt_T_20 = 71'h1001fffe0003fff800 & _res_3_T_7[70:0]; // @[ECC.scala 156:66]
  wire [70:0] _res_3_syndromeUInt_T_22 = 71'h2001fffffffc000000 & _res_3_T_7[70:0]; // @[ECC.scala 156:66]
  wire [70:0] _res_3_syndromeUInt_T_24 = 71'h40fe00000000000000 & _res_3_T_7[70:0]; // @[ECC.scala 156:66]
  wire [6:0] res_3_syndromeUInt_1 = {^_res_3_syndromeUInt_T_24,^_res_3_syndromeUInt_T_22,^_res_3_syndromeUInt_T_20,^
    _res_3_syndromeUInt_T_18,^_res_3_syndromeUInt_T_16,^_res_3_syndromeUInt_T_14,^_res_3_syndromeUInt_T_12}; // @[ECC.scala 156:78]
  wire  res_3_correctable_1 = |res_3_syndromeUInt_1; // @[ECC.scala 163:36]
  wire  res_3_uncorrectable_4 = ^_res_3_T_7; // @[ECC.scala 87:27]
  wire  res_3_uncorrectable_5 = ~res_3_uncorrectable_4 & res_3_correctable_1; // @[ECC.scala 195:47]
  wire  res_1_3 = res_3_uncorrectable_4 | res_3_uncorrectable_5; // @[ECC.scala 31:27]
  wire [45:0] _res_4_T_2 = {_T_218_ecc[38:32],data_4[294:256]}; // @[Cat.scala 31:58]
  wire [44:0] _res_4_syndromeUInt_T = 45'hd556aaad5b & _res_4_T_2[44:0]; // @[ECC.scala 156:66]
  wire [44:0] _res_4_syndromeUInt_T_2 = 45'h1199b33366d & _res_4_T_2[44:0]; // @[ECC.scala 156:66]
  wire [44:0] _res_4_syndromeUInt_T_4 = 45'h261e3c3c78e & _res_4_T_2[44:0]; // @[ECC.scala 156:66]
  wire [44:0] _res_4_syndromeUInt_T_6 = 45'h47e03fc07f0 & _res_4_T_2[44:0]; // @[ECC.scala 156:66]
  wire [44:0] _res_4_syndromeUInt_T_8 = 45'h80003fff800 & _res_4_T_2[44:0]; // @[ECC.scala 156:66]
  wire [44:0] _res_4_syndromeUInt_T_10 = 45'h107ffc000000 & _res_4_T_2[44:0]; // @[ECC.scala 156:66]
  wire [5:0] res_4_syndromeUInt = {^_res_4_syndromeUInt_T_10,^_res_4_syndromeUInt_T_8,^_res_4_syndromeUInt_T_6,^
    _res_4_syndromeUInt_T_4,^_res_4_syndromeUInt_T_2,^_res_4_syndromeUInt_T}; // @[ECC.scala 156:78]
  wire  res_4_correctable = |res_4_syndromeUInt; // @[ECC.scala 163:36]
  wire  res_4_uncorrectable_1 = ^_res_4_T_2; // @[ECC.scala 87:27]
  wire  res_4_uncorrectable_2 = ~res_4_uncorrectable_1 & res_4_correctable; // @[ECC.scala 195:47]
  wire  res_1_4 = res_4_uncorrectable_1 | res_4_uncorrectable_2; // @[ECC.scala 31:27]
  wire [4:0] _T_239 = {res_1_0,res_1_1,res_1_2,res_1_3,res_1_4}; // @[Cat.scala 31:58]
  wire  l3eccError = |_T_239; // @[MMUBundle.scala 727:14]
  wire  state_vec_set_left_older_1 = ~l3_hitWay[2]; // @[Replacement.scala 196:33]
  wire [6:0] _GEN_1507 = 2'h1 == data_1_req_info_vpn[4:3] ? state_vec_1_1 : state_vec_1_0; // @[package.scala 154:{13,13}]
  wire [6:0] _GEN_1508 = 2'h2 == data_1_req_info_vpn[4:3] ? state_vec_1_2 : _GEN_1507; // @[package.scala 154:{13,13}]
  wire [6:0] _GEN_1509 = 2'h3 == data_1_req_info_vpn[4:3] ? state_vec_1_3 : _GEN_1508; // @[package.scala 154:{13,13}]
  wire [2:0] state_vec_left_subtree_state_1 = _GEN_1509[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_right_subtree_state_1 = _GEN_1509[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_set_left_older_2 = ~l3_hitWay[1]; // @[Replacement.scala 196:33]
  wire  state_vec_left_subtree_state_2 = state_vec_left_subtree_state_1[1]; // @[package.scala 154:13]
  wire  state_vec_right_subtree_state_2 = state_vec_left_subtree_state_1[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_T_12 = ~l3_hitWay[0]; // @[Replacement.scala 218:7]
  wire  _state_vec_T_13 = state_vec_set_left_older_2 ? state_vec_left_subtree_state_2 : _state_vec_T_12; // @[Replacement.scala 203:16]
  wire  _state_vec_T_17 = state_vec_set_left_older_2 ? _state_vec_T_12 : state_vec_right_subtree_state_2; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_T_18 = {state_vec_set_left_older_2,_state_vec_T_13,_state_vec_T_17}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_T_19 = state_vec_set_left_older_1 ? state_vec_left_subtree_state_1 : _state_vec_T_18; // @[Replacement.scala 203:16]
  wire  state_vec_left_subtree_state_3 = state_vec_right_subtree_state_1[1]; // @[package.scala 154:13]
  wire  state_vec_right_subtree_state_3 = state_vec_right_subtree_state_1[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_T_24 = state_vec_set_left_older_2 ? state_vec_left_subtree_state_3 : _state_vec_T_12; // @[Replacement.scala 203:16]
  wire  _state_vec_T_28 = state_vec_set_left_older_2 ? _state_vec_T_12 : state_vec_right_subtree_state_3; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_T_29 = {state_vec_set_left_older_2,_state_vec_T_24,_state_vec_T_28}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_T_30 = state_vec_set_left_older_1 ? _state_vec_T_29 : state_vec_right_subtree_state_1; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_T_31 = {state_vec_set_left_older_1,_state_vec_T_19,_state_vec_T_30}; // @[Cat.scala 31:58]
  wire [6:0] _GEN_1510 = 2'h0 == data_1_req_info_vpn[4:3] ? _state_vec_T_31 : state_vec_1_0; // @[Replacement.scala 305:17 308:{20,20}]
  wire [6:0] _GEN_1511 = 2'h1 == data_1_req_info_vpn[4:3] ? _state_vec_T_31 : state_vec_1_1; // @[Replacement.scala 305:17 308:{20,20}]
  wire [6:0] _GEN_1512 = 2'h2 == data_1_req_info_vpn[4:3] ? _state_vec_T_31 : state_vec_1_2; // @[Replacement.scala 305:17 308:{20,20}]
  wire [6:0] _GEN_1513 = 2'h3 == data_1_req_info_vpn[4:3] ? _state_vec_T_31 : state_vec_1_3; // @[Replacement.scala 305:17 308:{20,20}]
  wire [6:0] _GEN_1514 = _T_217 & stageCheck_valid_1cycle ? _GEN_1510 : state_vec_1_0; // @[PageTableCache.scala 330:43 Replacement.scala 305:17]
  wire [6:0] _GEN_1515 = _T_217 & stageCheck_valid_1cycle ? _GEN_1511 : state_vec_1_1; // @[PageTableCache.scala 330:43 Replacement.scala 305:17]
  wire [6:0] _GEN_1516 = _T_217 & stageCheck_valid_1cycle ? _GEN_1512 : state_vec_1_2; // @[PageTableCache.scala 330:43 Replacement.scala 305:17]
  wire [6:0] _GEN_1517 = _T_217 & stageCheck_valid_1cycle ? _GEN_1513 : state_vec_1_3; // @[PageTableCache.scala 330:43 Replacement.scala 305:17]
  reg  state_reg_3; // @[Replacement.scala 168:70]
  wire  asid_hit_20 = sp_0_asid == io_csr_dup_0_satp_asid; // @[MMUBundle.scala 578:59]
  wire  hit0 = sp_0_tag[17:9] == io_req_bits_req_info_vpn[26:18]; // @[MMUBundle.scala 587:52]
  wire  hit1 = sp_0_tag[8:0] == io_req_bits_req_info_vpn[17:9]; // @[MMUBundle.scala 588:66]
  wire  _T_256 = sp_0_level == 2'h0 ? hit0 : hit0 & hit1; // @[MMUBundle.scala 590:22]
  wire  _T_257 = asid_hit_20 & _T_256; // @[MMUBundle.scala 590:16]
  wire  sp_hitVecT_0 = _T_257 & spv[0]; // @[PageTableCache.scala 353:115]
  wire  asid_hit_21 = sp_1_asid == io_csr_dup_0_satp_asid; // @[MMUBundle.scala 578:59]
  wire  hit0_1 = sp_1_tag[17:9] == io_req_bits_req_info_vpn[26:18]; // @[MMUBundle.scala 587:52]
  wire  hit1_1 = sp_1_tag[8:0] == io_req_bits_req_info_vpn[17:9]; // @[MMUBundle.scala 588:66]
  wire  _T_262 = sp_1_level == 2'h0 ? hit0_1 : hit0_1 & hit1_1; // @[MMUBundle.scala 590:22]
  wire  _T_263 = asid_hit_21 & _T_262; // @[MMUBundle.scala 590:16]
  wire  sp_hitVecT_1 = _T_263 & spv[1]; // @[PageTableCache.scala 353:115]
  reg  r_13; // @[Reg.scala 16:16]
  reg  r_14; // @[Reg.scala 16:16]
  wire  _T_268 = r_13 | r_14; // @[ParallelMux.scala 90:65]
  wire [1:0] _T_272 = {r_14,r_13}; // @[Cat.scala 31:58]
  wire  state_reg_touch_way_sized_1 = _T_272[1]; // @[CircuitMath.scala 30:8]
  wire  _state_reg_T_10 = ~state_reg_touch_way_sized_1; // @[Replacement.scala 218:7]
  reg  spHit; // @[Reg.scala 16:16]
  reg [23:0] spHitData_ppn; // @[Reg.scala 16:16]
  reg  spHitData_perm_d; // @[Reg.scala 16:16]
  reg  spHitData_perm_a; // @[Reg.scala 16:16]
  reg  spHitData_perm_g; // @[Reg.scala 16:16]
  reg  spHitData_perm_u; // @[Reg.scala 16:16]
  reg  spHitData_perm_x; // @[Reg.scala 16:16]
  reg  spHitData_perm_w; // @[Reg.scala 16:16]
  reg  spHitData_perm_r; // @[Reg.scala 16:16]
  reg [1:0] spHitData_level; // @[Reg.scala 16:16]
  reg  spPre; // @[Reg.scala 16:16]
  reg  spValid; // @[Reg.scala 16:16]
  wire  check_res_l2_hit = _T_117 & ~l2eccError; // @[PageTableCache.scala 47:21]
  wire [23:0] _GEN_1538 = 3'h1 == data_1_req_info_vpn[11:9] ? _T_118_entries_ppns_1 : _T_118_entries_ppns_0; // @[PageTableCache.scala 49:{14,14}]
  wire [23:0] _GEN_1539 = 3'h2 == data_1_req_info_vpn[11:9] ? _T_118_entries_ppns_2 : _GEN_1538; // @[PageTableCache.scala 49:{14,14}]
  wire [23:0] _GEN_1540 = 3'h3 == data_1_req_info_vpn[11:9] ? _T_118_entries_ppns_3 : _GEN_1539; // @[PageTableCache.scala 49:{14,14}]
  wire [23:0] _GEN_1541 = 3'h4 == data_1_req_info_vpn[11:9] ? _T_118_entries_ppns_4 : _GEN_1540; // @[PageTableCache.scala 49:{14,14}]
  wire  check_res_l2_ecc = l2eccError & _T_117; // @[PageTableCache.scala 51:21]
  wire  check_res_l3_hit = _T_217 & ~l3eccError; // @[PageTableCache.scala 47:21]
  wire [23:0] _GEN_1546 = 3'h1 == data_1_req_info_vpn[2:0] ? _T_218_entries_ppns_1 : _T_218_entries_ppns_0; // @[PageTableCache.scala 49:{14,14}]
  wire [23:0] _GEN_1547 = 3'h2 == data_1_req_info_vpn[2:0] ? _T_218_entries_ppns_2 : _GEN_1546; // @[PageTableCache.scala 49:{14,14}]
  wire [23:0] _GEN_1548 = 3'h3 == data_1_req_info_vpn[2:0] ? _T_218_entries_ppns_3 : _GEN_1547; // @[PageTableCache.scala 49:{14,14}]
  wire [23:0] _GEN_1549 = 3'h4 == data_1_req_info_vpn[2:0] ? _T_218_entries_ppns_4 : _GEN_1548; // @[PageTableCache.scala 49:{14,14}]
  wire  _GEN_1554 = 3'h1 == data_1_req_info_vpn[2:0] ? _T_218_entries_perms_1_d : _T_218_entries_perms_0_d; // @[PageTableCache.scala 50:{15,15}]
  wire  _GEN_1555 = 3'h2 == data_1_req_info_vpn[2:0] ? _T_218_entries_perms_2_d : _GEN_1554; // @[PageTableCache.scala 50:{15,15}]
  wire  _GEN_1556 = 3'h3 == data_1_req_info_vpn[2:0] ? _T_218_entries_perms_3_d : _GEN_1555; // @[PageTableCache.scala 50:{15,15}]
  wire  _GEN_1557 = 3'h4 == data_1_req_info_vpn[2:0] ? _T_218_entries_perms_4_d : _GEN_1556; // @[PageTableCache.scala 50:{15,15}]
  wire  _GEN_1562 = 3'h1 == data_1_req_info_vpn[2:0] ? _T_218_entries_perms_1_a : _T_218_entries_perms_0_a; // @[PageTableCache.scala 50:{15,15}]
  wire  _GEN_1563 = 3'h2 == data_1_req_info_vpn[2:0] ? _T_218_entries_perms_2_a : _GEN_1562; // @[PageTableCache.scala 50:{15,15}]
  wire  _GEN_1564 = 3'h3 == data_1_req_info_vpn[2:0] ? _T_218_entries_perms_3_a : _GEN_1563; // @[PageTableCache.scala 50:{15,15}]
  wire  _GEN_1565 = 3'h4 == data_1_req_info_vpn[2:0] ? _T_218_entries_perms_4_a : _GEN_1564; // @[PageTableCache.scala 50:{15,15}]
  wire  _GEN_1570 = 3'h1 == data_1_req_info_vpn[2:0] ? _T_218_entries_perms_1_g : _T_218_entries_perms_0_g; // @[PageTableCache.scala 50:{15,15}]
  wire  _GEN_1571 = 3'h2 == data_1_req_info_vpn[2:0] ? _T_218_entries_perms_2_g : _GEN_1570; // @[PageTableCache.scala 50:{15,15}]
  wire  _GEN_1572 = 3'h3 == data_1_req_info_vpn[2:0] ? _T_218_entries_perms_3_g : _GEN_1571; // @[PageTableCache.scala 50:{15,15}]
  wire  _GEN_1573 = 3'h4 == data_1_req_info_vpn[2:0] ? _T_218_entries_perms_4_g : _GEN_1572; // @[PageTableCache.scala 50:{15,15}]
  wire  _GEN_1578 = 3'h1 == data_1_req_info_vpn[2:0] ? _T_218_entries_perms_1_u : _T_218_entries_perms_0_u; // @[PageTableCache.scala 50:{15,15}]
  wire  _GEN_1579 = 3'h2 == data_1_req_info_vpn[2:0] ? _T_218_entries_perms_2_u : _GEN_1578; // @[PageTableCache.scala 50:{15,15}]
  wire  _GEN_1580 = 3'h3 == data_1_req_info_vpn[2:0] ? _T_218_entries_perms_3_u : _GEN_1579; // @[PageTableCache.scala 50:{15,15}]
  wire  _GEN_1581 = 3'h4 == data_1_req_info_vpn[2:0] ? _T_218_entries_perms_4_u : _GEN_1580; // @[PageTableCache.scala 50:{15,15}]
  wire  _GEN_1586 = 3'h1 == data_1_req_info_vpn[2:0] ? _T_218_entries_perms_1_x : _T_218_entries_perms_0_x; // @[PageTableCache.scala 50:{15,15}]
  wire  _GEN_1587 = 3'h2 == data_1_req_info_vpn[2:0] ? _T_218_entries_perms_2_x : _GEN_1586; // @[PageTableCache.scala 50:{15,15}]
  wire  _GEN_1588 = 3'h3 == data_1_req_info_vpn[2:0] ? _T_218_entries_perms_3_x : _GEN_1587; // @[PageTableCache.scala 50:{15,15}]
  wire  _GEN_1589 = 3'h4 == data_1_req_info_vpn[2:0] ? _T_218_entries_perms_4_x : _GEN_1588; // @[PageTableCache.scala 50:{15,15}]
  wire  _GEN_1594 = 3'h1 == data_1_req_info_vpn[2:0] ? _T_218_entries_perms_1_w : _T_218_entries_perms_0_w; // @[PageTableCache.scala 50:{15,15}]
  wire  _GEN_1595 = 3'h2 == data_1_req_info_vpn[2:0] ? _T_218_entries_perms_2_w : _GEN_1594; // @[PageTableCache.scala 50:{15,15}]
  wire  _GEN_1596 = 3'h3 == data_1_req_info_vpn[2:0] ? _T_218_entries_perms_3_w : _GEN_1595; // @[PageTableCache.scala 50:{15,15}]
  wire  _GEN_1597 = 3'h4 == data_1_req_info_vpn[2:0] ? _T_218_entries_perms_4_w : _GEN_1596; // @[PageTableCache.scala 50:{15,15}]
  wire  _GEN_1602 = 3'h1 == data_1_req_info_vpn[2:0] ? _T_218_entries_perms_1_r : _T_218_entries_perms_0_r; // @[PageTableCache.scala 50:{15,15}]
  wire  _GEN_1603 = 3'h2 == data_1_req_info_vpn[2:0] ? _T_218_entries_perms_2_r : _GEN_1602; // @[PageTableCache.scala 50:{15,15}]
  wire  _GEN_1604 = 3'h3 == data_1_req_info_vpn[2:0] ? _T_218_entries_perms_3_r : _GEN_1603; // @[PageTableCache.scala 50:{15,15}]
  wire  _GEN_1605 = 3'h4 == data_1_req_info_vpn[2:0] ? _T_218_entries_perms_4_r : _GEN_1604; // @[PageTableCache.scala 50:{15,15}]
  wire  check_res_l3_ecc = l3eccError & _T_217; // @[PageTableCache.scala 51:21]
  wire  _GEN_1610 = 3'h1 == data_1_req_info_vpn[2:0] ? _T_218_entries_vs_1 : _T_218_entries_vs_0; // @[PageTableCache.scala 53:{12,12}]
  wire  _GEN_1611 = 3'h2 == data_1_req_info_vpn[2:0] ? _T_218_entries_vs_2 : _GEN_1610; // @[PageTableCache.scala 53:{12,12}]
  wire  _GEN_1612 = 3'h3 == data_1_req_info_vpn[2:0] ? _T_218_entries_vs_3 : _GEN_1611; // @[PageTableCache.scala 53:{12,12}]
  wire  _GEN_1613 = 3'h4 == data_1_req_info_vpn[2:0] ? _T_218_entries_vs_4 : _GEN_1612; // @[PageTableCache.scala 53:{12,12}]
  reg  resp_res_l1_hit; // @[PageTableCache.scala 383:21]
  reg [23:0] resp_res_l1_ppn; // @[PageTableCache.scala 383:21]
  reg  resp_res_l2_hit; // @[PageTableCache.scala 383:21]
  reg [23:0] resp_res_l2_ppn; // @[PageTableCache.scala 383:21]
  reg  resp_res_l2_ecc; // @[PageTableCache.scala 383:21]
  reg  resp_res_l3_hit; // @[PageTableCache.scala 383:21]
  reg  resp_res_l3_pre; // @[PageTableCache.scala 383:21]
  reg [23:0] resp_res_l3_ppn; // @[PageTableCache.scala 383:21]
  reg  resp_res_l3_perm_d; // @[PageTableCache.scala 383:21]
  reg  resp_res_l3_perm_a; // @[PageTableCache.scala 383:21]
  reg  resp_res_l3_perm_g; // @[PageTableCache.scala 383:21]
  reg  resp_res_l3_perm_u; // @[PageTableCache.scala 383:21]
  reg  resp_res_l3_perm_x; // @[PageTableCache.scala 383:21]
  reg  resp_res_l3_perm_w; // @[PageTableCache.scala 383:21]
  reg  resp_res_l3_perm_r; // @[PageTableCache.scala 383:21]
  reg  resp_res_l3_ecc; // @[PageTableCache.scala 383:21]
  reg  resp_res_l3_v; // @[PageTableCache.scala 383:21]
  reg  resp_res_sp_hit; // @[PageTableCache.scala 383:21]
  reg  resp_res_sp_pre; // @[PageTableCache.scala 383:21]
  reg [23:0] resp_res_sp_ppn; // @[PageTableCache.scala 383:21]
  reg  resp_res_sp_perm_d; // @[PageTableCache.scala 383:21]
  reg  resp_res_sp_perm_a; // @[PageTableCache.scala 383:21]
  reg  resp_res_sp_perm_g; // @[PageTableCache.scala 383:21]
  reg  resp_res_sp_perm_u; // @[PageTableCache.scala 383:21]
  reg  resp_res_sp_perm_x; // @[PageTableCache.scala 383:21]
  reg  resp_res_sp_perm_w; // @[PageTableCache.scala 383:21]
  reg  resp_res_sp_perm_r; // @[PageTableCache.scala 383:21]
  reg [1:0] resp_res_sp_level; // @[PageTableCache.scala 383:21]
  reg  resp_res_sp_v; // @[PageTableCache.scala 383:21]
  wire  _bypassed_0_T_4 = io_refill_bits_req_info_dup_0_vpn[26:21] == data_2_req_info_vpn[26:21]; // @[PageTableCache.scala 221:44]
  wire  _bypassed_0_T_5 = io_refill_valid & 2'h0 == io_refill_bits_level_dup_0 & _bypassed_0_T_4; // @[PageTableCache.scala 225:66]
  reg  bypassed_0_valid; // @[Hold.scala 54:24]
  wire  _GEN_1669 = bypassed_0_valid ? 1'h0 : bypassed_0_valid; // @[Hold.scala 55:18 54:24 55:26]
  wire  _bypassed_0_T_7 = bypassed_0_valid | io_refill_valid; // @[PageTableCache.scala 391:52]
  reg  bypassed_0_valid_1; // @[MMUBundle.scala 796:24]
  wire  _GEN_1672 = _bypassed_0_T_5 | bypassed_0_valid_1; // @[MMUBundle.scala 797:19 796:24 797:27]
  wire  _bypassed_0_T_8 = bypassed_0_valid_1 | _bypassed_0_T_5; // @[MMUBundle.scala 800:11]
  wire  bypassed_0 = data_2_bypassed_0 | _bypassed_0_T_8; // @[PageTableCache.scala 389:47]
  wire  _bypassed_1_T_4 = io_refill_bits_req_info_dup_0_vpn[26:12] == data_2_req_info_vpn[26:12]; // @[PageTableCache.scala 221:44]
  wire  _bypassed_1_T_5 = io_refill_valid & 2'h1 == io_refill_bits_level_dup_0 & _bypassed_1_T_4; // @[PageTableCache.scala 225:66]
  reg  bypassed_1_valid; // @[Hold.scala 54:24]
  wire  _GEN_1675 = bypassed_1_valid ? 1'h0 : bypassed_1_valid; // @[Hold.scala 55:18 54:24 55:26]
  wire  _bypassed_1_T_7 = bypassed_1_valid | io_refill_valid; // @[PageTableCache.scala 391:52]
  reg  bypassed_1_valid_1; // @[MMUBundle.scala 796:24]
  wire  _GEN_1678 = _bypassed_1_T_5 | bypassed_1_valid_1; // @[MMUBundle.scala 797:19 796:24 797:27]
  wire  _bypassed_1_T_8 = bypassed_1_valid_1 | _bypassed_1_T_5; // @[MMUBundle.scala 800:11]
  wire  bypassed_1 = data_2_bypassed_1 | _bypassed_1_T_8; // @[PageTableCache.scala 389:47]
  wire  _bypassed_2_T_4 = io_refill_bits_req_info_dup_0_vpn[26:3] == data_2_req_info_vpn[26:3]; // @[PageTableCache.scala 221:44]
  wire  _bypassed_2_T_5 = io_refill_valid & 2'h2 == io_refill_bits_level_dup_0 & _bypassed_2_T_4; // @[PageTableCache.scala 225:66]
  reg  bypassed_2_valid; // @[Hold.scala 54:24]
  wire  _GEN_1681 = bypassed_2_valid ? 1'h0 : bypassed_2_valid; // @[Hold.scala 55:18 54:24 55:26]
  wire  _bypassed_2_T_7 = bypassed_2_valid | io_refill_valid; // @[PageTableCache.scala 391:52]
  reg  bypassed_2_valid_1; // @[MMUBundle.scala 796:24]
  wire  _GEN_1684 = _bypassed_2_T_5 | bypassed_2_valid_1; // @[MMUBundle.scala 797:19 796:24 797:27]
  wire  _bypassed_2_T_8 = bypassed_2_valid_1 | _bypassed_2_T_5; // @[MMUBundle.scala 800:11]
  wire  bypassed_2 = data_2_bypassed_2 | _bypassed_2_T_8; // @[PageTableCache.scala 389:47]
  wire  memPtes_0_perm_v = io_refill_bits_ptes[0]; // @[PageTableCache.scala 430:109]
  wire  memPtes_0_perm_r = io_refill_bits_ptes[1]; // @[PageTableCache.scala 430:109]
  wire  memPtes_0_perm_w = io_refill_bits_ptes[2]; // @[PageTableCache.scala 430:109]
  wire  memPtes_0_perm_x = io_refill_bits_ptes[3]; // @[PageTableCache.scala 430:109]
  wire  memPtes_0_perm_u = io_refill_bits_ptes[4]; // @[PageTableCache.scala 430:109]
  wire  memPtes_0_perm_g = io_refill_bits_ptes[5]; // @[PageTableCache.scala 430:109]
  wire  memPtes_0_perm_a = io_refill_bits_ptes[6]; // @[PageTableCache.scala 430:109]
  wire  memPtes_0_perm_d = io_refill_bits_ptes[7]; // @[PageTableCache.scala 430:109]
  wire [23:0] memPtes_0_ppn = io_refill_bits_ptes[33:10]; // @[PageTableCache.scala 430:109]
  wire  memPtes_1_perm_v = io_refill_bits_ptes[64]; // @[PageTableCache.scala 430:109]
  wire  memPtes_1_perm_r = io_refill_bits_ptes[65]; // @[PageTableCache.scala 430:109]
  wire  memPtes_1_perm_w = io_refill_bits_ptes[66]; // @[PageTableCache.scala 430:109]
  wire  memPtes_1_perm_x = io_refill_bits_ptes[67]; // @[PageTableCache.scala 430:109]
  wire  memPtes_1_perm_u = io_refill_bits_ptes[68]; // @[PageTableCache.scala 430:109]
  wire  memPtes_1_perm_g = io_refill_bits_ptes[69]; // @[PageTableCache.scala 430:109]
  wire  memPtes_1_perm_a = io_refill_bits_ptes[70]; // @[PageTableCache.scala 430:109]
  wire  memPtes_1_perm_d = io_refill_bits_ptes[71]; // @[PageTableCache.scala 430:109]
  wire [23:0] memPtes_1_ppn = io_refill_bits_ptes[97:74]; // @[PageTableCache.scala 430:109]
  wire  memPtes_2_perm_v = io_refill_bits_ptes[128]; // @[PageTableCache.scala 430:109]
  wire  memPtes_2_perm_r = io_refill_bits_ptes[129]; // @[PageTableCache.scala 430:109]
  wire  memPtes_2_perm_w = io_refill_bits_ptes[130]; // @[PageTableCache.scala 430:109]
  wire  memPtes_2_perm_x = io_refill_bits_ptes[131]; // @[PageTableCache.scala 430:109]
  wire  memPtes_2_perm_u = io_refill_bits_ptes[132]; // @[PageTableCache.scala 430:109]
  wire  memPtes_2_perm_g = io_refill_bits_ptes[133]; // @[PageTableCache.scala 430:109]
  wire  memPtes_2_perm_a = io_refill_bits_ptes[134]; // @[PageTableCache.scala 430:109]
  wire  memPtes_2_perm_d = io_refill_bits_ptes[135]; // @[PageTableCache.scala 430:109]
  wire [23:0] memPtes_2_ppn = io_refill_bits_ptes[161:138]; // @[PageTableCache.scala 430:109]
  wire  memPtes_3_perm_v = io_refill_bits_ptes[192]; // @[PageTableCache.scala 430:109]
  wire  memPtes_3_perm_r = io_refill_bits_ptes[193]; // @[PageTableCache.scala 430:109]
  wire  memPtes_3_perm_w = io_refill_bits_ptes[194]; // @[PageTableCache.scala 430:109]
  wire  memPtes_3_perm_x = io_refill_bits_ptes[195]; // @[PageTableCache.scala 430:109]
  wire  memPtes_3_perm_u = io_refill_bits_ptes[196]; // @[PageTableCache.scala 430:109]
  wire  memPtes_3_perm_g = io_refill_bits_ptes[197]; // @[PageTableCache.scala 430:109]
  wire  memPtes_3_perm_a = io_refill_bits_ptes[198]; // @[PageTableCache.scala 430:109]
  wire  memPtes_3_perm_d = io_refill_bits_ptes[199]; // @[PageTableCache.scala 430:109]
  wire [23:0] memPtes_3_ppn = io_refill_bits_ptes[225:202]; // @[PageTableCache.scala 430:109]
  wire  memPtes_4_perm_v = io_refill_bits_ptes[256]; // @[PageTableCache.scala 430:109]
  wire  memPtes_4_perm_r = io_refill_bits_ptes[257]; // @[PageTableCache.scala 430:109]
  wire  memPtes_4_perm_w = io_refill_bits_ptes[258]; // @[PageTableCache.scala 430:109]
  wire  memPtes_4_perm_x = io_refill_bits_ptes[259]; // @[PageTableCache.scala 430:109]
  wire  memPtes_4_perm_u = io_refill_bits_ptes[260]; // @[PageTableCache.scala 430:109]
  wire  memPtes_4_perm_g = io_refill_bits_ptes[261]; // @[PageTableCache.scala 430:109]
  wire  memPtes_4_perm_a = io_refill_bits_ptes[262]; // @[PageTableCache.scala 430:109]
  wire  memPtes_4_perm_d = io_refill_bits_ptes[263]; // @[PageTableCache.scala 430:109]
  wire [23:0] memPtes_4_ppn = io_refill_bits_ptes[289:266]; // @[PageTableCache.scala 430:109]
  wire  memPtes_5_perm_v = io_refill_bits_ptes[320]; // @[PageTableCache.scala 430:109]
  wire  memPtes_5_perm_r = io_refill_bits_ptes[321]; // @[PageTableCache.scala 430:109]
  wire  memPtes_5_perm_w = io_refill_bits_ptes[322]; // @[PageTableCache.scala 430:109]
  wire  memPtes_5_perm_x = io_refill_bits_ptes[323]; // @[PageTableCache.scala 430:109]
  wire  memPtes_5_perm_u = io_refill_bits_ptes[324]; // @[PageTableCache.scala 430:109]
  wire  memPtes_5_perm_g = io_refill_bits_ptes[325]; // @[PageTableCache.scala 430:109]
  wire  memPtes_5_perm_a = io_refill_bits_ptes[326]; // @[PageTableCache.scala 430:109]
  wire  memPtes_5_perm_d = io_refill_bits_ptes[327]; // @[PageTableCache.scala 430:109]
  wire [23:0] memPtes_5_ppn = io_refill_bits_ptes[353:330]; // @[PageTableCache.scala 430:109]
  wire  memPtes_6_perm_v = io_refill_bits_ptes[384]; // @[PageTableCache.scala 430:109]
  wire  memPtes_6_perm_r = io_refill_bits_ptes[385]; // @[PageTableCache.scala 430:109]
  wire  memPtes_6_perm_w = io_refill_bits_ptes[386]; // @[PageTableCache.scala 430:109]
  wire  memPtes_6_perm_x = io_refill_bits_ptes[387]; // @[PageTableCache.scala 430:109]
  wire  memPtes_6_perm_u = io_refill_bits_ptes[388]; // @[PageTableCache.scala 430:109]
  wire  memPtes_6_perm_g = io_refill_bits_ptes[389]; // @[PageTableCache.scala 430:109]
  wire  memPtes_6_perm_a = io_refill_bits_ptes[390]; // @[PageTableCache.scala 430:109]
  wire  memPtes_6_perm_d = io_refill_bits_ptes[391]; // @[PageTableCache.scala 430:109]
  wire [23:0] memPtes_6_ppn = io_refill_bits_ptes[417:394]; // @[PageTableCache.scala 430:109]
  wire  memPtes_7_perm_v = io_refill_bits_ptes[448]; // @[PageTableCache.scala 430:109]
  wire  memPtes_7_perm_r = io_refill_bits_ptes[449]; // @[PageTableCache.scala 430:109]
  wire  memPtes_7_perm_w = io_refill_bits_ptes[450]; // @[PageTableCache.scala 430:109]
  wire  memPtes_7_perm_x = io_refill_bits_ptes[451]; // @[PageTableCache.scala 430:109]
  wire  memPtes_7_perm_u = io_refill_bits_ptes[452]; // @[PageTableCache.scala 430:109]
  wire  memPtes_7_perm_g = io_refill_bits_ptes[453]; // @[PageTableCache.scala 430:109]
  wire  memPtes_7_perm_a = io_refill_bits_ptes[454]; // @[PageTableCache.scala 430:109]
  wire  memPtes_7_perm_d = io_refill_bits_ptes[455]; // @[PageTableCache.scala 430:109]
  wire [23:0] memPtes_7_ppn = io_refill_bits_ptes[481:458]; // @[PageTableCache.scala 430:109]
  wire  memPte_0_perm_v = io_refill_bits_sel_pte_dup_0[0]; // @[PageTableCache.scala 432:46]
  wire  memPte_0_perm_r = io_refill_bits_sel_pte_dup_0[1]; // @[PageTableCache.scala 432:46]
  wire  memPte_0_perm_w = io_refill_bits_sel_pte_dup_0[2]; // @[PageTableCache.scala 432:46]
  wire  memPte_0_perm_x = io_refill_bits_sel_pte_dup_0[3]; // @[PageTableCache.scala 432:46]
  wire  memPte_0_perm_u = io_refill_bits_sel_pte_dup_0[4]; // @[PageTableCache.scala 432:46]
  wire  memPte_0_perm_g = io_refill_bits_sel_pte_dup_0[5]; // @[PageTableCache.scala 432:46]
  wire  memPte_0_perm_a = io_refill_bits_sel_pte_dup_0[6]; // @[PageTableCache.scala 432:46]
  wire  memPte_0_perm_d = io_refill_bits_sel_pte_dup_0[7]; // @[PageTableCache.scala 432:46]
  wire [23:0] memPte_0_ppn = io_refill_bits_sel_pte_dup_0[33:10]; // @[PageTableCache.scala 432:46]
  wire [19:0] memPte_0_ppn_high = io_refill_bits_sel_pte_dup_0[53:34]; // @[PageTableCache.scala 432:46]
  wire  memPte_1_perm_v = io_refill_bits_sel_pte_dup_1[0]; // @[PageTableCache.scala 432:46]
  wire  memPte_1_perm_r = io_refill_bits_sel_pte_dup_1[1]; // @[PageTableCache.scala 432:46]
  wire  memPte_1_perm_w = io_refill_bits_sel_pte_dup_1[2]; // @[PageTableCache.scala 432:46]
  wire  memPte_1_perm_x = io_refill_bits_sel_pte_dup_1[3]; // @[PageTableCache.scala 432:46]
  wire [23:0] memPte_1_ppn = io_refill_bits_sel_pte_dup_1[33:10]; // @[PageTableCache.scala 432:46]
  wire [19:0] memPte_1_ppn_high = io_refill_bits_sel_pte_dup_1[53:34]; // @[PageTableCache.scala 432:46]
  wire [19:0] memPte_2_ppn_high = io_refill_bits_sel_pte_dup_2[53:34]; // @[PageTableCache.scala 432:46]
  wire  _T_296 = ~flush; // @[PageTableCache.scala 435:9]
  wire  _T_299 = memPte_0_perm_r | memPte_0_perm_x | memPte_0_perm_w; // @[MMUBundle.scala 532:22]
  wire  _T_312 = io_refill_bits_level_dup_0 == 2'h1 & memPte_0_ppn[8:0] == 9'h0; // @[MMUBundle.scala 517:33]
  wire  _T_313 = io_refill_bits_level_dup_0 == 2'h2 | _T_312; // @[MMUBundle.scala 516:33]
  wire  _T_317 = io_refill_bits_level_dup_0 == 2'h0 & memPte_0_ppn[17:0] == 18'h0; // @[MMUBundle.scala 518:33]
  wire  _T_318 = _T_313 | _T_317; // @[MMUBundle.scala 517:64]
  wire  _T_320 = _T_299 & ~_T_318; // @[MMUBundle.scala 516:14]
  wire  _T_321 = ~memPte_0_perm_v | ~memPte_0_perm_r & memPte_0_perm_w | _T_320; // @[MMUBundle.scala 522:36]
  wire  _T_322 = ~_T_321; // @[PageTableCache.scala 435:70]
  wire  _T_325 = ~(memPte_0_ppn_high == 20'h0); // @[MMUBundle.scala 528:5]
  wire  _T_326 = ~_T_325; // @[PageTableCache.scala 435:110]
  wire  refillIdx_left_subtree_older = state_reg[2]; // @[Replacement.scala 243:38]
  wire  _refillIdx_T_2 = refillIdx_left_subtree_older ? state_reg_left_subtree_state : state_reg_right_subtree_state; // @[Replacement.scala 250:16]
  wire [1:0] _refillIdx_T_3 = {refillIdx_left_subtree_older,_refillIdx_T_2}; // @[Cat.scala 31:58]
  wire  _refillIdx_emptyIdx_T_1 = ~l1v[0]; // @[MMUConst.scala 132:67]
  wire  _refillIdx_emptyIdx_T_3 = ~l1v[1]; // @[MMUConst.scala 132:67]
  wire  _refillIdx_emptyIdx_T_5 = ~l1v[2]; // @[MMUConst.scala 132:67]
  wire [1:0] _refillIdx_emptyIdx_T_9 = _refillIdx_emptyIdx_T_1 ? 2'h0 : 2'h1; // @[ParallelMux.scala 90:77]
  wire [1:0] _refillIdx_emptyIdx_T_11 = _refillIdx_emptyIdx_T_5 ? 2'h2 : 2'h3; // @[ParallelMux.scala 90:77]
  wire [1:0] refillIdx_emptyIdx = _refillIdx_emptyIdx_T_1 | _refillIdx_emptyIdx_T_3 ? _refillIdx_emptyIdx_T_9 :
    _refillIdx_emptyIdx_T_11; // @[ParallelMux.scala 90:77]
  wire  refillIdx_full = &l1v; // @[MMUConst.scala 133:23]
  wire [1:0] PtwL1RefillIdx = refillIdx_full ? _refillIdx_T_3 : refillIdx_emptyIdx; // @[MMUConst.scala 134:8]
  wire [3:0] l1_rfOH = 4'h1 << PtwL1RefillIdx; // @[OneHot.scala 57:35]
  wire  state_reg_set_left_older_1 = ~PtwL1RefillIdx[1]; // @[Replacement.scala 196:33]
  wire  _state_reg_T_13 = ~PtwL1RefillIdx[0]; // @[Replacement.scala 218:7]
  wire  _state_reg_T_14 = state_reg_set_left_older_1 ? state_reg_left_subtree_state : _state_reg_T_13; // @[Replacement.scala 203:16]
  wire  _state_reg_T_18 = state_reg_set_left_older_1 ? _state_reg_T_13 : state_reg_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_reg_T_19 = {state_reg_set_left_older_1,_state_reg_T_14,_state_reg_T_18}; // @[Cat.scala 31:58]
  wire [3:0] _l1v_T = l1v | l1_rfOH; // @[PageTableCache.scala 448:16]
  wire [3:0] _l1g_T = ~l1_rfOH; // @[PageTableCache.scala 449:19]
  wire [3:0] _l1g_T_1 = l1g & _l1g_T; // @[PageTableCache.scala 449:17]
  wire [3:0] _l1g_T_2 = memPte_0_perm_g ? l1_rfOH : 4'h0; // @[PageTableCache.scala 449:31]
  wire [3:0] _l1g_T_3 = _l1g_T_1 | _l1g_T_2; // @[PageTableCache.scala 449:26]
  wire [3:0] _GEN_1728 = ~flush & io_refill_bits_levelOH_l1 & ~_T_299 & ~_T_321 & ~_T_325 ? _l1v_T : l1v; // @[PageTableCache.scala 435:129 150:20 448:9]
  wire  _T_336 = memPte_1_perm_r | memPte_1_perm_x | memPte_1_perm_w; // @[MMUBundle.scala 532:22]
  wire  _T_349 = io_refill_bits_level_dup_1 == 2'h1 & memPte_1_ppn[8:0] == 9'h0; // @[MMUBundle.scala 517:33]
  wire  _T_350 = io_refill_bits_level_dup_1 == 2'h2 | _T_349; // @[MMUBundle.scala 516:33]
  wire  _T_354 = io_refill_bits_level_dup_1 == 2'h0 & memPte_1_ppn[17:0] == 18'h0; // @[MMUBundle.scala 518:33]
  wire  _T_355 = _T_350 | _T_354; // @[MMUBundle.scala 517:64]
  wire  _T_357 = _T_336 & ~_T_355; // @[MMUBundle.scala 516:14]
  wire  _T_358 = ~memPte_1_perm_v | ~memPte_1_perm_r & memPte_1_perm_w | _T_357; // @[MMUBundle.scala 522:36]
  wire  _T_362 = ~(memPte_1_ppn_high == 20'h0); // @[MMUBundle.scala 528:5]
  wire [1:0] l2_refillIdx = io_refill_bits_req_info_dup_1_vpn[13:12]; // @[MMUConst.scala 210:21]
  wire [2:0] _GEN_1735 = 2'h1 == l2_refillIdx ? state_vec__1 : state_vec__0; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1736 = 2'h2 == l2_refillIdx ? state_vec__2 : _GEN_1735; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1737 = 2'h3 == l2_refillIdx ? state_vec__3 : _GEN_1736; // @[Replacement.scala 243:{38,38}]
  wire  victimWay_left_subtree_older = _GEN_1737[2]; // @[Replacement.scala 243:38]
  wire  victimWay_left_subtree_state = _GEN_1737[1]; // @[package.scala 154:13]
  wire  victimWay_right_subtree_state = _GEN_1737[0]; // @[Replacement.scala 245:38]
  wire  _victimWay_T_2 = victimWay_left_subtree_older ? victimWay_left_subtree_state : victimWay_right_subtree_state; // @[Replacement.scala 250:16]
  wire [1:0] _victimWay_T_3 = {victimWay_left_subtree_older,_victimWay_T_2}; // @[Cat.scala 31:58]
  wire [3:0] _GEN_1739 = 2'h1 == l2_refillIdx ? l2vVec_1 : l2vVec_0; // @[MMUConst.scala 132:{69,69}]
  wire [3:0] _GEN_1740 = 2'h2 == l2_refillIdx ? l2vVec_2 : _GEN_1739; // @[MMUConst.scala 132:{69,69}]
  wire [3:0] _GEN_1741 = 2'h3 == l2_refillIdx ? l2vVec_3 : _GEN_1740; // @[MMUConst.scala 132:{69,69}]
  wire  _victimWay_emptyIdx_T_1 = ~_GEN_1741[0]; // @[MMUConst.scala 132:67]
  wire  _victimWay_emptyIdx_T_3 = ~_GEN_1741[1]; // @[MMUConst.scala 132:67]
  wire  _victimWay_emptyIdx_T_5 = ~_GEN_1741[2]; // @[MMUConst.scala 132:67]
  wire [1:0] _victimWay_emptyIdx_T_9 = _victimWay_emptyIdx_T_1 ? 2'h0 : 2'h1; // @[ParallelMux.scala 90:77]
  wire [1:0] _victimWay_emptyIdx_T_11 = _victimWay_emptyIdx_T_5 ? 2'h2 : 2'h3; // @[ParallelMux.scala 90:77]
  wire [1:0] victimWay_emptyIdx = _victimWay_emptyIdx_T_1 | _victimWay_emptyIdx_T_3 ? _victimWay_emptyIdx_T_9 :
    _victimWay_emptyIdx_T_11; // @[ParallelMux.scala 90:77]
  wire  victimWay_full = &_GEN_1741; // @[MMUConst.scala 133:23]
  wire [1:0] l2_victimWay = victimWay_full ? _victimWay_T_3 : victimWay_emptyIdx; // @[MMUConst.scala 134:8]
  wire [3:0] _rfvOH_T = {l2_refillIdx,l2_victimWay}; // @[Cat.scala 31:58]
  wire [15:0] l2_rfvOH = 16'h1 << _rfvOH_T; // @[OneHot.scala 57:35]
  wire [12:0] wdata_entries_ps_tag = io_refill_bits_req_info_dup_1_vpn[26:14]; // @[MMUBundle.scala 646:8]
  wire  _wdata_entries_ps_vs_0_T_3 = ~memPtes_0_perm_v | ~memPtes_0_perm_r & memPtes_0_perm_w; // @[MMUBundle.scala 522:13]
  wire  _wdata_entries_ps_vs_0_T_5 = memPtes_0_perm_r | memPtes_0_perm_x | memPtes_0_perm_w; // @[MMUBundle.scala 532:22]
  wire  _wdata_entries_ps_vs_0_T_9 = memPtes_0_ppn[8:0] == 9'h0; // @[MMUBundle.scala 517:56]
  wire  _wdata_entries_ps_vs_0_T_18 = _wdata_entries_ps_vs_0_T_5 & ~_wdata_entries_ps_vs_0_T_9; // @[MMUBundle.scala 516:14]
  wire  _wdata_entries_ps_vs_0_T_19 = ~memPtes_0_perm_v | ~memPtes_0_perm_r & memPtes_0_perm_w |
    _wdata_entries_ps_vs_0_T_18; // @[MMUBundle.scala 522:36]
  wire  wdata_entries_ps_vs_0 = ~_wdata_entries_ps_vs_0_T_19 & ~_wdata_entries_ps_vs_0_T_5; // @[MMUBundle.scala 669:42]
  wire  _wdata_entries_ps_vs_1_T_3 = ~memPtes_1_perm_v | ~memPtes_1_perm_r & memPtes_1_perm_w; // @[MMUBundle.scala 522:13]
  wire  _wdata_entries_ps_vs_1_T_5 = memPtes_1_perm_r | memPtes_1_perm_x | memPtes_1_perm_w; // @[MMUBundle.scala 532:22]
  wire  _wdata_entries_ps_vs_1_T_9 = memPtes_1_ppn[8:0] == 9'h0; // @[MMUBundle.scala 517:56]
  wire  _wdata_entries_ps_vs_1_T_18 = _wdata_entries_ps_vs_1_T_5 & ~_wdata_entries_ps_vs_1_T_9; // @[MMUBundle.scala 516:14]
  wire  _wdata_entries_ps_vs_1_T_19 = ~memPtes_1_perm_v | ~memPtes_1_perm_r & memPtes_1_perm_w |
    _wdata_entries_ps_vs_1_T_18; // @[MMUBundle.scala 522:36]
  wire  wdata_entries_ps_vs_1 = ~_wdata_entries_ps_vs_1_T_19 & ~_wdata_entries_ps_vs_1_T_5; // @[MMUBundle.scala 669:42]
  wire  _wdata_entries_ps_vs_2_T_3 = ~memPtes_2_perm_v | ~memPtes_2_perm_r & memPtes_2_perm_w; // @[MMUBundle.scala 522:13]
  wire  _wdata_entries_ps_vs_2_T_5 = memPtes_2_perm_r | memPtes_2_perm_x | memPtes_2_perm_w; // @[MMUBundle.scala 532:22]
  wire  _wdata_entries_ps_vs_2_T_9 = memPtes_2_ppn[8:0] == 9'h0; // @[MMUBundle.scala 517:56]
  wire  _wdata_entries_ps_vs_2_T_18 = _wdata_entries_ps_vs_2_T_5 & ~_wdata_entries_ps_vs_2_T_9; // @[MMUBundle.scala 516:14]
  wire  _wdata_entries_ps_vs_2_T_19 = ~memPtes_2_perm_v | ~memPtes_2_perm_r & memPtes_2_perm_w |
    _wdata_entries_ps_vs_2_T_18; // @[MMUBundle.scala 522:36]
  wire  wdata_entries_ps_vs_2 = ~_wdata_entries_ps_vs_2_T_19 & ~_wdata_entries_ps_vs_2_T_5; // @[MMUBundle.scala 669:42]
  wire  _wdata_entries_ps_vs_3_T_3 = ~memPtes_3_perm_v | ~memPtes_3_perm_r & memPtes_3_perm_w; // @[MMUBundle.scala 522:13]
  wire  _wdata_entries_ps_vs_3_T_5 = memPtes_3_perm_r | memPtes_3_perm_x | memPtes_3_perm_w; // @[MMUBundle.scala 532:22]
  wire  _wdata_entries_ps_vs_3_T_9 = memPtes_3_ppn[8:0] == 9'h0; // @[MMUBundle.scala 517:56]
  wire  _wdata_entries_ps_vs_3_T_18 = _wdata_entries_ps_vs_3_T_5 & ~_wdata_entries_ps_vs_3_T_9; // @[MMUBundle.scala 516:14]
  wire  _wdata_entries_ps_vs_3_T_19 = ~memPtes_3_perm_v | ~memPtes_3_perm_r & memPtes_3_perm_w |
    _wdata_entries_ps_vs_3_T_18; // @[MMUBundle.scala 522:36]
  wire  wdata_entries_ps_vs_3 = ~_wdata_entries_ps_vs_3_T_19 & ~_wdata_entries_ps_vs_3_T_5; // @[MMUBundle.scala 669:42]
  wire  _wdata_entries_ps_vs_4_T_3 = ~memPtes_4_perm_v | ~memPtes_4_perm_r & memPtes_4_perm_w; // @[MMUBundle.scala 522:13]
  wire  _wdata_entries_ps_vs_4_T_5 = memPtes_4_perm_r | memPtes_4_perm_x | memPtes_4_perm_w; // @[MMUBundle.scala 532:22]
  wire  _wdata_entries_ps_vs_4_T_9 = memPtes_4_ppn[8:0] == 9'h0; // @[MMUBundle.scala 517:56]
  wire  _wdata_entries_ps_vs_4_T_18 = _wdata_entries_ps_vs_4_T_5 & ~_wdata_entries_ps_vs_4_T_9; // @[MMUBundle.scala 516:14]
  wire  _wdata_entries_ps_vs_4_T_19 = ~memPtes_4_perm_v | ~memPtes_4_perm_r & memPtes_4_perm_w |
    _wdata_entries_ps_vs_4_T_18; // @[MMUBundle.scala 522:36]
  wire  wdata_entries_ps_vs_4 = ~_wdata_entries_ps_vs_4_T_19 & ~_wdata_entries_ps_vs_4_T_5; // @[MMUBundle.scala 669:42]
  wire  _wdata_entries_ps_vs_5_T_3 = ~memPtes_5_perm_v | ~memPtes_5_perm_r & memPtes_5_perm_w; // @[MMUBundle.scala 522:13]
  wire  _wdata_entries_ps_vs_5_T_5 = memPtes_5_perm_r | memPtes_5_perm_x | memPtes_5_perm_w; // @[MMUBundle.scala 532:22]
  wire  _wdata_entries_ps_vs_5_T_9 = memPtes_5_ppn[8:0] == 9'h0; // @[MMUBundle.scala 517:56]
  wire  _wdata_entries_ps_vs_5_T_18 = _wdata_entries_ps_vs_5_T_5 & ~_wdata_entries_ps_vs_5_T_9; // @[MMUBundle.scala 516:14]
  wire  _wdata_entries_ps_vs_5_T_19 = ~memPtes_5_perm_v | ~memPtes_5_perm_r & memPtes_5_perm_w |
    _wdata_entries_ps_vs_5_T_18; // @[MMUBundle.scala 522:36]
  wire  wdata_entries_ps_vs_5 = ~_wdata_entries_ps_vs_5_T_19 & ~_wdata_entries_ps_vs_5_T_5; // @[MMUBundle.scala 669:42]
  wire  _wdata_entries_ps_vs_6_T_3 = ~memPtes_6_perm_v | ~memPtes_6_perm_r & memPtes_6_perm_w; // @[MMUBundle.scala 522:13]
  wire  _wdata_entries_ps_vs_6_T_5 = memPtes_6_perm_r | memPtes_6_perm_x | memPtes_6_perm_w; // @[MMUBundle.scala 532:22]
  wire  _wdata_entries_ps_vs_6_T_9 = memPtes_6_ppn[8:0] == 9'h0; // @[MMUBundle.scala 517:56]
  wire  _wdata_entries_ps_vs_6_T_18 = _wdata_entries_ps_vs_6_T_5 & ~_wdata_entries_ps_vs_6_T_9; // @[MMUBundle.scala 516:14]
  wire  _wdata_entries_ps_vs_6_T_19 = ~memPtes_6_perm_v | ~memPtes_6_perm_r & memPtes_6_perm_w |
    _wdata_entries_ps_vs_6_T_18; // @[MMUBundle.scala 522:36]
  wire  wdata_entries_ps_vs_6 = ~_wdata_entries_ps_vs_6_T_19 & ~_wdata_entries_ps_vs_6_T_5; // @[MMUBundle.scala 669:42]
  wire  _wdata_entries_ps_vs_7_T_3 = ~memPtes_7_perm_v | ~memPtes_7_perm_r & memPtes_7_perm_w; // @[MMUBundle.scala 522:13]
  wire  _wdata_entries_ps_vs_7_T_5 = memPtes_7_perm_r | memPtes_7_perm_x | memPtes_7_perm_w; // @[MMUBundle.scala 532:22]
  wire  _wdata_entries_ps_vs_7_T_9 = memPtes_7_ppn[8:0] == 9'h0; // @[MMUBundle.scala 517:56]
  wire  _wdata_entries_ps_vs_7_T_18 = _wdata_entries_ps_vs_7_T_5 & ~_wdata_entries_ps_vs_7_T_9; // @[MMUBundle.scala 516:14]
  wire  _wdata_entries_ps_vs_7_T_19 = ~memPtes_7_perm_v | ~memPtes_7_perm_r & memPtes_7_perm_w |
    _wdata_entries_ps_vs_7_T_18; // @[MMUBundle.scala 522:36]
  wire  wdata_entries_ps_vs_7 = ~_wdata_entries_ps_vs_7_T_19 & ~_wdata_entries_ps_vs_7_T_5; // @[MMUBundle.scala 669:42]
  wire [220:0] data_hi_2 = {wdata_entries_ps_tag,io_csr_dup_1_satp_asid,memPtes_7_ppn,memPtes_6_ppn,memPtes_5_ppn,
    memPtes_4_ppn,memPtes_3_ppn,memPtes_2_ppn,memPtes_1_ppn,memPtes_0_ppn}; // @[MMUBundle.scala 705:30]
  wire [229:0] data_5 = {data_hi_2,wdata_entries_ps_vs_7,wdata_entries_ps_vs_6,wdata_entries_ps_vs_5,
    wdata_entries_ps_vs_4,wdata_entries_ps_vs_3,wdata_entries_ps_vs_2,wdata_entries_ps_vs_1,wdata_entries_ps_vs_0,
    refill_prefetch_dup_1}; // @[MMUBundle.scala 705:30]
  wire [63:0] _ecc_slices_0_syndromeUInt_T = 64'hab55555556aaad5b & data_5[63:0]; // @[ECC.scala 147:74]
  wire  _ecc_slices_0_syndromeUInt_T_1 = ^_ecc_slices_0_syndromeUInt_T; // @[ECC.scala 147:79]
  wire [63:0] _ecc_slices_0_syndromeUInt_T_3 = 64'hcd9999999b33366d & data_5[63:0]; // @[ECC.scala 147:74]
  wire  _ecc_slices_0_syndromeUInt_T_4 = ^_ecc_slices_0_syndromeUInt_T_3; // @[ECC.scala 147:79]
  wire [63:0] _ecc_slices_0_syndromeUInt_T_6 = 64'hf1e1e1e1e3c3c78e & data_5[63:0]; // @[ECC.scala 147:74]
  wire  _ecc_slices_0_syndromeUInt_T_7 = ^_ecc_slices_0_syndromeUInt_T_6; // @[ECC.scala 147:79]
  wire [63:0] _ecc_slices_0_syndromeUInt_T_9 = 64'h1fe01fe03fc07f0 & data_5[63:0]; // @[ECC.scala 147:74]
  wire  _ecc_slices_0_syndromeUInt_T_10 = ^_ecc_slices_0_syndromeUInt_T_9; // @[ECC.scala 147:79]
  wire [63:0] _ecc_slices_0_syndromeUInt_T_12 = 64'h1fffe0003fff800 & data_5[63:0]; // @[ECC.scala 147:74]
  wire  _ecc_slices_0_syndromeUInt_T_13 = ^_ecc_slices_0_syndromeUInt_T_12; // @[ECC.scala 147:79]
  wire [63:0] _ecc_slices_0_syndromeUInt_T_15 = 64'h1fffffffc000000 & data_5[63:0]; // @[ECC.scala 147:74]
  wire  _ecc_slices_0_syndromeUInt_T_16 = ^_ecc_slices_0_syndromeUInt_T_15; // @[ECC.scala 147:79]
  wire [63:0] _ecc_slices_0_syndromeUInt_T_18 = 64'hfe00000000000000 & data_5[63:0]; // @[ECC.scala 147:74]
  wire  _ecc_slices_0_syndromeUInt_T_19 = ^_ecc_slices_0_syndromeUInt_T_18; // @[ECC.scala 147:79]
  wire [70:0] _ecc_slices_0_T_1 = {_ecc_slices_0_syndromeUInt_T_19,_ecc_slices_0_syndromeUInt_T_16,
    _ecc_slices_0_syndromeUInt_T_13,_ecc_slices_0_syndromeUInt_T_10,_ecc_slices_0_syndromeUInt_T_7,
    _ecc_slices_0_syndromeUInt_T_4,_ecc_slices_0_syndromeUInt_T_1,data_5[63:0]}; // @[Cat.scala 31:58]
  wire  _ecc_slices_0_T_2 = ^_ecc_slices_0_T_1; // @[ECC.scala 81:55]
  wire [71:0] _ecc_slices_0_T_4 = {_ecc_slices_0_T_2,_ecc_slices_0_syndromeUInt_T_19,_ecc_slices_0_syndromeUInt_T_16,
    _ecc_slices_0_syndromeUInt_T_13,_ecc_slices_0_syndromeUInt_T_10,_ecc_slices_0_syndromeUInt_T_7,
    _ecc_slices_0_syndromeUInt_T_4,_ecc_slices_0_syndromeUInt_T_1,data_5[63:0]}; // @[Cat.scala 31:58]
  wire [7:0] ecc_slices__0 = _ecc_slices_0_T_4[71:64]; // @[MMUBundle.scala 708:77]
  wire [63:0] _ecc_slices_1_syndromeUInt_T = 64'hab55555556aaad5b & data_5[127:64]; // @[ECC.scala 147:74]
  wire  _ecc_slices_1_syndromeUInt_T_1 = ^_ecc_slices_1_syndromeUInt_T; // @[ECC.scala 147:79]
  wire [63:0] _ecc_slices_1_syndromeUInt_T_3 = 64'hcd9999999b33366d & data_5[127:64]; // @[ECC.scala 147:74]
  wire  _ecc_slices_1_syndromeUInt_T_4 = ^_ecc_slices_1_syndromeUInt_T_3; // @[ECC.scala 147:79]
  wire [63:0] _ecc_slices_1_syndromeUInt_T_6 = 64'hf1e1e1e1e3c3c78e & data_5[127:64]; // @[ECC.scala 147:74]
  wire  _ecc_slices_1_syndromeUInt_T_7 = ^_ecc_slices_1_syndromeUInt_T_6; // @[ECC.scala 147:79]
  wire [63:0] _ecc_slices_1_syndromeUInt_T_9 = 64'h1fe01fe03fc07f0 & data_5[127:64]; // @[ECC.scala 147:74]
  wire  _ecc_slices_1_syndromeUInt_T_10 = ^_ecc_slices_1_syndromeUInt_T_9; // @[ECC.scala 147:79]
  wire [63:0] _ecc_slices_1_syndromeUInt_T_12 = 64'h1fffe0003fff800 & data_5[127:64]; // @[ECC.scala 147:74]
  wire  _ecc_slices_1_syndromeUInt_T_13 = ^_ecc_slices_1_syndromeUInt_T_12; // @[ECC.scala 147:79]
  wire [63:0] _ecc_slices_1_syndromeUInt_T_15 = 64'h1fffffffc000000 & data_5[127:64]; // @[ECC.scala 147:74]
  wire  _ecc_slices_1_syndromeUInt_T_16 = ^_ecc_slices_1_syndromeUInt_T_15; // @[ECC.scala 147:79]
  wire [63:0] _ecc_slices_1_syndromeUInt_T_18 = 64'hfe00000000000000 & data_5[127:64]; // @[ECC.scala 147:74]
  wire  _ecc_slices_1_syndromeUInt_T_19 = ^_ecc_slices_1_syndromeUInt_T_18; // @[ECC.scala 147:79]
  wire [70:0] _ecc_slices_1_T_1 = {_ecc_slices_1_syndromeUInt_T_19,_ecc_slices_1_syndromeUInt_T_16,
    _ecc_slices_1_syndromeUInt_T_13,_ecc_slices_1_syndromeUInt_T_10,_ecc_slices_1_syndromeUInt_T_7,
    _ecc_slices_1_syndromeUInt_T_4,_ecc_slices_1_syndromeUInt_T_1,data_5[127:64]}; // @[Cat.scala 31:58]
  wire  _ecc_slices_1_T_2 = ^_ecc_slices_1_T_1; // @[ECC.scala 81:55]
  wire [71:0] _ecc_slices_1_T_4 = {_ecc_slices_1_T_2,_ecc_slices_1_syndromeUInt_T_19,_ecc_slices_1_syndromeUInt_T_16,
    _ecc_slices_1_syndromeUInt_T_13,_ecc_slices_1_syndromeUInt_T_10,_ecc_slices_1_syndromeUInt_T_7,
    _ecc_slices_1_syndromeUInt_T_4,_ecc_slices_1_syndromeUInt_T_1,data_5[127:64]}; // @[Cat.scala 31:58]
  wire [7:0] ecc_slices__1 = _ecc_slices_1_T_4[71:64]; // @[MMUBundle.scala 708:77]
  wire [63:0] _ecc_slices_2_syndromeUInt_T = 64'hab55555556aaad5b & data_5[191:128]; // @[ECC.scala 147:74]
  wire  _ecc_slices_2_syndromeUInt_T_1 = ^_ecc_slices_2_syndromeUInt_T; // @[ECC.scala 147:79]
  wire [63:0] _ecc_slices_2_syndromeUInt_T_3 = 64'hcd9999999b33366d & data_5[191:128]; // @[ECC.scala 147:74]
  wire  _ecc_slices_2_syndromeUInt_T_4 = ^_ecc_slices_2_syndromeUInt_T_3; // @[ECC.scala 147:79]
  wire [63:0] _ecc_slices_2_syndromeUInt_T_6 = 64'hf1e1e1e1e3c3c78e & data_5[191:128]; // @[ECC.scala 147:74]
  wire  _ecc_slices_2_syndromeUInt_T_7 = ^_ecc_slices_2_syndromeUInt_T_6; // @[ECC.scala 147:79]
  wire [63:0] _ecc_slices_2_syndromeUInt_T_9 = 64'h1fe01fe03fc07f0 & data_5[191:128]; // @[ECC.scala 147:74]
  wire  _ecc_slices_2_syndromeUInt_T_10 = ^_ecc_slices_2_syndromeUInt_T_9; // @[ECC.scala 147:79]
  wire [63:0] _ecc_slices_2_syndromeUInt_T_12 = 64'h1fffe0003fff800 & data_5[191:128]; // @[ECC.scala 147:74]
  wire  _ecc_slices_2_syndromeUInt_T_13 = ^_ecc_slices_2_syndromeUInt_T_12; // @[ECC.scala 147:79]
  wire [63:0] _ecc_slices_2_syndromeUInt_T_15 = 64'h1fffffffc000000 & data_5[191:128]; // @[ECC.scala 147:74]
  wire  _ecc_slices_2_syndromeUInt_T_16 = ^_ecc_slices_2_syndromeUInt_T_15; // @[ECC.scala 147:79]
  wire [63:0] _ecc_slices_2_syndromeUInt_T_18 = 64'hfe00000000000000 & data_5[191:128]; // @[ECC.scala 147:74]
  wire  _ecc_slices_2_syndromeUInt_T_19 = ^_ecc_slices_2_syndromeUInt_T_18; // @[ECC.scala 147:79]
  wire [70:0] _ecc_slices_2_T_1 = {_ecc_slices_2_syndromeUInt_T_19,_ecc_slices_2_syndromeUInt_T_16,
    _ecc_slices_2_syndromeUInt_T_13,_ecc_slices_2_syndromeUInt_T_10,_ecc_slices_2_syndromeUInt_T_7,
    _ecc_slices_2_syndromeUInt_T_4,_ecc_slices_2_syndromeUInt_T_1,data_5[191:128]}; // @[Cat.scala 31:58]
  wire  _ecc_slices_2_T_2 = ^_ecc_slices_2_T_1; // @[ECC.scala 81:55]
  wire [71:0] _ecc_slices_2_T_4 = {_ecc_slices_2_T_2,_ecc_slices_2_syndromeUInt_T_19,_ecc_slices_2_syndromeUInt_T_16,
    _ecc_slices_2_syndromeUInt_T_13,_ecc_slices_2_syndromeUInt_T_10,_ecc_slices_2_syndromeUInt_T_7,
    _ecc_slices_2_syndromeUInt_T_4,_ecc_slices_2_syndromeUInt_T_1,data_5[191:128]}; // @[Cat.scala 31:58]
  wire [7:0] ecc_slices__2 = _ecc_slices_2_T_4[71:64]; // @[MMUBundle.scala 708:77]
  wire [37:0] _ecc_unaligned_syndromeUInt_T = 38'h1556aaad5b & data_5[229:192]; // @[ECC.scala 147:74]
  wire  _ecc_unaligned_syndromeUInt_T_1 = ^_ecc_unaligned_syndromeUInt_T; // @[ECC.scala 147:79]
  wire [37:0] _ecc_unaligned_syndromeUInt_T_3 = 38'h199b33366d & data_5[229:192]; // @[ECC.scala 147:74]
  wire  _ecc_unaligned_syndromeUInt_T_4 = ^_ecc_unaligned_syndromeUInt_T_3; // @[ECC.scala 147:79]
  wire [37:0] _ecc_unaligned_syndromeUInt_T_6 = 38'h21e3c3c78e & data_5[229:192]; // @[ECC.scala 147:74]
  wire  _ecc_unaligned_syndromeUInt_T_7 = ^_ecc_unaligned_syndromeUInt_T_6; // @[ECC.scala 147:79]
  wire [37:0] _ecc_unaligned_syndromeUInt_T_9 = 38'h3e03fc07f0 & data_5[229:192]; // @[ECC.scala 147:74]
  wire  _ecc_unaligned_syndromeUInt_T_10 = ^_ecc_unaligned_syndromeUInt_T_9; // @[ECC.scala 147:79]
  wire [37:0] _ecc_unaligned_syndromeUInt_T_12 = 38'h3fff800 & data_5[229:192]; // @[ECC.scala 147:74]
  wire  _ecc_unaligned_syndromeUInt_T_13 = ^_ecc_unaligned_syndromeUInt_T_12; // @[ECC.scala 147:79]
  wire [37:0] _ecc_unaligned_syndromeUInt_T_15 = 38'h3ffc000000 & data_5[229:192]; // @[ECC.scala 147:74]
  wire  _ecc_unaligned_syndromeUInt_T_16 = ^_ecc_unaligned_syndromeUInt_T_15; // @[ECC.scala 147:79]
  wire [43:0] _ecc_unaligned_T_1 = {_ecc_unaligned_syndromeUInt_T_16,_ecc_unaligned_syndromeUInt_T_13,
    _ecc_unaligned_syndromeUInt_T_10,_ecc_unaligned_syndromeUInt_T_7,_ecc_unaligned_syndromeUInt_T_4,
    _ecc_unaligned_syndromeUInt_T_1,data_5[229:192]}; // @[Cat.scala 31:58]
  wire  _ecc_unaligned_T_2 = ^_ecc_unaligned_T_1; // @[ECC.scala 81:55]
  wire [44:0] _ecc_unaligned_T_4 = {_ecc_unaligned_T_2,_ecc_unaligned_syndromeUInt_T_16,_ecc_unaligned_syndromeUInt_T_13
    ,_ecc_unaligned_syndromeUInt_T_10,_ecc_unaligned_syndromeUInt_T_7,_ecc_unaligned_syndromeUInt_T_4,
    _ecc_unaligned_syndromeUInt_T_1,data_5[229:192]}; // @[Cat.scala 31:58]
  wire [6:0] ecc_unaligned = _ecc_unaligned_T_4[44:38]; // @[MMUBundle.scala 711:88]
  wire [23:0] _wdata_ecc_T = {ecc_slices__2,ecc_slices__1,ecc_slices__0}; // @[MMUBundle.scala 712:50]
  wire  state_vec_set_left_older_4 = ~l2_victimWay[1]; // @[Replacement.scala 196:33]
  wire  _state_vec_T_34 = ~l2_victimWay[0]; // @[Replacement.scala 218:7]
  wire  _state_vec_T_35 = state_vec_set_left_older_4 ? victimWay_left_subtree_state : _state_vec_T_34; // @[Replacement.scala 203:16]
  wire  _state_vec_T_39 = state_vec_set_left_older_4 ? _state_vec_T_34 : victimWay_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_T_40 = {state_vec_set_left_older_4,_state_vec_T_35,_state_vec_T_39}; // @[Cat.scala 31:58]
  wire [15:0] _l2v_T = l2v | l2_rfvOH; // @[PageTableCache.scala 482:16]
  wire [15:0] _l2g_T = ~l2_rfvOH; // @[PageTableCache.scala 483:18]
  wire [15:0] _l2g_T_1 = l2g & _l2g_T; // @[PageTableCache.scala 483:16]
  wire [7:0] _l2g_T_2 = {memPtes_0_perm_g,memPtes_1_perm_g,memPtes_2_perm_g,memPtes_3_perm_g,memPtes_4_perm_g,
    memPtes_5_perm_g,memPtes_6_perm_g,memPtes_7_perm_g}; // @[Cat.scala 31:58]
  wire  _l2g_T_3 = &_l2g_T_2; // @[PageTableCache.scala 483:58]
  wire [15:0] _l2g_T_4 = &_l2g_T_2 ? l2_rfvOH : 16'h0; // @[PageTableCache.scala 483:30]
  wire [15:0] _l2g_T_5 = _l2g_T_1 | _l2g_T_4; // @[PageTableCache.scala 483:25]
  wire [15:0] _GEN_1833 = ~flush_dup_1 & io_refill_bits_levelOH_l2 & ~_T_336 & ~_T_358 & ~_T_362 ? _l2v_T : l2v; // @[PageTableCache.scala 462:129 161:20 482:9]
  wire  _T_377 = ~(memPte_2_ppn_high == 20'h0); // @[MMUBundle.scala 528:5]
  wire [1:0] l3_refillIdx = io_refill_bits_req_info_dup_2_vpn[4:3]; // @[MMUConst.scala 226:21]
  wire [6:0] _GEN_1840 = 2'h1 == l3_refillIdx ? state_vec_1_1 : state_vec_1_0; // @[Replacement.scala 243:{38,38}]
  wire [6:0] _GEN_1841 = 2'h2 == l3_refillIdx ? state_vec_1_2 : _GEN_1840; // @[Replacement.scala 243:{38,38}]
  wire [6:0] _GEN_1842 = 2'h3 == l3_refillIdx ? state_vec_1_3 : _GEN_1841; // @[Replacement.scala 243:{38,38}]
  wire  victimWay_left_subtree_older_1 = _GEN_1842[6]; // @[Replacement.scala 243:38]
  wire [2:0] victimWay_left_subtree_state_1 = _GEN_1842[5:3]; // @[package.scala 154:13]
  wire [2:0] victimWay_right_subtree_state_1 = _GEN_1842[2:0]; // @[Replacement.scala 245:38]
  wire  victimWay_left_subtree_older_2 = victimWay_left_subtree_state_1[2]; // @[Replacement.scala 243:38]
  wire  victimWay_left_subtree_state_2 = victimWay_left_subtree_state_1[1]; // @[package.scala 154:13]
  wire  victimWay_right_subtree_state_2 = victimWay_left_subtree_state_1[0]; // @[Replacement.scala 245:38]
  wire  _victimWay_T_6 = victimWay_left_subtree_older_2 ? victimWay_left_subtree_state_2 :
    victimWay_right_subtree_state_2; // @[Replacement.scala 250:16]
  wire [1:0] _victimWay_T_7 = {victimWay_left_subtree_older_2,_victimWay_T_6}; // @[Cat.scala 31:58]
  wire  victimWay_left_subtree_older_3 = victimWay_right_subtree_state_1[2]; // @[Replacement.scala 243:38]
  wire  victimWay_left_subtree_state_3 = victimWay_right_subtree_state_1[1]; // @[package.scala 154:13]
  wire  victimWay_right_subtree_state_3 = victimWay_right_subtree_state_1[0]; // @[Replacement.scala 245:38]
  wire  _victimWay_T_10 = victimWay_left_subtree_older_3 ? victimWay_left_subtree_state_3 :
    victimWay_right_subtree_state_3; // @[Replacement.scala 250:16]
  wire [1:0] _victimWay_T_11 = {victimWay_left_subtree_older_3,_victimWay_T_10}; // @[Cat.scala 31:58]
  wire [1:0] _victimWay_T_12 = victimWay_left_subtree_older_1 ? _victimWay_T_7 : _victimWay_T_11; // @[Replacement.scala 250:16]
  wire [2:0] _victimWay_T_13 = {victimWay_left_subtree_older_1,_victimWay_T_12}; // @[Cat.scala 31:58]
  wire [7:0] _GEN_1844 = 2'h1 == l3_refillIdx ? l3vVec_1 : l3vVec_0; // @[MMUConst.scala 132:{69,69}]
  wire [7:0] _GEN_1845 = 2'h2 == l3_refillIdx ? l3vVec_2 : _GEN_1844; // @[MMUConst.scala 132:{69,69}]
  wire [7:0] _GEN_1846 = 2'h3 == l3_refillIdx ? l3vVec_3 : _GEN_1845; // @[MMUConst.scala 132:{69,69}]
  wire  _victimWay_emptyIdx_T_14 = ~_GEN_1846[0]; // @[MMUConst.scala 132:67]
  wire  _victimWay_emptyIdx_T_16 = ~_GEN_1846[1]; // @[MMUConst.scala 132:67]
  wire  _victimWay_emptyIdx_T_18 = ~_GEN_1846[2]; // @[MMUConst.scala 132:67]
  wire  _victimWay_emptyIdx_T_20 = ~_GEN_1846[3]; // @[MMUConst.scala 132:67]
  wire  _victimWay_emptyIdx_T_22 = ~_GEN_1846[4]; // @[MMUConst.scala 132:67]
  wire  _victimWay_emptyIdx_T_24 = ~_GEN_1846[5]; // @[MMUConst.scala 132:67]
  wire  _victimWay_emptyIdx_T_26 = ~_GEN_1846[6]; // @[MMUConst.scala 132:67]
  wire [2:0] _victimWay_emptyIdx_T_30 = _victimWay_emptyIdx_T_14 ? 3'h0 : 3'h1; // @[ParallelMux.scala 90:77]
  wire [2:0] _victimWay_emptyIdx_T_32 = _victimWay_emptyIdx_T_18 ? 3'h2 : 3'h3; // @[ParallelMux.scala 90:77]
  wire [2:0] _victimWay_emptyIdx_T_34 = _victimWay_emptyIdx_T_14 | _victimWay_emptyIdx_T_16 ? _victimWay_emptyIdx_T_30
     : _victimWay_emptyIdx_T_32; // @[ParallelMux.scala 90:77]
  wire [2:0] _victimWay_emptyIdx_T_36 = _victimWay_emptyIdx_T_22 ? 3'h4 : 3'h5; // @[ParallelMux.scala 90:77]
  wire [2:0] _victimWay_emptyIdx_T_38 = _victimWay_emptyIdx_T_26 ? 3'h6 : 3'h7; // @[ParallelMux.scala 90:77]
  wire [2:0] _victimWay_emptyIdx_T_40 = _victimWay_emptyIdx_T_22 | _victimWay_emptyIdx_T_24 ? _victimWay_emptyIdx_T_36
     : _victimWay_emptyIdx_T_38; // @[ParallelMux.scala 90:77]
  wire [2:0] victimWay_emptyIdx_1 = _victimWay_emptyIdx_T_14 | _victimWay_emptyIdx_T_16 | (_victimWay_emptyIdx_T_18 |
    _victimWay_emptyIdx_T_20) ? _victimWay_emptyIdx_T_34 : _victimWay_emptyIdx_T_40; // @[ParallelMux.scala 90:77]
  wire  victimWay_full_1 = &_GEN_1846; // @[MMUConst.scala 133:23]
  wire [2:0] l3_victimWay = victimWay_full_1 ? _victimWay_T_13 : victimWay_emptyIdx_1; // @[MMUConst.scala 134:8]
  wire [4:0] _rfvOH_T_1 = {l3_refillIdx,l3_victimWay}; // @[Cat.scala 31:58]
  wire [31:0] l3_rfvOH = 32'h1 << _rfvOH_T_1; // @[OneHot.scala 57:35]
  wire [21:0] wdata_entries_ps_1_tag = io_refill_bits_req_info_dup_2_vpn[26:5]; // @[MMUBundle.scala 646:8]
  wire  wdata_entries_ps_1_vs_0 = ~_wdata_entries_ps_vs_0_T_3 & _wdata_entries_ps_vs_0_T_5; // @[MMUBundle.scala 669:42]
  wire  wdata_entries_ps_1_vs_1 = ~_wdata_entries_ps_vs_1_T_3 & _wdata_entries_ps_vs_1_T_5; // @[MMUBundle.scala 669:42]
  wire  wdata_entries_ps_1_vs_2 = ~_wdata_entries_ps_vs_2_T_3 & _wdata_entries_ps_vs_2_T_5; // @[MMUBundle.scala 669:42]
  wire  wdata_entries_ps_1_vs_3 = ~_wdata_entries_ps_vs_3_T_3 & _wdata_entries_ps_vs_3_T_5; // @[MMUBundle.scala 669:42]
  wire  wdata_entries_ps_1_vs_4 = ~_wdata_entries_ps_vs_4_T_3 & _wdata_entries_ps_vs_4_T_5; // @[MMUBundle.scala 669:42]
  wire  wdata_entries_ps_1_vs_5 = ~_wdata_entries_ps_vs_5_T_3 & _wdata_entries_ps_vs_5_T_5; // @[MMUBundle.scala 669:42]
  wire  wdata_entries_ps_1_vs_6 = ~_wdata_entries_ps_vs_6_T_3 & _wdata_entries_ps_vs_6_T_5; // @[MMUBundle.scala 669:42]
  wire  wdata_entries_ps_1_vs_7 = ~_wdata_entries_ps_vs_7_T_3 & _wdata_entries_ps_vs_7_T_5; // @[MMUBundle.scala 669:42]
  wire [8:0] data_lo_lo_lo_3 = {memPtes_1_perm_r,memPtes_0_perm_d,memPtes_0_perm_a,memPtes_0_perm_g,memPtes_0_perm_u,
    memPtes_0_perm_x,memPtes_0_perm_w,memPtes_0_perm_r,refill_prefetch_dup_2}; // @[MMUBundle.scala 705:30]
  wire [17:0] data_lo_lo_3 = {memPtes_2_perm_x,memPtes_2_perm_w,memPtes_2_perm_r,memPtes_1_perm_d,memPtes_1_perm_a,
    memPtes_1_perm_g,memPtes_1_perm_u,memPtes_1_perm_x,memPtes_1_perm_w,data_lo_lo_lo_3}; // @[MMUBundle.scala 705:30]
  wire [9:0] data_lo_hi_hi_3 = {memPtes_5_perm_r,memPtes_4_perm_d,memPtes_4_perm_a,memPtes_4_perm_g,memPtes_4_perm_u,
    memPtes_4_perm_x,memPtes_4_perm_w,memPtes_4_perm_r,memPtes_3_perm_d,memPtes_3_perm_a}; // @[MMUBundle.scala 705:30]
  wire [18:0] data_lo_hi_3 = {data_lo_hi_hi_3,memPtes_3_perm_g,memPtes_3_perm_u,memPtes_3_perm_x,memPtes_3_perm_w,
    memPtes_3_perm_r,memPtes_2_perm_d,memPtes_2_perm_a,memPtes_2_perm_g,memPtes_2_perm_u}; // @[MMUBundle.scala 705:30]
  wire [9:0] data_hi_lo_hi_3 = {memPtes_7_perm_a,memPtes_7_perm_g,memPtes_7_perm_u,memPtes_7_perm_x,memPtes_7_perm_w,
    memPtes_7_perm_r,memPtes_6_perm_d,memPtes_6_perm_a,memPtes_6_perm_g,memPtes_6_perm_u}; // @[MMUBundle.scala 705:30]
  wire [18:0] data_hi_lo_3 = {data_hi_lo_hi_3,memPtes_6_perm_x,memPtes_6_perm_w,memPtes_6_perm_r,memPtes_5_perm_d,
    memPtes_5_perm_a,memPtes_5_perm_g,memPtes_5_perm_u,memPtes_5_perm_x,memPtes_5_perm_w}; // @[MMUBundle.scala 705:30]
  wire [229:0] data_hi_hi_hi_3 = {wdata_entries_ps_1_tag,io_csr_dup_2_satp_asid,memPtes_7_ppn,memPtes_6_ppn,
    memPtes_5_ppn,memPtes_4_ppn,memPtes_3_ppn,memPtes_2_ppn,memPtes_1_ppn,memPtes_0_ppn}; // @[MMUBundle.scala 705:30]
  wire [238:0] data_hi_hi_3 = {data_hi_hi_hi_3,wdata_entries_ps_1_vs_7,wdata_entries_ps_1_vs_6,wdata_entries_ps_1_vs_5,
    wdata_entries_ps_1_vs_4,wdata_entries_ps_1_vs_3,wdata_entries_ps_1_vs_2,wdata_entries_ps_1_vs_1,
    wdata_entries_ps_1_vs_0,memPtes_7_perm_d}; // @[MMUBundle.scala 705:30]
  wire [294:0] data_6 = {data_hi_hi_3,data_hi_lo_3,data_lo_hi_3,data_lo_lo_3}; // @[MMUBundle.scala 705:30]
  wire [63:0] _ecc_slices_0_syndromeUInt_T_21 = 64'hab55555556aaad5b & data_6[63:0]; // @[ECC.scala 147:74]
  wire  _ecc_slices_0_syndromeUInt_T_22 = ^_ecc_slices_0_syndromeUInt_T_21; // @[ECC.scala 147:79]
  wire [63:0] _ecc_slices_0_syndromeUInt_T_24 = 64'hcd9999999b33366d & data_6[63:0]; // @[ECC.scala 147:74]
  wire  _ecc_slices_0_syndromeUInt_T_25 = ^_ecc_slices_0_syndromeUInt_T_24; // @[ECC.scala 147:79]
  wire [63:0] _ecc_slices_0_syndromeUInt_T_27 = 64'hf1e1e1e1e3c3c78e & data_6[63:0]; // @[ECC.scala 147:74]
  wire  _ecc_slices_0_syndromeUInt_T_28 = ^_ecc_slices_0_syndromeUInt_T_27; // @[ECC.scala 147:79]
  wire [63:0] _ecc_slices_0_syndromeUInt_T_30 = 64'h1fe01fe03fc07f0 & data_6[63:0]; // @[ECC.scala 147:74]
  wire  _ecc_slices_0_syndromeUInt_T_31 = ^_ecc_slices_0_syndromeUInt_T_30; // @[ECC.scala 147:79]
  wire [63:0] _ecc_slices_0_syndromeUInt_T_33 = 64'h1fffe0003fff800 & data_6[63:0]; // @[ECC.scala 147:74]
  wire  _ecc_slices_0_syndromeUInt_T_34 = ^_ecc_slices_0_syndromeUInt_T_33; // @[ECC.scala 147:79]
  wire [63:0] _ecc_slices_0_syndromeUInt_T_36 = 64'h1fffffffc000000 & data_6[63:0]; // @[ECC.scala 147:74]
  wire  _ecc_slices_0_syndromeUInt_T_37 = ^_ecc_slices_0_syndromeUInt_T_36; // @[ECC.scala 147:79]
  wire [63:0] _ecc_slices_0_syndromeUInt_T_39 = 64'hfe00000000000000 & data_6[63:0]; // @[ECC.scala 147:74]
  wire  _ecc_slices_0_syndromeUInt_T_40 = ^_ecc_slices_0_syndromeUInt_T_39; // @[ECC.scala 147:79]
  wire [70:0] _ecc_slices_0_T_8 = {_ecc_slices_0_syndromeUInt_T_40,_ecc_slices_0_syndromeUInt_T_37,
    _ecc_slices_0_syndromeUInt_T_34,_ecc_slices_0_syndromeUInt_T_31,_ecc_slices_0_syndromeUInt_T_28,
    _ecc_slices_0_syndromeUInt_T_25,_ecc_slices_0_syndromeUInt_T_22,data_6[63:0]}; // @[Cat.scala 31:58]
  wire  _ecc_slices_0_T_9 = ^_ecc_slices_0_T_8; // @[ECC.scala 81:55]
  wire [71:0] _ecc_slices_0_T_11 = {_ecc_slices_0_T_9,_ecc_slices_0_syndromeUInt_T_40,_ecc_slices_0_syndromeUInt_T_37,
    _ecc_slices_0_syndromeUInt_T_34,_ecc_slices_0_syndromeUInt_T_31,_ecc_slices_0_syndromeUInt_T_28,
    _ecc_slices_0_syndromeUInt_T_25,_ecc_slices_0_syndromeUInt_T_22,data_6[63:0]}; // @[Cat.scala 31:58]
  wire [7:0] ecc_slices_1_0 = _ecc_slices_0_T_11[71:64]; // @[MMUBundle.scala 708:77]
  wire [63:0] _ecc_slices_1_syndromeUInt_T_21 = 64'hab55555556aaad5b & data_6[127:64]; // @[ECC.scala 147:74]
  wire  _ecc_slices_1_syndromeUInt_T_22 = ^_ecc_slices_1_syndromeUInt_T_21; // @[ECC.scala 147:79]
  wire [63:0] _ecc_slices_1_syndromeUInt_T_24 = 64'hcd9999999b33366d & data_6[127:64]; // @[ECC.scala 147:74]
  wire  _ecc_slices_1_syndromeUInt_T_25 = ^_ecc_slices_1_syndromeUInt_T_24; // @[ECC.scala 147:79]
  wire [63:0] _ecc_slices_1_syndromeUInt_T_27 = 64'hf1e1e1e1e3c3c78e & data_6[127:64]; // @[ECC.scala 147:74]
  wire  _ecc_slices_1_syndromeUInt_T_28 = ^_ecc_slices_1_syndromeUInt_T_27; // @[ECC.scala 147:79]
  wire [63:0] _ecc_slices_1_syndromeUInt_T_30 = 64'h1fe01fe03fc07f0 & data_6[127:64]; // @[ECC.scala 147:74]
  wire  _ecc_slices_1_syndromeUInt_T_31 = ^_ecc_slices_1_syndromeUInt_T_30; // @[ECC.scala 147:79]
  wire [63:0] _ecc_slices_1_syndromeUInt_T_33 = 64'h1fffe0003fff800 & data_6[127:64]; // @[ECC.scala 147:74]
  wire  _ecc_slices_1_syndromeUInt_T_34 = ^_ecc_slices_1_syndromeUInt_T_33; // @[ECC.scala 147:79]
  wire [63:0] _ecc_slices_1_syndromeUInt_T_36 = 64'h1fffffffc000000 & data_6[127:64]; // @[ECC.scala 147:74]
  wire  _ecc_slices_1_syndromeUInt_T_37 = ^_ecc_slices_1_syndromeUInt_T_36; // @[ECC.scala 147:79]
  wire [63:0] _ecc_slices_1_syndromeUInt_T_39 = 64'hfe00000000000000 & data_6[127:64]; // @[ECC.scala 147:74]
  wire  _ecc_slices_1_syndromeUInt_T_40 = ^_ecc_slices_1_syndromeUInt_T_39; // @[ECC.scala 147:79]
  wire [70:0] _ecc_slices_1_T_8 = {_ecc_slices_1_syndromeUInt_T_40,_ecc_slices_1_syndromeUInt_T_37,
    _ecc_slices_1_syndromeUInt_T_34,_ecc_slices_1_syndromeUInt_T_31,_ecc_slices_1_syndromeUInt_T_28,
    _ecc_slices_1_syndromeUInt_T_25,_ecc_slices_1_syndromeUInt_T_22,data_6[127:64]}; // @[Cat.scala 31:58]
  wire  _ecc_slices_1_T_9 = ^_ecc_slices_1_T_8; // @[ECC.scala 81:55]
  wire [71:0] _ecc_slices_1_T_11 = {_ecc_slices_1_T_9,_ecc_slices_1_syndromeUInt_T_40,_ecc_slices_1_syndromeUInt_T_37,
    _ecc_slices_1_syndromeUInt_T_34,_ecc_slices_1_syndromeUInt_T_31,_ecc_slices_1_syndromeUInt_T_28,
    _ecc_slices_1_syndromeUInt_T_25,_ecc_slices_1_syndromeUInt_T_22,data_6[127:64]}; // @[Cat.scala 31:58]
  wire [7:0] ecc_slices_1_1 = _ecc_slices_1_T_11[71:64]; // @[MMUBundle.scala 708:77]
  wire [63:0] _ecc_slices_2_syndromeUInt_T_21 = 64'hab55555556aaad5b & data_6[191:128]; // @[ECC.scala 147:74]
  wire  _ecc_slices_2_syndromeUInt_T_22 = ^_ecc_slices_2_syndromeUInt_T_21; // @[ECC.scala 147:79]
  wire [63:0] _ecc_slices_2_syndromeUInt_T_24 = 64'hcd9999999b33366d & data_6[191:128]; // @[ECC.scala 147:74]
  wire  _ecc_slices_2_syndromeUInt_T_25 = ^_ecc_slices_2_syndromeUInt_T_24; // @[ECC.scala 147:79]
  wire [63:0] _ecc_slices_2_syndromeUInt_T_27 = 64'hf1e1e1e1e3c3c78e & data_6[191:128]; // @[ECC.scala 147:74]
  wire  _ecc_slices_2_syndromeUInt_T_28 = ^_ecc_slices_2_syndromeUInt_T_27; // @[ECC.scala 147:79]
  wire [63:0] _ecc_slices_2_syndromeUInt_T_30 = 64'h1fe01fe03fc07f0 & data_6[191:128]; // @[ECC.scala 147:74]
  wire  _ecc_slices_2_syndromeUInt_T_31 = ^_ecc_slices_2_syndromeUInt_T_30; // @[ECC.scala 147:79]
  wire [63:0] _ecc_slices_2_syndromeUInt_T_33 = 64'h1fffe0003fff800 & data_6[191:128]; // @[ECC.scala 147:74]
  wire  _ecc_slices_2_syndromeUInt_T_34 = ^_ecc_slices_2_syndromeUInt_T_33; // @[ECC.scala 147:79]
  wire [63:0] _ecc_slices_2_syndromeUInt_T_36 = 64'h1fffffffc000000 & data_6[191:128]; // @[ECC.scala 147:74]
  wire  _ecc_slices_2_syndromeUInt_T_37 = ^_ecc_slices_2_syndromeUInt_T_36; // @[ECC.scala 147:79]
  wire [63:0] _ecc_slices_2_syndromeUInt_T_39 = 64'hfe00000000000000 & data_6[191:128]; // @[ECC.scala 147:74]
  wire  _ecc_slices_2_syndromeUInt_T_40 = ^_ecc_slices_2_syndromeUInt_T_39; // @[ECC.scala 147:79]
  wire [70:0] _ecc_slices_2_T_8 = {_ecc_slices_2_syndromeUInt_T_40,_ecc_slices_2_syndromeUInt_T_37,
    _ecc_slices_2_syndromeUInt_T_34,_ecc_slices_2_syndromeUInt_T_31,_ecc_slices_2_syndromeUInt_T_28,
    _ecc_slices_2_syndromeUInt_T_25,_ecc_slices_2_syndromeUInt_T_22,data_6[191:128]}; // @[Cat.scala 31:58]
  wire  _ecc_slices_2_T_9 = ^_ecc_slices_2_T_8; // @[ECC.scala 81:55]
  wire [71:0] _ecc_slices_2_T_11 = {_ecc_slices_2_T_9,_ecc_slices_2_syndromeUInt_T_40,_ecc_slices_2_syndromeUInt_T_37,
    _ecc_slices_2_syndromeUInt_T_34,_ecc_slices_2_syndromeUInt_T_31,_ecc_slices_2_syndromeUInt_T_28,
    _ecc_slices_2_syndromeUInt_T_25,_ecc_slices_2_syndromeUInt_T_22,data_6[191:128]}; // @[Cat.scala 31:58]
  wire [7:0] ecc_slices_1_2 = _ecc_slices_2_T_11[71:64]; // @[MMUBundle.scala 708:77]
  wire [63:0] _ecc_slices_3_syndromeUInt_T = 64'hab55555556aaad5b & data_6[255:192]; // @[ECC.scala 147:74]
  wire  _ecc_slices_3_syndromeUInt_T_1 = ^_ecc_slices_3_syndromeUInt_T; // @[ECC.scala 147:79]
  wire [63:0] _ecc_slices_3_syndromeUInt_T_3 = 64'hcd9999999b33366d & data_6[255:192]; // @[ECC.scala 147:74]
  wire  _ecc_slices_3_syndromeUInt_T_4 = ^_ecc_slices_3_syndromeUInt_T_3; // @[ECC.scala 147:79]
  wire [63:0] _ecc_slices_3_syndromeUInt_T_6 = 64'hf1e1e1e1e3c3c78e & data_6[255:192]; // @[ECC.scala 147:74]
  wire  _ecc_slices_3_syndromeUInt_T_7 = ^_ecc_slices_3_syndromeUInt_T_6; // @[ECC.scala 147:79]
  wire [63:0] _ecc_slices_3_syndromeUInt_T_9 = 64'h1fe01fe03fc07f0 & data_6[255:192]; // @[ECC.scala 147:74]
  wire  _ecc_slices_3_syndromeUInt_T_10 = ^_ecc_slices_3_syndromeUInt_T_9; // @[ECC.scala 147:79]
  wire [63:0] _ecc_slices_3_syndromeUInt_T_12 = 64'h1fffe0003fff800 & data_6[255:192]; // @[ECC.scala 147:74]
  wire  _ecc_slices_3_syndromeUInt_T_13 = ^_ecc_slices_3_syndromeUInt_T_12; // @[ECC.scala 147:79]
  wire [63:0] _ecc_slices_3_syndromeUInt_T_15 = 64'h1fffffffc000000 & data_6[255:192]; // @[ECC.scala 147:74]
  wire  _ecc_slices_3_syndromeUInt_T_16 = ^_ecc_slices_3_syndromeUInt_T_15; // @[ECC.scala 147:79]
  wire [63:0] _ecc_slices_3_syndromeUInt_T_18 = 64'hfe00000000000000 & data_6[255:192]; // @[ECC.scala 147:74]
  wire  _ecc_slices_3_syndromeUInt_T_19 = ^_ecc_slices_3_syndromeUInt_T_18; // @[ECC.scala 147:79]
  wire [70:0] _ecc_slices_3_T_1 = {_ecc_slices_3_syndromeUInt_T_19,_ecc_slices_3_syndromeUInt_T_16,
    _ecc_slices_3_syndromeUInt_T_13,_ecc_slices_3_syndromeUInt_T_10,_ecc_slices_3_syndromeUInt_T_7,
    _ecc_slices_3_syndromeUInt_T_4,_ecc_slices_3_syndromeUInt_T_1,data_6[255:192]}; // @[Cat.scala 31:58]
  wire  _ecc_slices_3_T_2 = ^_ecc_slices_3_T_1; // @[ECC.scala 81:55]
  wire [71:0] _ecc_slices_3_T_4 = {_ecc_slices_3_T_2,_ecc_slices_3_syndromeUInt_T_19,_ecc_slices_3_syndromeUInt_T_16,
    _ecc_slices_3_syndromeUInt_T_13,_ecc_slices_3_syndromeUInt_T_10,_ecc_slices_3_syndromeUInt_T_7,
    _ecc_slices_3_syndromeUInt_T_4,_ecc_slices_3_syndromeUInt_T_1,data_6[255:192]}; // @[Cat.scala 31:58]
  wire [7:0] ecc_slices_1_3 = _ecc_slices_3_T_4[71:64]; // @[MMUBundle.scala 708:77]
  wire [38:0] _ecc_unaligned_syndromeUInt_T_18 = 39'h5556aaad5b & data_6[294:256]; // @[ECC.scala 147:74]
  wire  _ecc_unaligned_syndromeUInt_T_19 = ^_ecc_unaligned_syndromeUInt_T_18; // @[ECC.scala 147:79]
  wire [38:0] _ecc_unaligned_syndromeUInt_T_21 = 39'h199b33366d & data_6[294:256]; // @[ECC.scala 147:74]
  wire  _ecc_unaligned_syndromeUInt_T_22 = ^_ecc_unaligned_syndromeUInt_T_21; // @[ECC.scala 147:79]
  wire [38:0] _ecc_unaligned_syndromeUInt_T_24 = 39'h61e3c3c78e & data_6[294:256]; // @[ECC.scala 147:74]
  wire  _ecc_unaligned_syndromeUInt_T_25 = ^_ecc_unaligned_syndromeUInt_T_24; // @[ECC.scala 147:79]
  wire [38:0] _ecc_unaligned_syndromeUInt_T_27 = 39'h7e03fc07f0 & data_6[294:256]; // @[ECC.scala 147:74]
  wire  _ecc_unaligned_syndromeUInt_T_28 = ^_ecc_unaligned_syndromeUInt_T_27; // @[ECC.scala 147:79]
  wire [38:0] _ecc_unaligned_syndromeUInt_T_30 = 39'h3fff800 & data_6[294:256]; // @[ECC.scala 147:74]
  wire  _ecc_unaligned_syndromeUInt_T_31 = ^_ecc_unaligned_syndromeUInt_T_30; // @[ECC.scala 147:79]
  wire [38:0] _ecc_unaligned_syndromeUInt_T_33 = 39'h7ffc000000 & data_6[294:256]; // @[ECC.scala 147:74]
  wire  _ecc_unaligned_syndromeUInt_T_34 = ^_ecc_unaligned_syndromeUInt_T_33; // @[ECC.scala 147:79]
  wire [44:0] _ecc_unaligned_T_7 = {_ecc_unaligned_syndromeUInt_T_34,_ecc_unaligned_syndromeUInt_T_31,
    _ecc_unaligned_syndromeUInt_T_28,_ecc_unaligned_syndromeUInt_T_25,_ecc_unaligned_syndromeUInt_T_22,
    _ecc_unaligned_syndromeUInt_T_19,data_6[294:256]}; // @[Cat.scala 31:58]
  wire  _ecc_unaligned_T_8 = ^_ecc_unaligned_T_7; // @[ECC.scala 81:55]
  wire [45:0] _ecc_unaligned_T_10 = {_ecc_unaligned_T_8,_ecc_unaligned_syndromeUInt_T_34,
    _ecc_unaligned_syndromeUInt_T_31,_ecc_unaligned_syndromeUInt_T_28,_ecc_unaligned_syndromeUInt_T_25,
    _ecc_unaligned_syndromeUInt_T_22,_ecc_unaligned_syndromeUInt_T_19,data_6[294:256]}; // @[Cat.scala 31:58]
  wire [6:0] ecc_unaligned_1 = _ecc_unaligned_T_10[45:39]; // @[MMUBundle.scala 711:88]
  wire [31:0] _wdata_ecc_T_2 = {ecc_slices_1_3,ecc_slices_1_2,ecc_slices_1_1,ecc_slices_1_0}; // @[MMUBundle.scala 712:50]
  wire  state_vec_set_left_older_5 = ~l3_victimWay[2]; // @[Replacement.scala 196:33]
  wire  state_vec_set_left_older_6 = ~l3_victimWay[1]; // @[Replacement.scala 196:33]
  wire  _state_vec_T_44 = ~l3_victimWay[0]; // @[Replacement.scala 218:7]
  wire  _state_vec_T_45 = state_vec_set_left_older_6 ? victimWay_left_subtree_state_2 : _state_vec_T_44; // @[Replacement.scala 203:16]
  wire  _state_vec_T_49 = state_vec_set_left_older_6 ? _state_vec_T_44 : victimWay_right_subtree_state_2; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_T_50 = {state_vec_set_left_older_6,_state_vec_T_45,_state_vec_T_49}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_T_51 = state_vec_set_left_older_5 ? victimWay_left_subtree_state_1 : _state_vec_T_50; // @[Replacement.scala 203:16]
  wire  _state_vec_T_56 = state_vec_set_left_older_6 ? victimWay_left_subtree_state_3 : _state_vec_T_44; // @[Replacement.scala 203:16]
  wire  _state_vec_T_60 = state_vec_set_left_older_6 ? _state_vec_T_44 : victimWay_right_subtree_state_3; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_T_61 = {state_vec_set_left_older_6,_state_vec_T_56,_state_vec_T_60}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_T_62 = state_vec_set_left_older_5 ? _state_vec_T_61 : victimWay_right_subtree_state_1; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_T_63 = {state_vec_set_left_older_5,_state_vec_T_51,_state_vec_T_62}; // @[Cat.scala 31:58]
  wire [31:0] _l3v_T = l3v | l3_rfvOH; // @[PageTableCache.scala 520:16]
  wire [31:0] _l3g_T = ~l3_rfvOH; // @[PageTableCache.scala 521:18]
  wire [31:0] _l3g_T_1 = l3g & _l3g_T; // @[PageTableCache.scala 521:16]
  wire [31:0] _l3g_T_4 = _l2g_T_3 ? l3_rfvOH : 32'h0; // @[PageTableCache.scala 521:30]
  wire [31:0] _l3g_T_5 = _l3g_T_1 | _l3g_T_4; // @[PageTableCache.scala 521:25]
  wire [1:0] sp_rfOH = 2'h1 << state_reg_3; // @[OneHot.scala 57:35]
  wire  _state_reg_T_21 = ~state_reg_3; // @[Replacement.scala 218:7]
  wire [1:0] _spv_T = spv | sp_rfOH; // @[PageTableCache.scala 552:16]
  wire [1:0] _spg_T = ~sp_rfOH; // @[PageTableCache.scala 553:18]
  wire [1:0] _spg_T_1 = spg & _spg_T; // @[PageTableCache.scala 553:16]
  wire [1:0] _spg_T_2 = memPte_0_perm_g ? sp_rfOH : 2'h0; // @[PageTableCache.scala 553:29]
  wire [1:0] _spg_T_3 = _spg_T_1 | _spg_T_2; // @[PageTableCache.scala 553:24]
  wire  l2eccFlush = resp_res_l2_ecc & stageResp_valid_1cycle_dup_0_valid; // @[PageTableCache.scala 566:36]
  wire  l3eccFlush = resp_res_l3_ecc & stageResp_valid_1cycle_dup_1_valid; // @[PageTableCache.scala 567:36]
  wire [3:0] flushSetIdxOH = 4'h1 << data_2_req_info_vpn[13:12]; // @[OneHot.scala 57:35]
  wire [3:0] _flushMask_T_5 = flushSetIdxOH[0] ? 4'hf : 4'h0; // @[Bitwise.scala 74:12]
  wire [3:0] _flushMask_T_7 = flushSetIdxOH[1] ? 4'hf : 4'h0; // @[Bitwise.scala 74:12]
  wire [3:0] _flushMask_T_9 = flushSetIdxOH[2] ? 4'hf : 4'h0; // @[Bitwise.scala 74:12]
  wire [3:0] _flushMask_T_11 = flushSetIdxOH[3] ? 4'hf : 4'h0; // @[Bitwise.scala 74:12]
  wire [15:0] flushMask = {_flushMask_T_11,_flushMask_T_9,_flushMask_T_7,_flushMask_T_5}; // @[PageTableCache.scala 574:101]
  wire [15:0] _l2v_T_1 = ~flushMask; // @[PageTableCache.scala 575:18]
  wire [15:0] _l2v_T_2 = l2v & _l2v_T_1; // @[PageTableCache.scala 575:16]
  wire [15:0] _l2g_T_7 = l2g & _l2v_T_1; // @[PageTableCache.scala 576:16]
  wire [15:0] _GEN_2533 = l2eccFlush ? _l2v_T_2 : _GEN_1833; // @[PageTableCache.scala 572:21 575:9]
  wire [3:0] flushSetIdxOH_1 = 4'h1 << data_2_req_info_vpn[4:3]; // @[OneHot.scala 57:35]
  wire [7:0] _flushMask_T_17 = flushSetIdxOH_1[0] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _flushMask_T_19 = flushSetIdxOH_1[1] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _flushMask_T_21 = flushSetIdxOH_1[2] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _flushMask_T_23 = flushSetIdxOH_1[3] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [31:0] flushMask_1 = {_flushMask_T_23,_flushMask_T_21,_flushMask_T_19,_flushMask_T_17}; // @[PageTableCache.scala 581:101]
  wire [31:0] _l3v_T_1 = ~flushMask_1; // @[PageTableCache.scala 582:18]
  wire [31:0] _l3v_T_2 = l3v & _l3v_T_1; // @[PageTableCache.scala 582:16]
  wire [31:0] _l3g_T_7 = l3g & _l3v_T_1; // @[PageTableCache.scala 583:16]
  wire [26:0] sfence_vpn = io_sfence_dup_3_bits_addr[38:12]; // @[PageTableCache.scala 588:45]
  wire [31:0] _l3v_T_3 = l3v & l3g; // @[PageTableCache.scala 596:20]
  wire [3:0] sfence_nrs1_flushSetIdxOH = 4'h1 << sfence_vpn[4:3]; // @[OneHot.scala 57:35]
  wire [7:0] _flushMask_T_29 = sfence_nrs1_flushSetIdxOH[0] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _flushMask_T_31 = sfence_nrs1_flushSetIdxOH[1] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _flushMask_T_33 = sfence_nrs1_flushSetIdxOH[2] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [7:0] _flushMask_T_35 = sfence_nrs1_flushSetIdxOH[3] ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [31:0] sfence_nrs1_flushMask = {_flushMask_T_35,_flushMask_T_33,_flushMask_T_31,_flushMask_T_29}; // @[PageTableCache.scala 602:103]
  wire [31:0] _l3v_T_4 = ~sfence_nrs1_flushMask; // @[PageTableCache.scala 608:22]
  wire [31:0] _l3v_T_5 = l3v & _l3v_T_4; // @[PageTableCache.scala 608:20]
  wire [31:0] _l3v_T_7 = _l3v_T_4 | l3g; // @[PageTableCache.scala 611:34]
  wire [31:0] _l3v_T_8 = l3v & _l3v_T_7; // @[PageTableCache.scala 611:20]
  wire [3:0] l1asidhit = {l1_3_asid == io_sfence_dup_0_bits_asid,l1_2_asid == io_sfence_dup_0_bits_asid,l1_1_asid ==
    io_sfence_dup_0_bits_asid,l1_0_asid == io_sfence_dup_0_bits_asid}; // @[PageTableCache.scala 617:73]
  wire  _spasidhit_T = sp_0_asid == io_sfence_dup_0_bits_asid; // @[PageTableCache.scala 618:43]
  wire  _spasidhit_T_1 = sp_1_asid == io_sfence_dup_0_bits_asid; // @[PageTableCache.scala 618:43]
  wire [1:0] spasidhit = {sp_1_asid == io_sfence_dup_0_bits_asid,sp_0_asid == io_sfence_dup_0_bits_asid}; // @[PageTableCache.scala 618:73]
  wire [26:0] sfence_vpn_1 = io_sfence_dup_0_bits_addr[38:12]; // @[PageTableCache.scala 619:45]
  wire [3:0] _l1v_T_1 = ~l1asidhit; // @[PageTableCache.scala 630:23]
  wire [3:0] _l1v_T_2 = _l1v_T_1 | l1g; // @[PageTableCache.scala 630:34]
  wire [3:0] _l1v_T_3 = l1v & _l1v_T_2; // @[PageTableCache.scala 630:20]
  wire [15:0] _l2v_T_3 = l2v & l2g; // @[PageTableCache.scala 631:20]
  wire [1:0] _spv_T_1 = ~spasidhit; // @[PageTableCache.scala 632:23]
  wire [1:0] _spv_T_2 = _spv_T_1 | spg; // @[PageTableCache.scala 632:34]
  wire [1:0] _spv_T_3 = spv & _spv_T_2; // @[PageTableCache.scala 632:20]
  wire  spv_hit0 = sp_0_tag[17:9] == sfence_vpn_1[26:18]; // @[MMUBundle.scala 587:52]
  wire  spv_hit1 = sp_0_tag[8:0] == sfence_vpn_1[17:9]; // @[MMUBundle.scala 588:66]
  wire  _spv_T_6 = sp_0_level == 2'h0 ? spv_hit0 : spv_hit0 & spv_hit1; // @[MMUBundle.scala 590:22]
  wire  spv_hit0_1 = sp_1_tag[17:9] == sfence_vpn_1[26:18]; // @[MMUBundle.scala 587:52]
  wire  spv_hit1_1 = sp_1_tag[8:0] == sfence_vpn_1[17:9]; // @[MMUBundle.scala 588:66]
  wire  _spv_T_10 = sp_1_level == 2'h0 ? spv_hit0_1 : spv_hit0_1 & spv_hit1_1; // @[MMUBundle.scala 590:22]
  wire [1:0] _spv_T_12 = {_spv_T_10,_spv_T_6}; // @[PageTableCache.scala 644:103]
  wire [1:0] _spv_T_13 = ~_spv_T_12; // @[PageTableCache.scala 644:23]
  wire [1:0] _spv_T_14 = spv & _spv_T_13; // @[PageTableCache.scala 644:20]
  wire  _spv_T_18 = _spasidhit_T & _spv_T_6; // @[MMUBundle.scala 590:16]
  wire  _spv_T_22 = _spasidhit_T_1 & _spv_T_10; // @[MMUBundle.scala 590:16]
  wire [1:0] _spv_T_23 = {_spv_T_22,_spv_T_18}; // @[PageTableCache.scala 647:84]
  wire [1:0] _spv_T_24 = ~_spv_T_23; // @[PageTableCache.scala 647:23]
  wire [1:0] _spv_T_25 = _spv_T_24 | spg; // @[PageTableCache.scala 647:91]
  wire [1:0] _spv_T_26 = spv & _spv_T_25; // @[PageTableCache.scala 647:20]
  wire  _base_valid_access_0_T = io_resp_bits_req_info_source == 2'h2; // @[MMUConst.scala 254:13]
  wire  _base_valid_access_0_T_2 = io_resp_ready & io_resp_valid; // @[Decoupled.scala 50:35]
  wire  _T_565 = ~io_req_ready; // @[PageTableCache.scala 729:48]
  wire  _T_567 = ~io_resp_ready; // @[PageTableCache.scala 730:52]
  reg  io_perf_0_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg  io_perf_0_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg  io_perf_1_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg  io_perf_1_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg  io_perf_2_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg  io_perf_2_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg  io_perf_3_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg  io_perf_3_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg  io_perf_4_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg  io_perf_4_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg  io_perf_5_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg  io_perf_5_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg  io_perf_6_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg  io_perf_6_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg  io_perf_7_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg  io_perf_7_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  SRAMTemplate_68 l2 ( // @[PageTableCache.scala 155:18]
    .clock(l2_clock),
    .io_rreq_valid(l2_io_rreq_valid),
    .io_rreq_bits_setIdx(l2_io_rreq_bits_setIdx),
    .io_rresp_data_0_entries_tag(l2_io_rresp_data_0_entries_tag),
    .io_rresp_data_0_entries_asid(l2_io_rresp_data_0_entries_asid),
    .io_rresp_data_0_entries_ppns_0(l2_io_rresp_data_0_entries_ppns_0),
    .io_rresp_data_0_entries_ppns_1(l2_io_rresp_data_0_entries_ppns_1),
    .io_rresp_data_0_entries_ppns_2(l2_io_rresp_data_0_entries_ppns_2),
    .io_rresp_data_0_entries_ppns_3(l2_io_rresp_data_0_entries_ppns_3),
    .io_rresp_data_0_entries_ppns_4(l2_io_rresp_data_0_entries_ppns_4),
    .io_rresp_data_0_entries_ppns_5(l2_io_rresp_data_0_entries_ppns_5),
    .io_rresp_data_0_entries_ppns_6(l2_io_rresp_data_0_entries_ppns_6),
    .io_rresp_data_0_entries_ppns_7(l2_io_rresp_data_0_entries_ppns_7),
    .io_rresp_data_0_entries_vs_0(l2_io_rresp_data_0_entries_vs_0),
    .io_rresp_data_0_entries_vs_1(l2_io_rresp_data_0_entries_vs_1),
    .io_rresp_data_0_entries_vs_2(l2_io_rresp_data_0_entries_vs_2),
    .io_rresp_data_0_entries_vs_3(l2_io_rresp_data_0_entries_vs_3),
    .io_rresp_data_0_entries_vs_4(l2_io_rresp_data_0_entries_vs_4),
    .io_rresp_data_0_entries_vs_5(l2_io_rresp_data_0_entries_vs_5),
    .io_rresp_data_0_entries_vs_6(l2_io_rresp_data_0_entries_vs_6),
    .io_rresp_data_0_entries_vs_7(l2_io_rresp_data_0_entries_vs_7),
    .io_rresp_data_0_entries_prefetch(l2_io_rresp_data_0_entries_prefetch),
    .io_rresp_data_0_ecc(l2_io_rresp_data_0_ecc),
    .io_rresp_data_1_entries_tag(l2_io_rresp_data_1_entries_tag),
    .io_rresp_data_1_entries_asid(l2_io_rresp_data_1_entries_asid),
    .io_rresp_data_1_entries_ppns_0(l2_io_rresp_data_1_entries_ppns_0),
    .io_rresp_data_1_entries_ppns_1(l2_io_rresp_data_1_entries_ppns_1),
    .io_rresp_data_1_entries_ppns_2(l2_io_rresp_data_1_entries_ppns_2),
    .io_rresp_data_1_entries_ppns_3(l2_io_rresp_data_1_entries_ppns_3),
    .io_rresp_data_1_entries_ppns_4(l2_io_rresp_data_1_entries_ppns_4),
    .io_rresp_data_1_entries_ppns_5(l2_io_rresp_data_1_entries_ppns_5),
    .io_rresp_data_1_entries_ppns_6(l2_io_rresp_data_1_entries_ppns_6),
    .io_rresp_data_1_entries_ppns_7(l2_io_rresp_data_1_entries_ppns_7),
    .io_rresp_data_1_entries_vs_0(l2_io_rresp_data_1_entries_vs_0),
    .io_rresp_data_1_entries_vs_1(l2_io_rresp_data_1_entries_vs_1),
    .io_rresp_data_1_entries_vs_2(l2_io_rresp_data_1_entries_vs_2),
    .io_rresp_data_1_entries_vs_3(l2_io_rresp_data_1_entries_vs_3),
    .io_rresp_data_1_entries_vs_4(l2_io_rresp_data_1_entries_vs_4),
    .io_rresp_data_1_entries_vs_5(l2_io_rresp_data_1_entries_vs_5),
    .io_rresp_data_1_entries_vs_6(l2_io_rresp_data_1_entries_vs_6),
    .io_rresp_data_1_entries_vs_7(l2_io_rresp_data_1_entries_vs_7),
    .io_rresp_data_1_entries_prefetch(l2_io_rresp_data_1_entries_prefetch),
    .io_rresp_data_1_ecc(l2_io_rresp_data_1_ecc),
    .io_rresp_data_2_entries_tag(l2_io_rresp_data_2_entries_tag),
    .io_rresp_data_2_entries_asid(l2_io_rresp_data_2_entries_asid),
    .io_rresp_data_2_entries_ppns_0(l2_io_rresp_data_2_entries_ppns_0),
    .io_rresp_data_2_entries_ppns_1(l2_io_rresp_data_2_entries_ppns_1),
    .io_rresp_data_2_entries_ppns_2(l2_io_rresp_data_2_entries_ppns_2),
    .io_rresp_data_2_entries_ppns_3(l2_io_rresp_data_2_entries_ppns_3),
    .io_rresp_data_2_entries_ppns_4(l2_io_rresp_data_2_entries_ppns_4),
    .io_rresp_data_2_entries_ppns_5(l2_io_rresp_data_2_entries_ppns_5),
    .io_rresp_data_2_entries_ppns_6(l2_io_rresp_data_2_entries_ppns_6),
    .io_rresp_data_2_entries_ppns_7(l2_io_rresp_data_2_entries_ppns_7),
    .io_rresp_data_2_entries_vs_0(l2_io_rresp_data_2_entries_vs_0),
    .io_rresp_data_2_entries_vs_1(l2_io_rresp_data_2_entries_vs_1),
    .io_rresp_data_2_entries_vs_2(l2_io_rresp_data_2_entries_vs_2),
    .io_rresp_data_2_entries_vs_3(l2_io_rresp_data_2_entries_vs_3),
    .io_rresp_data_2_entries_vs_4(l2_io_rresp_data_2_entries_vs_4),
    .io_rresp_data_2_entries_vs_5(l2_io_rresp_data_2_entries_vs_5),
    .io_rresp_data_2_entries_vs_6(l2_io_rresp_data_2_entries_vs_6),
    .io_rresp_data_2_entries_vs_7(l2_io_rresp_data_2_entries_vs_7),
    .io_rresp_data_2_entries_prefetch(l2_io_rresp_data_2_entries_prefetch),
    .io_rresp_data_2_ecc(l2_io_rresp_data_2_ecc),
    .io_rresp_data_3_entries_tag(l2_io_rresp_data_3_entries_tag),
    .io_rresp_data_3_entries_asid(l2_io_rresp_data_3_entries_asid),
    .io_rresp_data_3_entries_ppns_0(l2_io_rresp_data_3_entries_ppns_0),
    .io_rresp_data_3_entries_ppns_1(l2_io_rresp_data_3_entries_ppns_1),
    .io_rresp_data_3_entries_ppns_2(l2_io_rresp_data_3_entries_ppns_2),
    .io_rresp_data_3_entries_ppns_3(l2_io_rresp_data_3_entries_ppns_3),
    .io_rresp_data_3_entries_ppns_4(l2_io_rresp_data_3_entries_ppns_4),
    .io_rresp_data_3_entries_ppns_5(l2_io_rresp_data_3_entries_ppns_5),
    .io_rresp_data_3_entries_ppns_6(l2_io_rresp_data_3_entries_ppns_6),
    .io_rresp_data_3_entries_ppns_7(l2_io_rresp_data_3_entries_ppns_7),
    .io_rresp_data_3_entries_vs_0(l2_io_rresp_data_3_entries_vs_0),
    .io_rresp_data_3_entries_vs_1(l2_io_rresp_data_3_entries_vs_1),
    .io_rresp_data_3_entries_vs_2(l2_io_rresp_data_3_entries_vs_2),
    .io_rresp_data_3_entries_vs_3(l2_io_rresp_data_3_entries_vs_3),
    .io_rresp_data_3_entries_vs_4(l2_io_rresp_data_3_entries_vs_4),
    .io_rresp_data_3_entries_vs_5(l2_io_rresp_data_3_entries_vs_5),
    .io_rresp_data_3_entries_vs_6(l2_io_rresp_data_3_entries_vs_6),
    .io_rresp_data_3_entries_vs_7(l2_io_rresp_data_3_entries_vs_7),
    .io_rresp_data_3_entries_prefetch(l2_io_rresp_data_3_entries_prefetch),
    .io_rresp_data_3_ecc(l2_io_rresp_data_3_ecc),
    .io_wreq_valid(l2_io_wreq_valid),
    .io_wreq_bits_setIdx(l2_io_wreq_bits_setIdx),
    .io_wreq_bits_data_0_entries_tag(l2_io_wreq_bits_data_0_entries_tag),
    .io_wreq_bits_data_0_entries_asid(l2_io_wreq_bits_data_0_entries_asid),
    .io_wreq_bits_data_0_entries_ppns_0(l2_io_wreq_bits_data_0_entries_ppns_0),
    .io_wreq_bits_data_0_entries_ppns_1(l2_io_wreq_bits_data_0_entries_ppns_1),
    .io_wreq_bits_data_0_entries_ppns_2(l2_io_wreq_bits_data_0_entries_ppns_2),
    .io_wreq_bits_data_0_entries_ppns_3(l2_io_wreq_bits_data_0_entries_ppns_3),
    .io_wreq_bits_data_0_entries_ppns_4(l2_io_wreq_bits_data_0_entries_ppns_4),
    .io_wreq_bits_data_0_entries_ppns_5(l2_io_wreq_bits_data_0_entries_ppns_5),
    .io_wreq_bits_data_0_entries_ppns_6(l2_io_wreq_bits_data_0_entries_ppns_6),
    .io_wreq_bits_data_0_entries_ppns_7(l2_io_wreq_bits_data_0_entries_ppns_7),
    .io_wreq_bits_data_0_entries_vs_0(l2_io_wreq_bits_data_0_entries_vs_0),
    .io_wreq_bits_data_0_entries_vs_1(l2_io_wreq_bits_data_0_entries_vs_1),
    .io_wreq_bits_data_0_entries_vs_2(l2_io_wreq_bits_data_0_entries_vs_2),
    .io_wreq_bits_data_0_entries_vs_3(l2_io_wreq_bits_data_0_entries_vs_3),
    .io_wreq_bits_data_0_entries_vs_4(l2_io_wreq_bits_data_0_entries_vs_4),
    .io_wreq_bits_data_0_entries_vs_5(l2_io_wreq_bits_data_0_entries_vs_5),
    .io_wreq_bits_data_0_entries_vs_6(l2_io_wreq_bits_data_0_entries_vs_6),
    .io_wreq_bits_data_0_entries_vs_7(l2_io_wreq_bits_data_0_entries_vs_7),
    .io_wreq_bits_data_0_entries_prefetch(l2_io_wreq_bits_data_0_entries_prefetch),
    .io_wreq_bits_data_0_ecc(l2_io_wreq_bits_data_0_ecc),
    .io_wreq_bits_data_1_entries_tag(l2_io_wreq_bits_data_1_entries_tag),
    .io_wreq_bits_data_1_entries_asid(l2_io_wreq_bits_data_1_entries_asid),
    .io_wreq_bits_data_1_entries_ppns_0(l2_io_wreq_bits_data_1_entries_ppns_0),
    .io_wreq_bits_data_1_entries_ppns_1(l2_io_wreq_bits_data_1_entries_ppns_1),
    .io_wreq_bits_data_1_entries_ppns_2(l2_io_wreq_bits_data_1_entries_ppns_2),
    .io_wreq_bits_data_1_entries_ppns_3(l2_io_wreq_bits_data_1_entries_ppns_3),
    .io_wreq_bits_data_1_entries_ppns_4(l2_io_wreq_bits_data_1_entries_ppns_4),
    .io_wreq_bits_data_1_entries_ppns_5(l2_io_wreq_bits_data_1_entries_ppns_5),
    .io_wreq_bits_data_1_entries_ppns_6(l2_io_wreq_bits_data_1_entries_ppns_6),
    .io_wreq_bits_data_1_entries_ppns_7(l2_io_wreq_bits_data_1_entries_ppns_7),
    .io_wreq_bits_data_1_entries_vs_0(l2_io_wreq_bits_data_1_entries_vs_0),
    .io_wreq_bits_data_1_entries_vs_1(l2_io_wreq_bits_data_1_entries_vs_1),
    .io_wreq_bits_data_1_entries_vs_2(l2_io_wreq_bits_data_1_entries_vs_2),
    .io_wreq_bits_data_1_entries_vs_3(l2_io_wreq_bits_data_1_entries_vs_3),
    .io_wreq_bits_data_1_entries_vs_4(l2_io_wreq_bits_data_1_entries_vs_4),
    .io_wreq_bits_data_1_entries_vs_5(l2_io_wreq_bits_data_1_entries_vs_5),
    .io_wreq_bits_data_1_entries_vs_6(l2_io_wreq_bits_data_1_entries_vs_6),
    .io_wreq_bits_data_1_entries_vs_7(l2_io_wreq_bits_data_1_entries_vs_7),
    .io_wreq_bits_data_1_entries_prefetch(l2_io_wreq_bits_data_1_entries_prefetch),
    .io_wreq_bits_data_1_ecc(l2_io_wreq_bits_data_1_ecc),
    .io_wreq_bits_data_2_entries_tag(l2_io_wreq_bits_data_2_entries_tag),
    .io_wreq_bits_data_2_entries_asid(l2_io_wreq_bits_data_2_entries_asid),
    .io_wreq_bits_data_2_entries_ppns_0(l2_io_wreq_bits_data_2_entries_ppns_0),
    .io_wreq_bits_data_2_entries_ppns_1(l2_io_wreq_bits_data_2_entries_ppns_1),
    .io_wreq_bits_data_2_entries_ppns_2(l2_io_wreq_bits_data_2_entries_ppns_2),
    .io_wreq_bits_data_2_entries_ppns_3(l2_io_wreq_bits_data_2_entries_ppns_3),
    .io_wreq_bits_data_2_entries_ppns_4(l2_io_wreq_bits_data_2_entries_ppns_4),
    .io_wreq_bits_data_2_entries_ppns_5(l2_io_wreq_bits_data_2_entries_ppns_5),
    .io_wreq_bits_data_2_entries_ppns_6(l2_io_wreq_bits_data_2_entries_ppns_6),
    .io_wreq_bits_data_2_entries_ppns_7(l2_io_wreq_bits_data_2_entries_ppns_7),
    .io_wreq_bits_data_2_entries_vs_0(l2_io_wreq_bits_data_2_entries_vs_0),
    .io_wreq_bits_data_2_entries_vs_1(l2_io_wreq_bits_data_2_entries_vs_1),
    .io_wreq_bits_data_2_entries_vs_2(l2_io_wreq_bits_data_2_entries_vs_2),
    .io_wreq_bits_data_2_entries_vs_3(l2_io_wreq_bits_data_2_entries_vs_3),
    .io_wreq_bits_data_2_entries_vs_4(l2_io_wreq_bits_data_2_entries_vs_4),
    .io_wreq_bits_data_2_entries_vs_5(l2_io_wreq_bits_data_2_entries_vs_5),
    .io_wreq_bits_data_2_entries_vs_6(l2_io_wreq_bits_data_2_entries_vs_6),
    .io_wreq_bits_data_2_entries_vs_7(l2_io_wreq_bits_data_2_entries_vs_7),
    .io_wreq_bits_data_2_entries_prefetch(l2_io_wreq_bits_data_2_entries_prefetch),
    .io_wreq_bits_data_2_ecc(l2_io_wreq_bits_data_2_ecc),
    .io_wreq_bits_data_3_entries_tag(l2_io_wreq_bits_data_3_entries_tag),
    .io_wreq_bits_data_3_entries_asid(l2_io_wreq_bits_data_3_entries_asid),
    .io_wreq_bits_data_3_entries_ppns_0(l2_io_wreq_bits_data_3_entries_ppns_0),
    .io_wreq_bits_data_3_entries_ppns_1(l2_io_wreq_bits_data_3_entries_ppns_1),
    .io_wreq_bits_data_3_entries_ppns_2(l2_io_wreq_bits_data_3_entries_ppns_2),
    .io_wreq_bits_data_3_entries_ppns_3(l2_io_wreq_bits_data_3_entries_ppns_3),
    .io_wreq_bits_data_3_entries_ppns_4(l2_io_wreq_bits_data_3_entries_ppns_4),
    .io_wreq_bits_data_3_entries_ppns_5(l2_io_wreq_bits_data_3_entries_ppns_5),
    .io_wreq_bits_data_3_entries_ppns_6(l2_io_wreq_bits_data_3_entries_ppns_6),
    .io_wreq_bits_data_3_entries_ppns_7(l2_io_wreq_bits_data_3_entries_ppns_7),
    .io_wreq_bits_data_3_entries_vs_0(l2_io_wreq_bits_data_3_entries_vs_0),
    .io_wreq_bits_data_3_entries_vs_1(l2_io_wreq_bits_data_3_entries_vs_1),
    .io_wreq_bits_data_3_entries_vs_2(l2_io_wreq_bits_data_3_entries_vs_2),
    .io_wreq_bits_data_3_entries_vs_3(l2_io_wreq_bits_data_3_entries_vs_3),
    .io_wreq_bits_data_3_entries_vs_4(l2_io_wreq_bits_data_3_entries_vs_4),
    .io_wreq_bits_data_3_entries_vs_5(l2_io_wreq_bits_data_3_entries_vs_5),
    .io_wreq_bits_data_3_entries_vs_6(l2_io_wreq_bits_data_3_entries_vs_6),
    .io_wreq_bits_data_3_entries_vs_7(l2_io_wreq_bits_data_3_entries_vs_7),
    .io_wreq_bits_data_3_entries_prefetch(l2_io_wreq_bits_data_3_entries_prefetch),
    .io_wreq_bits_data_3_ecc(l2_io_wreq_bits_data_3_ecc),
    .io_wreq_bits_waymask(l2_io_wreq_bits_waymask)
  );
  SRAMTemplate_69 l3 ( // @[PageTableCache.scala 179:18]
    .clock(l3_clock),
    .io_rreq_valid(l3_io_rreq_valid),
    .io_rreq_bits_setIdx(l3_io_rreq_bits_setIdx),
    .io_rresp_data_0_entries_tag(l3_io_rresp_data_0_entries_tag),
    .io_rresp_data_0_entries_asid(l3_io_rresp_data_0_entries_asid),
    .io_rresp_data_0_entries_ppns_0(l3_io_rresp_data_0_entries_ppns_0),
    .io_rresp_data_0_entries_ppns_1(l3_io_rresp_data_0_entries_ppns_1),
    .io_rresp_data_0_entries_ppns_2(l3_io_rresp_data_0_entries_ppns_2),
    .io_rresp_data_0_entries_ppns_3(l3_io_rresp_data_0_entries_ppns_3),
    .io_rresp_data_0_entries_ppns_4(l3_io_rresp_data_0_entries_ppns_4),
    .io_rresp_data_0_entries_ppns_5(l3_io_rresp_data_0_entries_ppns_5),
    .io_rresp_data_0_entries_ppns_6(l3_io_rresp_data_0_entries_ppns_6),
    .io_rresp_data_0_entries_ppns_7(l3_io_rresp_data_0_entries_ppns_7),
    .io_rresp_data_0_entries_vs_0(l3_io_rresp_data_0_entries_vs_0),
    .io_rresp_data_0_entries_vs_1(l3_io_rresp_data_0_entries_vs_1),
    .io_rresp_data_0_entries_vs_2(l3_io_rresp_data_0_entries_vs_2),
    .io_rresp_data_0_entries_vs_3(l3_io_rresp_data_0_entries_vs_3),
    .io_rresp_data_0_entries_vs_4(l3_io_rresp_data_0_entries_vs_4),
    .io_rresp_data_0_entries_vs_5(l3_io_rresp_data_0_entries_vs_5),
    .io_rresp_data_0_entries_vs_6(l3_io_rresp_data_0_entries_vs_6),
    .io_rresp_data_0_entries_vs_7(l3_io_rresp_data_0_entries_vs_7),
    .io_rresp_data_0_entries_perms_0_d(l3_io_rresp_data_0_entries_perms_0_d),
    .io_rresp_data_0_entries_perms_0_a(l3_io_rresp_data_0_entries_perms_0_a),
    .io_rresp_data_0_entries_perms_0_g(l3_io_rresp_data_0_entries_perms_0_g),
    .io_rresp_data_0_entries_perms_0_u(l3_io_rresp_data_0_entries_perms_0_u),
    .io_rresp_data_0_entries_perms_0_x(l3_io_rresp_data_0_entries_perms_0_x),
    .io_rresp_data_0_entries_perms_0_w(l3_io_rresp_data_0_entries_perms_0_w),
    .io_rresp_data_0_entries_perms_0_r(l3_io_rresp_data_0_entries_perms_0_r),
    .io_rresp_data_0_entries_perms_1_d(l3_io_rresp_data_0_entries_perms_1_d),
    .io_rresp_data_0_entries_perms_1_a(l3_io_rresp_data_0_entries_perms_1_a),
    .io_rresp_data_0_entries_perms_1_g(l3_io_rresp_data_0_entries_perms_1_g),
    .io_rresp_data_0_entries_perms_1_u(l3_io_rresp_data_0_entries_perms_1_u),
    .io_rresp_data_0_entries_perms_1_x(l3_io_rresp_data_0_entries_perms_1_x),
    .io_rresp_data_0_entries_perms_1_w(l3_io_rresp_data_0_entries_perms_1_w),
    .io_rresp_data_0_entries_perms_1_r(l3_io_rresp_data_0_entries_perms_1_r),
    .io_rresp_data_0_entries_perms_2_d(l3_io_rresp_data_0_entries_perms_2_d),
    .io_rresp_data_0_entries_perms_2_a(l3_io_rresp_data_0_entries_perms_2_a),
    .io_rresp_data_0_entries_perms_2_g(l3_io_rresp_data_0_entries_perms_2_g),
    .io_rresp_data_0_entries_perms_2_u(l3_io_rresp_data_0_entries_perms_2_u),
    .io_rresp_data_0_entries_perms_2_x(l3_io_rresp_data_0_entries_perms_2_x),
    .io_rresp_data_0_entries_perms_2_w(l3_io_rresp_data_0_entries_perms_2_w),
    .io_rresp_data_0_entries_perms_2_r(l3_io_rresp_data_0_entries_perms_2_r),
    .io_rresp_data_0_entries_perms_3_d(l3_io_rresp_data_0_entries_perms_3_d),
    .io_rresp_data_0_entries_perms_3_a(l3_io_rresp_data_0_entries_perms_3_a),
    .io_rresp_data_0_entries_perms_3_g(l3_io_rresp_data_0_entries_perms_3_g),
    .io_rresp_data_0_entries_perms_3_u(l3_io_rresp_data_0_entries_perms_3_u),
    .io_rresp_data_0_entries_perms_3_x(l3_io_rresp_data_0_entries_perms_3_x),
    .io_rresp_data_0_entries_perms_3_w(l3_io_rresp_data_0_entries_perms_3_w),
    .io_rresp_data_0_entries_perms_3_r(l3_io_rresp_data_0_entries_perms_3_r),
    .io_rresp_data_0_entries_perms_4_d(l3_io_rresp_data_0_entries_perms_4_d),
    .io_rresp_data_0_entries_perms_4_a(l3_io_rresp_data_0_entries_perms_4_a),
    .io_rresp_data_0_entries_perms_4_g(l3_io_rresp_data_0_entries_perms_4_g),
    .io_rresp_data_0_entries_perms_4_u(l3_io_rresp_data_0_entries_perms_4_u),
    .io_rresp_data_0_entries_perms_4_x(l3_io_rresp_data_0_entries_perms_4_x),
    .io_rresp_data_0_entries_perms_4_w(l3_io_rresp_data_0_entries_perms_4_w),
    .io_rresp_data_0_entries_perms_4_r(l3_io_rresp_data_0_entries_perms_4_r),
    .io_rresp_data_0_entries_perms_5_d(l3_io_rresp_data_0_entries_perms_5_d),
    .io_rresp_data_0_entries_perms_5_a(l3_io_rresp_data_0_entries_perms_5_a),
    .io_rresp_data_0_entries_perms_5_g(l3_io_rresp_data_0_entries_perms_5_g),
    .io_rresp_data_0_entries_perms_5_u(l3_io_rresp_data_0_entries_perms_5_u),
    .io_rresp_data_0_entries_perms_5_x(l3_io_rresp_data_0_entries_perms_5_x),
    .io_rresp_data_0_entries_perms_5_w(l3_io_rresp_data_0_entries_perms_5_w),
    .io_rresp_data_0_entries_perms_5_r(l3_io_rresp_data_0_entries_perms_5_r),
    .io_rresp_data_0_entries_perms_6_d(l3_io_rresp_data_0_entries_perms_6_d),
    .io_rresp_data_0_entries_perms_6_a(l3_io_rresp_data_0_entries_perms_6_a),
    .io_rresp_data_0_entries_perms_6_g(l3_io_rresp_data_0_entries_perms_6_g),
    .io_rresp_data_0_entries_perms_6_u(l3_io_rresp_data_0_entries_perms_6_u),
    .io_rresp_data_0_entries_perms_6_x(l3_io_rresp_data_0_entries_perms_6_x),
    .io_rresp_data_0_entries_perms_6_w(l3_io_rresp_data_0_entries_perms_6_w),
    .io_rresp_data_0_entries_perms_6_r(l3_io_rresp_data_0_entries_perms_6_r),
    .io_rresp_data_0_entries_perms_7_d(l3_io_rresp_data_0_entries_perms_7_d),
    .io_rresp_data_0_entries_perms_7_a(l3_io_rresp_data_0_entries_perms_7_a),
    .io_rresp_data_0_entries_perms_7_g(l3_io_rresp_data_0_entries_perms_7_g),
    .io_rresp_data_0_entries_perms_7_u(l3_io_rresp_data_0_entries_perms_7_u),
    .io_rresp_data_0_entries_perms_7_x(l3_io_rresp_data_0_entries_perms_7_x),
    .io_rresp_data_0_entries_perms_7_w(l3_io_rresp_data_0_entries_perms_7_w),
    .io_rresp_data_0_entries_perms_7_r(l3_io_rresp_data_0_entries_perms_7_r),
    .io_rresp_data_0_entries_prefetch(l3_io_rresp_data_0_entries_prefetch),
    .io_rresp_data_0_ecc(l3_io_rresp_data_0_ecc),
    .io_rresp_data_1_entries_tag(l3_io_rresp_data_1_entries_tag),
    .io_rresp_data_1_entries_asid(l3_io_rresp_data_1_entries_asid),
    .io_rresp_data_1_entries_ppns_0(l3_io_rresp_data_1_entries_ppns_0),
    .io_rresp_data_1_entries_ppns_1(l3_io_rresp_data_1_entries_ppns_1),
    .io_rresp_data_1_entries_ppns_2(l3_io_rresp_data_1_entries_ppns_2),
    .io_rresp_data_1_entries_ppns_3(l3_io_rresp_data_1_entries_ppns_3),
    .io_rresp_data_1_entries_ppns_4(l3_io_rresp_data_1_entries_ppns_4),
    .io_rresp_data_1_entries_ppns_5(l3_io_rresp_data_1_entries_ppns_5),
    .io_rresp_data_1_entries_ppns_6(l3_io_rresp_data_1_entries_ppns_6),
    .io_rresp_data_1_entries_ppns_7(l3_io_rresp_data_1_entries_ppns_7),
    .io_rresp_data_1_entries_vs_0(l3_io_rresp_data_1_entries_vs_0),
    .io_rresp_data_1_entries_vs_1(l3_io_rresp_data_1_entries_vs_1),
    .io_rresp_data_1_entries_vs_2(l3_io_rresp_data_1_entries_vs_2),
    .io_rresp_data_1_entries_vs_3(l3_io_rresp_data_1_entries_vs_3),
    .io_rresp_data_1_entries_vs_4(l3_io_rresp_data_1_entries_vs_4),
    .io_rresp_data_1_entries_vs_5(l3_io_rresp_data_1_entries_vs_5),
    .io_rresp_data_1_entries_vs_6(l3_io_rresp_data_1_entries_vs_6),
    .io_rresp_data_1_entries_vs_7(l3_io_rresp_data_1_entries_vs_7),
    .io_rresp_data_1_entries_perms_0_d(l3_io_rresp_data_1_entries_perms_0_d),
    .io_rresp_data_1_entries_perms_0_a(l3_io_rresp_data_1_entries_perms_0_a),
    .io_rresp_data_1_entries_perms_0_g(l3_io_rresp_data_1_entries_perms_0_g),
    .io_rresp_data_1_entries_perms_0_u(l3_io_rresp_data_1_entries_perms_0_u),
    .io_rresp_data_1_entries_perms_0_x(l3_io_rresp_data_1_entries_perms_0_x),
    .io_rresp_data_1_entries_perms_0_w(l3_io_rresp_data_1_entries_perms_0_w),
    .io_rresp_data_1_entries_perms_0_r(l3_io_rresp_data_1_entries_perms_0_r),
    .io_rresp_data_1_entries_perms_1_d(l3_io_rresp_data_1_entries_perms_1_d),
    .io_rresp_data_1_entries_perms_1_a(l3_io_rresp_data_1_entries_perms_1_a),
    .io_rresp_data_1_entries_perms_1_g(l3_io_rresp_data_1_entries_perms_1_g),
    .io_rresp_data_1_entries_perms_1_u(l3_io_rresp_data_1_entries_perms_1_u),
    .io_rresp_data_1_entries_perms_1_x(l3_io_rresp_data_1_entries_perms_1_x),
    .io_rresp_data_1_entries_perms_1_w(l3_io_rresp_data_1_entries_perms_1_w),
    .io_rresp_data_1_entries_perms_1_r(l3_io_rresp_data_1_entries_perms_1_r),
    .io_rresp_data_1_entries_perms_2_d(l3_io_rresp_data_1_entries_perms_2_d),
    .io_rresp_data_1_entries_perms_2_a(l3_io_rresp_data_1_entries_perms_2_a),
    .io_rresp_data_1_entries_perms_2_g(l3_io_rresp_data_1_entries_perms_2_g),
    .io_rresp_data_1_entries_perms_2_u(l3_io_rresp_data_1_entries_perms_2_u),
    .io_rresp_data_1_entries_perms_2_x(l3_io_rresp_data_1_entries_perms_2_x),
    .io_rresp_data_1_entries_perms_2_w(l3_io_rresp_data_1_entries_perms_2_w),
    .io_rresp_data_1_entries_perms_2_r(l3_io_rresp_data_1_entries_perms_2_r),
    .io_rresp_data_1_entries_perms_3_d(l3_io_rresp_data_1_entries_perms_3_d),
    .io_rresp_data_1_entries_perms_3_a(l3_io_rresp_data_1_entries_perms_3_a),
    .io_rresp_data_1_entries_perms_3_g(l3_io_rresp_data_1_entries_perms_3_g),
    .io_rresp_data_1_entries_perms_3_u(l3_io_rresp_data_1_entries_perms_3_u),
    .io_rresp_data_1_entries_perms_3_x(l3_io_rresp_data_1_entries_perms_3_x),
    .io_rresp_data_1_entries_perms_3_w(l3_io_rresp_data_1_entries_perms_3_w),
    .io_rresp_data_1_entries_perms_3_r(l3_io_rresp_data_1_entries_perms_3_r),
    .io_rresp_data_1_entries_perms_4_d(l3_io_rresp_data_1_entries_perms_4_d),
    .io_rresp_data_1_entries_perms_4_a(l3_io_rresp_data_1_entries_perms_4_a),
    .io_rresp_data_1_entries_perms_4_g(l3_io_rresp_data_1_entries_perms_4_g),
    .io_rresp_data_1_entries_perms_4_u(l3_io_rresp_data_1_entries_perms_4_u),
    .io_rresp_data_1_entries_perms_4_x(l3_io_rresp_data_1_entries_perms_4_x),
    .io_rresp_data_1_entries_perms_4_w(l3_io_rresp_data_1_entries_perms_4_w),
    .io_rresp_data_1_entries_perms_4_r(l3_io_rresp_data_1_entries_perms_4_r),
    .io_rresp_data_1_entries_perms_5_d(l3_io_rresp_data_1_entries_perms_5_d),
    .io_rresp_data_1_entries_perms_5_a(l3_io_rresp_data_1_entries_perms_5_a),
    .io_rresp_data_1_entries_perms_5_g(l3_io_rresp_data_1_entries_perms_5_g),
    .io_rresp_data_1_entries_perms_5_u(l3_io_rresp_data_1_entries_perms_5_u),
    .io_rresp_data_1_entries_perms_5_x(l3_io_rresp_data_1_entries_perms_5_x),
    .io_rresp_data_1_entries_perms_5_w(l3_io_rresp_data_1_entries_perms_5_w),
    .io_rresp_data_1_entries_perms_5_r(l3_io_rresp_data_1_entries_perms_5_r),
    .io_rresp_data_1_entries_perms_6_d(l3_io_rresp_data_1_entries_perms_6_d),
    .io_rresp_data_1_entries_perms_6_a(l3_io_rresp_data_1_entries_perms_6_a),
    .io_rresp_data_1_entries_perms_6_g(l3_io_rresp_data_1_entries_perms_6_g),
    .io_rresp_data_1_entries_perms_6_u(l3_io_rresp_data_1_entries_perms_6_u),
    .io_rresp_data_1_entries_perms_6_x(l3_io_rresp_data_1_entries_perms_6_x),
    .io_rresp_data_1_entries_perms_6_w(l3_io_rresp_data_1_entries_perms_6_w),
    .io_rresp_data_1_entries_perms_6_r(l3_io_rresp_data_1_entries_perms_6_r),
    .io_rresp_data_1_entries_perms_7_d(l3_io_rresp_data_1_entries_perms_7_d),
    .io_rresp_data_1_entries_perms_7_a(l3_io_rresp_data_1_entries_perms_7_a),
    .io_rresp_data_1_entries_perms_7_g(l3_io_rresp_data_1_entries_perms_7_g),
    .io_rresp_data_1_entries_perms_7_u(l3_io_rresp_data_1_entries_perms_7_u),
    .io_rresp_data_1_entries_perms_7_x(l3_io_rresp_data_1_entries_perms_7_x),
    .io_rresp_data_1_entries_perms_7_w(l3_io_rresp_data_1_entries_perms_7_w),
    .io_rresp_data_1_entries_perms_7_r(l3_io_rresp_data_1_entries_perms_7_r),
    .io_rresp_data_1_entries_prefetch(l3_io_rresp_data_1_entries_prefetch),
    .io_rresp_data_1_ecc(l3_io_rresp_data_1_ecc),
    .io_rresp_data_2_entries_tag(l3_io_rresp_data_2_entries_tag),
    .io_rresp_data_2_entries_asid(l3_io_rresp_data_2_entries_asid),
    .io_rresp_data_2_entries_ppns_0(l3_io_rresp_data_2_entries_ppns_0),
    .io_rresp_data_2_entries_ppns_1(l3_io_rresp_data_2_entries_ppns_1),
    .io_rresp_data_2_entries_ppns_2(l3_io_rresp_data_2_entries_ppns_2),
    .io_rresp_data_2_entries_ppns_3(l3_io_rresp_data_2_entries_ppns_3),
    .io_rresp_data_2_entries_ppns_4(l3_io_rresp_data_2_entries_ppns_4),
    .io_rresp_data_2_entries_ppns_5(l3_io_rresp_data_2_entries_ppns_5),
    .io_rresp_data_2_entries_ppns_6(l3_io_rresp_data_2_entries_ppns_6),
    .io_rresp_data_2_entries_ppns_7(l3_io_rresp_data_2_entries_ppns_7),
    .io_rresp_data_2_entries_vs_0(l3_io_rresp_data_2_entries_vs_0),
    .io_rresp_data_2_entries_vs_1(l3_io_rresp_data_2_entries_vs_1),
    .io_rresp_data_2_entries_vs_2(l3_io_rresp_data_2_entries_vs_2),
    .io_rresp_data_2_entries_vs_3(l3_io_rresp_data_2_entries_vs_3),
    .io_rresp_data_2_entries_vs_4(l3_io_rresp_data_2_entries_vs_4),
    .io_rresp_data_2_entries_vs_5(l3_io_rresp_data_2_entries_vs_5),
    .io_rresp_data_2_entries_vs_6(l3_io_rresp_data_2_entries_vs_6),
    .io_rresp_data_2_entries_vs_7(l3_io_rresp_data_2_entries_vs_7),
    .io_rresp_data_2_entries_perms_0_d(l3_io_rresp_data_2_entries_perms_0_d),
    .io_rresp_data_2_entries_perms_0_a(l3_io_rresp_data_2_entries_perms_0_a),
    .io_rresp_data_2_entries_perms_0_g(l3_io_rresp_data_2_entries_perms_0_g),
    .io_rresp_data_2_entries_perms_0_u(l3_io_rresp_data_2_entries_perms_0_u),
    .io_rresp_data_2_entries_perms_0_x(l3_io_rresp_data_2_entries_perms_0_x),
    .io_rresp_data_2_entries_perms_0_w(l3_io_rresp_data_2_entries_perms_0_w),
    .io_rresp_data_2_entries_perms_0_r(l3_io_rresp_data_2_entries_perms_0_r),
    .io_rresp_data_2_entries_perms_1_d(l3_io_rresp_data_2_entries_perms_1_d),
    .io_rresp_data_2_entries_perms_1_a(l3_io_rresp_data_2_entries_perms_1_a),
    .io_rresp_data_2_entries_perms_1_g(l3_io_rresp_data_2_entries_perms_1_g),
    .io_rresp_data_2_entries_perms_1_u(l3_io_rresp_data_2_entries_perms_1_u),
    .io_rresp_data_2_entries_perms_1_x(l3_io_rresp_data_2_entries_perms_1_x),
    .io_rresp_data_2_entries_perms_1_w(l3_io_rresp_data_2_entries_perms_1_w),
    .io_rresp_data_2_entries_perms_1_r(l3_io_rresp_data_2_entries_perms_1_r),
    .io_rresp_data_2_entries_perms_2_d(l3_io_rresp_data_2_entries_perms_2_d),
    .io_rresp_data_2_entries_perms_2_a(l3_io_rresp_data_2_entries_perms_2_a),
    .io_rresp_data_2_entries_perms_2_g(l3_io_rresp_data_2_entries_perms_2_g),
    .io_rresp_data_2_entries_perms_2_u(l3_io_rresp_data_2_entries_perms_2_u),
    .io_rresp_data_2_entries_perms_2_x(l3_io_rresp_data_2_entries_perms_2_x),
    .io_rresp_data_2_entries_perms_2_w(l3_io_rresp_data_2_entries_perms_2_w),
    .io_rresp_data_2_entries_perms_2_r(l3_io_rresp_data_2_entries_perms_2_r),
    .io_rresp_data_2_entries_perms_3_d(l3_io_rresp_data_2_entries_perms_3_d),
    .io_rresp_data_2_entries_perms_3_a(l3_io_rresp_data_2_entries_perms_3_a),
    .io_rresp_data_2_entries_perms_3_g(l3_io_rresp_data_2_entries_perms_3_g),
    .io_rresp_data_2_entries_perms_3_u(l3_io_rresp_data_2_entries_perms_3_u),
    .io_rresp_data_2_entries_perms_3_x(l3_io_rresp_data_2_entries_perms_3_x),
    .io_rresp_data_2_entries_perms_3_w(l3_io_rresp_data_2_entries_perms_3_w),
    .io_rresp_data_2_entries_perms_3_r(l3_io_rresp_data_2_entries_perms_3_r),
    .io_rresp_data_2_entries_perms_4_d(l3_io_rresp_data_2_entries_perms_4_d),
    .io_rresp_data_2_entries_perms_4_a(l3_io_rresp_data_2_entries_perms_4_a),
    .io_rresp_data_2_entries_perms_4_g(l3_io_rresp_data_2_entries_perms_4_g),
    .io_rresp_data_2_entries_perms_4_u(l3_io_rresp_data_2_entries_perms_4_u),
    .io_rresp_data_2_entries_perms_4_x(l3_io_rresp_data_2_entries_perms_4_x),
    .io_rresp_data_2_entries_perms_4_w(l3_io_rresp_data_2_entries_perms_4_w),
    .io_rresp_data_2_entries_perms_4_r(l3_io_rresp_data_2_entries_perms_4_r),
    .io_rresp_data_2_entries_perms_5_d(l3_io_rresp_data_2_entries_perms_5_d),
    .io_rresp_data_2_entries_perms_5_a(l3_io_rresp_data_2_entries_perms_5_a),
    .io_rresp_data_2_entries_perms_5_g(l3_io_rresp_data_2_entries_perms_5_g),
    .io_rresp_data_2_entries_perms_5_u(l3_io_rresp_data_2_entries_perms_5_u),
    .io_rresp_data_2_entries_perms_5_x(l3_io_rresp_data_2_entries_perms_5_x),
    .io_rresp_data_2_entries_perms_5_w(l3_io_rresp_data_2_entries_perms_5_w),
    .io_rresp_data_2_entries_perms_5_r(l3_io_rresp_data_2_entries_perms_5_r),
    .io_rresp_data_2_entries_perms_6_d(l3_io_rresp_data_2_entries_perms_6_d),
    .io_rresp_data_2_entries_perms_6_a(l3_io_rresp_data_2_entries_perms_6_a),
    .io_rresp_data_2_entries_perms_6_g(l3_io_rresp_data_2_entries_perms_6_g),
    .io_rresp_data_2_entries_perms_6_u(l3_io_rresp_data_2_entries_perms_6_u),
    .io_rresp_data_2_entries_perms_6_x(l3_io_rresp_data_2_entries_perms_6_x),
    .io_rresp_data_2_entries_perms_6_w(l3_io_rresp_data_2_entries_perms_6_w),
    .io_rresp_data_2_entries_perms_6_r(l3_io_rresp_data_2_entries_perms_6_r),
    .io_rresp_data_2_entries_perms_7_d(l3_io_rresp_data_2_entries_perms_7_d),
    .io_rresp_data_2_entries_perms_7_a(l3_io_rresp_data_2_entries_perms_7_a),
    .io_rresp_data_2_entries_perms_7_g(l3_io_rresp_data_2_entries_perms_7_g),
    .io_rresp_data_2_entries_perms_7_u(l3_io_rresp_data_2_entries_perms_7_u),
    .io_rresp_data_2_entries_perms_7_x(l3_io_rresp_data_2_entries_perms_7_x),
    .io_rresp_data_2_entries_perms_7_w(l3_io_rresp_data_2_entries_perms_7_w),
    .io_rresp_data_2_entries_perms_7_r(l3_io_rresp_data_2_entries_perms_7_r),
    .io_rresp_data_2_entries_prefetch(l3_io_rresp_data_2_entries_prefetch),
    .io_rresp_data_2_ecc(l3_io_rresp_data_2_ecc),
    .io_rresp_data_3_entries_tag(l3_io_rresp_data_3_entries_tag),
    .io_rresp_data_3_entries_asid(l3_io_rresp_data_3_entries_asid),
    .io_rresp_data_3_entries_ppns_0(l3_io_rresp_data_3_entries_ppns_0),
    .io_rresp_data_3_entries_ppns_1(l3_io_rresp_data_3_entries_ppns_1),
    .io_rresp_data_3_entries_ppns_2(l3_io_rresp_data_3_entries_ppns_2),
    .io_rresp_data_3_entries_ppns_3(l3_io_rresp_data_3_entries_ppns_3),
    .io_rresp_data_3_entries_ppns_4(l3_io_rresp_data_3_entries_ppns_4),
    .io_rresp_data_3_entries_ppns_5(l3_io_rresp_data_3_entries_ppns_5),
    .io_rresp_data_3_entries_ppns_6(l3_io_rresp_data_3_entries_ppns_6),
    .io_rresp_data_3_entries_ppns_7(l3_io_rresp_data_3_entries_ppns_7),
    .io_rresp_data_3_entries_vs_0(l3_io_rresp_data_3_entries_vs_0),
    .io_rresp_data_3_entries_vs_1(l3_io_rresp_data_3_entries_vs_1),
    .io_rresp_data_3_entries_vs_2(l3_io_rresp_data_3_entries_vs_2),
    .io_rresp_data_3_entries_vs_3(l3_io_rresp_data_3_entries_vs_3),
    .io_rresp_data_3_entries_vs_4(l3_io_rresp_data_3_entries_vs_4),
    .io_rresp_data_3_entries_vs_5(l3_io_rresp_data_3_entries_vs_5),
    .io_rresp_data_3_entries_vs_6(l3_io_rresp_data_3_entries_vs_6),
    .io_rresp_data_3_entries_vs_7(l3_io_rresp_data_3_entries_vs_7),
    .io_rresp_data_3_entries_perms_0_d(l3_io_rresp_data_3_entries_perms_0_d),
    .io_rresp_data_3_entries_perms_0_a(l3_io_rresp_data_3_entries_perms_0_a),
    .io_rresp_data_3_entries_perms_0_g(l3_io_rresp_data_3_entries_perms_0_g),
    .io_rresp_data_3_entries_perms_0_u(l3_io_rresp_data_3_entries_perms_0_u),
    .io_rresp_data_3_entries_perms_0_x(l3_io_rresp_data_3_entries_perms_0_x),
    .io_rresp_data_3_entries_perms_0_w(l3_io_rresp_data_3_entries_perms_0_w),
    .io_rresp_data_3_entries_perms_0_r(l3_io_rresp_data_3_entries_perms_0_r),
    .io_rresp_data_3_entries_perms_1_d(l3_io_rresp_data_3_entries_perms_1_d),
    .io_rresp_data_3_entries_perms_1_a(l3_io_rresp_data_3_entries_perms_1_a),
    .io_rresp_data_3_entries_perms_1_g(l3_io_rresp_data_3_entries_perms_1_g),
    .io_rresp_data_3_entries_perms_1_u(l3_io_rresp_data_3_entries_perms_1_u),
    .io_rresp_data_3_entries_perms_1_x(l3_io_rresp_data_3_entries_perms_1_x),
    .io_rresp_data_3_entries_perms_1_w(l3_io_rresp_data_3_entries_perms_1_w),
    .io_rresp_data_3_entries_perms_1_r(l3_io_rresp_data_3_entries_perms_1_r),
    .io_rresp_data_3_entries_perms_2_d(l3_io_rresp_data_3_entries_perms_2_d),
    .io_rresp_data_3_entries_perms_2_a(l3_io_rresp_data_3_entries_perms_2_a),
    .io_rresp_data_3_entries_perms_2_g(l3_io_rresp_data_3_entries_perms_2_g),
    .io_rresp_data_3_entries_perms_2_u(l3_io_rresp_data_3_entries_perms_2_u),
    .io_rresp_data_3_entries_perms_2_x(l3_io_rresp_data_3_entries_perms_2_x),
    .io_rresp_data_3_entries_perms_2_w(l3_io_rresp_data_3_entries_perms_2_w),
    .io_rresp_data_3_entries_perms_2_r(l3_io_rresp_data_3_entries_perms_2_r),
    .io_rresp_data_3_entries_perms_3_d(l3_io_rresp_data_3_entries_perms_3_d),
    .io_rresp_data_3_entries_perms_3_a(l3_io_rresp_data_3_entries_perms_3_a),
    .io_rresp_data_3_entries_perms_3_g(l3_io_rresp_data_3_entries_perms_3_g),
    .io_rresp_data_3_entries_perms_3_u(l3_io_rresp_data_3_entries_perms_3_u),
    .io_rresp_data_3_entries_perms_3_x(l3_io_rresp_data_3_entries_perms_3_x),
    .io_rresp_data_3_entries_perms_3_w(l3_io_rresp_data_3_entries_perms_3_w),
    .io_rresp_data_3_entries_perms_3_r(l3_io_rresp_data_3_entries_perms_3_r),
    .io_rresp_data_3_entries_perms_4_d(l3_io_rresp_data_3_entries_perms_4_d),
    .io_rresp_data_3_entries_perms_4_a(l3_io_rresp_data_3_entries_perms_4_a),
    .io_rresp_data_3_entries_perms_4_g(l3_io_rresp_data_3_entries_perms_4_g),
    .io_rresp_data_3_entries_perms_4_u(l3_io_rresp_data_3_entries_perms_4_u),
    .io_rresp_data_3_entries_perms_4_x(l3_io_rresp_data_3_entries_perms_4_x),
    .io_rresp_data_3_entries_perms_4_w(l3_io_rresp_data_3_entries_perms_4_w),
    .io_rresp_data_3_entries_perms_4_r(l3_io_rresp_data_3_entries_perms_4_r),
    .io_rresp_data_3_entries_perms_5_d(l3_io_rresp_data_3_entries_perms_5_d),
    .io_rresp_data_3_entries_perms_5_a(l3_io_rresp_data_3_entries_perms_5_a),
    .io_rresp_data_3_entries_perms_5_g(l3_io_rresp_data_3_entries_perms_5_g),
    .io_rresp_data_3_entries_perms_5_u(l3_io_rresp_data_3_entries_perms_5_u),
    .io_rresp_data_3_entries_perms_5_x(l3_io_rresp_data_3_entries_perms_5_x),
    .io_rresp_data_3_entries_perms_5_w(l3_io_rresp_data_3_entries_perms_5_w),
    .io_rresp_data_3_entries_perms_5_r(l3_io_rresp_data_3_entries_perms_5_r),
    .io_rresp_data_3_entries_perms_6_d(l3_io_rresp_data_3_entries_perms_6_d),
    .io_rresp_data_3_entries_perms_6_a(l3_io_rresp_data_3_entries_perms_6_a),
    .io_rresp_data_3_entries_perms_6_g(l3_io_rresp_data_3_entries_perms_6_g),
    .io_rresp_data_3_entries_perms_6_u(l3_io_rresp_data_3_entries_perms_6_u),
    .io_rresp_data_3_entries_perms_6_x(l3_io_rresp_data_3_entries_perms_6_x),
    .io_rresp_data_3_entries_perms_6_w(l3_io_rresp_data_3_entries_perms_6_w),
    .io_rresp_data_3_entries_perms_6_r(l3_io_rresp_data_3_entries_perms_6_r),
    .io_rresp_data_3_entries_perms_7_d(l3_io_rresp_data_3_entries_perms_7_d),
    .io_rresp_data_3_entries_perms_7_a(l3_io_rresp_data_3_entries_perms_7_a),
    .io_rresp_data_3_entries_perms_7_g(l3_io_rresp_data_3_entries_perms_7_g),
    .io_rresp_data_3_entries_perms_7_u(l3_io_rresp_data_3_entries_perms_7_u),
    .io_rresp_data_3_entries_perms_7_x(l3_io_rresp_data_3_entries_perms_7_x),
    .io_rresp_data_3_entries_perms_7_w(l3_io_rresp_data_3_entries_perms_7_w),
    .io_rresp_data_3_entries_perms_7_r(l3_io_rresp_data_3_entries_perms_7_r),
    .io_rresp_data_3_entries_prefetch(l3_io_rresp_data_3_entries_prefetch),
    .io_rresp_data_3_ecc(l3_io_rresp_data_3_ecc),
    .io_rresp_data_4_entries_tag(l3_io_rresp_data_4_entries_tag),
    .io_rresp_data_4_entries_asid(l3_io_rresp_data_4_entries_asid),
    .io_rresp_data_4_entries_ppns_0(l3_io_rresp_data_4_entries_ppns_0),
    .io_rresp_data_4_entries_ppns_1(l3_io_rresp_data_4_entries_ppns_1),
    .io_rresp_data_4_entries_ppns_2(l3_io_rresp_data_4_entries_ppns_2),
    .io_rresp_data_4_entries_ppns_3(l3_io_rresp_data_4_entries_ppns_3),
    .io_rresp_data_4_entries_ppns_4(l3_io_rresp_data_4_entries_ppns_4),
    .io_rresp_data_4_entries_ppns_5(l3_io_rresp_data_4_entries_ppns_5),
    .io_rresp_data_4_entries_ppns_6(l3_io_rresp_data_4_entries_ppns_6),
    .io_rresp_data_4_entries_ppns_7(l3_io_rresp_data_4_entries_ppns_7),
    .io_rresp_data_4_entries_vs_0(l3_io_rresp_data_4_entries_vs_0),
    .io_rresp_data_4_entries_vs_1(l3_io_rresp_data_4_entries_vs_1),
    .io_rresp_data_4_entries_vs_2(l3_io_rresp_data_4_entries_vs_2),
    .io_rresp_data_4_entries_vs_3(l3_io_rresp_data_4_entries_vs_3),
    .io_rresp_data_4_entries_vs_4(l3_io_rresp_data_4_entries_vs_4),
    .io_rresp_data_4_entries_vs_5(l3_io_rresp_data_4_entries_vs_5),
    .io_rresp_data_4_entries_vs_6(l3_io_rresp_data_4_entries_vs_6),
    .io_rresp_data_4_entries_vs_7(l3_io_rresp_data_4_entries_vs_7),
    .io_rresp_data_4_entries_perms_0_d(l3_io_rresp_data_4_entries_perms_0_d),
    .io_rresp_data_4_entries_perms_0_a(l3_io_rresp_data_4_entries_perms_0_a),
    .io_rresp_data_4_entries_perms_0_g(l3_io_rresp_data_4_entries_perms_0_g),
    .io_rresp_data_4_entries_perms_0_u(l3_io_rresp_data_4_entries_perms_0_u),
    .io_rresp_data_4_entries_perms_0_x(l3_io_rresp_data_4_entries_perms_0_x),
    .io_rresp_data_4_entries_perms_0_w(l3_io_rresp_data_4_entries_perms_0_w),
    .io_rresp_data_4_entries_perms_0_r(l3_io_rresp_data_4_entries_perms_0_r),
    .io_rresp_data_4_entries_perms_1_d(l3_io_rresp_data_4_entries_perms_1_d),
    .io_rresp_data_4_entries_perms_1_a(l3_io_rresp_data_4_entries_perms_1_a),
    .io_rresp_data_4_entries_perms_1_g(l3_io_rresp_data_4_entries_perms_1_g),
    .io_rresp_data_4_entries_perms_1_u(l3_io_rresp_data_4_entries_perms_1_u),
    .io_rresp_data_4_entries_perms_1_x(l3_io_rresp_data_4_entries_perms_1_x),
    .io_rresp_data_4_entries_perms_1_w(l3_io_rresp_data_4_entries_perms_1_w),
    .io_rresp_data_4_entries_perms_1_r(l3_io_rresp_data_4_entries_perms_1_r),
    .io_rresp_data_4_entries_perms_2_d(l3_io_rresp_data_4_entries_perms_2_d),
    .io_rresp_data_4_entries_perms_2_a(l3_io_rresp_data_4_entries_perms_2_a),
    .io_rresp_data_4_entries_perms_2_g(l3_io_rresp_data_4_entries_perms_2_g),
    .io_rresp_data_4_entries_perms_2_u(l3_io_rresp_data_4_entries_perms_2_u),
    .io_rresp_data_4_entries_perms_2_x(l3_io_rresp_data_4_entries_perms_2_x),
    .io_rresp_data_4_entries_perms_2_w(l3_io_rresp_data_4_entries_perms_2_w),
    .io_rresp_data_4_entries_perms_2_r(l3_io_rresp_data_4_entries_perms_2_r),
    .io_rresp_data_4_entries_perms_3_d(l3_io_rresp_data_4_entries_perms_3_d),
    .io_rresp_data_4_entries_perms_3_a(l3_io_rresp_data_4_entries_perms_3_a),
    .io_rresp_data_4_entries_perms_3_g(l3_io_rresp_data_4_entries_perms_3_g),
    .io_rresp_data_4_entries_perms_3_u(l3_io_rresp_data_4_entries_perms_3_u),
    .io_rresp_data_4_entries_perms_3_x(l3_io_rresp_data_4_entries_perms_3_x),
    .io_rresp_data_4_entries_perms_3_w(l3_io_rresp_data_4_entries_perms_3_w),
    .io_rresp_data_4_entries_perms_3_r(l3_io_rresp_data_4_entries_perms_3_r),
    .io_rresp_data_4_entries_perms_4_d(l3_io_rresp_data_4_entries_perms_4_d),
    .io_rresp_data_4_entries_perms_4_a(l3_io_rresp_data_4_entries_perms_4_a),
    .io_rresp_data_4_entries_perms_4_g(l3_io_rresp_data_4_entries_perms_4_g),
    .io_rresp_data_4_entries_perms_4_u(l3_io_rresp_data_4_entries_perms_4_u),
    .io_rresp_data_4_entries_perms_4_x(l3_io_rresp_data_4_entries_perms_4_x),
    .io_rresp_data_4_entries_perms_4_w(l3_io_rresp_data_4_entries_perms_4_w),
    .io_rresp_data_4_entries_perms_4_r(l3_io_rresp_data_4_entries_perms_4_r),
    .io_rresp_data_4_entries_perms_5_d(l3_io_rresp_data_4_entries_perms_5_d),
    .io_rresp_data_4_entries_perms_5_a(l3_io_rresp_data_4_entries_perms_5_a),
    .io_rresp_data_4_entries_perms_5_g(l3_io_rresp_data_4_entries_perms_5_g),
    .io_rresp_data_4_entries_perms_5_u(l3_io_rresp_data_4_entries_perms_5_u),
    .io_rresp_data_4_entries_perms_5_x(l3_io_rresp_data_4_entries_perms_5_x),
    .io_rresp_data_4_entries_perms_5_w(l3_io_rresp_data_4_entries_perms_5_w),
    .io_rresp_data_4_entries_perms_5_r(l3_io_rresp_data_4_entries_perms_5_r),
    .io_rresp_data_4_entries_perms_6_d(l3_io_rresp_data_4_entries_perms_6_d),
    .io_rresp_data_4_entries_perms_6_a(l3_io_rresp_data_4_entries_perms_6_a),
    .io_rresp_data_4_entries_perms_6_g(l3_io_rresp_data_4_entries_perms_6_g),
    .io_rresp_data_4_entries_perms_6_u(l3_io_rresp_data_4_entries_perms_6_u),
    .io_rresp_data_4_entries_perms_6_x(l3_io_rresp_data_4_entries_perms_6_x),
    .io_rresp_data_4_entries_perms_6_w(l3_io_rresp_data_4_entries_perms_6_w),
    .io_rresp_data_4_entries_perms_6_r(l3_io_rresp_data_4_entries_perms_6_r),
    .io_rresp_data_4_entries_perms_7_d(l3_io_rresp_data_4_entries_perms_7_d),
    .io_rresp_data_4_entries_perms_7_a(l3_io_rresp_data_4_entries_perms_7_a),
    .io_rresp_data_4_entries_perms_7_g(l3_io_rresp_data_4_entries_perms_7_g),
    .io_rresp_data_4_entries_perms_7_u(l3_io_rresp_data_4_entries_perms_7_u),
    .io_rresp_data_4_entries_perms_7_x(l3_io_rresp_data_4_entries_perms_7_x),
    .io_rresp_data_4_entries_perms_7_w(l3_io_rresp_data_4_entries_perms_7_w),
    .io_rresp_data_4_entries_perms_7_r(l3_io_rresp_data_4_entries_perms_7_r),
    .io_rresp_data_4_entries_prefetch(l3_io_rresp_data_4_entries_prefetch),
    .io_rresp_data_4_ecc(l3_io_rresp_data_4_ecc),
    .io_rresp_data_5_entries_tag(l3_io_rresp_data_5_entries_tag),
    .io_rresp_data_5_entries_asid(l3_io_rresp_data_5_entries_asid),
    .io_rresp_data_5_entries_ppns_0(l3_io_rresp_data_5_entries_ppns_0),
    .io_rresp_data_5_entries_ppns_1(l3_io_rresp_data_5_entries_ppns_1),
    .io_rresp_data_5_entries_ppns_2(l3_io_rresp_data_5_entries_ppns_2),
    .io_rresp_data_5_entries_ppns_3(l3_io_rresp_data_5_entries_ppns_3),
    .io_rresp_data_5_entries_ppns_4(l3_io_rresp_data_5_entries_ppns_4),
    .io_rresp_data_5_entries_ppns_5(l3_io_rresp_data_5_entries_ppns_5),
    .io_rresp_data_5_entries_ppns_6(l3_io_rresp_data_5_entries_ppns_6),
    .io_rresp_data_5_entries_ppns_7(l3_io_rresp_data_5_entries_ppns_7),
    .io_rresp_data_5_entries_vs_0(l3_io_rresp_data_5_entries_vs_0),
    .io_rresp_data_5_entries_vs_1(l3_io_rresp_data_5_entries_vs_1),
    .io_rresp_data_5_entries_vs_2(l3_io_rresp_data_5_entries_vs_2),
    .io_rresp_data_5_entries_vs_3(l3_io_rresp_data_5_entries_vs_3),
    .io_rresp_data_5_entries_vs_4(l3_io_rresp_data_5_entries_vs_4),
    .io_rresp_data_5_entries_vs_5(l3_io_rresp_data_5_entries_vs_5),
    .io_rresp_data_5_entries_vs_6(l3_io_rresp_data_5_entries_vs_6),
    .io_rresp_data_5_entries_vs_7(l3_io_rresp_data_5_entries_vs_7),
    .io_rresp_data_5_entries_perms_0_d(l3_io_rresp_data_5_entries_perms_0_d),
    .io_rresp_data_5_entries_perms_0_a(l3_io_rresp_data_5_entries_perms_0_a),
    .io_rresp_data_5_entries_perms_0_g(l3_io_rresp_data_5_entries_perms_0_g),
    .io_rresp_data_5_entries_perms_0_u(l3_io_rresp_data_5_entries_perms_0_u),
    .io_rresp_data_5_entries_perms_0_x(l3_io_rresp_data_5_entries_perms_0_x),
    .io_rresp_data_5_entries_perms_0_w(l3_io_rresp_data_5_entries_perms_0_w),
    .io_rresp_data_5_entries_perms_0_r(l3_io_rresp_data_5_entries_perms_0_r),
    .io_rresp_data_5_entries_perms_1_d(l3_io_rresp_data_5_entries_perms_1_d),
    .io_rresp_data_5_entries_perms_1_a(l3_io_rresp_data_5_entries_perms_1_a),
    .io_rresp_data_5_entries_perms_1_g(l3_io_rresp_data_5_entries_perms_1_g),
    .io_rresp_data_5_entries_perms_1_u(l3_io_rresp_data_5_entries_perms_1_u),
    .io_rresp_data_5_entries_perms_1_x(l3_io_rresp_data_5_entries_perms_1_x),
    .io_rresp_data_5_entries_perms_1_w(l3_io_rresp_data_5_entries_perms_1_w),
    .io_rresp_data_5_entries_perms_1_r(l3_io_rresp_data_5_entries_perms_1_r),
    .io_rresp_data_5_entries_perms_2_d(l3_io_rresp_data_5_entries_perms_2_d),
    .io_rresp_data_5_entries_perms_2_a(l3_io_rresp_data_5_entries_perms_2_a),
    .io_rresp_data_5_entries_perms_2_g(l3_io_rresp_data_5_entries_perms_2_g),
    .io_rresp_data_5_entries_perms_2_u(l3_io_rresp_data_5_entries_perms_2_u),
    .io_rresp_data_5_entries_perms_2_x(l3_io_rresp_data_5_entries_perms_2_x),
    .io_rresp_data_5_entries_perms_2_w(l3_io_rresp_data_5_entries_perms_2_w),
    .io_rresp_data_5_entries_perms_2_r(l3_io_rresp_data_5_entries_perms_2_r),
    .io_rresp_data_5_entries_perms_3_d(l3_io_rresp_data_5_entries_perms_3_d),
    .io_rresp_data_5_entries_perms_3_a(l3_io_rresp_data_5_entries_perms_3_a),
    .io_rresp_data_5_entries_perms_3_g(l3_io_rresp_data_5_entries_perms_3_g),
    .io_rresp_data_5_entries_perms_3_u(l3_io_rresp_data_5_entries_perms_3_u),
    .io_rresp_data_5_entries_perms_3_x(l3_io_rresp_data_5_entries_perms_3_x),
    .io_rresp_data_5_entries_perms_3_w(l3_io_rresp_data_5_entries_perms_3_w),
    .io_rresp_data_5_entries_perms_3_r(l3_io_rresp_data_5_entries_perms_3_r),
    .io_rresp_data_5_entries_perms_4_d(l3_io_rresp_data_5_entries_perms_4_d),
    .io_rresp_data_5_entries_perms_4_a(l3_io_rresp_data_5_entries_perms_4_a),
    .io_rresp_data_5_entries_perms_4_g(l3_io_rresp_data_5_entries_perms_4_g),
    .io_rresp_data_5_entries_perms_4_u(l3_io_rresp_data_5_entries_perms_4_u),
    .io_rresp_data_5_entries_perms_4_x(l3_io_rresp_data_5_entries_perms_4_x),
    .io_rresp_data_5_entries_perms_4_w(l3_io_rresp_data_5_entries_perms_4_w),
    .io_rresp_data_5_entries_perms_4_r(l3_io_rresp_data_5_entries_perms_4_r),
    .io_rresp_data_5_entries_perms_5_d(l3_io_rresp_data_5_entries_perms_5_d),
    .io_rresp_data_5_entries_perms_5_a(l3_io_rresp_data_5_entries_perms_5_a),
    .io_rresp_data_5_entries_perms_5_g(l3_io_rresp_data_5_entries_perms_5_g),
    .io_rresp_data_5_entries_perms_5_u(l3_io_rresp_data_5_entries_perms_5_u),
    .io_rresp_data_5_entries_perms_5_x(l3_io_rresp_data_5_entries_perms_5_x),
    .io_rresp_data_5_entries_perms_5_w(l3_io_rresp_data_5_entries_perms_5_w),
    .io_rresp_data_5_entries_perms_5_r(l3_io_rresp_data_5_entries_perms_5_r),
    .io_rresp_data_5_entries_perms_6_d(l3_io_rresp_data_5_entries_perms_6_d),
    .io_rresp_data_5_entries_perms_6_a(l3_io_rresp_data_5_entries_perms_6_a),
    .io_rresp_data_5_entries_perms_6_g(l3_io_rresp_data_5_entries_perms_6_g),
    .io_rresp_data_5_entries_perms_6_u(l3_io_rresp_data_5_entries_perms_6_u),
    .io_rresp_data_5_entries_perms_6_x(l3_io_rresp_data_5_entries_perms_6_x),
    .io_rresp_data_5_entries_perms_6_w(l3_io_rresp_data_5_entries_perms_6_w),
    .io_rresp_data_5_entries_perms_6_r(l3_io_rresp_data_5_entries_perms_6_r),
    .io_rresp_data_5_entries_perms_7_d(l3_io_rresp_data_5_entries_perms_7_d),
    .io_rresp_data_5_entries_perms_7_a(l3_io_rresp_data_5_entries_perms_7_a),
    .io_rresp_data_5_entries_perms_7_g(l3_io_rresp_data_5_entries_perms_7_g),
    .io_rresp_data_5_entries_perms_7_u(l3_io_rresp_data_5_entries_perms_7_u),
    .io_rresp_data_5_entries_perms_7_x(l3_io_rresp_data_5_entries_perms_7_x),
    .io_rresp_data_5_entries_perms_7_w(l3_io_rresp_data_5_entries_perms_7_w),
    .io_rresp_data_5_entries_perms_7_r(l3_io_rresp_data_5_entries_perms_7_r),
    .io_rresp_data_5_entries_prefetch(l3_io_rresp_data_5_entries_prefetch),
    .io_rresp_data_5_ecc(l3_io_rresp_data_5_ecc),
    .io_rresp_data_6_entries_tag(l3_io_rresp_data_6_entries_tag),
    .io_rresp_data_6_entries_asid(l3_io_rresp_data_6_entries_asid),
    .io_rresp_data_6_entries_ppns_0(l3_io_rresp_data_6_entries_ppns_0),
    .io_rresp_data_6_entries_ppns_1(l3_io_rresp_data_6_entries_ppns_1),
    .io_rresp_data_6_entries_ppns_2(l3_io_rresp_data_6_entries_ppns_2),
    .io_rresp_data_6_entries_ppns_3(l3_io_rresp_data_6_entries_ppns_3),
    .io_rresp_data_6_entries_ppns_4(l3_io_rresp_data_6_entries_ppns_4),
    .io_rresp_data_6_entries_ppns_5(l3_io_rresp_data_6_entries_ppns_5),
    .io_rresp_data_6_entries_ppns_6(l3_io_rresp_data_6_entries_ppns_6),
    .io_rresp_data_6_entries_ppns_7(l3_io_rresp_data_6_entries_ppns_7),
    .io_rresp_data_6_entries_vs_0(l3_io_rresp_data_6_entries_vs_0),
    .io_rresp_data_6_entries_vs_1(l3_io_rresp_data_6_entries_vs_1),
    .io_rresp_data_6_entries_vs_2(l3_io_rresp_data_6_entries_vs_2),
    .io_rresp_data_6_entries_vs_3(l3_io_rresp_data_6_entries_vs_3),
    .io_rresp_data_6_entries_vs_4(l3_io_rresp_data_6_entries_vs_4),
    .io_rresp_data_6_entries_vs_5(l3_io_rresp_data_6_entries_vs_5),
    .io_rresp_data_6_entries_vs_6(l3_io_rresp_data_6_entries_vs_6),
    .io_rresp_data_6_entries_vs_7(l3_io_rresp_data_6_entries_vs_7),
    .io_rresp_data_6_entries_perms_0_d(l3_io_rresp_data_6_entries_perms_0_d),
    .io_rresp_data_6_entries_perms_0_a(l3_io_rresp_data_6_entries_perms_0_a),
    .io_rresp_data_6_entries_perms_0_g(l3_io_rresp_data_6_entries_perms_0_g),
    .io_rresp_data_6_entries_perms_0_u(l3_io_rresp_data_6_entries_perms_0_u),
    .io_rresp_data_6_entries_perms_0_x(l3_io_rresp_data_6_entries_perms_0_x),
    .io_rresp_data_6_entries_perms_0_w(l3_io_rresp_data_6_entries_perms_0_w),
    .io_rresp_data_6_entries_perms_0_r(l3_io_rresp_data_6_entries_perms_0_r),
    .io_rresp_data_6_entries_perms_1_d(l3_io_rresp_data_6_entries_perms_1_d),
    .io_rresp_data_6_entries_perms_1_a(l3_io_rresp_data_6_entries_perms_1_a),
    .io_rresp_data_6_entries_perms_1_g(l3_io_rresp_data_6_entries_perms_1_g),
    .io_rresp_data_6_entries_perms_1_u(l3_io_rresp_data_6_entries_perms_1_u),
    .io_rresp_data_6_entries_perms_1_x(l3_io_rresp_data_6_entries_perms_1_x),
    .io_rresp_data_6_entries_perms_1_w(l3_io_rresp_data_6_entries_perms_1_w),
    .io_rresp_data_6_entries_perms_1_r(l3_io_rresp_data_6_entries_perms_1_r),
    .io_rresp_data_6_entries_perms_2_d(l3_io_rresp_data_6_entries_perms_2_d),
    .io_rresp_data_6_entries_perms_2_a(l3_io_rresp_data_6_entries_perms_2_a),
    .io_rresp_data_6_entries_perms_2_g(l3_io_rresp_data_6_entries_perms_2_g),
    .io_rresp_data_6_entries_perms_2_u(l3_io_rresp_data_6_entries_perms_2_u),
    .io_rresp_data_6_entries_perms_2_x(l3_io_rresp_data_6_entries_perms_2_x),
    .io_rresp_data_6_entries_perms_2_w(l3_io_rresp_data_6_entries_perms_2_w),
    .io_rresp_data_6_entries_perms_2_r(l3_io_rresp_data_6_entries_perms_2_r),
    .io_rresp_data_6_entries_perms_3_d(l3_io_rresp_data_6_entries_perms_3_d),
    .io_rresp_data_6_entries_perms_3_a(l3_io_rresp_data_6_entries_perms_3_a),
    .io_rresp_data_6_entries_perms_3_g(l3_io_rresp_data_6_entries_perms_3_g),
    .io_rresp_data_6_entries_perms_3_u(l3_io_rresp_data_6_entries_perms_3_u),
    .io_rresp_data_6_entries_perms_3_x(l3_io_rresp_data_6_entries_perms_3_x),
    .io_rresp_data_6_entries_perms_3_w(l3_io_rresp_data_6_entries_perms_3_w),
    .io_rresp_data_6_entries_perms_3_r(l3_io_rresp_data_6_entries_perms_3_r),
    .io_rresp_data_6_entries_perms_4_d(l3_io_rresp_data_6_entries_perms_4_d),
    .io_rresp_data_6_entries_perms_4_a(l3_io_rresp_data_6_entries_perms_4_a),
    .io_rresp_data_6_entries_perms_4_g(l3_io_rresp_data_6_entries_perms_4_g),
    .io_rresp_data_6_entries_perms_4_u(l3_io_rresp_data_6_entries_perms_4_u),
    .io_rresp_data_6_entries_perms_4_x(l3_io_rresp_data_6_entries_perms_4_x),
    .io_rresp_data_6_entries_perms_4_w(l3_io_rresp_data_6_entries_perms_4_w),
    .io_rresp_data_6_entries_perms_4_r(l3_io_rresp_data_6_entries_perms_4_r),
    .io_rresp_data_6_entries_perms_5_d(l3_io_rresp_data_6_entries_perms_5_d),
    .io_rresp_data_6_entries_perms_5_a(l3_io_rresp_data_6_entries_perms_5_a),
    .io_rresp_data_6_entries_perms_5_g(l3_io_rresp_data_6_entries_perms_5_g),
    .io_rresp_data_6_entries_perms_5_u(l3_io_rresp_data_6_entries_perms_5_u),
    .io_rresp_data_6_entries_perms_5_x(l3_io_rresp_data_6_entries_perms_5_x),
    .io_rresp_data_6_entries_perms_5_w(l3_io_rresp_data_6_entries_perms_5_w),
    .io_rresp_data_6_entries_perms_5_r(l3_io_rresp_data_6_entries_perms_5_r),
    .io_rresp_data_6_entries_perms_6_d(l3_io_rresp_data_6_entries_perms_6_d),
    .io_rresp_data_6_entries_perms_6_a(l3_io_rresp_data_6_entries_perms_6_a),
    .io_rresp_data_6_entries_perms_6_g(l3_io_rresp_data_6_entries_perms_6_g),
    .io_rresp_data_6_entries_perms_6_u(l3_io_rresp_data_6_entries_perms_6_u),
    .io_rresp_data_6_entries_perms_6_x(l3_io_rresp_data_6_entries_perms_6_x),
    .io_rresp_data_6_entries_perms_6_w(l3_io_rresp_data_6_entries_perms_6_w),
    .io_rresp_data_6_entries_perms_6_r(l3_io_rresp_data_6_entries_perms_6_r),
    .io_rresp_data_6_entries_perms_7_d(l3_io_rresp_data_6_entries_perms_7_d),
    .io_rresp_data_6_entries_perms_7_a(l3_io_rresp_data_6_entries_perms_7_a),
    .io_rresp_data_6_entries_perms_7_g(l3_io_rresp_data_6_entries_perms_7_g),
    .io_rresp_data_6_entries_perms_7_u(l3_io_rresp_data_6_entries_perms_7_u),
    .io_rresp_data_6_entries_perms_7_x(l3_io_rresp_data_6_entries_perms_7_x),
    .io_rresp_data_6_entries_perms_7_w(l3_io_rresp_data_6_entries_perms_7_w),
    .io_rresp_data_6_entries_perms_7_r(l3_io_rresp_data_6_entries_perms_7_r),
    .io_rresp_data_6_entries_prefetch(l3_io_rresp_data_6_entries_prefetch),
    .io_rresp_data_6_ecc(l3_io_rresp_data_6_ecc),
    .io_rresp_data_7_entries_tag(l3_io_rresp_data_7_entries_tag),
    .io_rresp_data_7_entries_asid(l3_io_rresp_data_7_entries_asid),
    .io_rresp_data_7_entries_ppns_0(l3_io_rresp_data_7_entries_ppns_0),
    .io_rresp_data_7_entries_ppns_1(l3_io_rresp_data_7_entries_ppns_1),
    .io_rresp_data_7_entries_ppns_2(l3_io_rresp_data_7_entries_ppns_2),
    .io_rresp_data_7_entries_ppns_3(l3_io_rresp_data_7_entries_ppns_3),
    .io_rresp_data_7_entries_ppns_4(l3_io_rresp_data_7_entries_ppns_4),
    .io_rresp_data_7_entries_ppns_5(l3_io_rresp_data_7_entries_ppns_5),
    .io_rresp_data_7_entries_ppns_6(l3_io_rresp_data_7_entries_ppns_6),
    .io_rresp_data_7_entries_ppns_7(l3_io_rresp_data_7_entries_ppns_7),
    .io_rresp_data_7_entries_vs_0(l3_io_rresp_data_7_entries_vs_0),
    .io_rresp_data_7_entries_vs_1(l3_io_rresp_data_7_entries_vs_1),
    .io_rresp_data_7_entries_vs_2(l3_io_rresp_data_7_entries_vs_2),
    .io_rresp_data_7_entries_vs_3(l3_io_rresp_data_7_entries_vs_3),
    .io_rresp_data_7_entries_vs_4(l3_io_rresp_data_7_entries_vs_4),
    .io_rresp_data_7_entries_vs_5(l3_io_rresp_data_7_entries_vs_5),
    .io_rresp_data_7_entries_vs_6(l3_io_rresp_data_7_entries_vs_6),
    .io_rresp_data_7_entries_vs_7(l3_io_rresp_data_7_entries_vs_7),
    .io_rresp_data_7_entries_perms_0_d(l3_io_rresp_data_7_entries_perms_0_d),
    .io_rresp_data_7_entries_perms_0_a(l3_io_rresp_data_7_entries_perms_0_a),
    .io_rresp_data_7_entries_perms_0_g(l3_io_rresp_data_7_entries_perms_0_g),
    .io_rresp_data_7_entries_perms_0_u(l3_io_rresp_data_7_entries_perms_0_u),
    .io_rresp_data_7_entries_perms_0_x(l3_io_rresp_data_7_entries_perms_0_x),
    .io_rresp_data_7_entries_perms_0_w(l3_io_rresp_data_7_entries_perms_0_w),
    .io_rresp_data_7_entries_perms_0_r(l3_io_rresp_data_7_entries_perms_0_r),
    .io_rresp_data_7_entries_perms_1_d(l3_io_rresp_data_7_entries_perms_1_d),
    .io_rresp_data_7_entries_perms_1_a(l3_io_rresp_data_7_entries_perms_1_a),
    .io_rresp_data_7_entries_perms_1_g(l3_io_rresp_data_7_entries_perms_1_g),
    .io_rresp_data_7_entries_perms_1_u(l3_io_rresp_data_7_entries_perms_1_u),
    .io_rresp_data_7_entries_perms_1_x(l3_io_rresp_data_7_entries_perms_1_x),
    .io_rresp_data_7_entries_perms_1_w(l3_io_rresp_data_7_entries_perms_1_w),
    .io_rresp_data_7_entries_perms_1_r(l3_io_rresp_data_7_entries_perms_1_r),
    .io_rresp_data_7_entries_perms_2_d(l3_io_rresp_data_7_entries_perms_2_d),
    .io_rresp_data_7_entries_perms_2_a(l3_io_rresp_data_7_entries_perms_2_a),
    .io_rresp_data_7_entries_perms_2_g(l3_io_rresp_data_7_entries_perms_2_g),
    .io_rresp_data_7_entries_perms_2_u(l3_io_rresp_data_7_entries_perms_2_u),
    .io_rresp_data_7_entries_perms_2_x(l3_io_rresp_data_7_entries_perms_2_x),
    .io_rresp_data_7_entries_perms_2_w(l3_io_rresp_data_7_entries_perms_2_w),
    .io_rresp_data_7_entries_perms_2_r(l3_io_rresp_data_7_entries_perms_2_r),
    .io_rresp_data_7_entries_perms_3_d(l3_io_rresp_data_7_entries_perms_3_d),
    .io_rresp_data_7_entries_perms_3_a(l3_io_rresp_data_7_entries_perms_3_a),
    .io_rresp_data_7_entries_perms_3_g(l3_io_rresp_data_7_entries_perms_3_g),
    .io_rresp_data_7_entries_perms_3_u(l3_io_rresp_data_7_entries_perms_3_u),
    .io_rresp_data_7_entries_perms_3_x(l3_io_rresp_data_7_entries_perms_3_x),
    .io_rresp_data_7_entries_perms_3_w(l3_io_rresp_data_7_entries_perms_3_w),
    .io_rresp_data_7_entries_perms_3_r(l3_io_rresp_data_7_entries_perms_3_r),
    .io_rresp_data_7_entries_perms_4_d(l3_io_rresp_data_7_entries_perms_4_d),
    .io_rresp_data_7_entries_perms_4_a(l3_io_rresp_data_7_entries_perms_4_a),
    .io_rresp_data_7_entries_perms_4_g(l3_io_rresp_data_7_entries_perms_4_g),
    .io_rresp_data_7_entries_perms_4_u(l3_io_rresp_data_7_entries_perms_4_u),
    .io_rresp_data_7_entries_perms_4_x(l3_io_rresp_data_7_entries_perms_4_x),
    .io_rresp_data_7_entries_perms_4_w(l3_io_rresp_data_7_entries_perms_4_w),
    .io_rresp_data_7_entries_perms_4_r(l3_io_rresp_data_7_entries_perms_4_r),
    .io_rresp_data_7_entries_perms_5_d(l3_io_rresp_data_7_entries_perms_5_d),
    .io_rresp_data_7_entries_perms_5_a(l3_io_rresp_data_7_entries_perms_5_a),
    .io_rresp_data_7_entries_perms_5_g(l3_io_rresp_data_7_entries_perms_5_g),
    .io_rresp_data_7_entries_perms_5_u(l3_io_rresp_data_7_entries_perms_5_u),
    .io_rresp_data_7_entries_perms_5_x(l3_io_rresp_data_7_entries_perms_5_x),
    .io_rresp_data_7_entries_perms_5_w(l3_io_rresp_data_7_entries_perms_5_w),
    .io_rresp_data_7_entries_perms_5_r(l3_io_rresp_data_7_entries_perms_5_r),
    .io_rresp_data_7_entries_perms_6_d(l3_io_rresp_data_7_entries_perms_6_d),
    .io_rresp_data_7_entries_perms_6_a(l3_io_rresp_data_7_entries_perms_6_a),
    .io_rresp_data_7_entries_perms_6_g(l3_io_rresp_data_7_entries_perms_6_g),
    .io_rresp_data_7_entries_perms_6_u(l3_io_rresp_data_7_entries_perms_6_u),
    .io_rresp_data_7_entries_perms_6_x(l3_io_rresp_data_7_entries_perms_6_x),
    .io_rresp_data_7_entries_perms_6_w(l3_io_rresp_data_7_entries_perms_6_w),
    .io_rresp_data_7_entries_perms_6_r(l3_io_rresp_data_7_entries_perms_6_r),
    .io_rresp_data_7_entries_perms_7_d(l3_io_rresp_data_7_entries_perms_7_d),
    .io_rresp_data_7_entries_perms_7_a(l3_io_rresp_data_7_entries_perms_7_a),
    .io_rresp_data_7_entries_perms_7_g(l3_io_rresp_data_7_entries_perms_7_g),
    .io_rresp_data_7_entries_perms_7_u(l3_io_rresp_data_7_entries_perms_7_u),
    .io_rresp_data_7_entries_perms_7_x(l3_io_rresp_data_7_entries_perms_7_x),
    .io_rresp_data_7_entries_perms_7_w(l3_io_rresp_data_7_entries_perms_7_w),
    .io_rresp_data_7_entries_perms_7_r(l3_io_rresp_data_7_entries_perms_7_r),
    .io_rresp_data_7_entries_prefetch(l3_io_rresp_data_7_entries_prefetch),
    .io_rresp_data_7_ecc(l3_io_rresp_data_7_ecc),
    .io_wreq_valid(l3_io_wreq_valid),
    .io_wreq_bits_setIdx(l3_io_wreq_bits_setIdx),
    .io_wreq_bits_data_0_entries_tag(l3_io_wreq_bits_data_0_entries_tag),
    .io_wreq_bits_data_0_entries_asid(l3_io_wreq_bits_data_0_entries_asid),
    .io_wreq_bits_data_0_entries_ppns_0(l3_io_wreq_bits_data_0_entries_ppns_0),
    .io_wreq_bits_data_0_entries_ppns_1(l3_io_wreq_bits_data_0_entries_ppns_1),
    .io_wreq_bits_data_0_entries_ppns_2(l3_io_wreq_bits_data_0_entries_ppns_2),
    .io_wreq_bits_data_0_entries_ppns_3(l3_io_wreq_bits_data_0_entries_ppns_3),
    .io_wreq_bits_data_0_entries_ppns_4(l3_io_wreq_bits_data_0_entries_ppns_4),
    .io_wreq_bits_data_0_entries_ppns_5(l3_io_wreq_bits_data_0_entries_ppns_5),
    .io_wreq_bits_data_0_entries_ppns_6(l3_io_wreq_bits_data_0_entries_ppns_6),
    .io_wreq_bits_data_0_entries_ppns_7(l3_io_wreq_bits_data_0_entries_ppns_7),
    .io_wreq_bits_data_0_entries_vs_0(l3_io_wreq_bits_data_0_entries_vs_0),
    .io_wreq_bits_data_0_entries_vs_1(l3_io_wreq_bits_data_0_entries_vs_1),
    .io_wreq_bits_data_0_entries_vs_2(l3_io_wreq_bits_data_0_entries_vs_2),
    .io_wreq_bits_data_0_entries_vs_3(l3_io_wreq_bits_data_0_entries_vs_3),
    .io_wreq_bits_data_0_entries_vs_4(l3_io_wreq_bits_data_0_entries_vs_4),
    .io_wreq_bits_data_0_entries_vs_5(l3_io_wreq_bits_data_0_entries_vs_5),
    .io_wreq_bits_data_0_entries_vs_6(l3_io_wreq_bits_data_0_entries_vs_6),
    .io_wreq_bits_data_0_entries_vs_7(l3_io_wreq_bits_data_0_entries_vs_7),
    .io_wreq_bits_data_0_entries_perms_0_d(l3_io_wreq_bits_data_0_entries_perms_0_d),
    .io_wreq_bits_data_0_entries_perms_0_a(l3_io_wreq_bits_data_0_entries_perms_0_a),
    .io_wreq_bits_data_0_entries_perms_0_g(l3_io_wreq_bits_data_0_entries_perms_0_g),
    .io_wreq_bits_data_0_entries_perms_0_u(l3_io_wreq_bits_data_0_entries_perms_0_u),
    .io_wreq_bits_data_0_entries_perms_0_x(l3_io_wreq_bits_data_0_entries_perms_0_x),
    .io_wreq_bits_data_0_entries_perms_0_w(l3_io_wreq_bits_data_0_entries_perms_0_w),
    .io_wreq_bits_data_0_entries_perms_0_r(l3_io_wreq_bits_data_0_entries_perms_0_r),
    .io_wreq_bits_data_0_entries_perms_1_d(l3_io_wreq_bits_data_0_entries_perms_1_d),
    .io_wreq_bits_data_0_entries_perms_1_a(l3_io_wreq_bits_data_0_entries_perms_1_a),
    .io_wreq_bits_data_0_entries_perms_1_g(l3_io_wreq_bits_data_0_entries_perms_1_g),
    .io_wreq_bits_data_0_entries_perms_1_u(l3_io_wreq_bits_data_0_entries_perms_1_u),
    .io_wreq_bits_data_0_entries_perms_1_x(l3_io_wreq_bits_data_0_entries_perms_1_x),
    .io_wreq_bits_data_0_entries_perms_1_w(l3_io_wreq_bits_data_0_entries_perms_1_w),
    .io_wreq_bits_data_0_entries_perms_1_r(l3_io_wreq_bits_data_0_entries_perms_1_r),
    .io_wreq_bits_data_0_entries_perms_2_d(l3_io_wreq_bits_data_0_entries_perms_2_d),
    .io_wreq_bits_data_0_entries_perms_2_a(l3_io_wreq_bits_data_0_entries_perms_2_a),
    .io_wreq_bits_data_0_entries_perms_2_g(l3_io_wreq_bits_data_0_entries_perms_2_g),
    .io_wreq_bits_data_0_entries_perms_2_u(l3_io_wreq_bits_data_0_entries_perms_2_u),
    .io_wreq_bits_data_0_entries_perms_2_x(l3_io_wreq_bits_data_0_entries_perms_2_x),
    .io_wreq_bits_data_0_entries_perms_2_w(l3_io_wreq_bits_data_0_entries_perms_2_w),
    .io_wreq_bits_data_0_entries_perms_2_r(l3_io_wreq_bits_data_0_entries_perms_2_r),
    .io_wreq_bits_data_0_entries_perms_3_d(l3_io_wreq_bits_data_0_entries_perms_3_d),
    .io_wreq_bits_data_0_entries_perms_3_a(l3_io_wreq_bits_data_0_entries_perms_3_a),
    .io_wreq_bits_data_0_entries_perms_3_g(l3_io_wreq_bits_data_0_entries_perms_3_g),
    .io_wreq_bits_data_0_entries_perms_3_u(l3_io_wreq_bits_data_0_entries_perms_3_u),
    .io_wreq_bits_data_0_entries_perms_3_x(l3_io_wreq_bits_data_0_entries_perms_3_x),
    .io_wreq_bits_data_0_entries_perms_3_w(l3_io_wreq_bits_data_0_entries_perms_3_w),
    .io_wreq_bits_data_0_entries_perms_3_r(l3_io_wreq_bits_data_0_entries_perms_3_r),
    .io_wreq_bits_data_0_entries_perms_4_d(l3_io_wreq_bits_data_0_entries_perms_4_d),
    .io_wreq_bits_data_0_entries_perms_4_a(l3_io_wreq_bits_data_0_entries_perms_4_a),
    .io_wreq_bits_data_0_entries_perms_4_g(l3_io_wreq_bits_data_0_entries_perms_4_g),
    .io_wreq_bits_data_0_entries_perms_4_u(l3_io_wreq_bits_data_0_entries_perms_4_u),
    .io_wreq_bits_data_0_entries_perms_4_x(l3_io_wreq_bits_data_0_entries_perms_4_x),
    .io_wreq_bits_data_0_entries_perms_4_w(l3_io_wreq_bits_data_0_entries_perms_4_w),
    .io_wreq_bits_data_0_entries_perms_4_r(l3_io_wreq_bits_data_0_entries_perms_4_r),
    .io_wreq_bits_data_0_entries_perms_5_d(l3_io_wreq_bits_data_0_entries_perms_5_d),
    .io_wreq_bits_data_0_entries_perms_5_a(l3_io_wreq_bits_data_0_entries_perms_5_a),
    .io_wreq_bits_data_0_entries_perms_5_g(l3_io_wreq_bits_data_0_entries_perms_5_g),
    .io_wreq_bits_data_0_entries_perms_5_u(l3_io_wreq_bits_data_0_entries_perms_5_u),
    .io_wreq_bits_data_0_entries_perms_5_x(l3_io_wreq_bits_data_0_entries_perms_5_x),
    .io_wreq_bits_data_0_entries_perms_5_w(l3_io_wreq_bits_data_0_entries_perms_5_w),
    .io_wreq_bits_data_0_entries_perms_5_r(l3_io_wreq_bits_data_0_entries_perms_5_r),
    .io_wreq_bits_data_0_entries_perms_6_d(l3_io_wreq_bits_data_0_entries_perms_6_d),
    .io_wreq_bits_data_0_entries_perms_6_a(l3_io_wreq_bits_data_0_entries_perms_6_a),
    .io_wreq_bits_data_0_entries_perms_6_g(l3_io_wreq_bits_data_0_entries_perms_6_g),
    .io_wreq_bits_data_0_entries_perms_6_u(l3_io_wreq_bits_data_0_entries_perms_6_u),
    .io_wreq_bits_data_0_entries_perms_6_x(l3_io_wreq_bits_data_0_entries_perms_6_x),
    .io_wreq_bits_data_0_entries_perms_6_w(l3_io_wreq_bits_data_0_entries_perms_6_w),
    .io_wreq_bits_data_0_entries_perms_6_r(l3_io_wreq_bits_data_0_entries_perms_6_r),
    .io_wreq_bits_data_0_entries_perms_7_d(l3_io_wreq_bits_data_0_entries_perms_7_d),
    .io_wreq_bits_data_0_entries_perms_7_a(l3_io_wreq_bits_data_0_entries_perms_7_a),
    .io_wreq_bits_data_0_entries_perms_7_g(l3_io_wreq_bits_data_0_entries_perms_7_g),
    .io_wreq_bits_data_0_entries_perms_7_u(l3_io_wreq_bits_data_0_entries_perms_7_u),
    .io_wreq_bits_data_0_entries_perms_7_x(l3_io_wreq_bits_data_0_entries_perms_7_x),
    .io_wreq_bits_data_0_entries_perms_7_w(l3_io_wreq_bits_data_0_entries_perms_7_w),
    .io_wreq_bits_data_0_entries_perms_7_r(l3_io_wreq_bits_data_0_entries_perms_7_r),
    .io_wreq_bits_data_0_entries_prefetch(l3_io_wreq_bits_data_0_entries_prefetch),
    .io_wreq_bits_data_0_ecc(l3_io_wreq_bits_data_0_ecc),
    .io_wreq_bits_data_1_entries_tag(l3_io_wreq_bits_data_1_entries_tag),
    .io_wreq_bits_data_1_entries_asid(l3_io_wreq_bits_data_1_entries_asid),
    .io_wreq_bits_data_1_entries_ppns_0(l3_io_wreq_bits_data_1_entries_ppns_0),
    .io_wreq_bits_data_1_entries_ppns_1(l3_io_wreq_bits_data_1_entries_ppns_1),
    .io_wreq_bits_data_1_entries_ppns_2(l3_io_wreq_bits_data_1_entries_ppns_2),
    .io_wreq_bits_data_1_entries_ppns_3(l3_io_wreq_bits_data_1_entries_ppns_3),
    .io_wreq_bits_data_1_entries_ppns_4(l3_io_wreq_bits_data_1_entries_ppns_4),
    .io_wreq_bits_data_1_entries_ppns_5(l3_io_wreq_bits_data_1_entries_ppns_5),
    .io_wreq_bits_data_1_entries_ppns_6(l3_io_wreq_bits_data_1_entries_ppns_6),
    .io_wreq_bits_data_1_entries_ppns_7(l3_io_wreq_bits_data_1_entries_ppns_7),
    .io_wreq_bits_data_1_entries_vs_0(l3_io_wreq_bits_data_1_entries_vs_0),
    .io_wreq_bits_data_1_entries_vs_1(l3_io_wreq_bits_data_1_entries_vs_1),
    .io_wreq_bits_data_1_entries_vs_2(l3_io_wreq_bits_data_1_entries_vs_2),
    .io_wreq_bits_data_1_entries_vs_3(l3_io_wreq_bits_data_1_entries_vs_3),
    .io_wreq_bits_data_1_entries_vs_4(l3_io_wreq_bits_data_1_entries_vs_4),
    .io_wreq_bits_data_1_entries_vs_5(l3_io_wreq_bits_data_1_entries_vs_5),
    .io_wreq_bits_data_1_entries_vs_6(l3_io_wreq_bits_data_1_entries_vs_6),
    .io_wreq_bits_data_1_entries_vs_7(l3_io_wreq_bits_data_1_entries_vs_7),
    .io_wreq_bits_data_1_entries_perms_0_d(l3_io_wreq_bits_data_1_entries_perms_0_d),
    .io_wreq_bits_data_1_entries_perms_0_a(l3_io_wreq_bits_data_1_entries_perms_0_a),
    .io_wreq_bits_data_1_entries_perms_0_g(l3_io_wreq_bits_data_1_entries_perms_0_g),
    .io_wreq_bits_data_1_entries_perms_0_u(l3_io_wreq_bits_data_1_entries_perms_0_u),
    .io_wreq_bits_data_1_entries_perms_0_x(l3_io_wreq_bits_data_1_entries_perms_0_x),
    .io_wreq_bits_data_1_entries_perms_0_w(l3_io_wreq_bits_data_1_entries_perms_0_w),
    .io_wreq_bits_data_1_entries_perms_0_r(l3_io_wreq_bits_data_1_entries_perms_0_r),
    .io_wreq_bits_data_1_entries_perms_1_d(l3_io_wreq_bits_data_1_entries_perms_1_d),
    .io_wreq_bits_data_1_entries_perms_1_a(l3_io_wreq_bits_data_1_entries_perms_1_a),
    .io_wreq_bits_data_1_entries_perms_1_g(l3_io_wreq_bits_data_1_entries_perms_1_g),
    .io_wreq_bits_data_1_entries_perms_1_u(l3_io_wreq_bits_data_1_entries_perms_1_u),
    .io_wreq_bits_data_1_entries_perms_1_x(l3_io_wreq_bits_data_1_entries_perms_1_x),
    .io_wreq_bits_data_1_entries_perms_1_w(l3_io_wreq_bits_data_1_entries_perms_1_w),
    .io_wreq_bits_data_1_entries_perms_1_r(l3_io_wreq_bits_data_1_entries_perms_1_r),
    .io_wreq_bits_data_1_entries_perms_2_d(l3_io_wreq_bits_data_1_entries_perms_2_d),
    .io_wreq_bits_data_1_entries_perms_2_a(l3_io_wreq_bits_data_1_entries_perms_2_a),
    .io_wreq_bits_data_1_entries_perms_2_g(l3_io_wreq_bits_data_1_entries_perms_2_g),
    .io_wreq_bits_data_1_entries_perms_2_u(l3_io_wreq_bits_data_1_entries_perms_2_u),
    .io_wreq_bits_data_1_entries_perms_2_x(l3_io_wreq_bits_data_1_entries_perms_2_x),
    .io_wreq_bits_data_1_entries_perms_2_w(l3_io_wreq_bits_data_1_entries_perms_2_w),
    .io_wreq_bits_data_1_entries_perms_2_r(l3_io_wreq_bits_data_1_entries_perms_2_r),
    .io_wreq_bits_data_1_entries_perms_3_d(l3_io_wreq_bits_data_1_entries_perms_3_d),
    .io_wreq_bits_data_1_entries_perms_3_a(l3_io_wreq_bits_data_1_entries_perms_3_a),
    .io_wreq_bits_data_1_entries_perms_3_g(l3_io_wreq_bits_data_1_entries_perms_3_g),
    .io_wreq_bits_data_1_entries_perms_3_u(l3_io_wreq_bits_data_1_entries_perms_3_u),
    .io_wreq_bits_data_1_entries_perms_3_x(l3_io_wreq_bits_data_1_entries_perms_3_x),
    .io_wreq_bits_data_1_entries_perms_3_w(l3_io_wreq_bits_data_1_entries_perms_3_w),
    .io_wreq_bits_data_1_entries_perms_3_r(l3_io_wreq_bits_data_1_entries_perms_3_r),
    .io_wreq_bits_data_1_entries_perms_4_d(l3_io_wreq_bits_data_1_entries_perms_4_d),
    .io_wreq_bits_data_1_entries_perms_4_a(l3_io_wreq_bits_data_1_entries_perms_4_a),
    .io_wreq_bits_data_1_entries_perms_4_g(l3_io_wreq_bits_data_1_entries_perms_4_g),
    .io_wreq_bits_data_1_entries_perms_4_u(l3_io_wreq_bits_data_1_entries_perms_4_u),
    .io_wreq_bits_data_1_entries_perms_4_x(l3_io_wreq_bits_data_1_entries_perms_4_x),
    .io_wreq_bits_data_1_entries_perms_4_w(l3_io_wreq_bits_data_1_entries_perms_4_w),
    .io_wreq_bits_data_1_entries_perms_4_r(l3_io_wreq_bits_data_1_entries_perms_4_r),
    .io_wreq_bits_data_1_entries_perms_5_d(l3_io_wreq_bits_data_1_entries_perms_5_d),
    .io_wreq_bits_data_1_entries_perms_5_a(l3_io_wreq_bits_data_1_entries_perms_5_a),
    .io_wreq_bits_data_1_entries_perms_5_g(l3_io_wreq_bits_data_1_entries_perms_5_g),
    .io_wreq_bits_data_1_entries_perms_5_u(l3_io_wreq_bits_data_1_entries_perms_5_u),
    .io_wreq_bits_data_1_entries_perms_5_x(l3_io_wreq_bits_data_1_entries_perms_5_x),
    .io_wreq_bits_data_1_entries_perms_5_w(l3_io_wreq_bits_data_1_entries_perms_5_w),
    .io_wreq_bits_data_1_entries_perms_5_r(l3_io_wreq_bits_data_1_entries_perms_5_r),
    .io_wreq_bits_data_1_entries_perms_6_d(l3_io_wreq_bits_data_1_entries_perms_6_d),
    .io_wreq_bits_data_1_entries_perms_6_a(l3_io_wreq_bits_data_1_entries_perms_6_a),
    .io_wreq_bits_data_1_entries_perms_6_g(l3_io_wreq_bits_data_1_entries_perms_6_g),
    .io_wreq_bits_data_1_entries_perms_6_u(l3_io_wreq_bits_data_1_entries_perms_6_u),
    .io_wreq_bits_data_1_entries_perms_6_x(l3_io_wreq_bits_data_1_entries_perms_6_x),
    .io_wreq_bits_data_1_entries_perms_6_w(l3_io_wreq_bits_data_1_entries_perms_6_w),
    .io_wreq_bits_data_1_entries_perms_6_r(l3_io_wreq_bits_data_1_entries_perms_6_r),
    .io_wreq_bits_data_1_entries_perms_7_d(l3_io_wreq_bits_data_1_entries_perms_7_d),
    .io_wreq_bits_data_1_entries_perms_7_a(l3_io_wreq_bits_data_1_entries_perms_7_a),
    .io_wreq_bits_data_1_entries_perms_7_g(l3_io_wreq_bits_data_1_entries_perms_7_g),
    .io_wreq_bits_data_1_entries_perms_7_u(l3_io_wreq_bits_data_1_entries_perms_7_u),
    .io_wreq_bits_data_1_entries_perms_7_x(l3_io_wreq_bits_data_1_entries_perms_7_x),
    .io_wreq_bits_data_1_entries_perms_7_w(l3_io_wreq_bits_data_1_entries_perms_7_w),
    .io_wreq_bits_data_1_entries_perms_7_r(l3_io_wreq_bits_data_1_entries_perms_7_r),
    .io_wreq_bits_data_1_entries_prefetch(l3_io_wreq_bits_data_1_entries_prefetch),
    .io_wreq_bits_data_1_ecc(l3_io_wreq_bits_data_1_ecc),
    .io_wreq_bits_data_2_entries_tag(l3_io_wreq_bits_data_2_entries_tag),
    .io_wreq_bits_data_2_entries_asid(l3_io_wreq_bits_data_2_entries_asid),
    .io_wreq_bits_data_2_entries_ppns_0(l3_io_wreq_bits_data_2_entries_ppns_0),
    .io_wreq_bits_data_2_entries_ppns_1(l3_io_wreq_bits_data_2_entries_ppns_1),
    .io_wreq_bits_data_2_entries_ppns_2(l3_io_wreq_bits_data_2_entries_ppns_2),
    .io_wreq_bits_data_2_entries_ppns_3(l3_io_wreq_bits_data_2_entries_ppns_3),
    .io_wreq_bits_data_2_entries_ppns_4(l3_io_wreq_bits_data_2_entries_ppns_4),
    .io_wreq_bits_data_2_entries_ppns_5(l3_io_wreq_bits_data_2_entries_ppns_5),
    .io_wreq_bits_data_2_entries_ppns_6(l3_io_wreq_bits_data_2_entries_ppns_6),
    .io_wreq_bits_data_2_entries_ppns_7(l3_io_wreq_bits_data_2_entries_ppns_7),
    .io_wreq_bits_data_2_entries_vs_0(l3_io_wreq_bits_data_2_entries_vs_0),
    .io_wreq_bits_data_2_entries_vs_1(l3_io_wreq_bits_data_2_entries_vs_1),
    .io_wreq_bits_data_2_entries_vs_2(l3_io_wreq_bits_data_2_entries_vs_2),
    .io_wreq_bits_data_2_entries_vs_3(l3_io_wreq_bits_data_2_entries_vs_3),
    .io_wreq_bits_data_2_entries_vs_4(l3_io_wreq_bits_data_2_entries_vs_4),
    .io_wreq_bits_data_2_entries_vs_5(l3_io_wreq_bits_data_2_entries_vs_5),
    .io_wreq_bits_data_2_entries_vs_6(l3_io_wreq_bits_data_2_entries_vs_6),
    .io_wreq_bits_data_2_entries_vs_7(l3_io_wreq_bits_data_2_entries_vs_7),
    .io_wreq_bits_data_2_entries_perms_0_d(l3_io_wreq_bits_data_2_entries_perms_0_d),
    .io_wreq_bits_data_2_entries_perms_0_a(l3_io_wreq_bits_data_2_entries_perms_0_a),
    .io_wreq_bits_data_2_entries_perms_0_g(l3_io_wreq_bits_data_2_entries_perms_0_g),
    .io_wreq_bits_data_2_entries_perms_0_u(l3_io_wreq_bits_data_2_entries_perms_0_u),
    .io_wreq_bits_data_2_entries_perms_0_x(l3_io_wreq_bits_data_2_entries_perms_0_x),
    .io_wreq_bits_data_2_entries_perms_0_w(l3_io_wreq_bits_data_2_entries_perms_0_w),
    .io_wreq_bits_data_2_entries_perms_0_r(l3_io_wreq_bits_data_2_entries_perms_0_r),
    .io_wreq_bits_data_2_entries_perms_1_d(l3_io_wreq_bits_data_2_entries_perms_1_d),
    .io_wreq_bits_data_2_entries_perms_1_a(l3_io_wreq_bits_data_2_entries_perms_1_a),
    .io_wreq_bits_data_2_entries_perms_1_g(l3_io_wreq_bits_data_2_entries_perms_1_g),
    .io_wreq_bits_data_2_entries_perms_1_u(l3_io_wreq_bits_data_2_entries_perms_1_u),
    .io_wreq_bits_data_2_entries_perms_1_x(l3_io_wreq_bits_data_2_entries_perms_1_x),
    .io_wreq_bits_data_2_entries_perms_1_w(l3_io_wreq_bits_data_2_entries_perms_1_w),
    .io_wreq_bits_data_2_entries_perms_1_r(l3_io_wreq_bits_data_2_entries_perms_1_r),
    .io_wreq_bits_data_2_entries_perms_2_d(l3_io_wreq_bits_data_2_entries_perms_2_d),
    .io_wreq_bits_data_2_entries_perms_2_a(l3_io_wreq_bits_data_2_entries_perms_2_a),
    .io_wreq_bits_data_2_entries_perms_2_g(l3_io_wreq_bits_data_2_entries_perms_2_g),
    .io_wreq_bits_data_2_entries_perms_2_u(l3_io_wreq_bits_data_2_entries_perms_2_u),
    .io_wreq_bits_data_2_entries_perms_2_x(l3_io_wreq_bits_data_2_entries_perms_2_x),
    .io_wreq_bits_data_2_entries_perms_2_w(l3_io_wreq_bits_data_2_entries_perms_2_w),
    .io_wreq_bits_data_2_entries_perms_2_r(l3_io_wreq_bits_data_2_entries_perms_2_r),
    .io_wreq_bits_data_2_entries_perms_3_d(l3_io_wreq_bits_data_2_entries_perms_3_d),
    .io_wreq_bits_data_2_entries_perms_3_a(l3_io_wreq_bits_data_2_entries_perms_3_a),
    .io_wreq_bits_data_2_entries_perms_3_g(l3_io_wreq_bits_data_2_entries_perms_3_g),
    .io_wreq_bits_data_2_entries_perms_3_u(l3_io_wreq_bits_data_2_entries_perms_3_u),
    .io_wreq_bits_data_2_entries_perms_3_x(l3_io_wreq_bits_data_2_entries_perms_3_x),
    .io_wreq_bits_data_2_entries_perms_3_w(l3_io_wreq_bits_data_2_entries_perms_3_w),
    .io_wreq_bits_data_2_entries_perms_3_r(l3_io_wreq_bits_data_2_entries_perms_3_r),
    .io_wreq_bits_data_2_entries_perms_4_d(l3_io_wreq_bits_data_2_entries_perms_4_d),
    .io_wreq_bits_data_2_entries_perms_4_a(l3_io_wreq_bits_data_2_entries_perms_4_a),
    .io_wreq_bits_data_2_entries_perms_4_g(l3_io_wreq_bits_data_2_entries_perms_4_g),
    .io_wreq_bits_data_2_entries_perms_4_u(l3_io_wreq_bits_data_2_entries_perms_4_u),
    .io_wreq_bits_data_2_entries_perms_4_x(l3_io_wreq_bits_data_2_entries_perms_4_x),
    .io_wreq_bits_data_2_entries_perms_4_w(l3_io_wreq_bits_data_2_entries_perms_4_w),
    .io_wreq_bits_data_2_entries_perms_4_r(l3_io_wreq_bits_data_2_entries_perms_4_r),
    .io_wreq_bits_data_2_entries_perms_5_d(l3_io_wreq_bits_data_2_entries_perms_5_d),
    .io_wreq_bits_data_2_entries_perms_5_a(l3_io_wreq_bits_data_2_entries_perms_5_a),
    .io_wreq_bits_data_2_entries_perms_5_g(l3_io_wreq_bits_data_2_entries_perms_5_g),
    .io_wreq_bits_data_2_entries_perms_5_u(l3_io_wreq_bits_data_2_entries_perms_5_u),
    .io_wreq_bits_data_2_entries_perms_5_x(l3_io_wreq_bits_data_2_entries_perms_5_x),
    .io_wreq_bits_data_2_entries_perms_5_w(l3_io_wreq_bits_data_2_entries_perms_5_w),
    .io_wreq_bits_data_2_entries_perms_5_r(l3_io_wreq_bits_data_2_entries_perms_5_r),
    .io_wreq_bits_data_2_entries_perms_6_d(l3_io_wreq_bits_data_2_entries_perms_6_d),
    .io_wreq_bits_data_2_entries_perms_6_a(l3_io_wreq_bits_data_2_entries_perms_6_a),
    .io_wreq_bits_data_2_entries_perms_6_g(l3_io_wreq_bits_data_2_entries_perms_6_g),
    .io_wreq_bits_data_2_entries_perms_6_u(l3_io_wreq_bits_data_2_entries_perms_6_u),
    .io_wreq_bits_data_2_entries_perms_6_x(l3_io_wreq_bits_data_2_entries_perms_6_x),
    .io_wreq_bits_data_2_entries_perms_6_w(l3_io_wreq_bits_data_2_entries_perms_6_w),
    .io_wreq_bits_data_2_entries_perms_6_r(l3_io_wreq_bits_data_2_entries_perms_6_r),
    .io_wreq_bits_data_2_entries_perms_7_d(l3_io_wreq_bits_data_2_entries_perms_7_d),
    .io_wreq_bits_data_2_entries_perms_7_a(l3_io_wreq_bits_data_2_entries_perms_7_a),
    .io_wreq_bits_data_2_entries_perms_7_g(l3_io_wreq_bits_data_2_entries_perms_7_g),
    .io_wreq_bits_data_2_entries_perms_7_u(l3_io_wreq_bits_data_2_entries_perms_7_u),
    .io_wreq_bits_data_2_entries_perms_7_x(l3_io_wreq_bits_data_2_entries_perms_7_x),
    .io_wreq_bits_data_2_entries_perms_7_w(l3_io_wreq_bits_data_2_entries_perms_7_w),
    .io_wreq_bits_data_2_entries_perms_7_r(l3_io_wreq_bits_data_2_entries_perms_7_r),
    .io_wreq_bits_data_2_entries_prefetch(l3_io_wreq_bits_data_2_entries_prefetch),
    .io_wreq_bits_data_2_ecc(l3_io_wreq_bits_data_2_ecc),
    .io_wreq_bits_data_3_entries_tag(l3_io_wreq_bits_data_3_entries_tag),
    .io_wreq_bits_data_3_entries_asid(l3_io_wreq_bits_data_3_entries_asid),
    .io_wreq_bits_data_3_entries_ppns_0(l3_io_wreq_bits_data_3_entries_ppns_0),
    .io_wreq_bits_data_3_entries_ppns_1(l3_io_wreq_bits_data_3_entries_ppns_1),
    .io_wreq_bits_data_3_entries_ppns_2(l3_io_wreq_bits_data_3_entries_ppns_2),
    .io_wreq_bits_data_3_entries_ppns_3(l3_io_wreq_bits_data_3_entries_ppns_3),
    .io_wreq_bits_data_3_entries_ppns_4(l3_io_wreq_bits_data_3_entries_ppns_4),
    .io_wreq_bits_data_3_entries_ppns_5(l3_io_wreq_bits_data_3_entries_ppns_5),
    .io_wreq_bits_data_3_entries_ppns_6(l3_io_wreq_bits_data_3_entries_ppns_6),
    .io_wreq_bits_data_3_entries_ppns_7(l3_io_wreq_bits_data_3_entries_ppns_7),
    .io_wreq_bits_data_3_entries_vs_0(l3_io_wreq_bits_data_3_entries_vs_0),
    .io_wreq_bits_data_3_entries_vs_1(l3_io_wreq_bits_data_3_entries_vs_1),
    .io_wreq_bits_data_3_entries_vs_2(l3_io_wreq_bits_data_3_entries_vs_2),
    .io_wreq_bits_data_3_entries_vs_3(l3_io_wreq_bits_data_3_entries_vs_3),
    .io_wreq_bits_data_3_entries_vs_4(l3_io_wreq_bits_data_3_entries_vs_4),
    .io_wreq_bits_data_3_entries_vs_5(l3_io_wreq_bits_data_3_entries_vs_5),
    .io_wreq_bits_data_3_entries_vs_6(l3_io_wreq_bits_data_3_entries_vs_6),
    .io_wreq_bits_data_3_entries_vs_7(l3_io_wreq_bits_data_3_entries_vs_7),
    .io_wreq_bits_data_3_entries_perms_0_d(l3_io_wreq_bits_data_3_entries_perms_0_d),
    .io_wreq_bits_data_3_entries_perms_0_a(l3_io_wreq_bits_data_3_entries_perms_0_a),
    .io_wreq_bits_data_3_entries_perms_0_g(l3_io_wreq_bits_data_3_entries_perms_0_g),
    .io_wreq_bits_data_3_entries_perms_0_u(l3_io_wreq_bits_data_3_entries_perms_0_u),
    .io_wreq_bits_data_3_entries_perms_0_x(l3_io_wreq_bits_data_3_entries_perms_0_x),
    .io_wreq_bits_data_3_entries_perms_0_w(l3_io_wreq_bits_data_3_entries_perms_0_w),
    .io_wreq_bits_data_3_entries_perms_0_r(l3_io_wreq_bits_data_3_entries_perms_0_r),
    .io_wreq_bits_data_3_entries_perms_1_d(l3_io_wreq_bits_data_3_entries_perms_1_d),
    .io_wreq_bits_data_3_entries_perms_1_a(l3_io_wreq_bits_data_3_entries_perms_1_a),
    .io_wreq_bits_data_3_entries_perms_1_g(l3_io_wreq_bits_data_3_entries_perms_1_g),
    .io_wreq_bits_data_3_entries_perms_1_u(l3_io_wreq_bits_data_3_entries_perms_1_u),
    .io_wreq_bits_data_3_entries_perms_1_x(l3_io_wreq_bits_data_3_entries_perms_1_x),
    .io_wreq_bits_data_3_entries_perms_1_w(l3_io_wreq_bits_data_3_entries_perms_1_w),
    .io_wreq_bits_data_3_entries_perms_1_r(l3_io_wreq_bits_data_3_entries_perms_1_r),
    .io_wreq_bits_data_3_entries_perms_2_d(l3_io_wreq_bits_data_3_entries_perms_2_d),
    .io_wreq_bits_data_3_entries_perms_2_a(l3_io_wreq_bits_data_3_entries_perms_2_a),
    .io_wreq_bits_data_3_entries_perms_2_g(l3_io_wreq_bits_data_3_entries_perms_2_g),
    .io_wreq_bits_data_3_entries_perms_2_u(l3_io_wreq_bits_data_3_entries_perms_2_u),
    .io_wreq_bits_data_3_entries_perms_2_x(l3_io_wreq_bits_data_3_entries_perms_2_x),
    .io_wreq_bits_data_3_entries_perms_2_w(l3_io_wreq_bits_data_3_entries_perms_2_w),
    .io_wreq_bits_data_3_entries_perms_2_r(l3_io_wreq_bits_data_3_entries_perms_2_r),
    .io_wreq_bits_data_3_entries_perms_3_d(l3_io_wreq_bits_data_3_entries_perms_3_d),
    .io_wreq_bits_data_3_entries_perms_3_a(l3_io_wreq_bits_data_3_entries_perms_3_a),
    .io_wreq_bits_data_3_entries_perms_3_g(l3_io_wreq_bits_data_3_entries_perms_3_g),
    .io_wreq_bits_data_3_entries_perms_3_u(l3_io_wreq_bits_data_3_entries_perms_3_u),
    .io_wreq_bits_data_3_entries_perms_3_x(l3_io_wreq_bits_data_3_entries_perms_3_x),
    .io_wreq_bits_data_3_entries_perms_3_w(l3_io_wreq_bits_data_3_entries_perms_3_w),
    .io_wreq_bits_data_3_entries_perms_3_r(l3_io_wreq_bits_data_3_entries_perms_3_r),
    .io_wreq_bits_data_3_entries_perms_4_d(l3_io_wreq_bits_data_3_entries_perms_4_d),
    .io_wreq_bits_data_3_entries_perms_4_a(l3_io_wreq_bits_data_3_entries_perms_4_a),
    .io_wreq_bits_data_3_entries_perms_4_g(l3_io_wreq_bits_data_3_entries_perms_4_g),
    .io_wreq_bits_data_3_entries_perms_4_u(l3_io_wreq_bits_data_3_entries_perms_4_u),
    .io_wreq_bits_data_3_entries_perms_4_x(l3_io_wreq_bits_data_3_entries_perms_4_x),
    .io_wreq_bits_data_3_entries_perms_4_w(l3_io_wreq_bits_data_3_entries_perms_4_w),
    .io_wreq_bits_data_3_entries_perms_4_r(l3_io_wreq_bits_data_3_entries_perms_4_r),
    .io_wreq_bits_data_3_entries_perms_5_d(l3_io_wreq_bits_data_3_entries_perms_5_d),
    .io_wreq_bits_data_3_entries_perms_5_a(l3_io_wreq_bits_data_3_entries_perms_5_a),
    .io_wreq_bits_data_3_entries_perms_5_g(l3_io_wreq_bits_data_3_entries_perms_5_g),
    .io_wreq_bits_data_3_entries_perms_5_u(l3_io_wreq_bits_data_3_entries_perms_5_u),
    .io_wreq_bits_data_3_entries_perms_5_x(l3_io_wreq_bits_data_3_entries_perms_5_x),
    .io_wreq_bits_data_3_entries_perms_5_w(l3_io_wreq_bits_data_3_entries_perms_5_w),
    .io_wreq_bits_data_3_entries_perms_5_r(l3_io_wreq_bits_data_3_entries_perms_5_r),
    .io_wreq_bits_data_3_entries_perms_6_d(l3_io_wreq_bits_data_3_entries_perms_6_d),
    .io_wreq_bits_data_3_entries_perms_6_a(l3_io_wreq_bits_data_3_entries_perms_6_a),
    .io_wreq_bits_data_3_entries_perms_6_g(l3_io_wreq_bits_data_3_entries_perms_6_g),
    .io_wreq_bits_data_3_entries_perms_6_u(l3_io_wreq_bits_data_3_entries_perms_6_u),
    .io_wreq_bits_data_3_entries_perms_6_x(l3_io_wreq_bits_data_3_entries_perms_6_x),
    .io_wreq_bits_data_3_entries_perms_6_w(l3_io_wreq_bits_data_3_entries_perms_6_w),
    .io_wreq_bits_data_3_entries_perms_6_r(l3_io_wreq_bits_data_3_entries_perms_6_r),
    .io_wreq_bits_data_3_entries_perms_7_d(l3_io_wreq_bits_data_3_entries_perms_7_d),
    .io_wreq_bits_data_3_entries_perms_7_a(l3_io_wreq_bits_data_3_entries_perms_7_a),
    .io_wreq_bits_data_3_entries_perms_7_g(l3_io_wreq_bits_data_3_entries_perms_7_g),
    .io_wreq_bits_data_3_entries_perms_7_u(l3_io_wreq_bits_data_3_entries_perms_7_u),
    .io_wreq_bits_data_3_entries_perms_7_x(l3_io_wreq_bits_data_3_entries_perms_7_x),
    .io_wreq_bits_data_3_entries_perms_7_w(l3_io_wreq_bits_data_3_entries_perms_7_w),
    .io_wreq_bits_data_3_entries_perms_7_r(l3_io_wreq_bits_data_3_entries_perms_7_r),
    .io_wreq_bits_data_3_entries_prefetch(l3_io_wreq_bits_data_3_entries_prefetch),
    .io_wreq_bits_data_3_ecc(l3_io_wreq_bits_data_3_ecc),
    .io_wreq_bits_data_4_entries_tag(l3_io_wreq_bits_data_4_entries_tag),
    .io_wreq_bits_data_4_entries_asid(l3_io_wreq_bits_data_4_entries_asid),
    .io_wreq_bits_data_4_entries_ppns_0(l3_io_wreq_bits_data_4_entries_ppns_0),
    .io_wreq_bits_data_4_entries_ppns_1(l3_io_wreq_bits_data_4_entries_ppns_1),
    .io_wreq_bits_data_4_entries_ppns_2(l3_io_wreq_bits_data_4_entries_ppns_2),
    .io_wreq_bits_data_4_entries_ppns_3(l3_io_wreq_bits_data_4_entries_ppns_3),
    .io_wreq_bits_data_4_entries_ppns_4(l3_io_wreq_bits_data_4_entries_ppns_4),
    .io_wreq_bits_data_4_entries_ppns_5(l3_io_wreq_bits_data_4_entries_ppns_5),
    .io_wreq_bits_data_4_entries_ppns_6(l3_io_wreq_bits_data_4_entries_ppns_6),
    .io_wreq_bits_data_4_entries_ppns_7(l3_io_wreq_bits_data_4_entries_ppns_7),
    .io_wreq_bits_data_4_entries_vs_0(l3_io_wreq_bits_data_4_entries_vs_0),
    .io_wreq_bits_data_4_entries_vs_1(l3_io_wreq_bits_data_4_entries_vs_1),
    .io_wreq_bits_data_4_entries_vs_2(l3_io_wreq_bits_data_4_entries_vs_2),
    .io_wreq_bits_data_4_entries_vs_3(l3_io_wreq_bits_data_4_entries_vs_3),
    .io_wreq_bits_data_4_entries_vs_4(l3_io_wreq_bits_data_4_entries_vs_4),
    .io_wreq_bits_data_4_entries_vs_5(l3_io_wreq_bits_data_4_entries_vs_5),
    .io_wreq_bits_data_4_entries_vs_6(l3_io_wreq_bits_data_4_entries_vs_6),
    .io_wreq_bits_data_4_entries_vs_7(l3_io_wreq_bits_data_4_entries_vs_7),
    .io_wreq_bits_data_4_entries_perms_0_d(l3_io_wreq_bits_data_4_entries_perms_0_d),
    .io_wreq_bits_data_4_entries_perms_0_a(l3_io_wreq_bits_data_4_entries_perms_0_a),
    .io_wreq_bits_data_4_entries_perms_0_g(l3_io_wreq_bits_data_4_entries_perms_0_g),
    .io_wreq_bits_data_4_entries_perms_0_u(l3_io_wreq_bits_data_4_entries_perms_0_u),
    .io_wreq_bits_data_4_entries_perms_0_x(l3_io_wreq_bits_data_4_entries_perms_0_x),
    .io_wreq_bits_data_4_entries_perms_0_w(l3_io_wreq_bits_data_4_entries_perms_0_w),
    .io_wreq_bits_data_4_entries_perms_0_r(l3_io_wreq_bits_data_4_entries_perms_0_r),
    .io_wreq_bits_data_4_entries_perms_1_d(l3_io_wreq_bits_data_4_entries_perms_1_d),
    .io_wreq_bits_data_4_entries_perms_1_a(l3_io_wreq_bits_data_4_entries_perms_1_a),
    .io_wreq_bits_data_4_entries_perms_1_g(l3_io_wreq_bits_data_4_entries_perms_1_g),
    .io_wreq_bits_data_4_entries_perms_1_u(l3_io_wreq_bits_data_4_entries_perms_1_u),
    .io_wreq_bits_data_4_entries_perms_1_x(l3_io_wreq_bits_data_4_entries_perms_1_x),
    .io_wreq_bits_data_4_entries_perms_1_w(l3_io_wreq_bits_data_4_entries_perms_1_w),
    .io_wreq_bits_data_4_entries_perms_1_r(l3_io_wreq_bits_data_4_entries_perms_1_r),
    .io_wreq_bits_data_4_entries_perms_2_d(l3_io_wreq_bits_data_4_entries_perms_2_d),
    .io_wreq_bits_data_4_entries_perms_2_a(l3_io_wreq_bits_data_4_entries_perms_2_a),
    .io_wreq_bits_data_4_entries_perms_2_g(l3_io_wreq_bits_data_4_entries_perms_2_g),
    .io_wreq_bits_data_4_entries_perms_2_u(l3_io_wreq_bits_data_4_entries_perms_2_u),
    .io_wreq_bits_data_4_entries_perms_2_x(l3_io_wreq_bits_data_4_entries_perms_2_x),
    .io_wreq_bits_data_4_entries_perms_2_w(l3_io_wreq_bits_data_4_entries_perms_2_w),
    .io_wreq_bits_data_4_entries_perms_2_r(l3_io_wreq_bits_data_4_entries_perms_2_r),
    .io_wreq_bits_data_4_entries_perms_3_d(l3_io_wreq_bits_data_4_entries_perms_3_d),
    .io_wreq_bits_data_4_entries_perms_3_a(l3_io_wreq_bits_data_4_entries_perms_3_a),
    .io_wreq_bits_data_4_entries_perms_3_g(l3_io_wreq_bits_data_4_entries_perms_3_g),
    .io_wreq_bits_data_4_entries_perms_3_u(l3_io_wreq_bits_data_4_entries_perms_3_u),
    .io_wreq_bits_data_4_entries_perms_3_x(l3_io_wreq_bits_data_4_entries_perms_3_x),
    .io_wreq_bits_data_4_entries_perms_3_w(l3_io_wreq_bits_data_4_entries_perms_3_w),
    .io_wreq_bits_data_4_entries_perms_3_r(l3_io_wreq_bits_data_4_entries_perms_3_r),
    .io_wreq_bits_data_4_entries_perms_4_d(l3_io_wreq_bits_data_4_entries_perms_4_d),
    .io_wreq_bits_data_4_entries_perms_4_a(l3_io_wreq_bits_data_4_entries_perms_4_a),
    .io_wreq_bits_data_4_entries_perms_4_g(l3_io_wreq_bits_data_4_entries_perms_4_g),
    .io_wreq_bits_data_4_entries_perms_4_u(l3_io_wreq_bits_data_4_entries_perms_4_u),
    .io_wreq_bits_data_4_entries_perms_4_x(l3_io_wreq_bits_data_4_entries_perms_4_x),
    .io_wreq_bits_data_4_entries_perms_4_w(l3_io_wreq_bits_data_4_entries_perms_4_w),
    .io_wreq_bits_data_4_entries_perms_4_r(l3_io_wreq_bits_data_4_entries_perms_4_r),
    .io_wreq_bits_data_4_entries_perms_5_d(l3_io_wreq_bits_data_4_entries_perms_5_d),
    .io_wreq_bits_data_4_entries_perms_5_a(l3_io_wreq_bits_data_4_entries_perms_5_a),
    .io_wreq_bits_data_4_entries_perms_5_g(l3_io_wreq_bits_data_4_entries_perms_5_g),
    .io_wreq_bits_data_4_entries_perms_5_u(l3_io_wreq_bits_data_4_entries_perms_5_u),
    .io_wreq_bits_data_4_entries_perms_5_x(l3_io_wreq_bits_data_4_entries_perms_5_x),
    .io_wreq_bits_data_4_entries_perms_5_w(l3_io_wreq_bits_data_4_entries_perms_5_w),
    .io_wreq_bits_data_4_entries_perms_5_r(l3_io_wreq_bits_data_4_entries_perms_5_r),
    .io_wreq_bits_data_4_entries_perms_6_d(l3_io_wreq_bits_data_4_entries_perms_6_d),
    .io_wreq_bits_data_4_entries_perms_6_a(l3_io_wreq_bits_data_4_entries_perms_6_a),
    .io_wreq_bits_data_4_entries_perms_6_g(l3_io_wreq_bits_data_4_entries_perms_6_g),
    .io_wreq_bits_data_4_entries_perms_6_u(l3_io_wreq_bits_data_4_entries_perms_6_u),
    .io_wreq_bits_data_4_entries_perms_6_x(l3_io_wreq_bits_data_4_entries_perms_6_x),
    .io_wreq_bits_data_4_entries_perms_6_w(l3_io_wreq_bits_data_4_entries_perms_6_w),
    .io_wreq_bits_data_4_entries_perms_6_r(l3_io_wreq_bits_data_4_entries_perms_6_r),
    .io_wreq_bits_data_4_entries_perms_7_d(l3_io_wreq_bits_data_4_entries_perms_7_d),
    .io_wreq_bits_data_4_entries_perms_7_a(l3_io_wreq_bits_data_4_entries_perms_7_a),
    .io_wreq_bits_data_4_entries_perms_7_g(l3_io_wreq_bits_data_4_entries_perms_7_g),
    .io_wreq_bits_data_4_entries_perms_7_u(l3_io_wreq_bits_data_4_entries_perms_7_u),
    .io_wreq_bits_data_4_entries_perms_7_x(l3_io_wreq_bits_data_4_entries_perms_7_x),
    .io_wreq_bits_data_4_entries_perms_7_w(l3_io_wreq_bits_data_4_entries_perms_7_w),
    .io_wreq_bits_data_4_entries_perms_7_r(l3_io_wreq_bits_data_4_entries_perms_7_r),
    .io_wreq_bits_data_4_entries_prefetch(l3_io_wreq_bits_data_4_entries_prefetch),
    .io_wreq_bits_data_4_ecc(l3_io_wreq_bits_data_4_ecc),
    .io_wreq_bits_data_5_entries_tag(l3_io_wreq_bits_data_5_entries_tag),
    .io_wreq_bits_data_5_entries_asid(l3_io_wreq_bits_data_5_entries_asid),
    .io_wreq_bits_data_5_entries_ppns_0(l3_io_wreq_bits_data_5_entries_ppns_0),
    .io_wreq_bits_data_5_entries_ppns_1(l3_io_wreq_bits_data_5_entries_ppns_1),
    .io_wreq_bits_data_5_entries_ppns_2(l3_io_wreq_bits_data_5_entries_ppns_2),
    .io_wreq_bits_data_5_entries_ppns_3(l3_io_wreq_bits_data_5_entries_ppns_3),
    .io_wreq_bits_data_5_entries_ppns_4(l3_io_wreq_bits_data_5_entries_ppns_4),
    .io_wreq_bits_data_5_entries_ppns_5(l3_io_wreq_bits_data_5_entries_ppns_5),
    .io_wreq_bits_data_5_entries_ppns_6(l3_io_wreq_bits_data_5_entries_ppns_6),
    .io_wreq_bits_data_5_entries_ppns_7(l3_io_wreq_bits_data_5_entries_ppns_7),
    .io_wreq_bits_data_5_entries_vs_0(l3_io_wreq_bits_data_5_entries_vs_0),
    .io_wreq_bits_data_5_entries_vs_1(l3_io_wreq_bits_data_5_entries_vs_1),
    .io_wreq_bits_data_5_entries_vs_2(l3_io_wreq_bits_data_5_entries_vs_2),
    .io_wreq_bits_data_5_entries_vs_3(l3_io_wreq_bits_data_5_entries_vs_3),
    .io_wreq_bits_data_5_entries_vs_4(l3_io_wreq_bits_data_5_entries_vs_4),
    .io_wreq_bits_data_5_entries_vs_5(l3_io_wreq_bits_data_5_entries_vs_5),
    .io_wreq_bits_data_5_entries_vs_6(l3_io_wreq_bits_data_5_entries_vs_6),
    .io_wreq_bits_data_5_entries_vs_7(l3_io_wreq_bits_data_5_entries_vs_7),
    .io_wreq_bits_data_5_entries_perms_0_d(l3_io_wreq_bits_data_5_entries_perms_0_d),
    .io_wreq_bits_data_5_entries_perms_0_a(l3_io_wreq_bits_data_5_entries_perms_0_a),
    .io_wreq_bits_data_5_entries_perms_0_g(l3_io_wreq_bits_data_5_entries_perms_0_g),
    .io_wreq_bits_data_5_entries_perms_0_u(l3_io_wreq_bits_data_5_entries_perms_0_u),
    .io_wreq_bits_data_5_entries_perms_0_x(l3_io_wreq_bits_data_5_entries_perms_0_x),
    .io_wreq_bits_data_5_entries_perms_0_w(l3_io_wreq_bits_data_5_entries_perms_0_w),
    .io_wreq_bits_data_5_entries_perms_0_r(l3_io_wreq_bits_data_5_entries_perms_0_r),
    .io_wreq_bits_data_5_entries_perms_1_d(l3_io_wreq_bits_data_5_entries_perms_1_d),
    .io_wreq_bits_data_5_entries_perms_1_a(l3_io_wreq_bits_data_5_entries_perms_1_a),
    .io_wreq_bits_data_5_entries_perms_1_g(l3_io_wreq_bits_data_5_entries_perms_1_g),
    .io_wreq_bits_data_5_entries_perms_1_u(l3_io_wreq_bits_data_5_entries_perms_1_u),
    .io_wreq_bits_data_5_entries_perms_1_x(l3_io_wreq_bits_data_5_entries_perms_1_x),
    .io_wreq_bits_data_5_entries_perms_1_w(l3_io_wreq_bits_data_5_entries_perms_1_w),
    .io_wreq_bits_data_5_entries_perms_1_r(l3_io_wreq_bits_data_5_entries_perms_1_r),
    .io_wreq_bits_data_5_entries_perms_2_d(l3_io_wreq_bits_data_5_entries_perms_2_d),
    .io_wreq_bits_data_5_entries_perms_2_a(l3_io_wreq_bits_data_5_entries_perms_2_a),
    .io_wreq_bits_data_5_entries_perms_2_g(l3_io_wreq_bits_data_5_entries_perms_2_g),
    .io_wreq_bits_data_5_entries_perms_2_u(l3_io_wreq_bits_data_5_entries_perms_2_u),
    .io_wreq_bits_data_5_entries_perms_2_x(l3_io_wreq_bits_data_5_entries_perms_2_x),
    .io_wreq_bits_data_5_entries_perms_2_w(l3_io_wreq_bits_data_5_entries_perms_2_w),
    .io_wreq_bits_data_5_entries_perms_2_r(l3_io_wreq_bits_data_5_entries_perms_2_r),
    .io_wreq_bits_data_5_entries_perms_3_d(l3_io_wreq_bits_data_5_entries_perms_3_d),
    .io_wreq_bits_data_5_entries_perms_3_a(l3_io_wreq_bits_data_5_entries_perms_3_a),
    .io_wreq_bits_data_5_entries_perms_3_g(l3_io_wreq_bits_data_5_entries_perms_3_g),
    .io_wreq_bits_data_5_entries_perms_3_u(l3_io_wreq_bits_data_5_entries_perms_3_u),
    .io_wreq_bits_data_5_entries_perms_3_x(l3_io_wreq_bits_data_5_entries_perms_3_x),
    .io_wreq_bits_data_5_entries_perms_3_w(l3_io_wreq_bits_data_5_entries_perms_3_w),
    .io_wreq_bits_data_5_entries_perms_3_r(l3_io_wreq_bits_data_5_entries_perms_3_r),
    .io_wreq_bits_data_5_entries_perms_4_d(l3_io_wreq_bits_data_5_entries_perms_4_d),
    .io_wreq_bits_data_5_entries_perms_4_a(l3_io_wreq_bits_data_5_entries_perms_4_a),
    .io_wreq_bits_data_5_entries_perms_4_g(l3_io_wreq_bits_data_5_entries_perms_4_g),
    .io_wreq_bits_data_5_entries_perms_4_u(l3_io_wreq_bits_data_5_entries_perms_4_u),
    .io_wreq_bits_data_5_entries_perms_4_x(l3_io_wreq_bits_data_5_entries_perms_4_x),
    .io_wreq_bits_data_5_entries_perms_4_w(l3_io_wreq_bits_data_5_entries_perms_4_w),
    .io_wreq_bits_data_5_entries_perms_4_r(l3_io_wreq_bits_data_5_entries_perms_4_r),
    .io_wreq_bits_data_5_entries_perms_5_d(l3_io_wreq_bits_data_5_entries_perms_5_d),
    .io_wreq_bits_data_5_entries_perms_5_a(l3_io_wreq_bits_data_5_entries_perms_5_a),
    .io_wreq_bits_data_5_entries_perms_5_g(l3_io_wreq_bits_data_5_entries_perms_5_g),
    .io_wreq_bits_data_5_entries_perms_5_u(l3_io_wreq_bits_data_5_entries_perms_5_u),
    .io_wreq_bits_data_5_entries_perms_5_x(l3_io_wreq_bits_data_5_entries_perms_5_x),
    .io_wreq_bits_data_5_entries_perms_5_w(l3_io_wreq_bits_data_5_entries_perms_5_w),
    .io_wreq_bits_data_5_entries_perms_5_r(l3_io_wreq_bits_data_5_entries_perms_5_r),
    .io_wreq_bits_data_5_entries_perms_6_d(l3_io_wreq_bits_data_5_entries_perms_6_d),
    .io_wreq_bits_data_5_entries_perms_6_a(l3_io_wreq_bits_data_5_entries_perms_6_a),
    .io_wreq_bits_data_5_entries_perms_6_g(l3_io_wreq_bits_data_5_entries_perms_6_g),
    .io_wreq_bits_data_5_entries_perms_6_u(l3_io_wreq_bits_data_5_entries_perms_6_u),
    .io_wreq_bits_data_5_entries_perms_6_x(l3_io_wreq_bits_data_5_entries_perms_6_x),
    .io_wreq_bits_data_5_entries_perms_6_w(l3_io_wreq_bits_data_5_entries_perms_6_w),
    .io_wreq_bits_data_5_entries_perms_6_r(l3_io_wreq_bits_data_5_entries_perms_6_r),
    .io_wreq_bits_data_5_entries_perms_7_d(l3_io_wreq_bits_data_5_entries_perms_7_d),
    .io_wreq_bits_data_5_entries_perms_7_a(l3_io_wreq_bits_data_5_entries_perms_7_a),
    .io_wreq_bits_data_5_entries_perms_7_g(l3_io_wreq_bits_data_5_entries_perms_7_g),
    .io_wreq_bits_data_5_entries_perms_7_u(l3_io_wreq_bits_data_5_entries_perms_7_u),
    .io_wreq_bits_data_5_entries_perms_7_x(l3_io_wreq_bits_data_5_entries_perms_7_x),
    .io_wreq_bits_data_5_entries_perms_7_w(l3_io_wreq_bits_data_5_entries_perms_7_w),
    .io_wreq_bits_data_5_entries_perms_7_r(l3_io_wreq_bits_data_5_entries_perms_7_r),
    .io_wreq_bits_data_5_entries_prefetch(l3_io_wreq_bits_data_5_entries_prefetch),
    .io_wreq_bits_data_5_ecc(l3_io_wreq_bits_data_5_ecc),
    .io_wreq_bits_data_6_entries_tag(l3_io_wreq_bits_data_6_entries_tag),
    .io_wreq_bits_data_6_entries_asid(l3_io_wreq_bits_data_6_entries_asid),
    .io_wreq_bits_data_6_entries_ppns_0(l3_io_wreq_bits_data_6_entries_ppns_0),
    .io_wreq_bits_data_6_entries_ppns_1(l3_io_wreq_bits_data_6_entries_ppns_1),
    .io_wreq_bits_data_6_entries_ppns_2(l3_io_wreq_bits_data_6_entries_ppns_2),
    .io_wreq_bits_data_6_entries_ppns_3(l3_io_wreq_bits_data_6_entries_ppns_3),
    .io_wreq_bits_data_6_entries_ppns_4(l3_io_wreq_bits_data_6_entries_ppns_4),
    .io_wreq_bits_data_6_entries_ppns_5(l3_io_wreq_bits_data_6_entries_ppns_5),
    .io_wreq_bits_data_6_entries_ppns_6(l3_io_wreq_bits_data_6_entries_ppns_6),
    .io_wreq_bits_data_6_entries_ppns_7(l3_io_wreq_bits_data_6_entries_ppns_7),
    .io_wreq_bits_data_6_entries_vs_0(l3_io_wreq_bits_data_6_entries_vs_0),
    .io_wreq_bits_data_6_entries_vs_1(l3_io_wreq_bits_data_6_entries_vs_1),
    .io_wreq_bits_data_6_entries_vs_2(l3_io_wreq_bits_data_6_entries_vs_2),
    .io_wreq_bits_data_6_entries_vs_3(l3_io_wreq_bits_data_6_entries_vs_3),
    .io_wreq_bits_data_6_entries_vs_4(l3_io_wreq_bits_data_6_entries_vs_4),
    .io_wreq_bits_data_6_entries_vs_5(l3_io_wreq_bits_data_6_entries_vs_5),
    .io_wreq_bits_data_6_entries_vs_6(l3_io_wreq_bits_data_6_entries_vs_6),
    .io_wreq_bits_data_6_entries_vs_7(l3_io_wreq_bits_data_6_entries_vs_7),
    .io_wreq_bits_data_6_entries_perms_0_d(l3_io_wreq_bits_data_6_entries_perms_0_d),
    .io_wreq_bits_data_6_entries_perms_0_a(l3_io_wreq_bits_data_6_entries_perms_0_a),
    .io_wreq_bits_data_6_entries_perms_0_g(l3_io_wreq_bits_data_6_entries_perms_0_g),
    .io_wreq_bits_data_6_entries_perms_0_u(l3_io_wreq_bits_data_6_entries_perms_0_u),
    .io_wreq_bits_data_6_entries_perms_0_x(l3_io_wreq_bits_data_6_entries_perms_0_x),
    .io_wreq_bits_data_6_entries_perms_0_w(l3_io_wreq_bits_data_6_entries_perms_0_w),
    .io_wreq_bits_data_6_entries_perms_0_r(l3_io_wreq_bits_data_6_entries_perms_0_r),
    .io_wreq_bits_data_6_entries_perms_1_d(l3_io_wreq_bits_data_6_entries_perms_1_d),
    .io_wreq_bits_data_6_entries_perms_1_a(l3_io_wreq_bits_data_6_entries_perms_1_a),
    .io_wreq_bits_data_6_entries_perms_1_g(l3_io_wreq_bits_data_6_entries_perms_1_g),
    .io_wreq_bits_data_6_entries_perms_1_u(l3_io_wreq_bits_data_6_entries_perms_1_u),
    .io_wreq_bits_data_6_entries_perms_1_x(l3_io_wreq_bits_data_6_entries_perms_1_x),
    .io_wreq_bits_data_6_entries_perms_1_w(l3_io_wreq_bits_data_6_entries_perms_1_w),
    .io_wreq_bits_data_6_entries_perms_1_r(l3_io_wreq_bits_data_6_entries_perms_1_r),
    .io_wreq_bits_data_6_entries_perms_2_d(l3_io_wreq_bits_data_6_entries_perms_2_d),
    .io_wreq_bits_data_6_entries_perms_2_a(l3_io_wreq_bits_data_6_entries_perms_2_a),
    .io_wreq_bits_data_6_entries_perms_2_g(l3_io_wreq_bits_data_6_entries_perms_2_g),
    .io_wreq_bits_data_6_entries_perms_2_u(l3_io_wreq_bits_data_6_entries_perms_2_u),
    .io_wreq_bits_data_6_entries_perms_2_x(l3_io_wreq_bits_data_6_entries_perms_2_x),
    .io_wreq_bits_data_6_entries_perms_2_w(l3_io_wreq_bits_data_6_entries_perms_2_w),
    .io_wreq_bits_data_6_entries_perms_2_r(l3_io_wreq_bits_data_6_entries_perms_2_r),
    .io_wreq_bits_data_6_entries_perms_3_d(l3_io_wreq_bits_data_6_entries_perms_3_d),
    .io_wreq_bits_data_6_entries_perms_3_a(l3_io_wreq_bits_data_6_entries_perms_3_a),
    .io_wreq_bits_data_6_entries_perms_3_g(l3_io_wreq_bits_data_6_entries_perms_3_g),
    .io_wreq_bits_data_6_entries_perms_3_u(l3_io_wreq_bits_data_6_entries_perms_3_u),
    .io_wreq_bits_data_6_entries_perms_3_x(l3_io_wreq_bits_data_6_entries_perms_3_x),
    .io_wreq_bits_data_6_entries_perms_3_w(l3_io_wreq_bits_data_6_entries_perms_3_w),
    .io_wreq_bits_data_6_entries_perms_3_r(l3_io_wreq_bits_data_6_entries_perms_3_r),
    .io_wreq_bits_data_6_entries_perms_4_d(l3_io_wreq_bits_data_6_entries_perms_4_d),
    .io_wreq_bits_data_6_entries_perms_4_a(l3_io_wreq_bits_data_6_entries_perms_4_a),
    .io_wreq_bits_data_6_entries_perms_4_g(l3_io_wreq_bits_data_6_entries_perms_4_g),
    .io_wreq_bits_data_6_entries_perms_4_u(l3_io_wreq_bits_data_6_entries_perms_4_u),
    .io_wreq_bits_data_6_entries_perms_4_x(l3_io_wreq_bits_data_6_entries_perms_4_x),
    .io_wreq_bits_data_6_entries_perms_4_w(l3_io_wreq_bits_data_6_entries_perms_4_w),
    .io_wreq_bits_data_6_entries_perms_4_r(l3_io_wreq_bits_data_6_entries_perms_4_r),
    .io_wreq_bits_data_6_entries_perms_5_d(l3_io_wreq_bits_data_6_entries_perms_5_d),
    .io_wreq_bits_data_6_entries_perms_5_a(l3_io_wreq_bits_data_6_entries_perms_5_a),
    .io_wreq_bits_data_6_entries_perms_5_g(l3_io_wreq_bits_data_6_entries_perms_5_g),
    .io_wreq_bits_data_6_entries_perms_5_u(l3_io_wreq_bits_data_6_entries_perms_5_u),
    .io_wreq_bits_data_6_entries_perms_5_x(l3_io_wreq_bits_data_6_entries_perms_5_x),
    .io_wreq_bits_data_6_entries_perms_5_w(l3_io_wreq_bits_data_6_entries_perms_5_w),
    .io_wreq_bits_data_6_entries_perms_5_r(l3_io_wreq_bits_data_6_entries_perms_5_r),
    .io_wreq_bits_data_6_entries_perms_6_d(l3_io_wreq_bits_data_6_entries_perms_6_d),
    .io_wreq_bits_data_6_entries_perms_6_a(l3_io_wreq_bits_data_6_entries_perms_6_a),
    .io_wreq_bits_data_6_entries_perms_6_g(l3_io_wreq_bits_data_6_entries_perms_6_g),
    .io_wreq_bits_data_6_entries_perms_6_u(l3_io_wreq_bits_data_6_entries_perms_6_u),
    .io_wreq_bits_data_6_entries_perms_6_x(l3_io_wreq_bits_data_6_entries_perms_6_x),
    .io_wreq_bits_data_6_entries_perms_6_w(l3_io_wreq_bits_data_6_entries_perms_6_w),
    .io_wreq_bits_data_6_entries_perms_6_r(l3_io_wreq_bits_data_6_entries_perms_6_r),
    .io_wreq_bits_data_6_entries_perms_7_d(l3_io_wreq_bits_data_6_entries_perms_7_d),
    .io_wreq_bits_data_6_entries_perms_7_a(l3_io_wreq_bits_data_6_entries_perms_7_a),
    .io_wreq_bits_data_6_entries_perms_7_g(l3_io_wreq_bits_data_6_entries_perms_7_g),
    .io_wreq_bits_data_6_entries_perms_7_u(l3_io_wreq_bits_data_6_entries_perms_7_u),
    .io_wreq_bits_data_6_entries_perms_7_x(l3_io_wreq_bits_data_6_entries_perms_7_x),
    .io_wreq_bits_data_6_entries_perms_7_w(l3_io_wreq_bits_data_6_entries_perms_7_w),
    .io_wreq_bits_data_6_entries_perms_7_r(l3_io_wreq_bits_data_6_entries_perms_7_r),
    .io_wreq_bits_data_6_entries_prefetch(l3_io_wreq_bits_data_6_entries_prefetch),
    .io_wreq_bits_data_6_ecc(l3_io_wreq_bits_data_6_ecc),
    .io_wreq_bits_data_7_entries_tag(l3_io_wreq_bits_data_7_entries_tag),
    .io_wreq_bits_data_7_entries_asid(l3_io_wreq_bits_data_7_entries_asid),
    .io_wreq_bits_data_7_entries_ppns_0(l3_io_wreq_bits_data_7_entries_ppns_0),
    .io_wreq_bits_data_7_entries_ppns_1(l3_io_wreq_bits_data_7_entries_ppns_1),
    .io_wreq_bits_data_7_entries_ppns_2(l3_io_wreq_bits_data_7_entries_ppns_2),
    .io_wreq_bits_data_7_entries_ppns_3(l3_io_wreq_bits_data_7_entries_ppns_3),
    .io_wreq_bits_data_7_entries_ppns_4(l3_io_wreq_bits_data_7_entries_ppns_4),
    .io_wreq_bits_data_7_entries_ppns_5(l3_io_wreq_bits_data_7_entries_ppns_5),
    .io_wreq_bits_data_7_entries_ppns_6(l3_io_wreq_bits_data_7_entries_ppns_6),
    .io_wreq_bits_data_7_entries_ppns_7(l3_io_wreq_bits_data_7_entries_ppns_7),
    .io_wreq_bits_data_7_entries_vs_0(l3_io_wreq_bits_data_7_entries_vs_0),
    .io_wreq_bits_data_7_entries_vs_1(l3_io_wreq_bits_data_7_entries_vs_1),
    .io_wreq_bits_data_7_entries_vs_2(l3_io_wreq_bits_data_7_entries_vs_2),
    .io_wreq_bits_data_7_entries_vs_3(l3_io_wreq_bits_data_7_entries_vs_3),
    .io_wreq_bits_data_7_entries_vs_4(l3_io_wreq_bits_data_7_entries_vs_4),
    .io_wreq_bits_data_7_entries_vs_5(l3_io_wreq_bits_data_7_entries_vs_5),
    .io_wreq_bits_data_7_entries_vs_6(l3_io_wreq_bits_data_7_entries_vs_6),
    .io_wreq_bits_data_7_entries_vs_7(l3_io_wreq_bits_data_7_entries_vs_7),
    .io_wreq_bits_data_7_entries_perms_0_d(l3_io_wreq_bits_data_7_entries_perms_0_d),
    .io_wreq_bits_data_7_entries_perms_0_a(l3_io_wreq_bits_data_7_entries_perms_0_a),
    .io_wreq_bits_data_7_entries_perms_0_g(l3_io_wreq_bits_data_7_entries_perms_0_g),
    .io_wreq_bits_data_7_entries_perms_0_u(l3_io_wreq_bits_data_7_entries_perms_0_u),
    .io_wreq_bits_data_7_entries_perms_0_x(l3_io_wreq_bits_data_7_entries_perms_0_x),
    .io_wreq_bits_data_7_entries_perms_0_w(l3_io_wreq_bits_data_7_entries_perms_0_w),
    .io_wreq_bits_data_7_entries_perms_0_r(l3_io_wreq_bits_data_7_entries_perms_0_r),
    .io_wreq_bits_data_7_entries_perms_1_d(l3_io_wreq_bits_data_7_entries_perms_1_d),
    .io_wreq_bits_data_7_entries_perms_1_a(l3_io_wreq_bits_data_7_entries_perms_1_a),
    .io_wreq_bits_data_7_entries_perms_1_g(l3_io_wreq_bits_data_7_entries_perms_1_g),
    .io_wreq_bits_data_7_entries_perms_1_u(l3_io_wreq_bits_data_7_entries_perms_1_u),
    .io_wreq_bits_data_7_entries_perms_1_x(l3_io_wreq_bits_data_7_entries_perms_1_x),
    .io_wreq_bits_data_7_entries_perms_1_w(l3_io_wreq_bits_data_7_entries_perms_1_w),
    .io_wreq_bits_data_7_entries_perms_1_r(l3_io_wreq_bits_data_7_entries_perms_1_r),
    .io_wreq_bits_data_7_entries_perms_2_d(l3_io_wreq_bits_data_7_entries_perms_2_d),
    .io_wreq_bits_data_7_entries_perms_2_a(l3_io_wreq_bits_data_7_entries_perms_2_a),
    .io_wreq_bits_data_7_entries_perms_2_g(l3_io_wreq_bits_data_7_entries_perms_2_g),
    .io_wreq_bits_data_7_entries_perms_2_u(l3_io_wreq_bits_data_7_entries_perms_2_u),
    .io_wreq_bits_data_7_entries_perms_2_x(l3_io_wreq_bits_data_7_entries_perms_2_x),
    .io_wreq_bits_data_7_entries_perms_2_w(l3_io_wreq_bits_data_7_entries_perms_2_w),
    .io_wreq_bits_data_7_entries_perms_2_r(l3_io_wreq_bits_data_7_entries_perms_2_r),
    .io_wreq_bits_data_7_entries_perms_3_d(l3_io_wreq_bits_data_7_entries_perms_3_d),
    .io_wreq_bits_data_7_entries_perms_3_a(l3_io_wreq_bits_data_7_entries_perms_3_a),
    .io_wreq_bits_data_7_entries_perms_3_g(l3_io_wreq_bits_data_7_entries_perms_3_g),
    .io_wreq_bits_data_7_entries_perms_3_u(l3_io_wreq_bits_data_7_entries_perms_3_u),
    .io_wreq_bits_data_7_entries_perms_3_x(l3_io_wreq_bits_data_7_entries_perms_3_x),
    .io_wreq_bits_data_7_entries_perms_3_w(l3_io_wreq_bits_data_7_entries_perms_3_w),
    .io_wreq_bits_data_7_entries_perms_3_r(l3_io_wreq_bits_data_7_entries_perms_3_r),
    .io_wreq_bits_data_7_entries_perms_4_d(l3_io_wreq_bits_data_7_entries_perms_4_d),
    .io_wreq_bits_data_7_entries_perms_4_a(l3_io_wreq_bits_data_7_entries_perms_4_a),
    .io_wreq_bits_data_7_entries_perms_4_g(l3_io_wreq_bits_data_7_entries_perms_4_g),
    .io_wreq_bits_data_7_entries_perms_4_u(l3_io_wreq_bits_data_7_entries_perms_4_u),
    .io_wreq_bits_data_7_entries_perms_4_x(l3_io_wreq_bits_data_7_entries_perms_4_x),
    .io_wreq_bits_data_7_entries_perms_4_w(l3_io_wreq_bits_data_7_entries_perms_4_w),
    .io_wreq_bits_data_7_entries_perms_4_r(l3_io_wreq_bits_data_7_entries_perms_4_r),
    .io_wreq_bits_data_7_entries_perms_5_d(l3_io_wreq_bits_data_7_entries_perms_5_d),
    .io_wreq_bits_data_7_entries_perms_5_a(l3_io_wreq_bits_data_7_entries_perms_5_a),
    .io_wreq_bits_data_7_entries_perms_5_g(l3_io_wreq_bits_data_7_entries_perms_5_g),
    .io_wreq_bits_data_7_entries_perms_5_u(l3_io_wreq_bits_data_7_entries_perms_5_u),
    .io_wreq_bits_data_7_entries_perms_5_x(l3_io_wreq_bits_data_7_entries_perms_5_x),
    .io_wreq_bits_data_7_entries_perms_5_w(l3_io_wreq_bits_data_7_entries_perms_5_w),
    .io_wreq_bits_data_7_entries_perms_5_r(l3_io_wreq_bits_data_7_entries_perms_5_r),
    .io_wreq_bits_data_7_entries_perms_6_d(l3_io_wreq_bits_data_7_entries_perms_6_d),
    .io_wreq_bits_data_7_entries_perms_6_a(l3_io_wreq_bits_data_7_entries_perms_6_a),
    .io_wreq_bits_data_7_entries_perms_6_g(l3_io_wreq_bits_data_7_entries_perms_6_g),
    .io_wreq_bits_data_7_entries_perms_6_u(l3_io_wreq_bits_data_7_entries_perms_6_u),
    .io_wreq_bits_data_7_entries_perms_6_x(l3_io_wreq_bits_data_7_entries_perms_6_x),
    .io_wreq_bits_data_7_entries_perms_6_w(l3_io_wreq_bits_data_7_entries_perms_6_w),
    .io_wreq_bits_data_7_entries_perms_6_r(l3_io_wreq_bits_data_7_entries_perms_6_r),
    .io_wreq_bits_data_7_entries_perms_7_d(l3_io_wreq_bits_data_7_entries_perms_7_d),
    .io_wreq_bits_data_7_entries_perms_7_a(l3_io_wreq_bits_data_7_entries_perms_7_a),
    .io_wreq_bits_data_7_entries_perms_7_g(l3_io_wreq_bits_data_7_entries_perms_7_g),
    .io_wreq_bits_data_7_entries_perms_7_u(l3_io_wreq_bits_data_7_entries_perms_7_u),
    .io_wreq_bits_data_7_entries_perms_7_x(l3_io_wreq_bits_data_7_entries_perms_7_x),
    .io_wreq_bits_data_7_entries_perms_7_w(l3_io_wreq_bits_data_7_entries_perms_7_w),
    .io_wreq_bits_data_7_entries_perms_7_r(l3_io_wreq_bits_data_7_entries_perms_7_r),
    .io_wreq_bits_data_7_entries_prefetch(l3_io_wreq_bits_data_7_entries_prefetch),
    .io_wreq_bits_data_7_ecc(l3_io_wreq_bits_data_7_ecc),
    .io_wreq_bits_waymask(l3_io_wreq_bits_waymask)
  );
  assign io_req_ready = stageDelay_0_ready & ~io_refill_valid; // @[PipelineConnect.scala 114:31]
  assign io_resp_valid = valid_2; // @[PageTableCache.scala 133:23 PipelineConnect.scala 117:17]
  assign io_resp_bits_req_info_vpn = data_2_req_info_vpn; // @[PageTableCache.scala 133:23 PipelineConnect.scala 116:16]
  assign io_resp_bits_req_info_source = data_2_req_info_source; // @[PageTableCache.scala 133:23 PipelineConnect.scala 116:16]
  assign io_resp_bits_isFirst = data_2_isFirst; // @[PageTableCache.scala 133:23 PipelineConnect.scala 116:16]
  assign io_resp_bits_hit = resp_res_l3_hit | resp_res_sp_hit; // @[PageTableCache.scala 396:44]
  assign io_resp_bits_prefetch = resp_res_l3_pre & resp_res_l3_hit | resp_res_sp_pre & resp_res_sp_hit; // @[PageTableCache.scala 398:63]
  assign io_resp_bits_bypassed = bypassed_2 | bypassed_1 & ~resp_res_l2_hit | bypassed_0 & ~resp_res_l1_hit; // @[PageTableCache.scala 397:77]
  assign io_resp_bits_toFsm_l1Hit = resp_res_l1_hit; // @[PageTableCache.scala 399:28]
  assign io_resp_bits_toFsm_l2Hit = resp_res_l2_hit; // @[PageTableCache.scala 400:28]
  assign io_resp_bits_toFsm_ppn = resp_res_l2_hit ? resp_res_l2_ppn : resp_res_l1_ppn; // @[PageTableCache.scala 401:34]
  assign io_resp_bits_toTlb_tag = data_2_req_info_vpn; // @[PageTableCache.scala 133:23 PipelineConnect.scala 116:16]
  assign io_resp_bits_toTlb_asid = io_csr_dup_0_satp_asid; // @[PageTableCache.scala 403:28]
  assign io_resp_bits_toTlb_ppn = resp_res_l3_hit ? resp_res_l3_ppn : resp_res_sp_ppn; // @[PageTableCache.scala 404:34]
  assign io_resp_bits_toTlb_perm_d = resp_res_l3_hit ? resp_res_l3_perm_d : resp_res_sp_perm_d; // @[PageTableCache.scala 405:39]
  assign io_resp_bits_toTlb_perm_a = resp_res_l3_hit ? resp_res_l3_perm_a : resp_res_sp_perm_a; // @[PageTableCache.scala 405:39]
  assign io_resp_bits_toTlb_perm_g = resp_res_l3_hit ? resp_res_l3_perm_g : resp_res_sp_perm_g; // @[PageTableCache.scala 405:39]
  assign io_resp_bits_toTlb_perm_u = resp_res_l3_hit ? resp_res_l3_perm_u : resp_res_sp_perm_u; // @[PageTableCache.scala 405:39]
  assign io_resp_bits_toTlb_perm_x = resp_res_l3_hit ? resp_res_l3_perm_x : resp_res_sp_perm_x; // @[PageTableCache.scala 405:39]
  assign io_resp_bits_toTlb_perm_w = resp_res_l3_hit ? resp_res_l3_perm_w : resp_res_sp_perm_w; // @[PageTableCache.scala 405:39]
  assign io_resp_bits_toTlb_perm_r = resp_res_l3_hit ? resp_res_l3_perm_r : resp_res_sp_perm_r; // @[PageTableCache.scala 405:39]
  assign io_resp_bits_toTlb_level = resp_res_l3_hit ? 2'h2 : resp_res_sp_level; // @[PageTableCache.scala 406:40]
  assign io_resp_bits_toTlb_prefetch = data_2_req_info_source == 2'h2; // @[MMUConst.scala 254:13]
  assign io_resp_bits_toTlb_v = resp_res_sp_hit ? resp_res_sp_v : resp_res_l3_v; // @[PageTableCache.scala 408:30]
  assign io_perf_0_value = {{5'd0}, io_perf_0_value_REG_1}; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_1_value = {{5'd0}, io_perf_1_value_REG_1}; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_2_value = {{5'd0}, io_perf_2_value_REG_1}; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_3_value = {{5'd0}, io_perf_3_value_REG_1}; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_4_value = {{5'd0}, io_perf_4_value_REG_1}; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_5_value = {{5'd0}, io_perf_5_value_REG_1}; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_6_value = {{5'd0}, io_perf_6_value_REG_1}; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_7_value = {{5'd0}, io_perf_7_value_REG_1}; // @[PerfCounterUtils.scala 188:17]
  assign l2_clock = clock;
  assign l2_io_rreq_valid = stageReq_ready & io_req_valid; // @[Decoupled.scala 50:35]
  assign l2_io_rreq_bits_setIdx = io_req_bits_req_info_vpn[13:12]; // @[MMUConst.scala 210:21]
  assign l2_io_wreq_valid = ~flush_dup_1 & io_refill_bits_levelOH_l2 & ~_T_336 & ~_T_358 & ~_T_362; // @[PageTableCache.scala 462:107]
  assign l2_io_wreq_bits_setIdx = io_refill_bits_req_info_dup_1_vpn[13:12]; // @[MMUConst.scala 210:21]
  assign l2_io_wreq_bits_data_0_entries_tag = io_refill_bits_req_info_dup_1_vpn[26:14]; // @[MMUBundle.scala 646:8]
  assign l2_io_wreq_bits_data_0_entries_asid = io_csr_dup_1_satp_asid; // @[MMUBundle.scala 662:18 664:13]
  assign l2_io_wreq_bits_data_0_entries_ppns_0 = io_refill_bits_ptes[33:10]; // @[MMUBundle.scala 667:52]
  assign l2_io_wreq_bits_data_0_entries_ppns_1 = io_refill_bits_ptes[97:74]; // @[MMUBundle.scala 667:52]
  assign l2_io_wreq_bits_data_0_entries_ppns_2 = io_refill_bits_ptes[161:138]; // @[MMUBundle.scala 667:52]
  assign l2_io_wreq_bits_data_0_entries_ppns_3 = io_refill_bits_ptes[225:202]; // @[MMUBundle.scala 667:52]
  assign l2_io_wreq_bits_data_0_entries_ppns_4 = io_refill_bits_ptes[289:266]; // @[MMUBundle.scala 667:52]
  assign l2_io_wreq_bits_data_0_entries_ppns_5 = io_refill_bits_ptes[353:330]; // @[MMUBundle.scala 667:52]
  assign l2_io_wreq_bits_data_0_entries_ppns_6 = io_refill_bits_ptes[417:394]; // @[MMUBundle.scala 667:52]
  assign l2_io_wreq_bits_data_0_entries_ppns_7 = io_refill_bits_ptes[481:458]; // @[MMUBundle.scala 667:52]
  assign l2_io_wreq_bits_data_0_entries_vs_0 = ~_wdata_entries_ps_vs_0_T_19 & ~_wdata_entries_ps_vs_0_T_5; // @[MMUBundle.scala 669:42]
  assign l2_io_wreq_bits_data_0_entries_vs_1 = ~_wdata_entries_ps_vs_1_T_19 & ~_wdata_entries_ps_vs_1_T_5; // @[MMUBundle.scala 669:42]
  assign l2_io_wreq_bits_data_0_entries_vs_2 = ~_wdata_entries_ps_vs_2_T_19 & ~_wdata_entries_ps_vs_2_T_5; // @[MMUBundle.scala 669:42]
  assign l2_io_wreq_bits_data_0_entries_vs_3 = ~_wdata_entries_ps_vs_3_T_19 & ~_wdata_entries_ps_vs_3_T_5; // @[MMUBundle.scala 669:42]
  assign l2_io_wreq_bits_data_0_entries_vs_4 = ~_wdata_entries_ps_vs_4_T_19 & ~_wdata_entries_ps_vs_4_T_5; // @[MMUBundle.scala 669:42]
  assign l2_io_wreq_bits_data_0_entries_vs_5 = ~_wdata_entries_ps_vs_5_T_19 & ~_wdata_entries_ps_vs_5_T_5; // @[MMUBundle.scala 669:42]
  assign l2_io_wreq_bits_data_0_entries_vs_6 = ~_wdata_entries_ps_vs_6_T_19 & ~_wdata_entries_ps_vs_6_T_5; // @[MMUBundle.scala 669:42]
  assign l2_io_wreq_bits_data_0_entries_vs_7 = ~_wdata_entries_ps_vs_7_T_19 & ~_wdata_entries_ps_vs_7_T_5; // @[MMUBundle.scala 669:42]
  assign l2_io_wreq_bits_data_0_entries_prefetch = io_refill_bits_req_info_dup_1_source == 2'h2; // @[MMUConst.scala 254:13]
  assign l2_io_wreq_bits_data_0_ecc = {ecc_unaligned,_wdata_ecc_T}; // @[Cat.scala 31:58]
  assign l2_io_wreq_bits_data_1_entries_tag = io_refill_bits_req_info_dup_1_vpn[26:14]; // @[MMUBundle.scala 646:8]
  assign l2_io_wreq_bits_data_1_entries_asid = io_csr_dup_1_satp_asid; // @[MMUBundle.scala 662:18 664:13]
  assign l2_io_wreq_bits_data_1_entries_ppns_0 = io_refill_bits_ptes[33:10]; // @[MMUBundle.scala 667:52]
  assign l2_io_wreq_bits_data_1_entries_ppns_1 = io_refill_bits_ptes[97:74]; // @[MMUBundle.scala 667:52]
  assign l2_io_wreq_bits_data_1_entries_ppns_2 = io_refill_bits_ptes[161:138]; // @[MMUBundle.scala 667:52]
  assign l2_io_wreq_bits_data_1_entries_ppns_3 = io_refill_bits_ptes[225:202]; // @[MMUBundle.scala 667:52]
  assign l2_io_wreq_bits_data_1_entries_ppns_4 = io_refill_bits_ptes[289:266]; // @[MMUBundle.scala 667:52]
  assign l2_io_wreq_bits_data_1_entries_ppns_5 = io_refill_bits_ptes[353:330]; // @[MMUBundle.scala 667:52]
  assign l2_io_wreq_bits_data_1_entries_ppns_6 = io_refill_bits_ptes[417:394]; // @[MMUBundle.scala 667:52]
  assign l2_io_wreq_bits_data_1_entries_ppns_7 = io_refill_bits_ptes[481:458]; // @[MMUBundle.scala 667:52]
  assign l2_io_wreq_bits_data_1_entries_vs_0 = ~_wdata_entries_ps_vs_0_T_19 & ~_wdata_entries_ps_vs_0_T_5; // @[MMUBundle.scala 669:42]
  assign l2_io_wreq_bits_data_1_entries_vs_1 = ~_wdata_entries_ps_vs_1_T_19 & ~_wdata_entries_ps_vs_1_T_5; // @[MMUBundle.scala 669:42]
  assign l2_io_wreq_bits_data_1_entries_vs_2 = ~_wdata_entries_ps_vs_2_T_19 & ~_wdata_entries_ps_vs_2_T_5; // @[MMUBundle.scala 669:42]
  assign l2_io_wreq_bits_data_1_entries_vs_3 = ~_wdata_entries_ps_vs_3_T_19 & ~_wdata_entries_ps_vs_3_T_5; // @[MMUBundle.scala 669:42]
  assign l2_io_wreq_bits_data_1_entries_vs_4 = ~_wdata_entries_ps_vs_4_T_19 & ~_wdata_entries_ps_vs_4_T_5; // @[MMUBundle.scala 669:42]
  assign l2_io_wreq_bits_data_1_entries_vs_5 = ~_wdata_entries_ps_vs_5_T_19 & ~_wdata_entries_ps_vs_5_T_5; // @[MMUBundle.scala 669:42]
  assign l2_io_wreq_bits_data_1_entries_vs_6 = ~_wdata_entries_ps_vs_6_T_19 & ~_wdata_entries_ps_vs_6_T_5; // @[MMUBundle.scala 669:42]
  assign l2_io_wreq_bits_data_1_entries_vs_7 = ~_wdata_entries_ps_vs_7_T_19 & ~_wdata_entries_ps_vs_7_T_5; // @[MMUBundle.scala 669:42]
  assign l2_io_wreq_bits_data_1_entries_prefetch = io_refill_bits_req_info_dup_1_source == 2'h2; // @[MMUConst.scala 254:13]
  assign l2_io_wreq_bits_data_1_ecc = {ecc_unaligned,_wdata_ecc_T}; // @[Cat.scala 31:58]
  assign l2_io_wreq_bits_data_2_entries_tag = io_refill_bits_req_info_dup_1_vpn[26:14]; // @[MMUBundle.scala 646:8]
  assign l2_io_wreq_bits_data_2_entries_asid = io_csr_dup_1_satp_asid; // @[MMUBundle.scala 662:18 664:13]
  assign l2_io_wreq_bits_data_2_entries_ppns_0 = io_refill_bits_ptes[33:10]; // @[MMUBundle.scala 667:52]
  assign l2_io_wreq_bits_data_2_entries_ppns_1 = io_refill_bits_ptes[97:74]; // @[MMUBundle.scala 667:52]
  assign l2_io_wreq_bits_data_2_entries_ppns_2 = io_refill_bits_ptes[161:138]; // @[MMUBundle.scala 667:52]
  assign l2_io_wreq_bits_data_2_entries_ppns_3 = io_refill_bits_ptes[225:202]; // @[MMUBundle.scala 667:52]
  assign l2_io_wreq_bits_data_2_entries_ppns_4 = io_refill_bits_ptes[289:266]; // @[MMUBundle.scala 667:52]
  assign l2_io_wreq_bits_data_2_entries_ppns_5 = io_refill_bits_ptes[353:330]; // @[MMUBundle.scala 667:52]
  assign l2_io_wreq_bits_data_2_entries_ppns_6 = io_refill_bits_ptes[417:394]; // @[MMUBundle.scala 667:52]
  assign l2_io_wreq_bits_data_2_entries_ppns_7 = io_refill_bits_ptes[481:458]; // @[MMUBundle.scala 667:52]
  assign l2_io_wreq_bits_data_2_entries_vs_0 = ~_wdata_entries_ps_vs_0_T_19 & ~_wdata_entries_ps_vs_0_T_5; // @[MMUBundle.scala 669:42]
  assign l2_io_wreq_bits_data_2_entries_vs_1 = ~_wdata_entries_ps_vs_1_T_19 & ~_wdata_entries_ps_vs_1_T_5; // @[MMUBundle.scala 669:42]
  assign l2_io_wreq_bits_data_2_entries_vs_2 = ~_wdata_entries_ps_vs_2_T_19 & ~_wdata_entries_ps_vs_2_T_5; // @[MMUBundle.scala 669:42]
  assign l2_io_wreq_bits_data_2_entries_vs_3 = ~_wdata_entries_ps_vs_3_T_19 & ~_wdata_entries_ps_vs_3_T_5; // @[MMUBundle.scala 669:42]
  assign l2_io_wreq_bits_data_2_entries_vs_4 = ~_wdata_entries_ps_vs_4_T_19 & ~_wdata_entries_ps_vs_4_T_5; // @[MMUBundle.scala 669:42]
  assign l2_io_wreq_bits_data_2_entries_vs_5 = ~_wdata_entries_ps_vs_5_T_19 & ~_wdata_entries_ps_vs_5_T_5; // @[MMUBundle.scala 669:42]
  assign l2_io_wreq_bits_data_2_entries_vs_6 = ~_wdata_entries_ps_vs_6_T_19 & ~_wdata_entries_ps_vs_6_T_5; // @[MMUBundle.scala 669:42]
  assign l2_io_wreq_bits_data_2_entries_vs_7 = ~_wdata_entries_ps_vs_7_T_19 & ~_wdata_entries_ps_vs_7_T_5; // @[MMUBundle.scala 669:42]
  assign l2_io_wreq_bits_data_2_entries_prefetch = io_refill_bits_req_info_dup_1_source == 2'h2; // @[MMUConst.scala 254:13]
  assign l2_io_wreq_bits_data_2_ecc = {ecc_unaligned,_wdata_ecc_T}; // @[Cat.scala 31:58]
  assign l2_io_wreq_bits_data_3_entries_tag = io_refill_bits_req_info_dup_1_vpn[26:14]; // @[MMUBundle.scala 646:8]
  assign l2_io_wreq_bits_data_3_entries_asid = io_csr_dup_1_satp_asid; // @[MMUBundle.scala 662:18 664:13]
  assign l2_io_wreq_bits_data_3_entries_ppns_0 = io_refill_bits_ptes[33:10]; // @[MMUBundle.scala 667:52]
  assign l2_io_wreq_bits_data_3_entries_ppns_1 = io_refill_bits_ptes[97:74]; // @[MMUBundle.scala 667:52]
  assign l2_io_wreq_bits_data_3_entries_ppns_2 = io_refill_bits_ptes[161:138]; // @[MMUBundle.scala 667:52]
  assign l2_io_wreq_bits_data_3_entries_ppns_3 = io_refill_bits_ptes[225:202]; // @[MMUBundle.scala 667:52]
  assign l2_io_wreq_bits_data_3_entries_ppns_4 = io_refill_bits_ptes[289:266]; // @[MMUBundle.scala 667:52]
  assign l2_io_wreq_bits_data_3_entries_ppns_5 = io_refill_bits_ptes[353:330]; // @[MMUBundle.scala 667:52]
  assign l2_io_wreq_bits_data_3_entries_ppns_6 = io_refill_bits_ptes[417:394]; // @[MMUBundle.scala 667:52]
  assign l2_io_wreq_bits_data_3_entries_ppns_7 = io_refill_bits_ptes[481:458]; // @[MMUBundle.scala 667:52]
  assign l2_io_wreq_bits_data_3_entries_vs_0 = ~_wdata_entries_ps_vs_0_T_19 & ~_wdata_entries_ps_vs_0_T_5; // @[MMUBundle.scala 669:42]
  assign l2_io_wreq_bits_data_3_entries_vs_1 = ~_wdata_entries_ps_vs_1_T_19 & ~_wdata_entries_ps_vs_1_T_5; // @[MMUBundle.scala 669:42]
  assign l2_io_wreq_bits_data_3_entries_vs_2 = ~_wdata_entries_ps_vs_2_T_19 & ~_wdata_entries_ps_vs_2_T_5; // @[MMUBundle.scala 669:42]
  assign l2_io_wreq_bits_data_3_entries_vs_3 = ~_wdata_entries_ps_vs_3_T_19 & ~_wdata_entries_ps_vs_3_T_5; // @[MMUBundle.scala 669:42]
  assign l2_io_wreq_bits_data_3_entries_vs_4 = ~_wdata_entries_ps_vs_4_T_19 & ~_wdata_entries_ps_vs_4_T_5; // @[MMUBundle.scala 669:42]
  assign l2_io_wreq_bits_data_3_entries_vs_5 = ~_wdata_entries_ps_vs_5_T_19 & ~_wdata_entries_ps_vs_5_T_5; // @[MMUBundle.scala 669:42]
  assign l2_io_wreq_bits_data_3_entries_vs_6 = ~_wdata_entries_ps_vs_6_T_19 & ~_wdata_entries_ps_vs_6_T_5; // @[MMUBundle.scala 669:42]
  assign l2_io_wreq_bits_data_3_entries_vs_7 = ~_wdata_entries_ps_vs_7_T_19 & ~_wdata_entries_ps_vs_7_T_5; // @[MMUBundle.scala 669:42]
  assign l2_io_wreq_bits_data_3_entries_prefetch = io_refill_bits_req_info_dup_1_source == 2'h2; // @[MMUConst.scala 254:13]
  assign l2_io_wreq_bits_data_3_ecc = {ecc_unaligned,_wdata_ecc_T}; // @[Cat.scala 31:58]
  assign l2_io_wreq_bits_waymask = 4'h1 << l2_victimWay; // @[OneHot.scala 57:35]
  assign l3_clock = clock;
  assign l3_io_rreq_valid = stageReq_ready & io_req_valid; // @[Decoupled.scala 50:35]
  assign l3_io_rreq_bits_setIdx = io_req_bits_req_info_vpn[4:3]; // @[MMUConst.scala 226:21]
  assign l3_io_wreq_valid = ~flush_dup_2 & io_refill_bits_levelOH_l3 & ~_T_377; // @[PageTableCache.scala 500:44]
  assign l3_io_wreq_bits_setIdx = io_refill_bits_req_info_dup_2_vpn[4:3]; // @[MMUConst.scala 226:21]
  assign l3_io_wreq_bits_data_0_entries_tag = io_refill_bits_req_info_dup_2_vpn[26:5]; // @[MMUBundle.scala 646:8]
  assign l3_io_wreq_bits_data_0_entries_asid = io_csr_dup_2_satp_asid; // @[MMUBundle.scala 662:18 664:13]
  assign l3_io_wreq_bits_data_0_entries_ppns_0 = io_refill_bits_ptes[33:10]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_0_entries_ppns_1 = io_refill_bits_ptes[97:74]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_0_entries_ppns_2 = io_refill_bits_ptes[161:138]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_0_entries_ppns_3 = io_refill_bits_ptes[225:202]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_0_entries_ppns_4 = io_refill_bits_ptes[289:266]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_0_entries_ppns_5 = io_refill_bits_ptes[353:330]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_0_entries_ppns_6 = io_refill_bits_ptes[417:394]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_0_entries_ppns_7 = io_refill_bits_ptes[481:458]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_0_entries_vs_0 = ~_wdata_entries_ps_vs_0_T_3 & _wdata_entries_ps_vs_0_T_5; // @[MMUBundle.scala 669:42]
  assign l3_io_wreq_bits_data_0_entries_vs_1 = ~_wdata_entries_ps_vs_1_T_3 & _wdata_entries_ps_vs_1_T_5; // @[MMUBundle.scala 669:42]
  assign l3_io_wreq_bits_data_0_entries_vs_2 = ~_wdata_entries_ps_vs_2_T_3 & _wdata_entries_ps_vs_2_T_5; // @[MMUBundle.scala 669:42]
  assign l3_io_wreq_bits_data_0_entries_vs_3 = ~_wdata_entries_ps_vs_3_T_3 & _wdata_entries_ps_vs_3_T_5; // @[MMUBundle.scala 669:42]
  assign l3_io_wreq_bits_data_0_entries_vs_4 = ~_wdata_entries_ps_vs_4_T_3 & _wdata_entries_ps_vs_4_T_5; // @[MMUBundle.scala 669:42]
  assign l3_io_wreq_bits_data_0_entries_vs_5 = ~_wdata_entries_ps_vs_5_T_3 & _wdata_entries_ps_vs_5_T_5; // @[MMUBundle.scala 669:42]
  assign l3_io_wreq_bits_data_0_entries_vs_6 = ~_wdata_entries_ps_vs_6_T_3 & _wdata_entries_ps_vs_6_T_5; // @[MMUBundle.scala 669:42]
  assign l3_io_wreq_bits_data_0_entries_vs_7 = ~_wdata_entries_ps_vs_7_T_3 & _wdata_entries_ps_vs_7_T_5; // @[MMUBundle.scala 669:42]
  assign l3_io_wreq_bits_data_0_entries_perms_0_d = io_refill_bits_ptes[7]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_0_entries_perms_0_a = io_refill_bits_ptes[6]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_0_entries_perms_0_g = io_refill_bits_ptes[5]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_0_entries_perms_0_u = io_refill_bits_ptes[4]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_0_entries_perms_0_x = io_refill_bits_ptes[3]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_0_entries_perms_0_w = io_refill_bits_ptes[2]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_0_entries_perms_0_r = io_refill_bits_ptes[1]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_0_entries_perms_1_d = io_refill_bits_ptes[71]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_0_entries_perms_1_a = io_refill_bits_ptes[70]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_0_entries_perms_1_g = io_refill_bits_ptes[69]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_0_entries_perms_1_u = io_refill_bits_ptes[68]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_0_entries_perms_1_x = io_refill_bits_ptes[67]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_0_entries_perms_1_w = io_refill_bits_ptes[66]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_0_entries_perms_1_r = io_refill_bits_ptes[65]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_0_entries_perms_2_d = io_refill_bits_ptes[135]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_0_entries_perms_2_a = io_refill_bits_ptes[134]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_0_entries_perms_2_g = io_refill_bits_ptes[133]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_0_entries_perms_2_u = io_refill_bits_ptes[132]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_0_entries_perms_2_x = io_refill_bits_ptes[131]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_0_entries_perms_2_w = io_refill_bits_ptes[130]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_0_entries_perms_2_r = io_refill_bits_ptes[129]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_0_entries_perms_3_d = io_refill_bits_ptes[199]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_0_entries_perms_3_a = io_refill_bits_ptes[198]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_0_entries_perms_3_g = io_refill_bits_ptes[197]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_0_entries_perms_3_u = io_refill_bits_ptes[196]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_0_entries_perms_3_x = io_refill_bits_ptes[195]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_0_entries_perms_3_w = io_refill_bits_ptes[194]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_0_entries_perms_3_r = io_refill_bits_ptes[193]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_0_entries_perms_4_d = io_refill_bits_ptes[263]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_0_entries_perms_4_a = io_refill_bits_ptes[262]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_0_entries_perms_4_g = io_refill_bits_ptes[261]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_0_entries_perms_4_u = io_refill_bits_ptes[260]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_0_entries_perms_4_x = io_refill_bits_ptes[259]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_0_entries_perms_4_w = io_refill_bits_ptes[258]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_0_entries_perms_4_r = io_refill_bits_ptes[257]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_0_entries_perms_5_d = io_refill_bits_ptes[327]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_0_entries_perms_5_a = io_refill_bits_ptes[326]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_0_entries_perms_5_g = io_refill_bits_ptes[325]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_0_entries_perms_5_u = io_refill_bits_ptes[324]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_0_entries_perms_5_x = io_refill_bits_ptes[323]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_0_entries_perms_5_w = io_refill_bits_ptes[322]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_0_entries_perms_5_r = io_refill_bits_ptes[321]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_0_entries_perms_6_d = io_refill_bits_ptes[391]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_0_entries_perms_6_a = io_refill_bits_ptes[390]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_0_entries_perms_6_g = io_refill_bits_ptes[389]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_0_entries_perms_6_u = io_refill_bits_ptes[388]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_0_entries_perms_6_x = io_refill_bits_ptes[387]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_0_entries_perms_6_w = io_refill_bits_ptes[386]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_0_entries_perms_6_r = io_refill_bits_ptes[385]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_0_entries_perms_7_d = io_refill_bits_ptes[455]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_0_entries_perms_7_a = io_refill_bits_ptes[454]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_0_entries_perms_7_g = io_refill_bits_ptes[453]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_0_entries_perms_7_u = io_refill_bits_ptes[452]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_0_entries_perms_7_x = io_refill_bits_ptes[451]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_0_entries_perms_7_w = io_refill_bits_ptes[450]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_0_entries_perms_7_r = io_refill_bits_ptes[449]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_0_entries_prefetch = io_refill_bits_req_info_dup_2_source == 2'h2; // @[MMUConst.scala 254:13]
  assign l3_io_wreq_bits_data_0_ecc = {ecc_unaligned_1,_wdata_ecc_T_2}; // @[Cat.scala 31:58]
  assign l3_io_wreq_bits_data_1_entries_tag = io_refill_bits_req_info_dup_2_vpn[26:5]; // @[MMUBundle.scala 646:8]
  assign l3_io_wreq_bits_data_1_entries_asid = io_csr_dup_2_satp_asid; // @[MMUBundle.scala 662:18 664:13]
  assign l3_io_wreq_bits_data_1_entries_ppns_0 = io_refill_bits_ptes[33:10]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_1_entries_ppns_1 = io_refill_bits_ptes[97:74]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_1_entries_ppns_2 = io_refill_bits_ptes[161:138]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_1_entries_ppns_3 = io_refill_bits_ptes[225:202]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_1_entries_ppns_4 = io_refill_bits_ptes[289:266]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_1_entries_ppns_5 = io_refill_bits_ptes[353:330]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_1_entries_ppns_6 = io_refill_bits_ptes[417:394]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_1_entries_ppns_7 = io_refill_bits_ptes[481:458]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_1_entries_vs_0 = ~_wdata_entries_ps_vs_0_T_3 & _wdata_entries_ps_vs_0_T_5; // @[MMUBundle.scala 669:42]
  assign l3_io_wreq_bits_data_1_entries_vs_1 = ~_wdata_entries_ps_vs_1_T_3 & _wdata_entries_ps_vs_1_T_5; // @[MMUBundle.scala 669:42]
  assign l3_io_wreq_bits_data_1_entries_vs_2 = ~_wdata_entries_ps_vs_2_T_3 & _wdata_entries_ps_vs_2_T_5; // @[MMUBundle.scala 669:42]
  assign l3_io_wreq_bits_data_1_entries_vs_3 = ~_wdata_entries_ps_vs_3_T_3 & _wdata_entries_ps_vs_3_T_5; // @[MMUBundle.scala 669:42]
  assign l3_io_wreq_bits_data_1_entries_vs_4 = ~_wdata_entries_ps_vs_4_T_3 & _wdata_entries_ps_vs_4_T_5; // @[MMUBundle.scala 669:42]
  assign l3_io_wreq_bits_data_1_entries_vs_5 = ~_wdata_entries_ps_vs_5_T_3 & _wdata_entries_ps_vs_5_T_5; // @[MMUBundle.scala 669:42]
  assign l3_io_wreq_bits_data_1_entries_vs_6 = ~_wdata_entries_ps_vs_6_T_3 & _wdata_entries_ps_vs_6_T_5; // @[MMUBundle.scala 669:42]
  assign l3_io_wreq_bits_data_1_entries_vs_7 = ~_wdata_entries_ps_vs_7_T_3 & _wdata_entries_ps_vs_7_T_5; // @[MMUBundle.scala 669:42]
  assign l3_io_wreq_bits_data_1_entries_perms_0_d = io_refill_bits_ptes[7]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_1_entries_perms_0_a = io_refill_bits_ptes[6]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_1_entries_perms_0_g = io_refill_bits_ptes[5]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_1_entries_perms_0_u = io_refill_bits_ptes[4]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_1_entries_perms_0_x = io_refill_bits_ptes[3]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_1_entries_perms_0_w = io_refill_bits_ptes[2]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_1_entries_perms_0_r = io_refill_bits_ptes[1]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_1_entries_perms_1_d = io_refill_bits_ptes[71]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_1_entries_perms_1_a = io_refill_bits_ptes[70]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_1_entries_perms_1_g = io_refill_bits_ptes[69]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_1_entries_perms_1_u = io_refill_bits_ptes[68]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_1_entries_perms_1_x = io_refill_bits_ptes[67]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_1_entries_perms_1_w = io_refill_bits_ptes[66]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_1_entries_perms_1_r = io_refill_bits_ptes[65]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_1_entries_perms_2_d = io_refill_bits_ptes[135]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_1_entries_perms_2_a = io_refill_bits_ptes[134]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_1_entries_perms_2_g = io_refill_bits_ptes[133]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_1_entries_perms_2_u = io_refill_bits_ptes[132]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_1_entries_perms_2_x = io_refill_bits_ptes[131]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_1_entries_perms_2_w = io_refill_bits_ptes[130]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_1_entries_perms_2_r = io_refill_bits_ptes[129]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_1_entries_perms_3_d = io_refill_bits_ptes[199]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_1_entries_perms_3_a = io_refill_bits_ptes[198]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_1_entries_perms_3_g = io_refill_bits_ptes[197]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_1_entries_perms_3_u = io_refill_bits_ptes[196]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_1_entries_perms_3_x = io_refill_bits_ptes[195]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_1_entries_perms_3_w = io_refill_bits_ptes[194]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_1_entries_perms_3_r = io_refill_bits_ptes[193]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_1_entries_perms_4_d = io_refill_bits_ptes[263]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_1_entries_perms_4_a = io_refill_bits_ptes[262]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_1_entries_perms_4_g = io_refill_bits_ptes[261]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_1_entries_perms_4_u = io_refill_bits_ptes[260]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_1_entries_perms_4_x = io_refill_bits_ptes[259]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_1_entries_perms_4_w = io_refill_bits_ptes[258]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_1_entries_perms_4_r = io_refill_bits_ptes[257]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_1_entries_perms_5_d = io_refill_bits_ptes[327]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_1_entries_perms_5_a = io_refill_bits_ptes[326]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_1_entries_perms_5_g = io_refill_bits_ptes[325]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_1_entries_perms_5_u = io_refill_bits_ptes[324]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_1_entries_perms_5_x = io_refill_bits_ptes[323]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_1_entries_perms_5_w = io_refill_bits_ptes[322]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_1_entries_perms_5_r = io_refill_bits_ptes[321]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_1_entries_perms_6_d = io_refill_bits_ptes[391]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_1_entries_perms_6_a = io_refill_bits_ptes[390]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_1_entries_perms_6_g = io_refill_bits_ptes[389]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_1_entries_perms_6_u = io_refill_bits_ptes[388]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_1_entries_perms_6_x = io_refill_bits_ptes[387]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_1_entries_perms_6_w = io_refill_bits_ptes[386]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_1_entries_perms_6_r = io_refill_bits_ptes[385]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_1_entries_perms_7_d = io_refill_bits_ptes[455]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_1_entries_perms_7_a = io_refill_bits_ptes[454]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_1_entries_perms_7_g = io_refill_bits_ptes[453]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_1_entries_perms_7_u = io_refill_bits_ptes[452]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_1_entries_perms_7_x = io_refill_bits_ptes[451]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_1_entries_perms_7_w = io_refill_bits_ptes[450]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_1_entries_perms_7_r = io_refill_bits_ptes[449]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_1_entries_prefetch = io_refill_bits_req_info_dup_2_source == 2'h2; // @[MMUConst.scala 254:13]
  assign l3_io_wreq_bits_data_1_ecc = {ecc_unaligned_1,_wdata_ecc_T_2}; // @[Cat.scala 31:58]
  assign l3_io_wreq_bits_data_2_entries_tag = io_refill_bits_req_info_dup_2_vpn[26:5]; // @[MMUBundle.scala 646:8]
  assign l3_io_wreq_bits_data_2_entries_asid = io_csr_dup_2_satp_asid; // @[MMUBundle.scala 662:18 664:13]
  assign l3_io_wreq_bits_data_2_entries_ppns_0 = io_refill_bits_ptes[33:10]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_2_entries_ppns_1 = io_refill_bits_ptes[97:74]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_2_entries_ppns_2 = io_refill_bits_ptes[161:138]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_2_entries_ppns_3 = io_refill_bits_ptes[225:202]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_2_entries_ppns_4 = io_refill_bits_ptes[289:266]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_2_entries_ppns_5 = io_refill_bits_ptes[353:330]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_2_entries_ppns_6 = io_refill_bits_ptes[417:394]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_2_entries_ppns_7 = io_refill_bits_ptes[481:458]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_2_entries_vs_0 = ~_wdata_entries_ps_vs_0_T_3 & _wdata_entries_ps_vs_0_T_5; // @[MMUBundle.scala 669:42]
  assign l3_io_wreq_bits_data_2_entries_vs_1 = ~_wdata_entries_ps_vs_1_T_3 & _wdata_entries_ps_vs_1_T_5; // @[MMUBundle.scala 669:42]
  assign l3_io_wreq_bits_data_2_entries_vs_2 = ~_wdata_entries_ps_vs_2_T_3 & _wdata_entries_ps_vs_2_T_5; // @[MMUBundle.scala 669:42]
  assign l3_io_wreq_bits_data_2_entries_vs_3 = ~_wdata_entries_ps_vs_3_T_3 & _wdata_entries_ps_vs_3_T_5; // @[MMUBundle.scala 669:42]
  assign l3_io_wreq_bits_data_2_entries_vs_4 = ~_wdata_entries_ps_vs_4_T_3 & _wdata_entries_ps_vs_4_T_5; // @[MMUBundle.scala 669:42]
  assign l3_io_wreq_bits_data_2_entries_vs_5 = ~_wdata_entries_ps_vs_5_T_3 & _wdata_entries_ps_vs_5_T_5; // @[MMUBundle.scala 669:42]
  assign l3_io_wreq_bits_data_2_entries_vs_6 = ~_wdata_entries_ps_vs_6_T_3 & _wdata_entries_ps_vs_6_T_5; // @[MMUBundle.scala 669:42]
  assign l3_io_wreq_bits_data_2_entries_vs_7 = ~_wdata_entries_ps_vs_7_T_3 & _wdata_entries_ps_vs_7_T_5; // @[MMUBundle.scala 669:42]
  assign l3_io_wreq_bits_data_2_entries_perms_0_d = io_refill_bits_ptes[7]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_2_entries_perms_0_a = io_refill_bits_ptes[6]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_2_entries_perms_0_g = io_refill_bits_ptes[5]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_2_entries_perms_0_u = io_refill_bits_ptes[4]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_2_entries_perms_0_x = io_refill_bits_ptes[3]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_2_entries_perms_0_w = io_refill_bits_ptes[2]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_2_entries_perms_0_r = io_refill_bits_ptes[1]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_2_entries_perms_1_d = io_refill_bits_ptes[71]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_2_entries_perms_1_a = io_refill_bits_ptes[70]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_2_entries_perms_1_g = io_refill_bits_ptes[69]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_2_entries_perms_1_u = io_refill_bits_ptes[68]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_2_entries_perms_1_x = io_refill_bits_ptes[67]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_2_entries_perms_1_w = io_refill_bits_ptes[66]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_2_entries_perms_1_r = io_refill_bits_ptes[65]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_2_entries_perms_2_d = io_refill_bits_ptes[135]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_2_entries_perms_2_a = io_refill_bits_ptes[134]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_2_entries_perms_2_g = io_refill_bits_ptes[133]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_2_entries_perms_2_u = io_refill_bits_ptes[132]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_2_entries_perms_2_x = io_refill_bits_ptes[131]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_2_entries_perms_2_w = io_refill_bits_ptes[130]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_2_entries_perms_2_r = io_refill_bits_ptes[129]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_2_entries_perms_3_d = io_refill_bits_ptes[199]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_2_entries_perms_3_a = io_refill_bits_ptes[198]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_2_entries_perms_3_g = io_refill_bits_ptes[197]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_2_entries_perms_3_u = io_refill_bits_ptes[196]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_2_entries_perms_3_x = io_refill_bits_ptes[195]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_2_entries_perms_3_w = io_refill_bits_ptes[194]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_2_entries_perms_3_r = io_refill_bits_ptes[193]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_2_entries_perms_4_d = io_refill_bits_ptes[263]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_2_entries_perms_4_a = io_refill_bits_ptes[262]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_2_entries_perms_4_g = io_refill_bits_ptes[261]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_2_entries_perms_4_u = io_refill_bits_ptes[260]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_2_entries_perms_4_x = io_refill_bits_ptes[259]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_2_entries_perms_4_w = io_refill_bits_ptes[258]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_2_entries_perms_4_r = io_refill_bits_ptes[257]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_2_entries_perms_5_d = io_refill_bits_ptes[327]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_2_entries_perms_5_a = io_refill_bits_ptes[326]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_2_entries_perms_5_g = io_refill_bits_ptes[325]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_2_entries_perms_5_u = io_refill_bits_ptes[324]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_2_entries_perms_5_x = io_refill_bits_ptes[323]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_2_entries_perms_5_w = io_refill_bits_ptes[322]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_2_entries_perms_5_r = io_refill_bits_ptes[321]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_2_entries_perms_6_d = io_refill_bits_ptes[391]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_2_entries_perms_6_a = io_refill_bits_ptes[390]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_2_entries_perms_6_g = io_refill_bits_ptes[389]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_2_entries_perms_6_u = io_refill_bits_ptes[388]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_2_entries_perms_6_x = io_refill_bits_ptes[387]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_2_entries_perms_6_w = io_refill_bits_ptes[386]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_2_entries_perms_6_r = io_refill_bits_ptes[385]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_2_entries_perms_7_d = io_refill_bits_ptes[455]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_2_entries_perms_7_a = io_refill_bits_ptes[454]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_2_entries_perms_7_g = io_refill_bits_ptes[453]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_2_entries_perms_7_u = io_refill_bits_ptes[452]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_2_entries_perms_7_x = io_refill_bits_ptes[451]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_2_entries_perms_7_w = io_refill_bits_ptes[450]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_2_entries_perms_7_r = io_refill_bits_ptes[449]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_2_entries_prefetch = io_refill_bits_req_info_dup_2_source == 2'h2; // @[MMUConst.scala 254:13]
  assign l3_io_wreq_bits_data_2_ecc = {ecc_unaligned_1,_wdata_ecc_T_2}; // @[Cat.scala 31:58]
  assign l3_io_wreq_bits_data_3_entries_tag = io_refill_bits_req_info_dup_2_vpn[26:5]; // @[MMUBundle.scala 646:8]
  assign l3_io_wreq_bits_data_3_entries_asid = io_csr_dup_2_satp_asid; // @[MMUBundle.scala 662:18 664:13]
  assign l3_io_wreq_bits_data_3_entries_ppns_0 = io_refill_bits_ptes[33:10]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_3_entries_ppns_1 = io_refill_bits_ptes[97:74]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_3_entries_ppns_2 = io_refill_bits_ptes[161:138]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_3_entries_ppns_3 = io_refill_bits_ptes[225:202]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_3_entries_ppns_4 = io_refill_bits_ptes[289:266]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_3_entries_ppns_5 = io_refill_bits_ptes[353:330]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_3_entries_ppns_6 = io_refill_bits_ptes[417:394]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_3_entries_ppns_7 = io_refill_bits_ptes[481:458]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_3_entries_vs_0 = ~_wdata_entries_ps_vs_0_T_3 & _wdata_entries_ps_vs_0_T_5; // @[MMUBundle.scala 669:42]
  assign l3_io_wreq_bits_data_3_entries_vs_1 = ~_wdata_entries_ps_vs_1_T_3 & _wdata_entries_ps_vs_1_T_5; // @[MMUBundle.scala 669:42]
  assign l3_io_wreq_bits_data_3_entries_vs_2 = ~_wdata_entries_ps_vs_2_T_3 & _wdata_entries_ps_vs_2_T_5; // @[MMUBundle.scala 669:42]
  assign l3_io_wreq_bits_data_3_entries_vs_3 = ~_wdata_entries_ps_vs_3_T_3 & _wdata_entries_ps_vs_3_T_5; // @[MMUBundle.scala 669:42]
  assign l3_io_wreq_bits_data_3_entries_vs_4 = ~_wdata_entries_ps_vs_4_T_3 & _wdata_entries_ps_vs_4_T_5; // @[MMUBundle.scala 669:42]
  assign l3_io_wreq_bits_data_3_entries_vs_5 = ~_wdata_entries_ps_vs_5_T_3 & _wdata_entries_ps_vs_5_T_5; // @[MMUBundle.scala 669:42]
  assign l3_io_wreq_bits_data_3_entries_vs_6 = ~_wdata_entries_ps_vs_6_T_3 & _wdata_entries_ps_vs_6_T_5; // @[MMUBundle.scala 669:42]
  assign l3_io_wreq_bits_data_3_entries_vs_7 = ~_wdata_entries_ps_vs_7_T_3 & _wdata_entries_ps_vs_7_T_5; // @[MMUBundle.scala 669:42]
  assign l3_io_wreq_bits_data_3_entries_perms_0_d = io_refill_bits_ptes[7]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_3_entries_perms_0_a = io_refill_bits_ptes[6]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_3_entries_perms_0_g = io_refill_bits_ptes[5]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_3_entries_perms_0_u = io_refill_bits_ptes[4]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_3_entries_perms_0_x = io_refill_bits_ptes[3]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_3_entries_perms_0_w = io_refill_bits_ptes[2]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_3_entries_perms_0_r = io_refill_bits_ptes[1]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_3_entries_perms_1_d = io_refill_bits_ptes[71]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_3_entries_perms_1_a = io_refill_bits_ptes[70]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_3_entries_perms_1_g = io_refill_bits_ptes[69]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_3_entries_perms_1_u = io_refill_bits_ptes[68]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_3_entries_perms_1_x = io_refill_bits_ptes[67]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_3_entries_perms_1_w = io_refill_bits_ptes[66]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_3_entries_perms_1_r = io_refill_bits_ptes[65]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_3_entries_perms_2_d = io_refill_bits_ptes[135]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_3_entries_perms_2_a = io_refill_bits_ptes[134]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_3_entries_perms_2_g = io_refill_bits_ptes[133]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_3_entries_perms_2_u = io_refill_bits_ptes[132]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_3_entries_perms_2_x = io_refill_bits_ptes[131]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_3_entries_perms_2_w = io_refill_bits_ptes[130]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_3_entries_perms_2_r = io_refill_bits_ptes[129]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_3_entries_perms_3_d = io_refill_bits_ptes[199]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_3_entries_perms_3_a = io_refill_bits_ptes[198]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_3_entries_perms_3_g = io_refill_bits_ptes[197]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_3_entries_perms_3_u = io_refill_bits_ptes[196]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_3_entries_perms_3_x = io_refill_bits_ptes[195]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_3_entries_perms_3_w = io_refill_bits_ptes[194]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_3_entries_perms_3_r = io_refill_bits_ptes[193]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_3_entries_perms_4_d = io_refill_bits_ptes[263]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_3_entries_perms_4_a = io_refill_bits_ptes[262]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_3_entries_perms_4_g = io_refill_bits_ptes[261]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_3_entries_perms_4_u = io_refill_bits_ptes[260]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_3_entries_perms_4_x = io_refill_bits_ptes[259]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_3_entries_perms_4_w = io_refill_bits_ptes[258]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_3_entries_perms_4_r = io_refill_bits_ptes[257]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_3_entries_perms_5_d = io_refill_bits_ptes[327]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_3_entries_perms_5_a = io_refill_bits_ptes[326]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_3_entries_perms_5_g = io_refill_bits_ptes[325]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_3_entries_perms_5_u = io_refill_bits_ptes[324]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_3_entries_perms_5_x = io_refill_bits_ptes[323]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_3_entries_perms_5_w = io_refill_bits_ptes[322]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_3_entries_perms_5_r = io_refill_bits_ptes[321]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_3_entries_perms_6_d = io_refill_bits_ptes[391]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_3_entries_perms_6_a = io_refill_bits_ptes[390]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_3_entries_perms_6_g = io_refill_bits_ptes[389]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_3_entries_perms_6_u = io_refill_bits_ptes[388]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_3_entries_perms_6_x = io_refill_bits_ptes[387]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_3_entries_perms_6_w = io_refill_bits_ptes[386]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_3_entries_perms_6_r = io_refill_bits_ptes[385]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_3_entries_perms_7_d = io_refill_bits_ptes[455]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_3_entries_perms_7_a = io_refill_bits_ptes[454]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_3_entries_perms_7_g = io_refill_bits_ptes[453]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_3_entries_perms_7_u = io_refill_bits_ptes[452]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_3_entries_perms_7_x = io_refill_bits_ptes[451]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_3_entries_perms_7_w = io_refill_bits_ptes[450]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_3_entries_perms_7_r = io_refill_bits_ptes[449]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_3_entries_prefetch = io_refill_bits_req_info_dup_2_source == 2'h2; // @[MMUConst.scala 254:13]
  assign l3_io_wreq_bits_data_3_ecc = {ecc_unaligned_1,_wdata_ecc_T_2}; // @[Cat.scala 31:58]
  assign l3_io_wreq_bits_data_4_entries_tag = io_refill_bits_req_info_dup_2_vpn[26:5]; // @[MMUBundle.scala 646:8]
  assign l3_io_wreq_bits_data_4_entries_asid = io_csr_dup_2_satp_asid; // @[MMUBundle.scala 662:18 664:13]
  assign l3_io_wreq_bits_data_4_entries_ppns_0 = io_refill_bits_ptes[33:10]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_4_entries_ppns_1 = io_refill_bits_ptes[97:74]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_4_entries_ppns_2 = io_refill_bits_ptes[161:138]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_4_entries_ppns_3 = io_refill_bits_ptes[225:202]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_4_entries_ppns_4 = io_refill_bits_ptes[289:266]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_4_entries_ppns_5 = io_refill_bits_ptes[353:330]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_4_entries_ppns_6 = io_refill_bits_ptes[417:394]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_4_entries_ppns_7 = io_refill_bits_ptes[481:458]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_4_entries_vs_0 = ~_wdata_entries_ps_vs_0_T_3 & _wdata_entries_ps_vs_0_T_5; // @[MMUBundle.scala 669:42]
  assign l3_io_wreq_bits_data_4_entries_vs_1 = ~_wdata_entries_ps_vs_1_T_3 & _wdata_entries_ps_vs_1_T_5; // @[MMUBundle.scala 669:42]
  assign l3_io_wreq_bits_data_4_entries_vs_2 = ~_wdata_entries_ps_vs_2_T_3 & _wdata_entries_ps_vs_2_T_5; // @[MMUBundle.scala 669:42]
  assign l3_io_wreq_bits_data_4_entries_vs_3 = ~_wdata_entries_ps_vs_3_T_3 & _wdata_entries_ps_vs_3_T_5; // @[MMUBundle.scala 669:42]
  assign l3_io_wreq_bits_data_4_entries_vs_4 = ~_wdata_entries_ps_vs_4_T_3 & _wdata_entries_ps_vs_4_T_5; // @[MMUBundle.scala 669:42]
  assign l3_io_wreq_bits_data_4_entries_vs_5 = ~_wdata_entries_ps_vs_5_T_3 & _wdata_entries_ps_vs_5_T_5; // @[MMUBundle.scala 669:42]
  assign l3_io_wreq_bits_data_4_entries_vs_6 = ~_wdata_entries_ps_vs_6_T_3 & _wdata_entries_ps_vs_6_T_5; // @[MMUBundle.scala 669:42]
  assign l3_io_wreq_bits_data_4_entries_vs_7 = ~_wdata_entries_ps_vs_7_T_3 & _wdata_entries_ps_vs_7_T_5; // @[MMUBundle.scala 669:42]
  assign l3_io_wreq_bits_data_4_entries_perms_0_d = io_refill_bits_ptes[7]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_4_entries_perms_0_a = io_refill_bits_ptes[6]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_4_entries_perms_0_g = io_refill_bits_ptes[5]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_4_entries_perms_0_u = io_refill_bits_ptes[4]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_4_entries_perms_0_x = io_refill_bits_ptes[3]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_4_entries_perms_0_w = io_refill_bits_ptes[2]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_4_entries_perms_0_r = io_refill_bits_ptes[1]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_4_entries_perms_1_d = io_refill_bits_ptes[71]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_4_entries_perms_1_a = io_refill_bits_ptes[70]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_4_entries_perms_1_g = io_refill_bits_ptes[69]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_4_entries_perms_1_u = io_refill_bits_ptes[68]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_4_entries_perms_1_x = io_refill_bits_ptes[67]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_4_entries_perms_1_w = io_refill_bits_ptes[66]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_4_entries_perms_1_r = io_refill_bits_ptes[65]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_4_entries_perms_2_d = io_refill_bits_ptes[135]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_4_entries_perms_2_a = io_refill_bits_ptes[134]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_4_entries_perms_2_g = io_refill_bits_ptes[133]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_4_entries_perms_2_u = io_refill_bits_ptes[132]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_4_entries_perms_2_x = io_refill_bits_ptes[131]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_4_entries_perms_2_w = io_refill_bits_ptes[130]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_4_entries_perms_2_r = io_refill_bits_ptes[129]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_4_entries_perms_3_d = io_refill_bits_ptes[199]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_4_entries_perms_3_a = io_refill_bits_ptes[198]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_4_entries_perms_3_g = io_refill_bits_ptes[197]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_4_entries_perms_3_u = io_refill_bits_ptes[196]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_4_entries_perms_3_x = io_refill_bits_ptes[195]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_4_entries_perms_3_w = io_refill_bits_ptes[194]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_4_entries_perms_3_r = io_refill_bits_ptes[193]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_4_entries_perms_4_d = io_refill_bits_ptes[263]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_4_entries_perms_4_a = io_refill_bits_ptes[262]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_4_entries_perms_4_g = io_refill_bits_ptes[261]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_4_entries_perms_4_u = io_refill_bits_ptes[260]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_4_entries_perms_4_x = io_refill_bits_ptes[259]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_4_entries_perms_4_w = io_refill_bits_ptes[258]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_4_entries_perms_4_r = io_refill_bits_ptes[257]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_4_entries_perms_5_d = io_refill_bits_ptes[327]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_4_entries_perms_5_a = io_refill_bits_ptes[326]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_4_entries_perms_5_g = io_refill_bits_ptes[325]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_4_entries_perms_5_u = io_refill_bits_ptes[324]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_4_entries_perms_5_x = io_refill_bits_ptes[323]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_4_entries_perms_5_w = io_refill_bits_ptes[322]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_4_entries_perms_5_r = io_refill_bits_ptes[321]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_4_entries_perms_6_d = io_refill_bits_ptes[391]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_4_entries_perms_6_a = io_refill_bits_ptes[390]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_4_entries_perms_6_g = io_refill_bits_ptes[389]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_4_entries_perms_6_u = io_refill_bits_ptes[388]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_4_entries_perms_6_x = io_refill_bits_ptes[387]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_4_entries_perms_6_w = io_refill_bits_ptes[386]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_4_entries_perms_6_r = io_refill_bits_ptes[385]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_4_entries_perms_7_d = io_refill_bits_ptes[455]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_4_entries_perms_7_a = io_refill_bits_ptes[454]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_4_entries_perms_7_g = io_refill_bits_ptes[453]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_4_entries_perms_7_u = io_refill_bits_ptes[452]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_4_entries_perms_7_x = io_refill_bits_ptes[451]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_4_entries_perms_7_w = io_refill_bits_ptes[450]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_4_entries_perms_7_r = io_refill_bits_ptes[449]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_4_entries_prefetch = io_refill_bits_req_info_dup_2_source == 2'h2; // @[MMUConst.scala 254:13]
  assign l3_io_wreq_bits_data_4_ecc = {ecc_unaligned_1,_wdata_ecc_T_2}; // @[Cat.scala 31:58]
  assign l3_io_wreq_bits_data_5_entries_tag = io_refill_bits_req_info_dup_2_vpn[26:5]; // @[MMUBundle.scala 646:8]
  assign l3_io_wreq_bits_data_5_entries_asid = io_csr_dup_2_satp_asid; // @[MMUBundle.scala 662:18 664:13]
  assign l3_io_wreq_bits_data_5_entries_ppns_0 = io_refill_bits_ptes[33:10]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_5_entries_ppns_1 = io_refill_bits_ptes[97:74]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_5_entries_ppns_2 = io_refill_bits_ptes[161:138]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_5_entries_ppns_3 = io_refill_bits_ptes[225:202]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_5_entries_ppns_4 = io_refill_bits_ptes[289:266]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_5_entries_ppns_5 = io_refill_bits_ptes[353:330]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_5_entries_ppns_6 = io_refill_bits_ptes[417:394]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_5_entries_ppns_7 = io_refill_bits_ptes[481:458]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_5_entries_vs_0 = ~_wdata_entries_ps_vs_0_T_3 & _wdata_entries_ps_vs_0_T_5; // @[MMUBundle.scala 669:42]
  assign l3_io_wreq_bits_data_5_entries_vs_1 = ~_wdata_entries_ps_vs_1_T_3 & _wdata_entries_ps_vs_1_T_5; // @[MMUBundle.scala 669:42]
  assign l3_io_wreq_bits_data_5_entries_vs_2 = ~_wdata_entries_ps_vs_2_T_3 & _wdata_entries_ps_vs_2_T_5; // @[MMUBundle.scala 669:42]
  assign l3_io_wreq_bits_data_5_entries_vs_3 = ~_wdata_entries_ps_vs_3_T_3 & _wdata_entries_ps_vs_3_T_5; // @[MMUBundle.scala 669:42]
  assign l3_io_wreq_bits_data_5_entries_vs_4 = ~_wdata_entries_ps_vs_4_T_3 & _wdata_entries_ps_vs_4_T_5; // @[MMUBundle.scala 669:42]
  assign l3_io_wreq_bits_data_5_entries_vs_5 = ~_wdata_entries_ps_vs_5_T_3 & _wdata_entries_ps_vs_5_T_5; // @[MMUBundle.scala 669:42]
  assign l3_io_wreq_bits_data_5_entries_vs_6 = ~_wdata_entries_ps_vs_6_T_3 & _wdata_entries_ps_vs_6_T_5; // @[MMUBundle.scala 669:42]
  assign l3_io_wreq_bits_data_5_entries_vs_7 = ~_wdata_entries_ps_vs_7_T_3 & _wdata_entries_ps_vs_7_T_5; // @[MMUBundle.scala 669:42]
  assign l3_io_wreq_bits_data_5_entries_perms_0_d = io_refill_bits_ptes[7]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_5_entries_perms_0_a = io_refill_bits_ptes[6]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_5_entries_perms_0_g = io_refill_bits_ptes[5]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_5_entries_perms_0_u = io_refill_bits_ptes[4]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_5_entries_perms_0_x = io_refill_bits_ptes[3]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_5_entries_perms_0_w = io_refill_bits_ptes[2]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_5_entries_perms_0_r = io_refill_bits_ptes[1]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_5_entries_perms_1_d = io_refill_bits_ptes[71]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_5_entries_perms_1_a = io_refill_bits_ptes[70]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_5_entries_perms_1_g = io_refill_bits_ptes[69]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_5_entries_perms_1_u = io_refill_bits_ptes[68]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_5_entries_perms_1_x = io_refill_bits_ptes[67]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_5_entries_perms_1_w = io_refill_bits_ptes[66]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_5_entries_perms_1_r = io_refill_bits_ptes[65]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_5_entries_perms_2_d = io_refill_bits_ptes[135]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_5_entries_perms_2_a = io_refill_bits_ptes[134]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_5_entries_perms_2_g = io_refill_bits_ptes[133]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_5_entries_perms_2_u = io_refill_bits_ptes[132]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_5_entries_perms_2_x = io_refill_bits_ptes[131]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_5_entries_perms_2_w = io_refill_bits_ptes[130]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_5_entries_perms_2_r = io_refill_bits_ptes[129]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_5_entries_perms_3_d = io_refill_bits_ptes[199]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_5_entries_perms_3_a = io_refill_bits_ptes[198]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_5_entries_perms_3_g = io_refill_bits_ptes[197]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_5_entries_perms_3_u = io_refill_bits_ptes[196]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_5_entries_perms_3_x = io_refill_bits_ptes[195]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_5_entries_perms_3_w = io_refill_bits_ptes[194]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_5_entries_perms_3_r = io_refill_bits_ptes[193]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_5_entries_perms_4_d = io_refill_bits_ptes[263]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_5_entries_perms_4_a = io_refill_bits_ptes[262]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_5_entries_perms_4_g = io_refill_bits_ptes[261]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_5_entries_perms_4_u = io_refill_bits_ptes[260]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_5_entries_perms_4_x = io_refill_bits_ptes[259]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_5_entries_perms_4_w = io_refill_bits_ptes[258]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_5_entries_perms_4_r = io_refill_bits_ptes[257]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_5_entries_perms_5_d = io_refill_bits_ptes[327]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_5_entries_perms_5_a = io_refill_bits_ptes[326]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_5_entries_perms_5_g = io_refill_bits_ptes[325]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_5_entries_perms_5_u = io_refill_bits_ptes[324]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_5_entries_perms_5_x = io_refill_bits_ptes[323]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_5_entries_perms_5_w = io_refill_bits_ptes[322]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_5_entries_perms_5_r = io_refill_bits_ptes[321]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_5_entries_perms_6_d = io_refill_bits_ptes[391]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_5_entries_perms_6_a = io_refill_bits_ptes[390]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_5_entries_perms_6_g = io_refill_bits_ptes[389]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_5_entries_perms_6_u = io_refill_bits_ptes[388]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_5_entries_perms_6_x = io_refill_bits_ptes[387]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_5_entries_perms_6_w = io_refill_bits_ptes[386]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_5_entries_perms_6_r = io_refill_bits_ptes[385]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_5_entries_perms_7_d = io_refill_bits_ptes[455]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_5_entries_perms_7_a = io_refill_bits_ptes[454]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_5_entries_perms_7_g = io_refill_bits_ptes[453]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_5_entries_perms_7_u = io_refill_bits_ptes[452]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_5_entries_perms_7_x = io_refill_bits_ptes[451]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_5_entries_perms_7_w = io_refill_bits_ptes[450]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_5_entries_perms_7_r = io_refill_bits_ptes[449]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_5_entries_prefetch = io_refill_bits_req_info_dup_2_source == 2'h2; // @[MMUConst.scala 254:13]
  assign l3_io_wreq_bits_data_5_ecc = {ecc_unaligned_1,_wdata_ecc_T_2}; // @[Cat.scala 31:58]
  assign l3_io_wreq_bits_data_6_entries_tag = io_refill_bits_req_info_dup_2_vpn[26:5]; // @[MMUBundle.scala 646:8]
  assign l3_io_wreq_bits_data_6_entries_asid = io_csr_dup_2_satp_asid; // @[MMUBundle.scala 662:18 664:13]
  assign l3_io_wreq_bits_data_6_entries_ppns_0 = io_refill_bits_ptes[33:10]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_6_entries_ppns_1 = io_refill_bits_ptes[97:74]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_6_entries_ppns_2 = io_refill_bits_ptes[161:138]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_6_entries_ppns_3 = io_refill_bits_ptes[225:202]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_6_entries_ppns_4 = io_refill_bits_ptes[289:266]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_6_entries_ppns_5 = io_refill_bits_ptes[353:330]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_6_entries_ppns_6 = io_refill_bits_ptes[417:394]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_6_entries_ppns_7 = io_refill_bits_ptes[481:458]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_6_entries_vs_0 = ~_wdata_entries_ps_vs_0_T_3 & _wdata_entries_ps_vs_0_T_5; // @[MMUBundle.scala 669:42]
  assign l3_io_wreq_bits_data_6_entries_vs_1 = ~_wdata_entries_ps_vs_1_T_3 & _wdata_entries_ps_vs_1_T_5; // @[MMUBundle.scala 669:42]
  assign l3_io_wreq_bits_data_6_entries_vs_2 = ~_wdata_entries_ps_vs_2_T_3 & _wdata_entries_ps_vs_2_T_5; // @[MMUBundle.scala 669:42]
  assign l3_io_wreq_bits_data_6_entries_vs_3 = ~_wdata_entries_ps_vs_3_T_3 & _wdata_entries_ps_vs_3_T_5; // @[MMUBundle.scala 669:42]
  assign l3_io_wreq_bits_data_6_entries_vs_4 = ~_wdata_entries_ps_vs_4_T_3 & _wdata_entries_ps_vs_4_T_5; // @[MMUBundle.scala 669:42]
  assign l3_io_wreq_bits_data_6_entries_vs_5 = ~_wdata_entries_ps_vs_5_T_3 & _wdata_entries_ps_vs_5_T_5; // @[MMUBundle.scala 669:42]
  assign l3_io_wreq_bits_data_6_entries_vs_6 = ~_wdata_entries_ps_vs_6_T_3 & _wdata_entries_ps_vs_6_T_5; // @[MMUBundle.scala 669:42]
  assign l3_io_wreq_bits_data_6_entries_vs_7 = ~_wdata_entries_ps_vs_7_T_3 & _wdata_entries_ps_vs_7_T_5; // @[MMUBundle.scala 669:42]
  assign l3_io_wreq_bits_data_6_entries_perms_0_d = io_refill_bits_ptes[7]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_6_entries_perms_0_a = io_refill_bits_ptes[6]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_6_entries_perms_0_g = io_refill_bits_ptes[5]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_6_entries_perms_0_u = io_refill_bits_ptes[4]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_6_entries_perms_0_x = io_refill_bits_ptes[3]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_6_entries_perms_0_w = io_refill_bits_ptes[2]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_6_entries_perms_0_r = io_refill_bits_ptes[1]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_6_entries_perms_1_d = io_refill_bits_ptes[71]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_6_entries_perms_1_a = io_refill_bits_ptes[70]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_6_entries_perms_1_g = io_refill_bits_ptes[69]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_6_entries_perms_1_u = io_refill_bits_ptes[68]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_6_entries_perms_1_x = io_refill_bits_ptes[67]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_6_entries_perms_1_w = io_refill_bits_ptes[66]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_6_entries_perms_1_r = io_refill_bits_ptes[65]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_6_entries_perms_2_d = io_refill_bits_ptes[135]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_6_entries_perms_2_a = io_refill_bits_ptes[134]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_6_entries_perms_2_g = io_refill_bits_ptes[133]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_6_entries_perms_2_u = io_refill_bits_ptes[132]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_6_entries_perms_2_x = io_refill_bits_ptes[131]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_6_entries_perms_2_w = io_refill_bits_ptes[130]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_6_entries_perms_2_r = io_refill_bits_ptes[129]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_6_entries_perms_3_d = io_refill_bits_ptes[199]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_6_entries_perms_3_a = io_refill_bits_ptes[198]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_6_entries_perms_3_g = io_refill_bits_ptes[197]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_6_entries_perms_3_u = io_refill_bits_ptes[196]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_6_entries_perms_3_x = io_refill_bits_ptes[195]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_6_entries_perms_3_w = io_refill_bits_ptes[194]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_6_entries_perms_3_r = io_refill_bits_ptes[193]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_6_entries_perms_4_d = io_refill_bits_ptes[263]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_6_entries_perms_4_a = io_refill_bits_ptes[262]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_6_entries_perms_4_g = io_refill_bits_ptes[261]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_6_entries_perms_4_u = io_refill_bits_ptes[260]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_6_entries_perms_4_x = io_refill_bits_ptes[259]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_6_entries_perms_4_w = io_refill_bits_ptes[258]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_6_entries_perms_4_r = io_refill_bits_ptes[257]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_6_entries_perms_5_d = io_refill_bits_ptes[327]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_6_entries_perms_5_a = io_refill_bits_ptes[326]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_6_entries_perms_5_g = io_refill_bits_ptes[325]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_6_entries_perms_5_u = io_refill_bits_ptes[324]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_6_entries_perms_5_x = io_refill_bits_ptes[323]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_6_entries_perms_5_w = io_refill_bits_ptes[322]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_6_entries_perms_5_r = io_refill_bits_ptes[321]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_6_entries_perms_6_d = io_refill_bits_ptes[391]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_6_entries_perms_6_a = io_refill_bits_ptes[390]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_6_entries_perms_6_g = io_refill_bits_ptes[389]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_6_entries_perms_6_u = io_refill_bits_ptes[388]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_6_entries_perms_6_x = io_refill_bits_ptes[387]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_6_entries_perms_6_w = io_refill_bits_ptes[386]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_6_entries_perms_6_r = io_refill_bits_ptes[385]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_6_entries_perms_7_d = io_refill_bits_ptes[455]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_6_entries_perms_7_a = io_refill_bits_ptes[454]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_6_entries_perms_7_g = io_refill_bits_ptes[453]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_6_entries_perms_7_u = io_refill_bits_ptes[452]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_6_entries_perms_7_x = io_refill_bits_ptes[451]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_6_entries_perms_7_w = io_refill_bits_ptes[450]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_6_entries_perms_7_r = io_refill_bits_ptes[449]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_6_entries_prefetch = io_refill_bits_req_info_dup_2_source == 2'h2; // @[MMUConst.scala 254:13]
  assign l3_io_wreq_bits_data_6_ecc = {ecc_unaligned_1,_wdata_ecc_T_2}; // @[Cat.scala 31:58]
  assign l3_io_wreq_bits_data_7_entries_tag = io_refill_bits_req_info_dup_2_vpn[26:5]; // @[MMUBundle.scala 646:8]
  assign l3_io_wreq_bits_data_7_entries_asid = io_csr_dup_2_satp_asid; // @[MMUBundle.scala 662:18 664:13]
  assign l3_io_wreq_bits_data_7_entries_ppns_0 = io_refill_bits_ptes[33:10]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_7_entries_ppns_1 = io_refill_bits_ptes[97:74]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_7_entries_ppns_2 = io_refill_bits_ptes[161:138]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_7_entries_ppns_3 = io_refill_bits_ptes[225:202]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_7_entries_ppns_4 = io_refill_bits_ptes[289:266]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_7_entries_ppns_5 = io_refill_bits_ptes[353:330]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_7_entries_ppns_6 = io_refill_bits_ptes[417:394]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_7_entries_ppns_7 = io_refill_bits_ptes[481:458]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_7_entries_vs_0 = ~_wdata_entries_ps_vs_0_T_3 & _wdata_entries_ps_vs_0_T_5; // @[MMUBundle.scala 669:42]
  assign l3_io_wreq_bits_data_7_entries_vs_1 = ~_wdata_entries_ps_vs_1_T_3 & _wdata_entries_ps_vs_1_T_5; // @[MMUBundle.scala 669:42]
  assign l3_io_wreq_bits_data_7_entries_vs_2 = ~_wdata_entries_ps_vs_2_T_3 & _wdata_entries_ps_vs_2_T_5; // @[MMUBundle.scala 669:42]
  assign l3_io_wreq_bits_data_7_entries_vs_3 = ~_wdata_entries_ps_vs_3_T_3 & _wdata_entries_ps_vs_3_T_5; // @[MMUBundle.scala 669:42]
  assign l3_io_wreq_bits_data_7_entries_vs_4 = ~_wdata_entries_ps_vs_4_T_3 & _wdata_entries_ps_vs_4_T_5; // @[MMUBundle.scala 669:42]
  assign l3_io_wreq_bits_data_7_entries_vs_5 = ~_wdata_entries_ps_vs_5_T_3 & _wdata_entries_ps_vs_5_T_5; // @[MMUBundle.scala 669:42]
  assign l3_io_wreq_bits_data_7_entries_vs_6 = ~_wdata_entries_ps_vs_6_T_3 & _wdata_entries_ps_vs_6_T_5; // @[MMUBundle.scala 669:42]
  assign l3_io_wreq_bits_data_7_entries_vs_7 = ~_wdata_entries_ps_vs_7_T_3 & _wdata_entries_ps_vs_7_T_5; // @[MMUBundle.scala 669:42]
  assign l3_io_wreq_bits_data_7_entries_perms_0_d = io_refill_bits_ptes[7]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_7_entries_perms_0_a = io_refill_bits_ptes[6]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_7_entries_perms_0_g = io_refill_bits_ptes[5]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_7_entries_perms_0_u = io_refill_bits_ptes[4]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_7_entries_perms_0_x = io_refill_bits_ptes[3]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_7_entries_perms_0_w = io_refill_bits_ptes[2]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_7_entries_perms_0_r = io_refill_bits_ptes[1]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_7_entries_perms_1_d = io_refill_bits_ptes[71]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_7_entries_perms_1_a = io_refill_bits_ptes[70]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_7_entries_perms_1_g = io_refill_bits_ptes[69]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_7_entries_perms_1_u = io_refill_bits_ptes[68]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_7_entries_perms_1_x = io_refill_bits_ptes[67]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_7_entries_perms_1_w = io_refill_bits_ptes[66]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_7_entries_perms_1_r = io_refill_bits_ptes[65]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_7_entries_perms_2_d = io_refill_bits_ptes[135]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_7_entries_perms_2_a = io_refill_bits_ptes[134]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_7_entries_perms_2_g = io_refill_bits_ptes[133]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_7_entries_perms_2_u = io_refill_bits_ptes[132]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_7_entries_perms_2_x = io_refill_bits_ptes[131]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_7_entries_perms_2_w = io_refill_bits_ptes[130]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_7_entries_perms_2_r = io_refill_bits_ptes[129]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_7_entries_perms_3_d = io_refill_bits_ptes[199]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_7_entries_perms_3_a = io_refill_bits_ptes[198]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_7_entries_perms_3_g = io_refill_bits_ptes[197]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_7_entries_perms_3_u = io_refill_bits_ptes[196]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_7_entries_perms_3_x = io_refill_bits_ptes[195]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_7_entries_perms_3_w = io_refill_bits_ptes[194]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_7_entries_perms_3_r = io_refill_bits_ptes[193]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_7_entries_perms_4_d = io_refill_bits_ptes[263]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_7_entries_perms_4_a = io_refill_bits_ptes[262]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_7_entries_perms_4_g = io_refill_bits_ptes[261]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_7_entries_perms_4_u = io_refill_bits_ptes[260]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_7_entries_perms_4_x = io_refill_bits_ptes[259]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_7_entries_perms_4_w = io_refill_bits_ptes[258]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_7_entries_perms_4_r = io_refill_bits_ptes[257]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_7_entries_perms_5_d = io_refill_bits_ptes[327]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_7_entries_perms_5_a = io_refill_bits_ptes[326]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_7_entries_perms_5_g = io_refill_bits_ptes[325]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_7_entries_perms_5_u = io_refill_bits_ptes[324]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_7_entries_perms_5_x = io_refill_bits_ptes[323]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_7_entries_perms_5_w = io_refill_bits_ptes[322]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_7_entries_perms_5_r = io_refill_bits_ptes[321]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_7_entries_perms_6_d = io_refill_bits_ptes[391]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_7_entries_perms_6_a = io_refill_bits_ptes[390]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_7_entries_perms_6_g = io_refill_bits_ptes[389]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_7_entries_perms_6_u = io_refill_bits_ptes[388]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_7_entries_perms_6_x = io_refill_bits_ptes[387]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_7_entries_perms_6_w = io_refill_bits_ptes[386]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_7_entries_perms_6_r = io_refill_bits_ptes[385]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_7_entries_perms_7_d = io_refill_bits_ptes[455]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_7_entries_perms_7_a = io_refill_bits_ptes[454]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_7_entries_perms_7_g = io_refill_bits_ptes[453]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_7_entries_perms_7_u = io_refill_bits_ptes[452]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_7_entries_perms_7_x = io_refill_bits_ptes[451]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_7_entries_perms_7_w = io_refill_bits_ptes[450]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_7_entries_perms_7_r = io_refill_bits_ptes[449]; // @[MMUBundle.scala 667:52]
  assign l3_io_wreq_bits_data_7_entries_prefetch = io_refill_bits_req_info_dup_2_source == 2'h2; // @[MMUConst.scala 254:13]
  assign l3_io_wreq_bits_data_7_ecc = {ecc_unaligned_1,_wdata_ecc_T_2}; // @[Cat.scala 31:58]
  assign l3_io_wreq_bits_waymask = 8'h1 << l3_victimWay; // @[OneHot.scala 57:35]
  always @(posedge clock) begin
    if (leftFire) begin // @[Reg.scala 17:18]
      data_req_info_vpn <= io_req_bits_req_info_vpn; // @[Reg.scala 17:22]
    end
    if (leftFire) begin // @[Reg.scala 17:18]
      data_req_info_source <= io_req_bits_req_info_source; // @[Reg.scala 17:22]
    end
    if (leftFire) begin // @[Reg.scala 17:18]
      data_isFirst <= io_req_bits_isFirst; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[PageTableCache.scala 659:21]
      bypassed_reg <= bypassed_wire; // @[PageTableCache.scala 659:36]
    end else if (io_refill_valid) begin // @[PageTableCache.scala 660:35]
      bypassed_reg <= bypassed_reg | bypassed_wire; // @[PageTableCache.scala 660:50]
    end
    if (stageDelay_valid_1cycle) begin // @[PageTableCache.scala 659:21]
      bypassed_reg_1 <= bypassed_wire_1; // @[PageTableCache.scala 659:36]
    end else if (io_refill_valid) begin // @[PageTableCache.scala 660:35]
      bypassed_reg_1 <= bypassed_reg_1 | bypassed_wire_1; // @[PageTableCache.scala 660:50]
    end
    if (stageDelay_valid_1cycle) begin // @[PageTableCache.scala 659:21]
      bypassed_reg_2 <= bypassed_wire_2; // @[PageTableCache.scala 659:36]
    end else if (io_refill_valid) begin // @[PageTableCache.scala 660:35]
      bypassed_reg_2 <= bypassed_reg_2 | bypassed_wire_2; // @[PageTableCache.scala 660:50]
    end
    if (leftFire_1) begin // @[Reg.scala 17:18]
      data_1_req_info_vpn <= data_req_info_vpn; // @[Reg.scala 17:22]
    end
    if (leftFire_1) begin // @[Reg.scala 17:18]
      data_1_req_info_source <= data_req_info_source; // @[Reg.scala 17:22]
    end
    if (leftFire_1) begin // @[Reg.scala 17:18]
      data_1_isFirst <= data_isFirst; // @[Reg.scala 17:22]
    end
    if (leftFire_1) begin // @[Reg.scala 17:18]
      data_1_bypassed_0 <= stageDelay_1_bits_bypassed_0; // @[Reg.scala 17:22]
    end
    if (leftFire_1) begin // @[Reg.scala 17:18]
      data_1_bypassed_1 <= stageDelay_1_bits_bypassed_1; // @[Reg.scala 17:22]
    end
    if (leftFire_1) begin // @[Reg.scala 17:18]
      data_1_bypassed_2 <= stageDelay_1_bits_bypassed_2; // @[Reg.scala 17:22]
    end
    if (stageCheck_valid_1cycle) begin // @[PageTableCache.scala 659:21]
      bypassed_reg_3 <= bypassed_wire_3; // @[PageTableCache.scala 659:36]
    end else if (io_refill_valid) begin // @[PageTableCache.scala 660:35]
      bypassed_reg_3 <= bypassed_reg_3 | bypassed_wire_3; // @[PageTableCache.scala 660:50]
    end
    if (stageCheck_valid_1cycle) begin // @[PageTableCache.scala 659:21]
      bypassed_reg_4 <= bypassed_wire_4; // @[PageTableCache.scala 659:36]
    end else if (io_refill_valid) begin // @[PageTableCache.scala 660:35]
      bypassed_reg_4 <= bypassed_reg_4 | bypassed_wire_4; // @[PageTableCache.scala 660:50]
    end
    if (stageCheck_valid_1cycle) begin // @[PageTableCache.scala 659:21]
      bypassed_reg_5 <= bypassed_wire_5; // @[PageTableCache.scala 659:36]
    end else if (io_refill_valid) begin // @[PageTableCache.scala 660:35]
      bypassed_reg_5 <= bypassed_reg_5 | bypassed_wire_5; // @[PageTableCache.scala 660:50]
    end
    if (leftFire_2) begin // @[Reg.scala 17:18]
      data_2_req_info_vpn <= data_1_req_info_vpn; // @[Reg.scala 17:22]
    end
    if (leftFire_2) begin // @[Reg.scala 17:18]
      data_2_req_info_source <= data_1_req_info_source; // @[Reg.scala 17:22]
    end
    if (leftFire_2) begin // @[Reg.scala 17:18]
      data_2_isFirst <= data_1_isFirst; // @[Reg.scala 17:22]
    end
    if (leftFire_2) begin // @[Reg.scala 17:18]
      data_2_bypassed_0 <= stageCheck_1_bits_bypassed_0; // @[Reg.scala 17:22]
    end
    if (leftFire_2) begin // @[Reg.scala 17:18]
      data_2_bypassed_1 <= stageCheck_1_bits_bypassed_1; // @[Reg.scala 17:22]
    end
    if (leftFire_2) begin // @[Reg.scala 17:18]
      data_2_bypassed_2 <= stageCheck_1_bits_bypassed_2; // @[Reg.scala 17:22]
    end
    if (~flush & io_refill_bits_levelOH_l1 & ~_T_299 & ~_T_321 & ~_T_325) begin // @[PageTableCache.scala 435:129]
      if (2'h0 == PtwL1RefillIdx) begin // @[MMUBundle.scala 599:9]
        l1_0_tag <= io_refill_bits_req_info_dup_0_vpn[26:18]; // @[MMUBundle.scala 599:9]
      end
    end
    if (~flush & io_refill_bits_levelOH_l1 & ~_T_299 & ~_T_321 & ~_T_325) begin // @[PageTableCache.scala 435:129]
      if (2'h0 == PtwL1RefillIdx) begin // @[MMUBundle.scala 602:15]
        l1_0_asid <= io_csr_dup_0_satp_asid; // @[MMUBundle.scala 602:15]
      end
    end
    if (~flush & io_refill_bits_levelOH_l1 & ~_T_299 & ~_T_321 & ~_T_325) begin // @[PageTableCache.scala 435:129]
      if (2'h0 == PtwL1RefillIdx) begin // @[MMUBundle.scala 600:9]
        l1_0_ppn <= memPte_0_ppn; // @[MMUBundle.scala 600:9]
      end
    end
    if (~flush & io_refill_bits_levelOH_l1 & ~_T_299 & ~_T_321 & ~_T_325) begin // @[PageTableCache.scala 435:129]
      if (2'h1 == PtwL1RefillIdx) begin // @[MMUBundle.scala 599:9]
        l1_1_tag <= io_refill_bits_req_info_dup_0_vpn[26:18]; // @[MMUBundle.scala 599:9]
      end
    end
    if (~flush & io_refill_bits_levelOH_l1 & ~_T_299 & ~_T_321 & ~_T_325) begin // @[PageTableCache.scala 435:129]
      if (2'h1 == PtwL1RefillIdx) begin // @[MMUBundle.scala 602:15]
        l1_1_asid <= io_csr_dup_0_satp_asid; // @[MMUBundle.scala 602:15]
      end
    end
    if (~flush & io_refill_bits_levelOH_l1 & ~_T_299 & ~_T_321 & ~_T_325) begin // @[PageTableCache.scala 435:129]
      if (2'h1 == PtwL1RefillIdx) begin // @[MMUBundle.scala 600:9]
        l1_1_ppn <= memPte_0_ppn; // @[MMUBundle.scala 600:9]
      end
    end
    if (~flush & io_refill_bits_levelOH_l1 & ~_T_299 & ~_T_321 & ~_T_325) begin // @[PageTableCache.scala 435:129]
      if (2'h2 == PtwL1RefillIdx) begin // @[MMUBundle.scala 599:9]
        l1_2_tag <= io_refill_bits_req_info_dup_0_vpn[26:18]; // @[MMUBundle.scala 599:9]
      end
    end
    if (~flush & io_refill_bits_levelOH_l1 & ~_T_299 & ~_T_321 & ~_T_325) begin // @[PageTableCache.scala 435:129]
      if (2'h2 == PtwL1RefillIdx) begin // @[MMUBundle.scala 602:15]
        l1_2_asid <= io_csr_dup_0_satp_asid; // @[MMUBundle.scala 602:15]
      end
    end
    if (~flush & io_refill_bits_levelOH_l1 & ~_T_299 & ~_T_321 & ~_T_325) begin // @[PageTableCache.scala 435:129]
      if (2'h2 == PtwL1RefillIdx) begin // @[MMUBundle.scala 600:9]
        l1_2_ppn <= memPte_0_ppn; // @[MMUBundle.scala 600:9]
      end
    end
    if (~flush & io_refill_bits_levelOH_l1 & ~_T_299 & ~_T_321 & ~_T_325) begin // @[PageTableCache.scala 435:129]
      if (2'h3 == PtwL1RefillIdx) begin // @[MMUBundle.scala 599:9]
        l1_3_tag <= io_refill_bits_req_info_dup_0_vpn[26:18]; // @[MMUBundle.scala 599:9]
      end
    end
    if (~flush & io_refill_bits_levelOH_l1 & ~_T_299 & ~_T_321 & ~_T_325) begin // @[PageTableCache.scala 435:129]
      if (2'h3 == PtwL1RefillIdx) begin // @[MMUBundle.scala 602:15]
        l1_3_asid <= io_csr_dup_0_satp_asid; // @[MMUBundle.scala 602:15]
      end
    end
    if (~flush & io_refill_bits_levelOH_l1 & ~_T_299 & ~_T_321 & ~_T_325) begin // @[PageTableCache.scala 435:129]
      if (2'h3 == PtwL1RefillIdx) begin // @[MMUBundle.scala 600:9]
        l1_3_ppn <= memPte_0_ppn; // @[MMUBundle.scala 600:9]
      end
    end
    if (~flush & io_refill_bits_levelOH_l1 & ~_T_299 & ~_T_321 & ~_T_325) begin // @[PageTableCache.scala 435:129]
      l1g <= _l1g_T_3; // @[PageTableCache.scala 449:9]
    end
    if (l2eccFlush) begin // @[PageTableCache.scala 572:21]
      l2g <= _l2g_T_7; // @[PageTableCache.scala 576:9]
    end else if (~flush_dup_1 & io_refill_bits_levelOH_l2 & ~_T_336 & ~_T_358 & ~_T_362) begin // @[PageTableCache.scala 462:129]
      l2g <= _l2g_T_5; // @[PageTableCache.scala 483:9]
    end
    if (l3eccFlush) begin // @[PageTableCache.scala 579:21]
      l3g <= _l3g_T_7; // @[PageTableCache.scala 583:9]
    end else if (~flush_dup_2 & io_refill_bits_levelOH_l3 & ~_T_377) begin // @[PageTableCache.scala 500:66]
      l3g <= _l3g_T_5; // @[PageTableCache.scala 521:9]
    end
    if (_T_296 & io_refill_bits_levelOH_sp & (_T_299 | _T_321) & _T_326) begin // @[PageTableCache.scala 540:129]
      if (~state_reg_3) begin // @[MMUBundle.scala 599:9]
        sp_0_tag <= io_refill_bits_req_info_dup_0_vpn[26:9]; // @[MMUBundle.scala 599:9]
      end
    end
    if (_T_296 & io_refill_bits_levelOH_sp & (_T_299 | _T_321) & _T_326) begin // @[PageTableCache.scala 540:129]
      if (~state_reg_3) begin // @[MMUBundle.scala 602:15]
        sp_0_asid <= io_csr_dup_0_satp_asid; // @[MMUBundle.scala 602:15]
      end
    end
    if (_T_296 & io_refill_bits_levelOH_sp & (_T_299 | _T_321) & _T_326) begin // @[PageTableCache.scala 540:129]
      if (~state_reg_3) begin // @[MMUBundle.scala 600:9]
        sp_0_ppn <= memPte_0_ppn; // @[MMUBundle.scala 600:9]
      end
    end
    if (_T_296 & io_refill_bits_levelOH_sp & (_T_299 | _T_321) & _T_326) begin // @[PageTableCache.scala 540:129]
      if (~state_reg_3) begin // @[MMUBundle.scala 601:16]
        sp_0_perm_d <= memPte_0_perm_d; // @[MMUBundle.scala 601:16]
      end
    end
    if (_T_296 & io_refill_bits_levelOH_sp & (_T_299 | _T_321) & _T_326) begin // @[PageTableCache.scala 540:129]
      if (~state_reg_3) begin // @[MMUBundle.scala 601:16]
        sp_0_perm_a <= memPte_0_perm_a; // @[MMUBundle.scala 601:16]
      end
    end
    if (_T_296 & io_refill_bits_levelOH_sp & (_T_299 | _T_321) & _T_326) begin // @[PageTableCache.scala 540:129]
      if (~state_reg_3) begin // @[MMUBundle.scala 601:16]
        sp_0_perm_g <= memPte_0_perm_g; // @[MMUBundle.scala 601:16]
      end
    end
    if (_T_296 & io_refill_bits_levelOH_sp & (_T_299 | _T_321) & _T_326) begin // @[PageTableCache.scala 540:129]
      if (~state_reg_3) begin // @[MMUBundle.scala 601:16]
        sp_0_perm_u <= memPte_0_perm_u; // @[MMUBundle.scala 601:16]
      end
    end
    if (_T_296 & io_refill_bits_levelOH_sp & (_T_299 | _T_321) & _T_326) begin // @[PageTableCache.scala 540:129]
      if (~state_reg_3) begin // @[MMUBundle.scala 601:16]
        sp_0_perm_x <= memPte_0_perm_x; // @[MMUBundle.scala 601:16]
      end
    end
    if (_T_296 & io_refill_bits_levelOH_sp & (_T_299 | _T_321) & _T_326) begin // @[PageTableCache.scala 540:129]
      if (~state_reg_3) begin // @[MMUBundle.scala 601:16]
        sp_0_perm_w <= memPte_0_perm_w; // @[MMUBundle.scala 601:16]
      end
    end
    if (_T_296 & io_refill_bits_levelOH_sp & (_T_299 | _T_321) & _T_326) begin // @[PageTableCache.scala 540:129]
      if (~state_reg_3) begin // @[MMUBundle.scala 601:16]
        sp_0_perm_r <= memPte_0_perm_r; // @[MMUBundle.scala 601:16]
      end
    end
    if (_T_296 & io_refill_bits_levelOH_sp & (_T_299 | _T_321) & _T_326) begin // @[PageTableCache.scala 540:129]
      if (~state_reg_3) begin // @[MMUBundle.scala 605:22]
        sp_0_level <= io_refill_bits_level_dup_2; // @[MMUBundle.scala 605:22]
      end
    end
    if (_T_296 & io_refill_bits_levelOH_sp & (_T_299 | _T_321) & _T_326) begin // @[PageTableCache.scala 540:129]
      if (~state_reg_3) begin // @[MMUBundle.scala 603:19]
        sp_0_prefetch <= refill_prefetch_dup_0; // @[MMUBundle.scala 603:19]
      end
    end
    if (_T_296 & io_refill_bits_levelOH_sp & (_T_299 | _T_321) & _T_326) begin // @[PageTableCache.scala 540:129]
      if (~state_reg_3) begin // @[MMUBundle.scala 604:12]
        sp_0_v <= _T_322; // @[MMUBundle.scala 604:12]
      end
    end
    if (_T_296 & io_refill_bits_levelOH_sp & (_T_299 | _T_321) & _T_326) begin // @[PageTableCache.scala 540:129]
      if (state_reg_3) begin // @[MMUBundle.scala 599:9]
        sp_1_tag <= io_refill_bits_req_info_dup_0_vpn[26:9]; // @[MMUBundle.scala 599:9]
      end
    end
    if (_T_296 & io_refill_bits_levelOH_sp & (_T_299 | _T_321) & _T_326) begin // @[PageTableCache.scala 540:129]
      if (state_reg_3) begin // @[MMUBundle.scala 602:15]
        sp_1_asid <= io_csr_dup_0_satp_asid; // @[MMUBundle.scala 602:15]
      end
    end
    if (_T_296 & io_refill_bits_levelOH_sp & (_T_299 | _T_321) & _T_326) begin // @[PageTableCache.scala 540:129]
      if (state_reg_3) begin // @[MMUBundle.scala 600:9]
        sp_1_ppn <= memPte_0_ppn; // @[MMUBundle.scala 600:9]
      end
    end
    if (_T_296 & io_refill_bits_levelOH_sp & (_T_299 | _T_321) & _T_326) begin // @[PageTableCache.scala 540:129]
      if (state_reg_3) begin // @[MMUBundle.scala 601:16]
        sp_1_perm_d <= memPte_0_perm_d; // @[MMUBundle.scala 601:16]
      end
    end
    if (_T_296 & io_refill_bits_levelOH_sp & (_T_299 | _T_321) & _T_326) begin // @[PageTableCache.scala 540:129]
      if (state_reg_3) begin // @[MMUBundle.scala 601:16]
        sp_1_perm_a <= memPte_0_perm_a; // @[MMUBundle.scala 601:16]
      end
    end
    if (_T_296 & io_refill_bits_levelOH_sp & (_T_299 | _T_321) & _T_326) begin // @[PageTableCache.scala 540:129]
      if (state_reg_3) begin // @[MMUBundle.scala 601:16]
        sp_1_perm_g <= memPte_0_perm_g; // @[MMUBundle.scala 601:16]
      end
    end
    if (_T_296 & io_refill_bits_levelOH_sp & (_T_299 | _T_321) & _T_326) begin // @[PageTableCache.scala 540:129]
      if (state_reg_3) begin // @[MMUBundle.scala 601:16]
        sp_1_perm_u <= memPte_0_perm_u; // @[MMUBundle.scala 601:16]
      end
    end
    if (_T_296 & io_refill_bits_levelOH_sp & (_T_299 | _T_321) & _T_326) begin // @[PageTableCache.scala 540:129]
      if (state_reg_3) begin // @[MMUBundle.scala 601:16]
        sp_1_perm_x <= memPte_0_perm_x; // @[MMUBundle.scala 601:16]
      end
    end
    if (_T_296 & io_refill_bits_levelOH_sp & (_T_299 | _T_321) & _T_326) begin // @[PageTableCache.scala 540:129]
      if (state_reg_3) begin // @[MMUBundle.scala 601:16]
        sp_1_perm_w <= memPte_0_perm_w; // @[MMUBundle.scala 601:16]
      end
    end
    if (_T_296 & io_refill_bits_levelOH_sp & (_T_299 | _T_321) & _T_326) begin // @[PageTableCache.scala 540:129]
      if (state_reg_3) begin // @[MMUBundle.scala 601:16]
        sp_1_perm_r <= memPte_0_perm_r; // @[MMUBundle.scala 601:16]
      end
    end
    if (_T_296 & io_refill_bits_levelOH_sp & (_T_299 | _T_321) & _T_326) begin // @[PageTableCache.scala 540:129]
      if (state_reg_3) begin // @[MMUBundle.scala 605:22]
        sp_1_level <= io_refill_bits_level_dup_2; // @[MMUBundle.scala 605:22]
      end
    end
    if (_T_296 & io_refill_bits_levelOH_sp & (_T_299 | _T_321) & _T_326) begin // @[PageTableCache.scala 540:129]
      if (state_reg_3) begin // @[MMUBundle.scala 603:19]
        sp_1_prefetch <= refill_prefetch_dup_0; // @[MMUBundle.scala 603:19]
      end
    end
    if (_T_296 & io_refill_bits_levelOH_sp & (_T_299 | _T_321) & _T_326) begin // @[PageTableCache.scala 540:129]
      if (state_reg_3) begin // @[MMUBundle.scala 604:12]
        sp_1_v <= _T_322; // @[MMUBundle.scala 604:12]
      end
    end
    if (_T_296 & io_refill_bits_levelOH_sp & (_T_299 | _T_321) & _T_326) begin // @[PageTableCache.scala 540:129]
      spg <= _spg_T_3; // @[PageTableCache.scala 553:9]
    end
    if (_stageDelay_valid_1cycle_T) begin // @[Reg.scala 17:18]
      r <= l1_hitVecT_0; // @[Reg.scala 17:22]
    end
    if (_stageDelay_valid_1cycle_T) begin // @[Reg.scala 17:18]
      r_1 <= l1_hitVecT_1; // @[Reg.scala 17:22]
    end
    if (_stageDelay_valid_1cycle_T) begin // @[Reg.scala 17:18]
      r_2 <= l1_hitVecT_2; // @[Reg.scala 17:22]
    end
    if (_stageDelay_valid_1cycle_T) begin // @[Reg.scala 17:18]
      r_3 <= l1_hitVecT_3; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      if (r | r_1) begin // @[ParallelMux.scala 90:77]
        if (r) begin // @[ParallelMux.scala 90:77]
          r_4 <= l1_0_ppn;
        end else begin
          r_4 <= l1_1_ppn;
        end
      end else if (r_2) begin // @[ParallelMux.scala 90:77]
        r_4 <= l1_2_ppn;
      end else begin
        r_4 <= l1_3_ppn;
      end
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_6 <= _T_28; // @[Reg.scala 17:22]
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l1Hit <= _T_28; // @[Reg.scala 17:22]
      end else begin
        l1Hit <= r_6; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        if (r | r_1) begin // @[ParallelMux.scala 90:77]
          if (r) begin // @[ParallelMux.scala 90:77]
            l1HitPPN <= l1_0_ppn;
          end else begin
            l1HitPPN <= l1_1_ppn;
          end
        end else if (r_2) begin // @[ParallelMux.scala 90:77]
          l1HitPPN <= l1_2_ppn;
        end else begin
          l1HitPPN <= l1_3_ppn;
        end
      end else begin
        l1HitPPN <= r_4; // @[Reg.scala 16:16]
      end
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_0_entries_tag <= l2_io_rresp_data_0_entries_tag; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_0_entries_asid <= l2_io_rresp_data_0_entries_asid; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_0_entries_ppns_0 <= l2_io_rresp_data_0_entries_ppns_0; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_0_entries_ppns_1 <= l2_io_rresp_data_0_entries_ppns_1; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_0_entries_ppns_2 <= l2_io_rresp_data_0_entries_ppns_2; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_0_entries_ppns_3 <= l2_io_rresp_data_0_entries_ppns_3; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_0_entries_ppns_4 <= l2_io_rresp_data_0_entries_ppns_4; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_0_entries_ppns_5 <= l2_io_rresp_data_0_entries_ppns_5; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_0_entries_ppns_6 <= l2_io_rresp_data_0_entries_ppns_6; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_0_entries_ppns_7 <= l2_io_rresp_data_0_entries_ppns_7; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_0_entries_vs_0 <= l2_io_rresp_data_0_entries_vs_0; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_0_entries_vs_1 <= l2_io_rresp_data_0_entries_vs_1; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_0_entries_vs_2 <= l2_io_rresp_data_0_entries_vs_2; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_0_entries_vs_3 <= l2_io_rresp_data_0_entries_vs_3; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_0_entries_vs_4 <= l2_io_rresp_data_0_entries_vs_4; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_0_entries_vs_5 <= l2_io_rresp_data_0_entries_vs_5; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_0_entries_vs_6 <= l2_io_rresp_data_0_entries_vs_6; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_0_entries_vs_7 <= l2_io_rresp_data_0_entries_vs_7; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_0_entries_prefetch <= l2_io_rresp_data_0_entries_prefetch; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_0_ecc <= l2_io_rresp_data_0_ecc; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_1_entries_tag <= l2_io_rresp_data_1_entries_tag; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_1_entries_asid <= l2_io_rresp_data_1_entries_asid; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_1_entries_ppns_0 <= l2_io_rresp_data_1_entries_ppns_0; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_1_entries_ppns_1 <= l2_io_rresp_data_1_entries_ppns_1; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_1_entries_ppns_2 <= l2_io_rresp_data_1_entries_ppns_2; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_1_entries_ppns_3 <= l2_io_rresp_data_1_entries_ppns_3; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_1_entries_ppns_4 <= l2_io_rresp_data_1_entries_ppns_4; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_1_entries_ppns_5 <= l2_io_rresp_data_1_entries_ppns_5; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_1_entries_ppns_6 <= l2_io_rresp_data_1_entries_ppns_6; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_1_entries_ppns_7 <= l2_io_rresp_data_1_entries_ppns_7; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_1_entries_vs_0 <= l2_io_rresp_data_1_entries_vs_0; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_1_entries_vs_1 <= l2_io_rresp_data_1_entries_vs_1; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_1_entries_vs_2 <= l2_io_rresp_data_1_entries_vs_2; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_1_entries_vs_3 <= l2_io_rresp_data_1_entries_vs_3; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_1_entries_vs_4 <= l2_io_rresp_data_1_entries_vs_4; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_1_entries_vs_5 <= l2_io_rresp_data_1_entries_vs_5; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_1_entries_vs_6 <= l2_io_rresp_data_1_entries_vs_6; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_1_entries_vs_7 <= l2_io_rresp_data_1_entries_vs_7; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_1_entries_prefetch <= l2_io_rresp_data_1_entries_prefetch; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_1_ecc <= l2_io_rresp_data_1_ecc; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_2_entries_tag <= l2_io_rresp_data_2_entries_tag; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_2_entries_asid <= l2_io_rresp_data_2_entries_asid; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_2_entries_ppns_0 <= l2_io_rresp_data_2_entries_ppns_0; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_2_entries_ppns_1 <= l2_io_rresp_data_2_entries_ppns_1; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_2_entries_ppns_2 <= l2_io_rresp_data_2_entries_ppns_2; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_2_entries_ppns_3 <= l2_io_rresp_data_2_entries_ppns_3; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_2_entries_ppns_4 <= l2_io_rresp_data_2_entries_ppns_4; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_2_entries_ppns_5 <= l2_io_rresp_data_2_entries_ppns_5; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_2_entries_ppns_6 <= l2_io_rresp_data_2_entries_ppns_6; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_2_entries_ppns_7 <= l2_io_rresp_data_2_entries_ppns_7; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_2_entries_vs_0 <= l2_io_rresp_data_2_entries_vs_0; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_2_entries_vs_1 <= l2_io_rresp_data_2_entries_vs_1; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_2_entries_vs_2 <= l2_io_rresp_data_2_entries_vs_2; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_2_entries_vs_3 <= l2_io_rresp_data_2_entries_vs_3; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_2_entries_vs_4 <= l2_io_rresp_data_2_entries_vs_4; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_2_entries_vs_5 <= l2_io_rresp_data_2_entries_vs_5; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_2_entries_vs_6 <= l2_io_rresp_data_2_entries_vs_6; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_2_entries_vs_7 <= l2_io_rresp_data_2_entries_vs_7; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_2_entries_prefetch <= l2_io_rresp_data_2_entries_prefetch; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_2_ecc <= l2_io_rresp_data_2_ecc; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_3_entries_tag <= l2_io_rresp_data_3_entries_tag; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_3_entries_asid <= l2_io_rresp_data_3_entries_asid; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_3_entries_ppns_0 <= l2_io_rresp_data_3_entries_ppns_0; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_3_entries_ppns_1 <= l2_io_rresp_data_3_entries_ppns_1; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_3_entries_ppns_2 <= l2_io_rresp_data_3_entries_ppns_2; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_3_entries_ppns_3 <= l2_io_rresp_data_3_entries_ppns_3; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_3_entries_ppns_4 <= l2_io_rresp_data_3_entries_ppns_4; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_3_entries_ppns_5 <= l2_io_rresp_data_3_entries_ppns_5; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_3_entries_ppns_6 <= l2_io_rresp_data_3_entries_ppns_6; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_3_entries_ppns_7 <= l2_io_rresp_data_3_entries_ppns_7; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_3_entries_vs_0 <= l2_io_rresp_data_3_entries_vs_0; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_3_entries_vs_1 <= l2_io_rresp_data_3_entries_vs_1; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_3_entries_vs_2 <= l2_io_rresp_data_3_entries_vs_2; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_3_entries_vs_3 <= l2_io_rresp_data_3_entries_vs_3; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_3_entries_vs_4 <= l2_io_rresp_data_3_entries_vs_4; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_3_entries_vs_5 <= l2_io_rresp_data_3_entries_vs_5; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_3_entries_vs_6 <= l2_io_rresp_data_3_entries_vs_6; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_3_entries_vs_7 <= l2_io_rresp_data_3_entries_vs_7; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_3_entries_prefetch <= l2_io_rresp_data_3_entries_prefetch; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_7_3_ecc <= l2_io_rresp_data_3_ecc; // @[Reg.scala 17:22]
    end
    if (_stageDelay_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (2'h3 == l2_ridx) begin // @[Reg.scala 17:22]
        r_8 <= l2vVec_3; // @[Reg.scala 17:22]
      end else if (2'h2 == l2_ridx) begin // @[Reg.scala 17:22]
        r_8 <= l2vVec_2; // @[Reg.scala 17:22]
      end else if (2'h1 == l2_ridx) begin // @[Reg.scala 17:22]
        r_8 <= l2vVec_1; // @[Reg.scala 17:22]
      end else begin
        r_8 <= l2vVec_0;
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_0_entries_tag <= l2_io_rresp_data_0_entries_tag; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_0_entries_tag <= r_7_0_entries_tag; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_0_entries_asid <= l2_io_rresp_data_0_entries_asid; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_0_entries_asid <= r_7_0_entries_asid; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_0_entries_ppns_0 <= l2_io_rresp_data_0_entries_ppns_0; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_0_entries_ppns_0 <= r_7_0_entries_ppns_0; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_0_entries_ppns_1 <= l2_io_rresp_data_0_entries_ppns_1; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_0_entries_ppns_1 <= r_7_0_entries_ppns_1; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_0_entries_ppns_2 <= l2_io_rresp_data_0_entries_ppns_2; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_0_entries_ppns_2 <= r_7_0_entries_ppns_2; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_0_entries_ppns_3 <= l2_io_rresp_data_0_entries_ppns_3; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_0_entries_ppns_3 <= r_7_0_entries_ppns_3; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_0_entries_ppns_4 <= l2_io_rresp_data_0_entries_ppns_4; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_0_entries_ppns_4 <= r_7_0_entries_ppns_4; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_0_entries_ppns_5 <= l2_io_rresp_data_0_entries_ppns_5; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_0_entries_ppns_5 <= r_7_0_entries_ppns_5; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_0_entries_ppns_6 <= l2_io_rresp_data_0_entries_ppns_6; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_0_entries_ppns_6 <= r_7_0_entries_ppns_6; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_0_entries_ppns_7 <= l2_io_rresp_data_0_entries_ppns_7; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_0_entries_ppns_7 <= r_7_0_entries_ppns_7; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_0_entries_vs_0 <= l2_io_rresp_data_0_entries_vs_0; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_0_entries_vs_0 <= r_7_0_entries_vs_0; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_0_entries_vs_1 <= l2_io_rresp_data_0_entries_vs_1; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_0_entries_vs_1 <= r_7_0_entries_vs_1; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_0_entries_vs_2 <= l2_io_rresp_data_0_entries_vs_2; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_0_entries_vs_2 <= r_7_0_entries_vs_2; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_0_entries_vs_3 <= l2_io_rresp_data_0_entries_vs_3; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_0_entries_vs_3 <= r_7_0_entries_vs_3; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_0_entries_vs_4 <= l2_io_rresp_data_0_entries_vs_4; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_0_entries_vs_4 <= r_7_0_entries_vs_4; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_0_entries_vs_5 <= l2_io_rresp_data_0_entries_vs_5; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_0_entries_vs_5 <= r_7_0_entries_vs_5; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_0_entries_vs_6 <= l2_io_rresp_data_0_entries_vs_6; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_0_entries_vs_6 <= r_7_0_entries_vs_6; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_0_entries_vs_7 <= l2_io_rresp_data_0_entries_vs_7; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_0_entries_vs_7 <= r_7_0_entries_vs_7; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_0_entries_prefetch <= l2_io_rresp_data_0_entries_prefetch; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_0_entries_prefetch <= r_7_0_entries_prefetch; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_0_ecc <= l2_io_rresp_data_0_ecc; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_0_ecc <= r_7_0_ecc; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_1_entries_tag <= l2_io_rresp_data_1_entries_tag; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_1_entries_tag <= r_7_1_entries_tag; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_1_entries_asid <= l2_io_rresp_data_1_entries_asid; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_1_entries_asid <= r_7_1_entries_asid; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_1_entries_ppns_0 <= l2_io_rresp_data_1_entries_ppns_0; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_1_entries_ppns_0 <= r_7_1_entries_ppns_0; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_1_entries_ppns_1 <= l2_io_rresp_data_1_entries_ppns_1; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_1_entries_ppns_1 <= r_7_1_entries_ppns_1; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_1_entries_ppns_2 <= l2_io_rresp_data_1_entries_ppns_2; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_1_entries_ppns_2 <= r_7_1_entries_ppns_2; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_1_entries_ppns_3 <= l2_io_rresp_data_1_entries_ppns_3; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_1_entries_ppns_3 <= r_7_1_entries_ppns_3; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_1_entries_ppns_4 <= l2_io_rresp_data_1_entries_ppns_4; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_1_entries_ppns_4 <= r_7_1_entries_ppns_4; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_1_entries_ppns_5 <= l2_io_rresp_data_1_entries_ppns_5; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_1_entries_ppns_5 <= r_7_1_entries_ppns_5; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_1_entries_ppns_6 <= l2_io_rresp_data_1_entries_ppns_6; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_1_entries_ppns_6 <= r_7_1_entries_ppns_6; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_1_entries_ppns_7 <= l2_io_rresp_data_1_entries_ppns_7; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_1_entries_ppns_7 <= r_7_1_entries_ppns_7; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_1_entries_vs_0 <= l2_io_rresp_data_1_entries_vs_0; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_1_entries_vs_0 <= r_7_1_entries_vs_0; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_1_entries_vs_1 <= l2_io_rresp_data_1_entries_vs_1; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_1_entries_vs_1 <= r_7_1_entries_vs_1; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_1_entries_vs_2 <= l2_io_rresp_data_1_entries_vs_2; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_1_entries_vs_2 <= r_7_1_entries_vs_2; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_1_entries_vs_3 <= l2_io_rresp_data_1_entries_vs_3; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_1_entries_vs_3 <= r_7_1_entries_vs_3; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_1_entries_vs_4 <= l2_io_rresp_data_1_entries_vs_4; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_1_entries_vs_4 <= r_7_1_entries_vs_4; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_1_entries_vs_5 <= l2_io_rresp_data_1_entries_vs_5; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_1_entries_vs_5 <= r_7_1_entries_vs_5; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_1_entries_vs_6 <= l2_io_rresp_data_1_entries_vs_6; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_1_entries_vs_6 <= r_7_1_entries_vs_6; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_1_entries_vs_7 <= l2_io_rresp_data_1_entries_vs_7; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_1_entries_vs_7 <= r_7_1_entries_vs_7; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_1_entries_prefetch <= l2_io_rresp_data_1_entries_prefetch; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_1_entries_prefetch <= r_7_1_entries_prefetch; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_1_ecc <= l2_io_rresp_data_1_ecc; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_1_ecc <= r_7_1_ecc; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_2_entries_tag <= l2_io_rresp_data_2_entries_tag; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_2_entries_tag <= r_7_2_entries_tag; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_2_entries_asid <= l2_io_rresp_data_2_entries_asid; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_2_entries_asid <= r_7_2_entries_asid; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_2_entries_ppns_0 <= l2_io_rresp_data_2_entries_ppns_0; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_2_entries_ppns_0 <= r_7_2_entries_ppns_0; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_2_entries_ppns_1 <= l2_io_rresp_data_2_entries_ppns_1; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_2_entries_ppns_1 <= r_7_2_entries_ppns_1; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_2_entries_ppns_2 <= l2_io_rresp_data_2_entries_ppns_2; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_2_entries_ppns_2 <= r_7_2_entries_ppns_2; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_2_entries_ppns_3 <= l2_io_rresp_data_2_entries_ppns_3; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_2_entries_ppns_3 <= r_7_2_entries_ppns_3; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_2_entries_ppns_4 <= l2_io_rresp_data_2_entries_ppns_4; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_2_entries_ppns_4 <= r_7_2_entries_ppns_4; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_2_entries_ppns_5 <= l2_io_rresp_data_2_entries_ppns_5; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_2_entries_ppns_5 <= r_7_2_entries_ppns_5; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_2_entries_ppns_6 <= l2_io_rresp_data_2_entries_ppns_6; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_2_entries_ppns_6 <= r_7_2_entries_ppns_6; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_2_entries_ppns_7 <= l2_io_rresp_data_2_entries_ppns_7; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_2_entries_ppns_7 <= r_7_2_entries_ppns_7; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_2_entries_vs_0 <= l2_io_rresp_data_2_entries_vs_0; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_2_entries_vs_0 <= r_7_2_entries_vs_0; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_2_entries_vs_1 <= l2_io_rresp_data_2_entries_vs_1; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_2_entries_vs_1 <= r_7_2_entries_vs_1; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_2_entries_vs_2 <= l2_io_rresp_data_2_entries_vs_2; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_2_entries_vs_2 <= r_7_2_entries_vs_2; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_2_entries_vs_3 <= l2_io_rresp_data_2_entries_vs_3; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_2_entries_vs_3 <= r_7_2_entries_vs_3; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_2_entries_vs_4 <= l2_io_rresp_data_2_entries_vs_4; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_2_entries_vs_4 <= r_7_2_entries_vs_4; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_2_entries_vs_5 <= l2_io_rresp_data_2_entries_vs_5; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_2_entries_vs_5 <= r_7_2_entries_vs_5; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_2_entries_vs_6 <= l2_io_rresp_data_2_entries_vs_6; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_2_entries_vs_6 <= r_7_2_entries_vs_6; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_2_entries_vs_7 <= l2_io_rresp_data_2_entries_vs_7; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_2_entries_vs_7 <= r_7_2_entries_vs_7; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_2_entries_prefetch <= l2_io_rresp_data_2_entries_prefetch; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_2_entries_prefetch <= r_7_2_entries_prefetch; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_2_ecc <= l2_io_rresp_data_2_ecc; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_2_ecc <= r_7_2_ecc; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_3_entries_tag <= l2_io_rresp_data_3_entries_tag; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_3_entries_tag <= r_7_3_entries_tag; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_3_entries_asid <= l2_io_rresp_data_3_entries_asid; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_3_entries_asid <= r_7_3_entries_asid; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_3_entries_ppns_0 <= l2_io_rresp_data_3_entries_ppns_0; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_3_entries_ppns_0 <= r_7_3_entries_ppns_0; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_3_entries_ppns_1 <= l2_io_rresp_data_3_entries_ppns_1; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_3_entries_ppns_1 <= r_7_3_entries_ppns_1; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_3_entries_ppns_2 <= l2_io_rresp_data_3_entries_ppns_2; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_3_entries_ppns_2 <= r_7_3_entries_ppns_2; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_3_entries_ppns_3 <= l2_io_rresp_data_3_entries_ppns_3; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_3_entries_ppns_3 <= r_7_3_entries_ppns_3; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_3_entries_ppns_4 <= l2_io_rresp_data_3_entries_ppns_4; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_3_entries_ppns_4 <= r_7_3_entries_ppns_4; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_3_entries_ppns_5 <= l2_io_rresp_data_3_entries_ppns_5; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_3_entries_ppns_5 <= r_7_3_entries_ppns_5; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_3_entries_ppns_6 <= l2_io_rresp_data_3_entries_ppns_6; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_3_entries_ppns_6 <= r_7_3_entries_ppns_6; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_3_entries_ppns_7 <= l2_io_rresp_data_3_entries_ppns_7; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_3_entries_ppns_7 <= r_7_3_entries_ppns_7; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_3_entries_vs_0 <= l2_io_rresp_data_3_entries_vs_0; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_3_entries_vs_0 <= r_7_3_entries_vs_0; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_3_entries_vs_1 <= l2_io_rresp_data_3_entries_vs_1; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_3_entries_vs_1 <= r_7_3_entries_vs_1; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_3_entries_vs_2 <= l2_io_rresp_data_3_entries_vs_2; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_3_entries_vs_2 <= r_7_3_entries_vs_2; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_3_entries_vs_3 <= l2_io_rresp_data_3_entries_vs_3; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_3_entries_vs_3 <= r_7_3_entries_vs_3; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_3_entries_vs_4 <= l2_io_rresp_data_3_entries_vs_4; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_3_entries_vs_4 <= r_7_3_entries_vs_4; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_3_entries_vs_5 <= l2_io_rresp_data_3_entries_vs_5; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_3_entries_vs_5 <= r_7_3_entries_vs_5; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_3_entries_vs_6 <= l2_io_rresp_data_3_entries_vs_6; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_3_entries_vs_6 <= r_7_3_entries_vs_6; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_3_entries_vs_7 <= l2_io_rresp_data_3_entries_vs_7; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_3_entries_vs_7 <= r_7_3_entries_vs_7; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_3_entries_prefetch <= l2_io_rresp_data_3_entries_prefetch; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_3_entries_prefetch <= r_7_3_entries_prefetch; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l2_ramDatas_3_ecc <= l2_io_rresp_data_3_ecc; // @[Reg.scala 17:22]
      end else begin
        l2_ramDatas_3_ecc <= r_7_3_ecc; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      l2_hitVec_0 <= _T_84; // @[Reg.scala 17:22]
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      l2_hitVec_1 <= _T_91; // @[Reg.scala 17:22]
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      l2_hitVec_2 <= _T_98; // @[Reg.scala 17:22]
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      l2_hitVec_3 <= _T_105; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_tag <= l3_io_rresp_data_0_entries_tag; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_asid <= l3_io_rresp_data_0_entries_asid; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_ppns_0 <= l3_io_rresp_data_0_entries_ppns_0; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_ppns_1 <= l3_io_rresp_data_0_entries_ppns_1; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_ppns_2 <= l3_io_rresp_data_0_entries_ppns_2; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_ppns_3 <= l3_io_rresp_data_0_entries_ppns_3; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_ppns_4 <= l3_io_rresp_data_0_entries_ppns_4; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_ppns_5 <= l3_io_rresp_data_0_entries_ppns_5; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_ppns_6 <= l3_io_rresp_data_0_entries_ppns_6; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_ppns_7 <= l3_io_rresp_data_0_entries_ppns_7; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_vs_0 <= l3_io_rresp_data_0_entries_vs_0; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_vs_1 <= l3_io_rresp_data_0_entries_vs_1; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_vs_2 <= l3_io_rresp_data_0_entries_vs_2; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_vs_3 <= l3_io_rresp_data_0_entries_vs_3; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_vs_4 <= l3_io_rresp_data_0_entries_vs_4; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_vs_5 <= l3_io_rresp_data_0_entries_vs_5; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_vs_6 <= l3_io_rresp_data_0_entries_vs_6; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_vs_7 <= l3_io_rresp_data_0_entries_vs_7; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_perms_0_d <= l3_io_rresp_data_0_entries_perms_0_d; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_perms_0_a <= l3_io_rresp_data_0_entries_perms_0_a; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_perms_0_g <= l3_io_rresp_data_0_entries_perms_0_g; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_perms_0_u <= l3_io_rresp_data_0_entries_perms_0_u; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_perms_0_x <= l3_io_rresp_data_0_entries_perms_0_x; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_perms_0_w <= l3_io_rresp_data_0_entries_perms_0_w; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_perms_0_r <= l3_io_rresp_data_0_entries_perms_0_r; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_perms_1_d <= l3_io_rresp_data_0_entries_perms_1_d; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_perms_1_a <= l3_io_rresp_data_0_entries_perms_1_a; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_perms_1_g <= l3_io_rresp_data_0_entries_perms_1_g; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_perms_1_u <= l3_io_rresp_data_0_entries_perms_1_u; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_perms_1_x <= l3_io_rresp_data_0_entries_perms_1_x; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_perms_1_w <= l3_io_rresp_data_0_entries_perms_1_w; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_perms_1_r <= l3_io_rresp_data_0_entries_perms_1_r; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_perms_2_d <= l3_io_rresp_data_0_entries_perms_2_d; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_perms_2_a <= l3_io_rresp_data_0_entries_perms_2_a; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_perms_2_g <= l3_io_rresp_data_0_entries_perms_2_g; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_perms_2_u <= l3_io_rresp_data_0_entries_perms_2_u; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_perms_2_x <= l3_io_rresp_data_0_entries_perms_2_x; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_perms_2_w <= l3_io_rresp_data_0_entries_perms_2_w; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_perms_2_r <= l3_io_rresp_data_0_entries_perms_2_r; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_perms_3_d <= l3_io_rresp_data_0_entries_perms_3_d; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_perms_3_a <= l3_io_rresp_data_0_entries_perms_3_a; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_perms_3_g <= l3_io_rresp_data_0_entries_perms_3_g; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_perms_3_u <= l3_io_rresp_data_0_entries_perms_3_u; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_perms_3_x <= l3_io_rresp_data_0_entries_perms_3_x; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_perms_3_w <= l3_io_rresp_data_0_entries_perms_3_w; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_perms_3_r <= l3_io_rresp_data_0_entries_perms_3_r; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_perms_4_d <= l3_io_rresp_data_0_entries_perms_4_d; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_perms_4_a <= l3_io_rresp_data_0_entries_perms_4_a; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_perms_4_g <= l3_io_rresp_data_0_entries_perms_4_g; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_perms_4_u <= l3_io_rresp_data_0_entries_perms_4_u; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_perms_4_x <= l3_io_rresp_data_0_entries_perms_4_x; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_perms_4_w <= l3_io_rresp_data_0_entries_perms_4_w; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_perms_4_r <= l3_io_rresp_data_0_entries_perms_4_r; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_perms_5_d <= l3_io_rresp_data_0_entries_perms_5_d; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_perms_5_a <= l3_io_rresp_data_0_entries_perms_5_a; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_perms_5_g <= l3_io_rresp_data_0_entries_perms_5_g; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_perms_5_u <= l3_io_rresp_data_0_entries_perms_5_u; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_perms_5_x <= l3_io_rresp_data_0_entries_perms_5_x; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_perms_5_w <= l3_io_rresp_data_0_entries_perms_5_w; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_perms_5_r <= l3_io_rresp_data_0_entries_perms_5_r; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_perms_6_d <= l3_io_rresp_data_0_entries_perms_6_d; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_perms_6_a <= l3_io_rresp_data_0_entries_perms_6_a; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_perms_6_g <= l3_io_rresp_data_0_entries_perms_6_g; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_perms_6_u <= l3_io_rresp_data_0_entries_perms_6_u; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_perms_6_x <= l3_io_rresp_data_0_entries_perms_6_x; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_perms_6_w <= l3_io_rresp_data_0_entries_perms_6_w; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_perms_6_r <= l3_io_rresp_data_0_entries_perms_6_r; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_perms_7_d <= l3_io_rresp_data_0_entries_perms_7_d; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_perms_7_a <= l3_io_rresp_data_0_entries_perms_7_a; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_perms_7_g <= l3_io_rresp_data_0_entries_perms_7_g; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_perms_7_u <= l3_io_rresp_data_0_entries_perms_7_u; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_perms_7_x <= l3_io_rresp_data_0_entries_perms_7_x; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_perms_7_w <= l3_io_rresp_data_0_entries_perms_7_w; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_perms_7_r <= l3_io_rresp_data_0_entries_perms_7_r; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_entries_prefetch <= l3_io_rresp_data_0_entries_prefetch; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_0_ecc <= l3_io_rresp_data_0_ecc; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_tag <= l3_io_rresp_data_1_entries_tag; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_asid <= l3_io_rresp_data_1_entries_asid; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_ppns_0 <= l3_io_rresp_data_1_entries_ppns_0; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_ppns_1 <= l3_io_rresp_data_1_entries_ppns_1; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_ppns_2 <= l3_io_rresp_data_1_entries_ppns_2; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_ppns_3 <= l3_io_rresp_data_1_entries_ppns_3; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_ppns_4 <= l3_io_rresp_data_1_entries_ppns_4; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_ppns_5 <= l3_io_rresp_data_1_entries_ppns_5; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_ppns_6 <= l3_io_rresp_data_1_entries_ppns_6; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_ppns_7 <= l3_io_rresp_data_1_entries_ppns_7; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_vs_0 <= l3_io_rresp_data_1_entries_vs_0; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_vs_1 <= l3_io_rresp_data_1_entries_vs_1; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_vs_2 <= l3_io_rresp_data_1_entries_vs_2; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_vs_3 <= l3_io_rresp_data_1_entries_vs_3; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_vs_4 <= l3_io_rresp_data_1_entries_vs_4; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_vs_5 <= l3_io_rresp_data_1_entries_vs_5; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_vs_6 <= l3_io_rresp_data_1_entries_vs_6; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_vs_7 <= l3_io_rresp_data_1_entries_vs_7; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_perms_0_d <= l3_io_rresp_data_1_entries_perms_0_d; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_perms_0_a <= l3_io_rresp_data_1_entries_perms_0_a; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_perms_0_g <= l3_io_rresp_data_1_entries_perms_0_g; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_perms_0_u <= l3_io_rresp_data_1_entries_perms_0_u; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_perms_0_x <= l3_io_rresp_data_1_entries_perms_0_x; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_perms_0_w <= l3_io_rresp_data_1_entries_perms_0_w; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_perms_0_r <= l3_io_rresp_data_1_entries_perms_0_r; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_perms_1_d <= l3_io_rresp_data_1_entries_perms_1_d; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_perms_1_a <= l3_io_rresp_data_1_entries_perms_1_a; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_perms_1_g <= l3_io_rresp_data_1_entries_perms_1_g; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_perms_1_u <= l3_io_rresp_data_1_entries_perms_1_u; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_perms_1_x <= l3_io_rresp_data_1_entries_perms_1_x; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_perms_1_w <= l3_io_rresp_data_1_entries_perms_1_w; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_perms_1_r <= l3_io_rresp_data_1_entries_perms_1_r; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_perms_2_d <= l3_io_rresp_data_1_entries_perms_2_d; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_perms_2_a <= l3_io_rresp_data_1_entries_perms_2_a; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_perms_2_g <= l3_io_rresp_data_1_entries_perms_2_g; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_perms_2_u <= l3_io_rresp_data_1_entries_perms_2_u; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_perms_2_x <= l3_io_rresp_data_1_entries_perms_2_x; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_perms_2_w <= l3_io_rresp_data_1_entries_perms_2_w; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_perms_2_r <= l3_io_rresp_data_1_entries_perms_2_r; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_perms_3_d <= l3_io_rresp_data_1_entries_perms_3_d; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_perms_3_a <= l3_io_rresp_data_1_entries_perms_3_a; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_perms_3_g <= l3_io_rresp_data_1_entries_perms_3_g; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_perms_3_u <= l3_io_rresp_data_1_entries_perms_3_u; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_perms_3_x <= l3_io_rresp_data_1_entries_perms_3_x; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_perms_3_w <= l3_io_rresp_data_1_entries_perms_3_w; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_perms_3_r <= l3_io_rresp_data_1_entries_perms_3_r; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_perms_4_d <= l3_io_rresp_data_1_entries_perms_4_d; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_perms_4_a <= l3_io_rresp_data_1_entries_perms_4_a; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_perms_4_g <= l3_io_rresp_data_1_entries_perms_4_g; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_perms_4_u <= l3_io_rresp_data_1_entries_perms_4_u; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_perms_4_x <= l3_io_rresp_data_1_entries_perms_4_x; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_perms_4_w <= l3_io_rresp_data_1_entries_perms_4_w; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_perms_4_r <= l3_io_rresp_data_1_entries_perms_4_r; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_perms_5_d <= l3_io_rresp_data_1_entries_perms_5_d; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_perms_5_a <= l3_io_rresp_data_1_entries_perms_5_a; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_perms_5_g <= l3_io_rresp_data_1_entries_perms_5_g; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_perms_5_u <= l3_io_rresp_data_1_entries_perms_5_u; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_perms_5_x <= l3_io_rresp_data_1_entries_perms_5_x; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_perms_5_w <= l3_io_rresp_data_1_entries_perms_5_w; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_perms_5_r <= l3_io_rresp_data_1_entries_perms_5_r; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_perms_6_d <= l3_io_rresp_data_1_entries_perms_6_d; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_perms_6_a <= l3_io_rresp_data_1_entries_perms_6_a; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_perms_6_g <= l3_io_rresp_data_1_entries_perms_6_g; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_perms_6_u <= l3_io_rresp_data_1_entries_perms_6_u; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_perms_6_x <= l3_io_rresp_data_1_entries_perms_6_x; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_perms_6_w <= l3_io_rresp_data_1_entries_perms_6_w; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_perms_6_r <= l3_io_rresp_data_1_entries_perms_6_r; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_perms_7_d <= l3_io_rresp_data_1_entries_perms_7_d; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_perms_7_a <= l3_io_rresp_data_1_entries_perms_7_a; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_perms_7_g <= l3_io_rresp_data_1_entries_perms_7_g; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_perms_7_u <= l3_io_rresp_data_1_entries_perms_7_u; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_perms_7_x <= l3_io_rresp_data_1_entries_perms_7_x; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_perms_7_w <= l3_io_rresp_data_1_entries_perms_7_w; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_perms_7_r <= l3_io_rresp_data_1_entries_perms_7_r; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_entries_prefetch <= l3_io_rresp_data_1_entries_prefetch; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_1_ecc <= l3_io_rresp_data_1_ecc; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_tag <= l3_io_rresp_data_2_entries_tag; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_asid <= l3_io_rresp_data_2_entries_asid; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_ppns_0 <= l3_io_rresp_data_2_entries_ppns_0; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_ppns_1 <= l3_io_rresp_data_2_entries_ppns_1; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_ppns_2 <= l3_io_rresp_data_2_entries_ppns_2; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_ppns_3 <= l3_io_rresp_data_2_entries_ppns_3; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_ppns_4 <= l3_io_rresp_data_2_entries_ppns_4; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_ppns_5 <= l3_io_rresp_data_2_entries_ppns_5; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_ppns_6 <= l3_io_rresp_data_2_entries_ppns_6; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_ppns_7 <= l3_io_rresp_data_2_entries_ppns_7; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_vs_0 <= l3_io_rresp_data_2_entries_vs_0; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_vs_1 <= l3_io_rresp_data_2_entries_vs_1; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_vs_2 <= l3_io_rresp_data_2_entries_vs_2; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_vs_3 <= l3_io_rresp_data_2_entries_vs_3; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_vs_4 <= l3_io_rresp_data_2_entries_vs_4; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_vs_5 <= l3_io_rresp_data_2_entries_vs_5; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_vs_6 <= l3_io_rresp_data_2_entries_vs_6; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_vs_7 <= l3_io_rresp_data_2_entries_vs_7; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_perms_0_d <= l3_io_rresp_data_2_entries_perms_0_d; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_perms_0_a <= l3_io_rresp_data_2_entries_perms_0_a; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_perms_0_g <= l3_io_rresp_data_2_entries_perms_0_g; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_perms_0_u <= l3_io_rresp_data_2_entries_perms_0_u; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_perms_0_x <= l3_io_rresp_data_2_entries_perms_0_x; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_perms_0_w <= l3_io_rresp_data_2_entries_perms_0_w; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_perms_0_r <= l3_io_rresp_data_2_entries_perms_0_r; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_perms_1_d <= l3_io_rresp_data_2_entries_perms_1_d; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_perms_1_a <= l3_io_rresp_data_2_entries_perms_1_a; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_perms_1_g <= l3_io_rresp_data_2_entries_perms_1_g; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_perms_1_u <= l3_io_rresp_data_2_entries_perms_1_u; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_perms_1_x <= l3_io_rresp_data_2_entries_perms_1_x; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_perms_1_w <= l3_io_rresp_data_2_entries_perms_1_w; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_perms_1_r <= l3_io_rresp_data_2_entries_perms_1_r; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_perms_2_d <= l3_io_rresp_data_2_entries_perms_2_d; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_perms_2_a <= l3_io_rresp_data_2_entries_perms_2_a; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_perms_2_g <= l3_io_rresp_data_2_entries_perms_2_g; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_perms_2_u <= l3_io_rresp_data_2_entries_perms_2_u; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_perms_2_x <= l3_io_rresp_data_2_entries_perms_2_x; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_perms_2_w <= l3_io_rresp_data_2_entries_perms_2_w; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_perms_2_r <= l3_io_rresp_data_2_entries_perms_2_r; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_perms_3_d <= l3_io_rresp_data_2_entries_perms_3_d; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_perms_3_a <= l3_io_rresp_data_2_entries_perms_3_a; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_perms_3_g <= l3_io_rresp_data_2_entries_perms_3_g; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_perms_3_u <= l3_io_rresp_data_2_entries_perms_3_u; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_perms_3_x <= l3_io_rresp_data_2_entries_perms_3_x; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_perms_3_w <= l3_io_rresp_data_2_entries_perms_3_w; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_perms_3_r <= l3_io_rresp_data_2_entries_perms_3_r; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_perms_4_d <= l3_io_rresp_data_2_entries_perms_4_d; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_perms_4_a <= l3_io_rresp_data_2_entries_perms_4_a; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_perms_4_g <= l3_io_rresp_data_2_entries_perms_4_g; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_perms_4_u <= l3_io_rresp_data_2_entries_perms_4_u; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_perms_4_x <= l3_io_rresp_data_2_entries_perms_4_x; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_perms_4_w <= l3_io_rresp_data_2_entries_perms_4_w; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_perms_4_r <= l3_io_rresp_data_2_entries_perms_4_r; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_perms_5_d <= l3_io_rresp_data_2_entries_perms_5_d; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_perms_5_a <= l3_io_rresp_data_2_entries_perms_5_a; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_perms_5_g <= l3_io_rresp_data_2_entries_perms_5_g; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_perms_5_u <= l3_io_rresp_data_2_entries_perms_5_u; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_perms_5_x <= l3_io_rresp_data_2_entries_perms_5_x; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_perms_5_w <= l3_io_rresp_data_2_entries_perms_5_w; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_perms_5_r <= l3_io_rresp_data_2_entries_perms_5_r; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_perms_6_d <= l3_io_rresp_data_2_entries_perms_6_d; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_perms_6_a <= l3_io_rresp_data_2_entries_perms_6_a; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_perms_6_g <= l3_io_rresp_data_2_entries_perms_6_g; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_perms_6_u <= l3_io_rresp_data_2_entries_perms_6_u; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_perms_6_x <= l3_io_rresp_data_2_entries_perms_6_x; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_perms_6_w <= l3_io_rresp_data_2_entries_perms_6_w; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_perms_6_r <= l3_io_rresp_data_2_entries_perms_6_r; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_perms_7_d <= l3_io_rresp_data_2_entries_perms_7_d; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_perms_7_a <= l3_io_rresp_data_2_entries_perms_7_a; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_perms_7_g <= l3_io_rresp_data_2_entries_perms_7_g; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_perms_7_u <= l3_io_rresp_data_2_entries_perms_7_u; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_perms_7_x <= l3_io_rresp_data_2_entries_perms_7_x; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_perms_7_w <= l3_io_rresp_data_2_entries_perms_7_w; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_perms_7_r <= l3_io_rresp_data_2_entries_perms_7_r; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_entries_prefetch <= l3_io_rresp_data_2_entries_prefetch; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_2_ecc <= l3_io_rresp_data_2_ecc; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_tag <= l3_io_rresp_data_3_entries_tag; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_asid <= l3_io_rresp_data_3_entries_asid; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_ppns_0 <= l3_io_rresp_data_3_entries_ppns_0; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_ppns_1 <= l3_io_rresp_data_3_entries_ppns_1; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_ppns_2 <= l3_io_rresp_data_3_entries_ppns_2; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_ppns_3 <= l3_io_rresp_data_3_entries_ppns_3; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_ppns_4 <= l3_io_rresp_data_3_entries_ppns_4; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_ppns_5 <= l3_io_rresp_data_3_entries_ppns_5; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_ppns_6 <= l3_io_rresp_data_3_entries_ppns_6; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_ppns_7 <= l3_io_rresp_data_3_entries_ppns_7; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_vs_0 <= l3_io_rresp_data_3_entries_vs_0; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_vs_1 <= l3_io_rresp_data_3_entries_vs_1; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_vs_2 <= l3_io_rresp_data_3_entries_vs_2; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_vs_3 <= l3_io_rresp_data_3_entries_vs_3; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_vs_4 <= l3_io_rresp_data_3_entries_vs_4; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_vs_5 <= l3_io_rresp_data_3_entries_vs_5; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_vs_6 <= l3_io_rresp_data_3_entries_vs_6; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_vs_7 <= l3_io_rresp_data_3_entries_vs_7; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_perms_0_d <= l3_io_rresp_data_3_entries_perms_0_d; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_perms_0_a <= l3_io_rresp_data_3_entries_perms_0_a; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_perms_0_g <= l3_io_rresp_data_3_entries_perms_0_g; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_perms_0_u <= l3_io_rresp_data_3_entries_perms_0_u; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_perms_0_x <= l3_io_rresp_data_3_entries_perms_0_x; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_perms_0_w <= l3_io_rresp_data_3_entries_perms_0_w; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_perms_0_r <= l3_io_rresp_data_3_entries_perms_0_r; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_perms_1_d <= l3_io_rresp_data_3_entries_perms_1_d; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_perms_1_a <= l3_io_rresp_data_3_entries_perms_1_a; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_perms_1_g <= l3_io_rresp_data_3_entries_perms_1_g; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_perms_1_u <= l3_io_rresp_data_3_entries_perms_1_u; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_perms_1_x <= l3_io_rresp_data_3_entries_perms_1_x; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_perms_1_w <= l3_io_rresp_data_3_entries_perms_1_w; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_perms_1_r <= l3_io_rresp_data_3_entries_perms_1_r; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_perms_2_d <= l3_io_rresp_data_3_entries_perms_2_d; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_perms_2_a <= l3_io_rresp_data_3_entries_perms_2_a; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_perms_2_g <= l3_io_rresp_data_3_entries_perms_2_g; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_perms_2_u <= l3_io_rresp_data_3_entries_perms_2_u; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_perms_2_x <= l3_io_rresp_data_3_entries_perms_2_x; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_perms_2_w <= l3_io_rresp_data_3_entries_perms_2_w; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_perms_2_r <= l3_io_rresp_data_3_entries_perms_2_r; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_perms_3_d <= l3_io_rresp_data_3_entries_perms_3_d; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_perms_3_a <= l3_io_rresp_data_3_entries_perms_3_a; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_perms_3_g <= l3_io_rresp_data_3_entries_perms_3_g; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_perms_3_u <= l3_io_rresp_data_3_entries_perms_3_u; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_perms_3_x <= l3_io_rresp_data_3_entries_perms_3_x; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_perms_3_w <= l3_io_rresp_data_3_entries_perms_3_w; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_perms_3_r <= l3_io_rresp_data_3_entries_perms_3_r; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_perms_4_d <= l3_io_rresp_data_3_entries_perms_4_d; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_perms_4_a <= l3_io_rresp_data_3_entries_perms_4_a; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_perms_4_g <= l3_io_rresp_data_3_entries_perms_4_g; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_perms_4_u <= l3_io_rresp_data_3_entries_perms_4_u; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_perms_4_x <= l3_io_rresp_data_3_entries_perms_4_x; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_perms_4_w <= l3_io_rresp_data_3_entries_perms_4_w; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_perms_4_r <= l3_io_rresp_data_3_entries_perms_4_r; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_perms_5_d <= l3_io_rresp_data_3_entries_perms_5_d; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_perms_5_a <= l3_io_rresp_data_3_entries_perms_5_a; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_perms_5_g <= l3_io_rresp_data_3_entries_perms_5_g; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_perms_5_u <= l3_io_rresp_data_3_entries_perms_5_u; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_perms_5_x <= l3_io_rresp_data_3_entries_perms_5_x; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_perms_5_w <= l3_io_rresp_data_3_entries_perms_5_w; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_perms_5_r <= l3_io_rresp_data_3_entries_perms_5_r; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_perms_6_d <= l3_io_rresp_data_3_entries_perms_6_d; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_perms_6_a <= l3_io_rresp_data_3_entries_perms_6_a; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_perms_6_g <= l3_io_rresp_data_3_entries_perms_6_g; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_perms_6_u <= l3_io_rresp_data_3_entries_perms_6_u; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_perms_6_x <= l3_io_rresp_data_3_entries_perms_6_x; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_perms_6_w <= l3_io_rresp_data_3_entries_perms_6_w; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_perms_6_r <= l3_io_rresp_data_3_entries_perms_6_r; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_perms_7_d <= l3_io_rresp_data_3_entries_perms_7_d; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_perms_7_a <= l3_io_rresp_data_3_entries_perms_7_a; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_perms_7_g <= l3_io_rresp_data_3_entries_perms_7_g; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_perms_7_u <= l3_io_rresp_data_3_entries_perms_7_u; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_perms_7_x <= l3_io_rresp_data_3_entries_perms_7_x; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_perms_7_w <= l3_io_rresp_data_3_entries_perms_7_w; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_perms_7_r <= l3_io_rresp_data_3_entries_perms_7_r; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_entries_prefetch <= l3_io_rresp_data_3_entries_prefetch; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_3_ecc <= l3_io_rresp_data_3_ecc; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_tag <= l3_io_rresp_data_4_entries_tag; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_asid <= l3_io_rresp_data_4_entries_asid; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_ppns_0 <= l3_io_rresp_data_4_entries_ppns_0; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_ppns_1 <= l3_io_rresp_data_4_entries_ppns_1; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_ppns_2 <= l3_io_rresp_data_4_entries_ppns_2; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_ppns_3 <= l3_io_rresp_data_4_entries_ppns_3; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_ppns_4 <= l3_io_rresp_data_4_entries_ppns_4; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_ppns_5 <= l3_io_rresp_data_4_entries_ppns_5; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_ppns_6 <= l3_io_rresp_data_4_entries_ppns_6; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_ppns_7 <= l3_io_rresp_data_4_entries_ppns_7; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_vs_0 <= l3_io_rresp_data_4_entries_vs_0; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_vs_1 <= l3_io_rresp_data_4_entries_vs_1; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_vs_2 <= l3_io_rresp_data_4_entries_vs_2; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_vs_3 <= l3_io_rresp_data_4_entries_vs_3; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_vs_4 <= l3_io_rresp_data_4_entries_vs_4; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_vs_5 <= l3_io_rresp_data_4_entries_vs_5; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_vs_6 <= l3_io_rresp_data_4_entries_vs_6; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_vs_7 <= l3_io_rresp_data_4_entries_vs_7; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_perms_0_d <= l3_io_rresp_data_4_entries_perms_0_d; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_perms_0_a <= l3_io_rresp_data_4_entries_perms_0_a; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_perms_0_g <= l3_io_rresp_data_4_entries_perms_0_g; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_perms_0_u <= l3_io_rresp_data_4_entries_perms_0_u; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_perms_0_x <= l3_io_rresp_data_4_entries_perms_0_x; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_perms_0_w <= l3_io_rresp_data_4_entries_perms_0_w; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_perms_0_r <= l3_io_rresp_data_4_entries_perms_0_r; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_perms_1_d <= l3_io_rresp_data_4_entries_perms_1_d; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_perms_1_a <= l3_io_rresp_data_4_entries_perms_1_a; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_perms_1_g <= l3_io_rresp_data_4_entries_perms_1_g; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_perms_1_u <= l3_io_rresp_data_4_entries_perms_1_u; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_perms_1_x <= l3_io_rresp_data_4_entries_perms_1_x; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_perms_1_w <= l3_io_rresp_data_4_entries_perms_1_w; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_perms_1_r <= l3_io_rresp_data_4_entries_perms_1_r; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_perms_2_d <= l3_io_rresp_data_4_entries_perms_2_d; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_perms_2_a <= l3_io_rresp_data_4_entries_perms_2_a; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_perms_2_g <= l3_io_rresp_data_4_entries_perms_2_g; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_perms_2_u <= l3_io_rresp_data_4_entries_perms_2_u; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_perms_2_x <= l3_io_rresp_data_4_entries_perms_2_x; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_perms_2_w <= l3_io_rresp_data_4_entries_perms_2_w; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_perms_2_r <= l3_io_rresp_data_4_entries_perms_2_r; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_perms_3_d <= l3_io_rresp_data_4_entries_perms_3_d; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_perms_3_a <= l3_io_rresp_data_4_entries_perms_3_a; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_perms_3_g <= l3_io_rresp_data_4_entries_perms_3_g; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_perms_3_u <= l3_io_rresp_data_4_entries_perms_3_u; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_perms_3_x <= l3_io_rresp_data_4_entries_perms_3_x; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_perms_3_w <= l3_io_rresp_data_4_entries_perms_3_w; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_perms_3_r <= l3_io_rresp_data_4_entries_perms_3_r; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_perms_4_d <= l3_io_rresp_data_4_entries_perms_4_d; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_perms_4_a <= l3_io_rresp_data_4_entries_perms_4_a; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_perms_4_g <= l3_io_rresp_data_4_entries_perms_4_g; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_perms_4_u <= l3_io_rresp_data_4_entries_perms_4_u; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_perms_4_x <= l3_io_rresp_data_4_entries_perms_4_x; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_perms_4_w <= l3_io_rresp_data_4_entries_perms_4_w; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_perms_4_r <= l3_io_rresp_data_4_entries_perms_4_r; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_perms_5_d <= l3_io_rresp_data_4_entries_perms_5_d; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_perms_5_a <= l3_io_rresp_data_4_entries_perms_5_a; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_perms_5_g <= l3_io_rresp_data_4_entries_perms_5_g; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_perms_5_u <= l3_io_rresp_data_4_entries_perms_5_u; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_perms_5_x <= l3_io_rresp_data_4_entries_perms_5_x; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_perms_5_w <= l3_io_rresp_data_4_entries_perms_5_w; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_perms_5_r <= l3_io_rresp_data_4_entries_perms_5_r; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_perms_6_d <= l3_io_rresp_data_4_entries_perms_6_d; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_perms_6_a <= l3_io_rresp_data_4_entries_perms_6_a; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_perms_6_g <= l3_io_rresp_data_4_entries_perms_6_g; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_perms_6_u <= l3_io_rresp_data_4_entries_perms_6_u; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_perms_6_x <= l3_io_rresp_data_4_entries_perms_6_x; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_perms_6_w <= l3_io_rresp_data_4_entries_perms_6_w; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_perms_6_r <= l3_io_rresp_data_4_entries_perms_6_r; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_perms_7_d <= l3_io_rresp_data_4_entries_perms_7_d; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_perms_7_a <= l3_io_rresp_data_4_entries_perms_7_a; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_perms_7_g <= l3_io_rresp_data_4_entries_perms_7_g; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_perms_7_u <= l3_io_rresp_data_4_entries_perms_7_u; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_perms_7_x <= l3_io_rresp_data_4_entries_perms_7_x; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_perms_7_w <= l3_io_rresp_data_4_entries_perms_7_w; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_perms_7_r <= l3_io_rresp_data_4_entries_perms_7_r; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_entries_prefetch <= l3_io_rresp_data_4_entries_prefetch; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_4_ecc <= l3_io_rresp_data_4_ecc; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_tag <= l3_io_rresp_data_5_entries_tag; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_asid <= l3_io_rresp_data_5_entries_asid; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_ppns_0 <= l3_io_rresp_data_5_entries_ppns_0; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_ppns_1 <= l3_io_rresp_data_5_entries_ppns_1; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_ppns_2 <= l3_io_rresp_data_5_entries_ppns_2; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_ppns_3 <= l3_io_rresp_data_5_entries_ppns_3; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_ppns_4 <= l3_io_rresp_data_5_entries_ppns_4; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_ppns_5 <= l3_io_rresp_data_5_entries_ppns_5; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_ppns_6 <= l3_io_rresp_data_5_entries_ppns_6; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_ppns_7 <= l3_io_rresp_data_5_entries_ppns_7; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_vs_0 <= l3_io_rresp_data_5_entries_vs_0; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_vs_1 <= l3_io_rresp_data_5_entries_vs_1; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_vs_2 <= l3_io_rresp_data_5_entries_vs_2; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_vs_3 <= l3_io_rresp_data_5_entries_vs_3; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_vs_4 <= l3_io_rresp_data_5_entries_vs_4; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_vs_5 <= l3_io_rresp_data_5_entries_vs_5; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_vs_6 <= l3_io_rresp_data_5_entries_vs_6; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_vs_7 <= l3_io_rresp_data_5_entries_vs_7; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_perms_0_d <= l3_io_rresp_data_5_entries_perms_0_d; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_perms_0_a <= l3_io_rresp_data_5_entries_perms_0_a; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_perms_0_g <= l3_io_rresp_data_5_entries_perms_0_g; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_perms_0_u <= l3_io_rresp_data_5_entries_perms_0_u; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_perms_0_x <= l3_io_rresp_data_5_entries_perms_0_x; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_perms_0_w <= l3_io_rresp_data_5_entries_perms_0_w; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_perms_0_r <= l3_io_rresp_data_5_entries_perms_0_r; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_perms_1_d <= l3_io_rresp_data_5_entries_perms_1_d; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_perms_1_a <= l3_io_rresp_data_5_entries_perms_1_a; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_perms_1_g <= l3_io_rresp_data_5_entries_perms_1_g; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_perms_1_u <= l3_io_rresp_data_5_entries_perms_1_u; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_perms_1_x <= l3_io_rresp_data_5_entries_perms_1_x; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_perms_1_w <= l3_io_rresp_data_5_entries_perms_1_w; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_perms_1_r <= l3_io_rresp_data_5_entries_perms_1_r; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_perms_2_d <= l3_io_rresp_data_5_entries_perms_2_d; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_perms_2_a <= l3_io_rresp_data_5_entries_perms_2_a; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_perms_2_g <= l3_io_rresp_data_5_entries_perms_2_g; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_perms_2_u <= l3_io_rresp_data_5_entries_perms_2_u; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_perms_2_x <= l3_io_rresp_data_5_entries_perms_2_x; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_perms_2_w <= l3_io_rresp_data_5_entries_perms_2_w; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_perms_2_r <= l3_io_rresp_data_5_entries_perms_2_r; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_perms_3_d <= l3_io_rresp_data_5_entries_perms_3_d; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_perms_3_a <= l3_io_rresp_data_5_entries_perms_3_a; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_perms_3_g <= l3_io_rresp_data_5_entries_perms_3_g; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_perms_3_u <= l3_io_rresp_data_5_entries_perms_3_u; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_perms_3_x <= l3_io_rresp_data_5_entries_perms_3_x; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_perms_3_w <= l3_io_rresp_data_5_entries_perms_3_w; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_perms_3_r <= l3_io_rresp_data_5_entries_perms_3_r; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_perms_4_d <= l3_io_rresp_data_5_entries_perms_4_d; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_perms_4_a <= l3_io_rresp_data_5_entries_perms_4_a; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_perms_4_g <= l3_io_rresp_data_5_entries_perms_4_g; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_perms_4_u <= l3_io_rresp_data_5_entries_perms_4_u; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_perms_4_x <= l3_io_rresp_data_5_entries_perms_4_x; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_perms_4_w <= l3_io_rresp_data_5_entries_perms_4_w; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_perms_4_r <= l3_io_rresp_data_5_entries_perms_4_r; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_perms_5_d <= l3_io_rresp_data_5_entries_perms_5_d; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_perms_5_a <= l3_io_rresp_data_5_entries_perms_5_a; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_perms_5_g <= l3_io_rresp_data_5_entries_perms_5_g; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_perms_5_u <= l3_io_rresp_data_5_entries_perms_5_u; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_perms_5_x <= l3_io_rresp_data_5_entries_perms_5_x; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_perms_5_w <= l3_io_rresp_data_5_entries_perms_5_w; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_perms_5_r <= l3_io_rresp_data_5_entries_perms_5_r; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_perms_6_d <= l3_io_rresp_data_5_entries_perms_6_d; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_perms_6_a <= l3_io_rresp_data_5_entries_perms_6_a; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_perms_6_g <= l3_io_rresp_data_5_entries_perms_6_g; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_perms_6_u <= l3_io_rresp_data_5_entries_perms_6_u; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_perms_6_x <= l3_io_rresp_data_5_entries_perms_6_x; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_perms_6_w <= l3_io_rresp_data_5_entries_perms_6_w; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_perms_6_r <= l3_io_rresp_data_5_entries_perms_6_r; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_perms_7_d <= l3_io_rresp_data_5_entries_perms_7_d; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_perms_7_a <= l3_io_rresp_data_5_entries_perms_7_a; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_perms_7_g <= l3_io_rresp_data_5_entries_perms_7_g; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_perms_7_u <= l3_io_rresp_data_5_entries_perms_7_u; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_perms_7_x <= l3_io_rresp_data_5_entries_perms_7_x; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_perms_7_w <= l3_io_rresp_data_5_entries_perms_7_w; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_perms_7_r <= l3_io_rresp_data_5_entries_perms_7_r; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_entries_prefetch <= l3_io_rresp_data_5_entries_prefetch; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_5_ecc <= l3_io_rresp_data_5_ecc; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_tag <= l3_io_rresp_data_6_entries_tag; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_asid <= l3_io_rresp_data_6_entries_asid; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_ppns_0 <= l3_io_rresp_data_6_entries_ppns_0; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_ppns_1 <= l3_io_rresp_data_6_entries_ppns_1; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_ppns_2 <= l3_io_rresp_data_6_entries_ppns_2; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_ppns_3 <= l3_io_rresp_data_6_entries_ppns_3; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_ppns_4 <= l3_io_rresp_data_6_entries_ppns_4; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_ppns_5 <= l3_io_rresp_data_6_entries_ppns_5; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_ppns_6 <= l3_io_rresp_data_6_entries_ppns_6; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_ppns_7 <= l3_io_rresp_data_6_entries_ppns_7; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_vs_0 <= l3_io_rresp_data_6_entries_vs_0; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_vs_1 <= l3_io_rresp_data_6_entries_vs_1; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_vs_2 <= l3_io_rresp_data_6_entries_vs_2; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_vs_3 <= l3_io_rresp_data_6_entries_vs_3; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_vs_4 <= l3_io_rresp_data_6_entries_vs_4; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_vs_5 <= l3_io_rresp_data_6_entries_vs_5; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_vs_6 <= l3_io_rresp_data_6_entries_vs_6; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_vs_7 <= l3_io_rresp_data_6_entries_vs_7; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_perms_0_d <= l3_io_rresp_data_6_entries_perms_0_d; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_perms_0_a <= l3_io_rresp_data_6_entries_perms_0_a; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_perms_0_g <= l3_io_rresp_data_6_entries_perms_0_g; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_perms_0_u <= l3_io_rresp_data_6_entries_perms_0_u; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_perms_0_x <= l3_io_rresp_data_6_entries_perms_0_x; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_perms_0_w <= l3_io_rresp_data_6_entries_perms_0_w; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_perms_0_r <= l3_io_rresp_data_6_entries_perms_0_r; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_perms_1_d <= l3_io_rresp_data_6_entries_perms_1_d; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_perms_1_a <= l3_io_rresp_data_6_entries_perms_1_a; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_perms_1_g <= l3_io_rresp_data_6_entries_perms_1_g; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_perms_1_u <= l3_io_rresp_data_6_entries_perms_1_u; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_perms_1_x <= l3_io_rresp_data_6_entries_perms_1_x; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_perms_1_w <= l3_io_rresp_data_6_entries_perms_1_w; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_perms_1_r <= l3_io_rresp_data_6_entries_perms_1_r; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_perms_2_d <= l3_io_rresp_data_6_entries_perms_2_d; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_perms_2_a <= l3_io_rresp_data_6_entries_perms_2_a; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_perms_2_g <= l3_io_rresp_data_6_entries_perms_2_g; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_perms_2_u <= l3_io_rresp_data_6_entries_perms_2_u; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_perms_2_x <= l3_io_rresp_data_6_entries_perms_2_x; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_perms_2_w <= l3_io_rresp_data_6_entries_perms_2_w; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_perms_2_r <= l3_io_rresp_data_6_entries_perms_2_r; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_perms_3_d <= l3_io_rresp_data_6_entries_perms_3_d; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_perms_3_a <= l3_io_rresp_data_6_entries_perms_3_a; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_perms_3_g <= l3_io_rresp_data_6_entries_perms_3_g; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_perms_3_u <= l3_io_rresp_data_6_entries_perms_3_u; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_perms_3_x <= l3_io_rresp_data_6_entries_perms_3_x; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_perms_3_w <= l3_io_rresp_data_6_entries_perms_3_w; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_perms_3_r <= l3_io_rresp_data_6_entries_perms_3_r; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_perms_4_d <= l3_io_rresp_data_6_entries_perms_4_d; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_perms_4_a <= l3_io_rresp_data_6_entries_perms_4_a; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_perms_4_g <= l3_io_rresp_data_6_entries_perms_4_g; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_perms_4_u <= l3_io_rresp_data_6_entries_perms_4_u; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_perms_4_x <= l3_io_rresp_data_6_entries_perms_4_x; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_perms_4_w <= l3_io_rresp_data_6_entries_perms_4_w; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_perms_4_r <= l3_io_rresp_data_6_entries_perms_4_r; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_perms_5_d <= l3_io_rresp_data_6_entries_perms_5_d; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_perms_5_a <= l3_io_rresp_data_6_entries_perms_5_a; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_perms_5_g <= l3_io_rresp_data_6_entries_perms_5_g; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_perms_5_u <= l3_io_rresp_data_6_entries_perms_5_u; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_perms_5_x <= l3_io_rresp_data_6_entries_perms_5_x; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_perms_5_w <= l3_io_rresp_data_6_entries_perms_5_w; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_perms_5_r <= l3_io_rresp_data_6_entries_perms_5_r; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_perms_6_d <= l3_io_rresp_data_6_entries_perms_6_d; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_perms_6_a <= l3_io_rresp_data_6_entries_perms_6_a; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_perms_6_g <= l3_io_rresp_data_6_entries_perms_6_g; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_perms_6_u <= l3_io_rresp_data_6_entries_perms_6_u; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_perms_6_x <= l3_io_rresp_data_6_entries_perms_6_x; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_perms_6_w <= l3_io_rresp_data_6_entries_perms_6_w; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_perms_6_r <= l3_io_rresp_data_6_entries_perms_6_r; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_perms_7_d <= l3_io_rresp_data_6_entries_perms_7_d; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_perms_7_a <= l3_io_rresp_data_6_entries_perms_7_a; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_perms_7_g <= l3_io_rresp_data_6_entries_perms_7_g; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_perms_7_u <= l3_io_rresp_data_6_entries_perms_7_u; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_perms_7_x <= l3_io_rresp_data_6_entries_perms_7_x; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_perms_7_w <= l3_io_rresp_data_6_entries_perms_7_w; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_perms_7_r <= l3_io_rresp_data_6_entries_perms_7_r; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_entries_prefetch <= l3_io_rresp_data_6_entries_prefetch; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_6_ecc <= l3_io_rresp_data_6_ecc; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_tag <= l3_io_rresp_data_7_entries_tag; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_asid <= l3_io_rresp_data_7_entries_asid; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_ppns_0 <= l3_io_rresp_data_7_entries_ppns_0; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_ppns_1 <= l3_io_rresp_data_7_entries_ppns_1; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_ppns_2 <= l3_io_rresp_data_7_entries_ppns_2; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_ppns_3 <= l3_io_rresp_data_7_entries_ppns_3; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_ppns_4 <= l3_io_rresp_data_7_entries_ppns_4; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_ppns_5 <= l3_io_rresp_data_7_entries_ppns_5; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_ppns_6 <= l3_io_rresp_data_7_entries_ppns_6; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_ppns_7 <= l3_io_rresp_data_7_entries_ppns_7; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_vs_0 <= l3_io_rresp_data_7_entries_vs_0; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_vs_1 <= l3_io_rresp_data_7_entries_vs_1; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_vs_2 <= l3_io_rresp_data_7_entries_vs_2; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_vs_3 <= l3_io_rresp_data_7_entries_vs_3; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_vs_4 <= l3_io_rresp_data_7_entries_vs_4; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_vs_5 <= l3_io_rresp_data_7_entries_vs_5; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_vs_6 <= l3_io_rresp_data_7_entries_vs_6; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_vs_7 <= l3_io_rresp_data_7_entries_vs_7; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_perms_0_d <= l3_io_rresp_data_7_entries_perms_0_d; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_perms_0_a <= l3_io_rresp_data_7_entries_perms_0_a; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_perms_0_g <= l3_io_rresp_data_7_entries_perms_0_g; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_perms_0_u <= l3_io_rresp_data_7_entries_perms_0_u; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_perms_0_x <= l3_io_rresp_data_7_entries_perms_0_x; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_perms_0_w <= l3_io_rresp_data_7_entries_perms_0_w; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_perms_0_r <= l3_io_rresp_data_7_entries_perms_0_r; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_perms_1_d <= l3_io_rresp_data_7_entries_perms_1_d; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_perms_1_a <= l3_io_rresp_data_7_entries_perms_1_a; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_perms_1_g <= l3_io_rresp_data_7_entries_perms_1_g; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_perms_1_u <= l3_io_rresp_data_7_entries_perms_1_u; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_perms_1_x <= l3_io_rresp_data_7_entries_perms_1_x; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_perms_1_w <= l3_io_rresp_data_7_entries_perms_1_w; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_perms_1_r <= l3_io_rresp_data_7_entries_perms_1_r; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_perms_2_d <= l3_io_rresp_data_7_entries_perms_2_d; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_perms_2_a <= l3_io_rresp_data_7_entries_perms_2_a; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_perms_2_g <= l3_io_rresp_data_7_entries_perms_2_g; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_perms_2_u <= l3_io_rresp_data_7_entries_perms_2_u; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_perms_2_x <= l3_io_rresp_data_7_entries_perms_2_x; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_perms_2_w <= l3_io_rresp_data_7_entries_perms_2_w; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_perms_2_r <= l3_io_rresp_data_7_entries_perms_2_r; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_perms_3_d <= l3_io_rresp_data_7_entries_perms_3_d; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_perms_3_a <= l3_io_rresp_data_7_entries_perms_3_a; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_perms_3_g <= l3_io_rresp_data_7_entries_perms_3_g; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_perms_3_u <= l3_io_rresp_data_7_entries_perms_3_u; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_perms_3_x <= l3_io_rresp_data_7_entries_perms_3_x; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_perms_3_w <= l3_io_rresp_data_7_entries_perms_3_w; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_perms_3_r <= l3_io_rresp_data_7_entries_perms_3_r; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_perms_4_d <= l3_io_rresp_data_7_entries_perms_4_d; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_perms_4_a <= l3_io_rresp_data_7_entries_perms_4_a; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_perms_4_g <= l3_io_rresp_data_7_entries_perms_4_g; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_perms_4_u <= l3_io_rresp_data_7_entries_perms_4_u; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_perms_4_x <= l3_io_rresp_data_7_entries_perms_4_x; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_perms_4_w <= l3_io_rresp_data_7_entries_perms_4_w; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_perms_4_r <= l3_io_rresp_data_7_entries_perms_4_r; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_perms_5_d <= l3_io_rresp_data_7_entries_perms_5_d; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_perms_5_a <= l3_io_rresp_data_7_entries_perms_5_a; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_perms_5_g <= l3_io_rresp_data_7_entries_perms_5_g; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_perms_5_u <= l3_io_rresp_data_7_entries_perms_5_u; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_perms_5_x <= l3_io_rresp_data_7_entries_perms_5_x; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_perms_5_w <= l3_io_rresp_data_7_entries_perms_5_w; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_perms_5_r <= l3_io_rresp_data_7_entries_perms_5_r; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_perms_6_d <= l3_io_rresp_data_7_entries_perms_6_d; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_perms_6_a <= l3_io_rresp_data_7_entries_perms_6_a; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_perms_6_g <= l3_io_rresp_data_7_entries_perms_6_g; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_perms_6_u <= l3_io_rresp_data_7_entries_perms_6_u; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_perms_6_x <= l3_io_rresp_data_7_entries_perms_6_x; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_perms_6_w <= l3_io_rresp_data_7_entries_perms_6_w; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_perms_6_r <= l3_io_rresp_data_7_entries_perms_6_r; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_perms_7_d <= l3_io_rresp_data_7_entries_perms_7_d; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_perms_7_a <= l3_io_rresp_data_7_entries_perms_7_a; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_perms_7_g <= l3_io_rresp_data_7_entries_perms_7_g; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_perms_7_u <= l3_io_rresp_data_7_entries_perms_7_u; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_perms_7_x <= l3_io_rresp_data_7_entries_perms_7_x; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_perms_7_w <= l3_io_rresp_data_7_entries_perms_7_w; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_perms_7_r <= l3_io_rresp_data_7_entries_perms_7_r; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_entries_prefetch <= l3_io_rresp_data_7_entries_prefetch; // @[Reg.scala 17:22]
    end
    if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
      r_10_7_ecc <= l3_io_rresp_data_7_ecc; // @[Reg.scala 17:22]
    end
    if (_stageDelay_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (2'h3 == l3_ridx) begin // @[Reg.scala 17:22]
        r_11 <= l3vVec_3; // @[Reg.scala 17:22]
      end else if (2'h2 == l3_ridx) begin // @[Reg.scala 17:22]
        r_11 <= l3vVec_2; // @[Reg.scala 17:22]
      end else if (2'h1 == l3_ridx) begin // @[Reg.scala 17:22]
        r_11 <= l3vVec_1; // @[Reg.scala 17:22]
      end else begin
        r_11 <= l3vVec_0;
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_tag <= l3_io_rresp_data_0_entries_tag; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_tag <= r_10_0_entries_tag; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_asid <= l3_io_rresp_data_0_entries_asid; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_asid <= r_10_0_entries_asid; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_ppns_0 <= l3_io_rresp_data_0_entries_ppns_0; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_ppns_0 <= r_10_0_entries_ppns_0; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_ppns_1 <= l3_io_rresp_data_0_entries_ppns_1; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_ppns_1 <= r_10_0_entries_ppns_1; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_ppns_2 <= l3_io_rresp_data_0_entries_ppns_2; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_ppns_2 <= r_10_0_entries_ppns_2; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_ppns_3 <= l3_io_rresp_data_0_entries_ppns_3; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_ppns_3 <= r_10_0_entries_ppns_3; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_ppns_4 <= l3_io_rresp_data_0_entries_ppns_4; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_ppns_4 <= r_10_0_entries_ppns_4; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_ppns_5 <= l3_io_rresp_data_0_entries_ppns_5; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_ppns_5 <= r_10_0_entries_ppns_5; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_ppns_6 <= l3_io_rresp_data_0_entries_ppns_6; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_ppns_6 <= r_10_0_entries_ppns_6; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_ppns_7 <= l3_io_rresp_data_0_entries_ppns_7; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_ppns_7 <= r_10_0_entries_ppns_7; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_vs_0 <= l3_io_rresp_data_0_entries_vs_0; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_vs_0 <= r_10_0_entries_vs_0; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_vs_1 <= l3_io_rresp_data_0_entries_vs_1; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_vs_1 <= r_10_0_entries_vs_1; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_vs_2 <= l3_io_rresp_data_0_entries_vs_2; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_vs_2 <= r_10_0_entries_vs_2; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_vs_3 <= l3_io_rresp_data_0_entries_vs_3; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_vs_3 <= r_10_0_entries_vs_3; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_vs_4 <= l3_io_rresp_data_0_entries_vs_4; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_vs_4 <= r_10_0_entries_vs_4; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_vs_5 <= l3_io_rresp_data_0_entries_vs_5; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_vs_5 <= r_10_0_entries_vs_5; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_vs_6 <= l3_io_rresp_data_0_entries_vs_6; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_vs_6 <= r_10_0_entries_vs_6; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_vs_7 <= l3_io_rresp_data_0_entries_vs_7; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_vs_7 <= r_10_0_entries_vs_7; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_perms_0_d <= l3_io_rresp_data_0_entries_perms_0_d; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_perms_0_d <= r_10_0_entries_perms_0_d; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_perms_0_a <= l3_io_rresp_data_0_entries_perms_0_a; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_perms_0_a <= r_10_0_entries_perms_0_a; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_perms_0_g <= l3_io_rresp_data_0_entries_perms_0_g; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_perms_0_g <= r_10_0_entries_perms_0_g; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_perms_0_u <= l3_io_rresp_data_0_entries_perms_0_u; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_perms_0_u <= r_10_0_entries_perms_0_u; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_perms_0_x <= l3_io_rresp_data_0_entries_perms_0_x; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_perms_0_x <= r_10_0_entries_perms_0_x; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_perms_0_w <= l3_io_rresp_data_0_entries_perms_0_w; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_perms_0_w <= r_10_0_entries_perms_0_w; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_perms_0_r <= l3_io_rresp_data_0_entries_perms_0_r; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_perms_0_r <= r_10_0_entries_perms_0_r; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_perms_1_d <= l3_io_rresp_data_0_entries_perms_1_d; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_perms_1_d <= r_10_0_entries_perms_1_d; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_perms_1_a <= l3_io_rresp_data_0_entries_perms_1_a; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_perms_1_a <= r_10_0_entries_perms_1_a; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_perms_1_g <= l3_io_rresp_data_0_entries_perms_1_g; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_perms_1_g <= r_10_0_entries_perms_1_g; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_perms_1_u <= l3_io_rresp_data_0_entries_perms_1_u; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_perms_1_u <= r_10_0_entries_perms_1_u; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_perms_1_x <= l3_io_rresp_data_0_entries_perms_1_x; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_perms_1_x <= r_10_0_entries_perms_1_x; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_perms_1_w <= l3_io_rresp_data_0_entries_perms_1_w; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_perms_1_w <= r_10_0_entries_perms_1_w; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_perms_1_r <= l3_io_rresp_data_0_entries_perms_1_r; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_perms_1_r <= r_10_0_entries_perms_1_r; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_perms_2_d <= l3_io_rresp_data_0_entries_perms_2_d; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_perms_2_d <= r_10_0_entries_perms_2_d; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_perms_2_a <= l3_io_rresp_data_0_entries_perms_2_a; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_perms_2_a <= r_10_0_entries_perms_2_a; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_perms_2_g <= l3_io_rresp_data_0_entries_perms_2_g; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_perms_2_g <= r_10_0_entries_perms_2_g; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_perms_2_u <= l3_io_rresp_data_0_entries_perms_2_u; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_perms_2_u <= r_10_0_entries_perms_2_u; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_perms_2_x <= l3_io_rresp_data_0_entries_perms_2_x; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_perms_2_x <= r_10_0_entries_perms_2_x; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_perms_2_w <= l3_io_rresp_data_0_entries_perms_2_w; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_perms_2_w <= r_10_0_entries_perms_2_w; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_perms_2_r <= l3_io_rresp_data_0_entries_perms_2_r; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_perms_2_r <= r_10_0_entries_perms_2_r; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_perms_3_d <= l3_io_rresp_data_0_entries_perms_3_d; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_perms_3_d <= r_10_0_entries_perms_3_d; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_perms_3_a <= l3_io_rresp_data_0_entries_perms_3_a; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_perms_3_a <= r_10_0_entries_perms_3_a; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_perms_3_g <= l3_io_rresp_data_0_entries_perms_3_g; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_perms_3_g <= r_10_0_entries_perms_3_g; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_perms_3_u <= l3_io_rresp_data_0_entries_perms_3_u; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_perms_3_u <= r_10_0_entries_perms_3_u; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_perms_3_x <= l3_io_rresp_data_0_entries_perms_3_x; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_perms_3_x <= r_10_0_entries_perms_3_x; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_perms_3_w <= l3_io_rresp_data_0_entries_perms_3_w; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_perms_3_w <= r_10_0_entries_perms_3_w; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_perms_3_r <= l3_io_rresp_data_0_entries_perms_3_r; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_perms_3_r <= r_10_0_entries_perms_3_r; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_perms_4_d <= l3_io_rresp_data_0_entries_perms_4_d; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_perms_4_d <= r_10_0_entries_perms_4_d; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_perms_4_a <= l3_io_rresp_data_0_entries_perms_4_a; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_perms_4_a <= r_10_0_entries_perms_4_a; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_perms_4_g <= l3_io_rresp_data_0_entries_perms_4_g; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_perms_4_g <= r_10_0_entries_perms_4_g; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_perms_4_u <= l3_io_rresp_data_0_entries_perms_4_u; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_perms_4_u <= r_10_0_entries_perms_4_u; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_perms_4_x <= l3_io_rresp_data_0_entries_perms_4_x; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_perms_4_x <= r_10_0_entries_perms_4_x; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_perms_4_w <= l3_io_rresp_data_0_entries_perms_4_w; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_perms_4_w <= r_10_0_entries_perms_4_w; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_perms_4_r <= l3_io_rresp_data_0_entries_perms_4_r; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_perms_4_r <= r_10_0_entries_perms_4_r; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_perms_5_d <= l3_io_rresp_data_0_entries_perms_5_d; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_perms_5_d <= r_10_0_entries_perms_5_d; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_perms_5_a <= l3_io_rresp_data_0_entries_perms_5_a; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_perms_5_a <= r_10_0_entries_perms_5_a; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_perms_5_g <= l3_io_rresp_data_0_entries_perms_5_g; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_perms_5_g <= r_10_0_entries_perms_5_g; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_perms_5_u <= l3_io_rresp_data_0_entries_perms_5_u; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_perms_5_u <= r_10_0_entries_perms_5_u; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_perms_5_x <= l3_io_rresp_data_0_entries_perms_5_x; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_perms_5_x <= r_10_0_entries_perms_5_x; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_perms_5_w <= l3_io_rresp_data_0_entries_perms_5_w; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_perms_5_w <= r_10_0_entries_perms_5_w; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_perms_5_r <= l3_io_rresp_data_0_entries_perms_5_r; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_perms_5_r <= r_10_0_entries_perms_5_r; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_perms_6_d <= l3_io_rresp_data_0_entries_perms_6_d; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_perms_6_d <= r_10_0_entries_perms_6_d; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_perms_6_a <= l3_io_rresp_data_0_entries_perms_6_a; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_perms_6_a <= r_10_0_entries_perms_6_a; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_perms_6_g <= l3_io_rresp_data_0_entries_perms_6_g; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_perms_6_g <= r_10_0_entries_perms_6_g; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_perms_6_u <= l3_io_rresp_data_0_entries_perms_6_u; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_perms_6_u <= r_10_0_entries_perms_6_u; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_perms_6_x <= l3_io_rresp_data_0_entries_perms_6_x; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_perms_6_x <= r_10_0_entries_perms_6_x; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_perms_6_w <= l3_io_rresp_data_0_entries_perms_6_w; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_perms_6_w <= r_10_0_entries_perms_6_w; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_perms_6_r <= l3_io_rresp_data_0_entries_perms_6_r; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_perms_6_r <= r_10_0_entries_perms_6_r; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_perms_7_d <= l3_io_rresp_data_0_entries_perms_7_d; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_perms_7_d <= r_10_0_entries_perms_7_d; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_perms_7_a <= l3_io_rresp_data_0_entries_perms_7_a; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_perms_7_a <= r_10_0_entries_perms_7_a; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_perms_7_g <= l3_io_rresp_data_0_entries_perms_7_g; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_perms_7_g <= r_10_0_entries_perms_7_g; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_perms_7_u <= l3_io_rresp_data_0_entries_perms_7_u; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_perms_7_u <= r_10_0_entries_perms_7_u; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_perms_7_x <= l3_io_rresp_data_0_entries_perms_7_x; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_perms_7_x <= r_10_0_entries_perms_7_x; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_perms_7_w <= l3_io_rresp_data_0_entries_perms_7_w; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_perms_7_w <= r_10_0_entries_perms_7_w; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_perms_7_r <= l3_io_rresp_data_0_entries_perms_7_r; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_perms_7_r <= r_10_0_entries_perms_7_r; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_entries_prefetch <= l3_io_rresp_data_0_entries_prefetch; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_entries_prefetch <= r_10_0_entries_prefetch; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_0_ecc <= l3_io_rresp_data_0_ecc; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_0_ecc <= r_10_0_ecc; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_tag <= l3_io_rresp_data_1_entries_tag; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_tag <= r_10_1_entries_tag; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_asid <= l3_io_rresp_data_1_entries_asid; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_asid <= r_10_1_entries_asid; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_ppns_0 <= l3_io_rresp_data_1_entries_ppns_0; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_ppns_0 <= r_10_1_entries_ppns_0; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_ppns_1 <= l3_io_rresp_data_1_entries_ppns_1; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_ppns_1 <= r_10_1_entries_ppns_1; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_ppns_2 <= l3_io_rresp_data_1_entries_ppns_2; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_ppns_2 <= r_10_1_entries_ppns_2; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_ppns_3 <= l3_io_rresp_data_1_entries_ppns_3; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_ppns_3 <= r_10_1_entries_ppns_3; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_ppns_4 <= l3_io_rresp_data_1_entries_ppns_4; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_ppns_4 <= r_10_1_entries_ppns_4; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_ppns_5 <= l3_io_rresp_data_1_entries_ppns_5; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_ppns_5 <= r_10_1_entries_ppns_5; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_ppns_6 <= l3_io_rresp_data_1_entries_ppns_6; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_ppns_6 <= r_10_1_entries_ppns_6; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_ppns_7 <= l3_io_rresp_data_1_entries_ppns_7; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_ppns_7 <= r_10_1_entries_ppns_7; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_vs_0 <= l3_io_rresp_data_1_entries_vs_0; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_vs_0 <= r_10_1_entries_vs_0; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_vs_1 <= l3_io_rresp_data_1_entries_vs_1; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_vs_1 <= r_10_1_entries_vs_1; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_vs_2 <= l3_io_rresp_data_1_entries_vs_2; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_vs_2 <= r_10_1_entries_vs_2; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_vs_3 <= l3_io_rresp_data_1_entries_vs_3; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_vs_3 <= r_10_1_entries_vs_3; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_vs_4 <= l3_io_rresp_data_1_entries_vs_4; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_vs_4 <= r_10_1_entries_vs_4; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_vs_5 <= l3_io_rresp_data_1_entries_vs_5; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_vs_5 <= r_10_1_entries_vs_5; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_vs_6 <= l3_io_rresp_data_1_entries_vs_6; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_vs_6 <= r_10_1_entries_vs_6; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_vs_7 <= l3_io_rresp_data_1_entries_vs_7; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_vs_7 <= r_10_1_entries_vs_7; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_perms_0_d <= l3_io_rresp_data_1_entries_perms_0_d; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_perms_0_d <= r_10_1_entries_perms_0_d; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_perms_0_a <= l3_io_rresp_data_1_entries_perms_0_a; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_perms_0_a <= r_10_1_entries_perms_0_a; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_perms_0_g <= l3_io_rresp_data_1_entries_perms_0_g; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_perms_0_g <= r_10_1_entries_perms_0_g; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_perms_0_u <= l3_io_rresp_data_1_entries_perms_0_u; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_perms_0_u <= r_10_1_entries_perms_0_u; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_perms_0_x <= l3_io_rresp_data_1_entries_perms_0_x; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_perms_0_x <= r_10_1_entries_perms_0_x; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_perms_0_w <= l3_io_rresp_data_1_entries_perms_0_w; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_perms_0_w <= r_10_1_entries_perms_0_w; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_perms_0_r <= l3_io_rresp_data_1_entries_perms_0_r; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_perms_0_r <= r_10_1_entries_perms_0_r; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_perms_1_d <= l3_io_rresp_data_1_entries_perms_1_d; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_perms_1_d <= r_10_1_entries_perms_1_d; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_perms_1_a <= l3_io_rresp_data_1_entries_perms_1_a; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_perms_1_a <= r_10_1_entries_perms_1_a; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_perms_1_g <= l3_io_rresp_data_1_entries_perms_1_g; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_perms_1_g <= r_10_1_entries_perms_1_g; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_perms_1_u <= l3_io_rresp_data_1_entries_perms_1_u; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_perms_1_u <= r_10_1_entries_perms_1_u; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_perms_1_x <= l3_io_rresp_data_1_entries_perms_1_x; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_perms_1_x <= r_10_1_entries_perms_1_x; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_perms_1_w <= l3_io_rresp_data_1_entries_perms_1_w; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_perms_1_w <= r_10_1_entries_perms_1_w; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_perms_1_r <= l3_io_rresp_data_1_entries_perms_1_r; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_perms_1_r <= r_10_1_entries_perms_1_r; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_perms_2_d <= l3_io_rresp_data_1_entries_perms_2_d; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_perms_2_d <= r_10_1_entries_perms_2_d; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_perms_2_a <= l3_io_rresp_data_1_entries_perms_2_a; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_perms_2_a <= r_10_1_entries_perms_2_a; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_perms_2_g <= l3_io_rresp_data_1_entries_perms_2_g; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_perms_2_g <= r_10_1_entries_perms_2_g; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_perms_2_u <= l3_io_rresp_data_1_entries_perms_2_u; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_perms_2_u <= r_10_1_entries_perms_2_u; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_perms_2_x <= l3_io_rresp_data_1_entries_perms_2_x; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_perms_2_x <= r_10_1_entries_perms_2_x; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_perms_2_w <= l3_io_rresp_data_1_entries_perms_2_w; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_perms_2_w <= r_10_1_entries_perms_2_w; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_perms_2_r <= l3_io_rresp_data_1_entries_perms_2_r; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_perms_2_r <= r_10_1_entries_perms_2_r; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_perms_3_d <= l3_io_rresp_data_1_entries_perms_3_d; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_perms_3_d <= r_10_1_entries_perms_3_d; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_perms_3_a <= l3_io_rresp_data_1_entries_perms_3_a; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_perms_3_a <= r_10_1_entries_perms_3_a; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_perms_3_g <= l3_io_rresp_data_1_entries_perms_3_g; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_perms_3_g <= r_10_1_entries_perms_3_g; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_perms_3_u <= l3_io_rresp_data_1_entries_perms_3_u; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_perms_3_u <= r_10_1_entries_perms_3_u; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_perms_3_x <= l3_io_rresp_data_1_entries_perms_3_x; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_perms_3_x <= r_10_1_entries_perms_3_x; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_perms_3_w <= l3_io_rresp_data_1_entries_perms_3_w; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_perms_3_w <= r_10_1_entries_perms_3_w; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_perms_3_r <= l3_io_rresp_data_1_entries_perms_3_r; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_perms_3_r <= r_10_1_entries_perms_3_r; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_perms_4_d <= l3_io_rresp_data_1_entries_perms_4_d; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_perms_4_d <= r_10_1_entries_perms_4_d; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_perms_4_a <= l3_io_rresp_data_1_entries_perms_4_a; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_perms_4_a <= r_10_1_entries_perms_4_a; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_perms_4_g <= l3_io_rresp_data_1_entries_perms_4_g; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_perms_4_g <= r_10_1_entries_perms_4_g; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_perms_4_u <= l3_io_rresp_data_1_entries_perms_4_u; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_perms_4_u <= r_10_1_entries_perms_4_u; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_perms_4_x <= l3_io_rresp_data_1_entries_perms_4_x; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_perms_4_x <= r_10_1_entries_perms_4_x; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_perms_4_w <= l3_io_rresp_data_1_entries_perms_4_w; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_perms_4_w <= r_10_1_entries_perms_4_w; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_perms_4_r <= l3_io_rresp_data_1_entries_perms_4_r; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_perms_4_r <= r_10_1_entries_perms_4_r; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_perms_5_d <= l3_io_rresp_data_1_entries_perms_5_d; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_perms_5_d <= r_10_1_entries_perms_5_d; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_perms_5_a <= l3_io_rresp_data_1_entries_perms_5_a; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_perms_5_a <= r_10_1_entries_perms_5_a; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_perms_5_g <= l3_io_rresp_data_1_entries_perms_5_g; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_perms_5_g <= r_10_1_entries_perms_5_g; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_perms_5_u <= l3_io_rresp_data_1_entries_perms_5_u; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_perms_5_u <= r_10_1_entries_perms_5_u; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_perms_5_x <= l3_io_rresp_data_1_entries_perms_5_x; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_perms_5_x <= r_10_1_entries_perms_5_x; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_perms_5_w <= l3_io_rresp_data_1_entries_perms_5_w; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_perms_5_w <= r_10_1_entries_perms_5_w; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_perms_5_r <= l3_io_rresp_data_1_entries_perms_5_r; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_perms_5_r <= r_10_1_entries_perms_5_r; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_perms_6_d <= l3_io_rresp_data_1_entries_perms_6_d; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_perms_6_d <= r_10_1_entries_perms_6_d; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_perms_6_a <= l3_io_rresp_data_1_entries_perms_6_a; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_perms_6_a <= r_10_1_entries_perms_6_a; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_perms_6_g <= l3_io_rresp_data_1_entries_perms_6_g; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_perms_6_g <= r_10_1_entries_perms_6_g; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_perms_6_u <= l3_io_rresp_data_1_entries_perms_6_u; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_perms_6_u <= r_10_1_entries_perms_6_u; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_perms_6_x <= l3_io_rresp_data_1_entries_perms_6_x; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_perms_6_x <= r_10_1_entries_perms_6_x; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_perms_6_w <= l3_io_rresp_data_1_entries_perms_6_w; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_perms_6_w <= r_10_1_entries_perms_6_w; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_perms_6_r <= l3_io_rresp_data_1_entries_perms_6_r; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_perms_6_r <= r_10_1_entries_perms_6_r; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_perms_7_d <= l3_io_rresp_data_1_entries_perms_7_d; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_perms_7_d <= r_10_1_entries_perms_7_d; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_perms_7_a <= l3_io_rresp_data_1_entries_perms_7_a; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_perms_7_a <= r_10_1_entries_perms_7_a; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_perms_7_g <= l3_io_rresp_data_1_entries_perms_7_g; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_perms_7_g <= r_10_1_entries_perms_7_g; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_perms_7_u <= l3_io_rresp_data_1_entries_perms_7_u; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_perms_7_u <= r_10_1_entries_perms_7_u; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_perms_7_x <= l3_io_rresp_data_1_entries_perms_7_x; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_perms_7_x <= r_10_1_entries_perms_7_x; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_perms_7_w <= l3_io_rresp_data_1_entries_perms_7_w; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_perms_7_w <= r_10_1_entries_perms_7_w; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_perms_7_r <= l3_io_rresp_data_1_entries_perms_7_r; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_perms_7_r <= r_10_1_entries_perms_7_r; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_entries_prefetch <= l3_io_rresp_data_1_entries_prefetch; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_entries_prefetch <= r_10_1_entries_prefetch; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_1_ecc <= l3_io_rresp_data_1_ecc; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_1_ecc <= r_10_1_ecc; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_tag <= l3_io_rresp_data_2_entries_tag; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_tag <= r_10_2_entries_tag; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_asid <= l3_io_rresp_data_2_entries_asid; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_asid <= r_10_2_entries_asid; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_ppns_0 <= l3_io_rresp_data_2_entries_ppns_0; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_ppns_0 <= r_10_2_entries_ppns_0; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_ppns_1 <= l3_io_rresp_data_2_entries_ppns_1; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_ppns_1 <= r_10_2_entries_ppns_1; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_ppns_2 <= l3_io_rresp_data_2_entries_ppns_2; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_ppns_2 <= r_10_2_entries_ppns_2; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_ppns_3 <= l3_io_rresp_data_2_entries_ppns_3; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_ppns_3 <= r_10_2_entries_ppns_3; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_ppns_4 <= l3_io_rresp_data_2_entries_ppns_4; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_ppns_4 <= r_10_2_entries_ppns_4; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_ppns_5 <= l3_io_rresp_data_2_entries_ppns_5; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_ppns_5 <= r_10_2_entries_ppns_5; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_ppns_6 <= l3_io_rresp_data_2_entries_ppns_6; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_ppns_6 <= r_10_2_entries_ppns_6; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_ppns_7 <= l3_io_rresp_data_2_entries_ppns_7; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_ppns_7 <= r_10_2_entries_ppns_7; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_vs_0 <= l3_io_rresp_data_2_entries_vs_0; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_vs_0 <= r_10_2_entries_vs_0; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_vs_1 <= l3_io_rresp_data_2_entries_vs_1; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_vs_1 <= r_10_2_entries_vs_1; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_vs_2 <= l3_io_rresp_data_2_entries_vs_2; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_vs_2 <= r_10_2_entries_vs_2; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_vs_3 <= l3_io_rresp_data_2_entries_vs_3; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_vs_3 <= r_10_2_entries_vs_3; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_vs_4 <= l3_io_rresp_data_2_entries_vs_4; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_vs_4 <= r_10_2_entries_vs_4; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_vs_5 <= l3_io_rresp_data_2_entries_vs_5; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_vs_5 <= r_10_2_entries_vs_5; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_vs_6 <= l3_io_rresp_data_2_entries_vs_6; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_vs_6 <= r_10_2_entries_vs_6; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_vs_7 <= l3_io_rresp_data_2_entries_vs_7; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_vs_7 <= r_10_2_entries_vs_7; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_perms_0_d <= l3_io_rresp_data_2_entries_perms_0_d; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_perms_0_d <= r_10_2_entries_perms_0_d; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_perms_0_a <= l3_io_rresp_data_2_entries_perms_0_a; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_perms_0_a <= r_10_2_entries_perms_0_a; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_perms_0_g <= l3_io_rresp_data_2_entries_perms_0_g; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_perms_0_g <= r_10_2_entries_perms_0_g; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_perms_0_u <= l3_io_rresp_data_2_entries_perms_0_u; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_perms_0_u <= r_10_2_entries_perms_0_u; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_perms_0_x <= l3_io_rresp_data_2_entries_perms_0_x; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_perms_0_x <= r_10_2_entries_perms_0_x; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_perms_0_w <= l3_io_rresp_data_2_entries_perms_0_w; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_perms_0_w <= r_10_2_entries_perms_0_w; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_perms_0_r <= l3_io_rresp_data_2_entries_perms_0_r; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_perms_0_r <= r_10_2_entries_perms_0_r; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_perms_1_d <= l3_io_rresp_data_2_entries_perms_1_d; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_perms_1_d <= r_10_2_entries_perms_1_d; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_perms_1_a <= l3_io_rresp_data_2_entries_perms_1_a; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_perms_1_a <= r_10_2_entries_perms_1_a; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_perms_1_g <= l3_io_rresp_data_2_entries_perms_1_g; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_perms_1_g <= r_10_2_entries_perms_1_g; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_perms_1_u <= l3_io_rresp_data_2_entries_perms_1_u; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_perms_1_u <= r_10_2_entries_perms_1_u; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_perms_1_x <= l3_io_rresp_data_2_entries_perms_1_x; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_perms_1_x <= r_10_2_entries_perms_1_x; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_perms_1_w <= l3_io_rresp_data_2_entries_perms_1_w; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_perms_1_w <= r_10_2_entries_perms_1_w; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_perms_1_r <= l3_io_rresp_data_2_entries_perms_1_r; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_perms_1_r <= r_10_2_entries_perms_1_r; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_perms_2_d <= l3_io_rresp_data_2_entries_perms_2_d; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_perms_2_d <= r_10_2_entries_perms_2_d; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_perms_2_a <= l3_io_rresp_data_2_entries_perms_2_a; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_perms_2_a <= r_10_2_entries_perms_2_a; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_perms_2_g <= l3_io_rresp_data_2_entries_perms_2_g; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_perms_2_g <= r_10_2_entries_perms_2_g; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_perms_2_u <= l3_io_rresp_data_2_entries_perms_2_u; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_perms_2_u <= r_10_2_entries_perms_2_u; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_perms_2_x <= l3_io_rresp_data_2_entries_perms_2_x; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_perms_2_x <= r_10_2_entries_perms_2_x; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_perms_2_w <= l3_io_rresp_data_2_entries_perms_2_w; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_perms_2_w <= r_10_2_entries_perms_2_w; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_perms_2_r <= l3_io_rresp_data_2_entries_perms_2_r; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_perms_2_r <= r_10_2_entries_perms_2_r; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_perms_3_d <= l3_io_rresp_data_2_entries_perms_3_d; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_perms_3_d <= r_10_2_entries_perms_3_d; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_perms_3_a <= l3_io_rresp_data_2_entries_perms_3_a; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_perms_3_a <= r_10_2_entries_perms_3_a; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_perms_3_g <= l3_io_rresp_data_2_entries_perms_3_g; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_perms_3_g <= r_10_2_entries_perms_3_g; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_perms_3_u <= l3_io_rresp_data_2_entries_perms_3_u; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_perms_3_u <= r_10_2_entries_perms_3_u; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_perms_3_x <= l3_io_rresp_data_2_entries_perms_3_x; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_perms_3_x <= r_10_2_entries_perms_3_x; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_perms_3_w <= l3_io_rresp_data_2_entries_perms_3_w; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_perms_3_w <= r_10_2_entries_perms_3_w; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_perms_3_r <= l3_io_rresp_data_2_entries_perms_3_r; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_perms_3_r <= r_10_2_entries_perms_3_r; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_perms_4_d <= l3_io_rresp_data_2_entries_perms_4_d; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_perms_4_d <= r_10_2_entries_perms_4_d; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_perms_4_a <= l3_io_rresp_data_2_entries_perms_4_a; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_perms_4_a <= r_10_2_entries_perms_4_a; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_perms_4_g <= l3_io_rresp_data_2_entries_perms_4_g; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_perms_4_g <= r_10_2_entries_perms_4_g; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_perms_4_u <= l3_io_rresp_data_2_entries_perms_4_u; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_perms_4_u <= r_10_2_entries_perms_4_u; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_perms_4_x <= l3_io_rresp_data_2_entries_perms_4_x; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_perms_4_x <= r_10_2_entries_perms_4_x; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_perms_4_w <= l3_io_rresp_data_2_entries_perms_4_w; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_perms_4_w <= r_10_2_entries_perms_4_w; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_perms_4_r <= l3_io_rresp_data_2_entries_perms_4_r; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_perms_4_r <= r_10_2_entries_perms_4_r; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_perms_5_d <= l3_io_rresp_data_2_entries_perms_5_d; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_perms_5_d <= r_10_2_entries_perms_5_d; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_perms_5_a <= l3_io_rresp_data_2_entries_perms_5_a; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_perms_5_a <= r_10_2_entries_perms_5_a; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_perms_5_g <= l3_io_rresp_data_2_entries_perms_5_g; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_perms_5_g <= r_10_2_entries_perms_5_g; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_perms_5_u <= l3_io_rresp_data_2_entries_perms_5_u; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_perms_5_u <= r_10_2_entries_perms_5_u; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_perms_5_x <= l3_io_rresp_data_2_entries_perms_5_x; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_perms_5_x <= r_10_2_entries_perms_5_x; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_perms_5_w <= l3_io_rresp_data_2_entries_perms_5_w; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_perms_5_w <= r_10_2_entries_perms_5_w; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_perms_5_r <= l3_io_rresp_data_2_entries_perms_5_r; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_perms_5_r <= r_10_2_entries_perms_5_r; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_perms_6_d <= l3_io_rresp_data_2_entries_perms_6_d; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_perms_6_d <= r_10_2_entries_perms_6_d; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_perms_6_a <= l3_io_rresp_data_2_entries_perms_6_a; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_perms_6_a <= r_10_2_entries_perms_6_a; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_perms_6_g <= l3_io_rresp_data_2_entries_perms_6_g; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_perms_6_g <= r_10_2_entries_perms_6_g; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_perms_6_u <= l3_io_rresp_data_2_entries_perms_6_u; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_perms_6_u <= r_10_2_entries_perms_6_u; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_perms_6_x <= l3_io_rresp_data_2_entries_perms_6_x; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_perms_6_x <= r_10_2_entries_perms_6_x; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_perms_6_w <= l3_io_rresp_data_2_entries_perms_6_w; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_perms_6_w <= r_10_2_entries_perms_6_w; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_perms_6_r <= l3_io_rresp_data_2_entries_perms_6_r; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_perms_6_r <= r_10_2_entries_perms_6_r; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_perms_7_d <= l3_io_rresp_data_2_entries_perms_7_d; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_perms_7_d <= r_10_2_entries_perms_7_d; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_perms_7_a <= l3_io_rresp_data_2_entries_perms_7_a; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_perms_7_a <= r_10_2_entries_perms_7_a; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_perms_7_g <= l3_io_rresp_data_2_entries_perms_7_g; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_perms_7_g <= r_10_2_entries_perms_7_g; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_perms_7_u <= l3_io_rresp_data_2_entries_perms_7_u; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_perms_7_u <= r_10_2_entries_perms_7_u; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_perms_7_x <= l3_io_rresp_data_2_entries_perms_7_x; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_perms_7_x <= r_10_2_entries_perms_7_x; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_perms_7_w <= l3_io_rresp_data_2_entries_perms_7_w; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_perms_7_w <= r_10_2_entries_perms_7_w; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_perms_7_r <= l3_io_rresp_data_2_entries_perms_7_r; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_perms_7_r <= r_10_2_entries_perms_7_r; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_entries_prefetch <= l3_io_rresp_data_2_entries_prefetch; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_entries_prefetch <= r_10_2_entries_prefetch; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_2_ecc <= l3_io_rresp_data_2_ecc; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_2_ecc <= r_10_2_ecc; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_tag <= l3_io_rresp_data_3_entries_tag; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_tag <= r_10_3_entries_tag; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_asid <= l3_io_rresp_data_3_entries_asid; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_asid <= r_10_3_entries_asid; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_ppns_0 <= l3_io_rresp_data_3_entries_ppns_0; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_ppns_0 <= r_10_3_entries_ppns_0; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_ppns_1 <= l3_io_rresp_data_3_entries_ppns_1; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_ppns_1 <= r_10_3_entries_ppns_1; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_ppns_2 <= l3_io_rresp_data_3_entries_ppns_2; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_ppns_2 <= r_10_3_entries_ppns_2; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_ppns_3 <= l3_io_rresp_data_3_entries_ppns_3; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_ppns_3 <= r_10_3_entries_ppns_3; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_ppns_4 <= l3_io_rresp_data_3_entries_ppns_4; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_ppns_4 <= r_10_3_entries_ppns_4; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_ppns_5 <= l3_io_rresp_data_3_entries_ppns_5; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_ppns_5 <= r_10_3_entries_ppns_5; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_ppns_6 <= l3_io_rresp_data_3_entries_ppns_6; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_ppns_6 <= r_10_3_entries_ppns_6; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_ppns_7 <= l3_io_rresp_data_3_entries_ppns_7; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_ppns_7 <= r_10_3_entries_ppns_7; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_vs_0 <= l3_io_rresp_data_3_entries_vs_0; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_vs_0 <= r_10_3_entries_vs_0; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_vs_1 <= l3_io_rresp_data_3_entries_vs_1; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_vs_1 <= r_10_3_entries_vs_1; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_vs_2 <= l3_io_rresp_data_3_entries_vs_2; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_vs_2 <= r_10_3_entries_vs_2; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_vs_3 <= l3_io_rresp_data_3_entries_vs_3; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_vs_3 <= r_10_3_entries_vs_3; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_vs_4 <= l3_io_rresp_data_3_entries_vs_4; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_vs_4 <= r_10_3_entries_vs_4; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_vs_5 <= l3_io_rresp_data_3_entries_vs_5; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_vs_5 <= r_10_3_entries_vs_5; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_vs_6 <= l3_io_rresp_data_3_entries_vs_6; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_vs_6 <= r_10_3_entries_vs_6; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_vs_7 <= l3_io_rresp_data_3_entries_vs_7; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_vs_7 <= r_10_3_entries_vs_7; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_perms_0_d <= l3_io_rresp_data_3_entries_perms_0_d; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_perms_0_d <= r_10_3_entries_perms_0_d; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_perms_0_a <= l3_io_rresp_data_3_entries_perms_0_a; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_perms_0_a <= r_10_3_entries_perms_0_a; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_perms_0_g <= l3_io_rresp_data_3_entries_perms_0_g; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_perms_0_g <= r_10_3_entries_perms_0_g; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_perms_0_u <= l3_io_rresp_data_3_entries_perms_0_u; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_perms_0_u <= r_10_3_entries_perms_0_u; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_perms_0_x <= l3_io_rresp_data_3_entries_perms_0_x; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_perms_0_x <= r_10_3_entries_perms_0_x; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_perms_0_w <= l3_io_rresp_data_3_entries_perms_0_w; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_perms_0_w <= r_10_3_entries_perms_0_w; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_perms_0_r <= l3_io_rresp_data_3_entries_perms_0_r; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_perms_0_r <= r_10_3_entries_perms_0_r; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_perms_1_d <= l3_io_rresp_data_3_entries_perms_1_d; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_perms_1_d <= r_10_3_entries_perms_1_d; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_perms_1_a <= l3_io_rresp_data_3_entries_perms_1_a; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_perms_1_a <= r_10_3_entries_perms_1_a; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_perms_1_g <= l3_io_rresp_data_3_entries_perms_1_g; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_perms_1_g <= r_10_3_entries_perms_1_g; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_perms_1_u <= l3_io_rresp_data_3_entries_perms_1_u; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_perms_1_u <= r_10_3_entries_perms_1_u; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_perms_1_x <= l3_io_rresp_data_3_entries_perms_1_x; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_perms_1_x <= r_10_3_entries_perms_1_x; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_perms_1_w <= l3_io_rresp_data_3_entries_perms_1_w; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_perms_1_w <= r_10_3_entries_perms_1_w; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_perms_1_r <= l3_io_rresp_data_3_entries_perms_1_r; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_perms_1_r <= r_10_3_entries_perms_1_r; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_perms_2_d <= l3_io_rresp_data_3_entries_perms_2_d; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_perms_2_d <= r_10_3_entries_perms_2_d; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_perms_2_a <= l3_io_rresp_data_3_entries_perms_2_a; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_perms_2_a <= r_10_3_entries_perms_2_a; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_perms_2_g <= l3_io_rresp_data_3_entries_perms_2_g; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_perms_2_g <= r_10_3_entries_perms_2_g; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_perms_2_u <= l3_io_rresp_data_3_entries_perms_2_u; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_perms_2_u <= r_10_3_entries_perms_2_u; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_perms_2_x <= l3_io_rresp_data_3_entries_perms_2_x; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_perms_2_x <= r_10_3_entries_perms_2_x; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_perms_2_w <= l3_io_rresp_data_3_entries_perms_2_w; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_perms_2_w <= r_10_3_entries_perms_2_w; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_perms_2_r <= l3_io_rresp_data_3_entries_perms_2_r; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_perms_2_r <= r_10_3_entries_perms_2_r; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_perms_3_d <= l3_io_rresp_data_3_entries_perms_3_d; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_perms_3_d <= r_10_3_entries_perms_3_d; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_perms_3_a <= l3_io_rresp_data_3_entries_perms_3_a; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_perms_3_a <= r_10_3_entries_perms_3_a; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_perms_3_g <= l3_io_rresp_data_3_entries_perms_3_g; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_perms_3_g <= r_10_3_entries_perms_3_g; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_perms_3_u <= l3_io_rresp_data_3_entries_perms_3_u; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_perms_3_u <= r_10_3_entries_perms_3_u; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_perms_3_x <= l3_io_rresp_data_3_entries_perms_3_x; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_perms_3_x <= r_10_3_entries_perms_3_x; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_perms_3_w <= l3_io_rresp_data_3_entries_perms_3_w; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_perms_3_w <= r_10_3_entries_perms_3_w; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_perms_3_r <= l3_io_rresp_data_3_entries_perms_3_r; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_perms_3_r <= r_10_3_entries_perms_3_r; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_perms_4_d <= l3_io_rresp_data_3_entries_perms_4_d; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_perms_4_d <= r_10_3_entries_perms_4_d; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_perms_4_a <= l3_io_rresp_data_3_entries_perms_4_a; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_perms_4_a <= r_10_3_entries_perms_4_a; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_perms_4_g <= l3_io_rresp_data_3_entries_perms_4_g; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_perms_4_g <= r_10_3_entries_perms_4_g; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_perms_4_u <= l3_io_rresp_data_3_entries_perms_4_u; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_perms_4_u <= r_10_3_entries_perms_4_u; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_perms_4_x <= l3_io_rresp_data_3_entries_perms_4_x; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_perms_4_x <= r_10_3_entries_perms_4_x; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_perms_4_w <= l3_io_rresp_data_3_entries_perms_4_w; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_perms_4_w <= r_10_3_entries_perms_4_w; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_perms_4_r <= l3_io_rresp_data_3_entries_perms_4_r; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_perms_4_r <= r_10_3_entries_perms_4_r; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_perms_5_d <= l3_io_rresp_data_3_entries_perms_5_d; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_perms_5_d <= r_10_3_entries_perms_5_d; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_perms_5_a <= l3_io_rresp_data_3_entries_perms_5_a; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_perms_5_a <= r_10_3_entries_perms_5_a; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_perms_5_g <= l3_io_rresp_data_3_entries_perms_5_g; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_perms_5_g <= r_10_3_entries_perms_5_g; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_perms_5_u <= l3_io_rresp_data_3_entries_perms_5_u; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_perms_5_u <= r_10_3_entries_perms_5_u; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_perms_5_x <= l3_io_rresp_data_3_entries_perms_5_x; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_perms_5_x <= r_10_3_entries_perms_5_x; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_perms_5_w <= l3_io_rresp_data_3_entries_perms_5_w; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_perms_5_w <= r_10_3_entries_perms_5_w; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_perms_5_r <= l3_io_rresp_data_3_entries_perms_5_r; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_perms_5_r <= r_10_3_entries_perms_5_r; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_perms_6_d <= l3_io_rresp_data_3_entries_perms_6_d; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_perms_6_d <= r_10_3_entries_perms_6_d; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_perms_6_a <= l3_io_rresp_data_3_entries_perms_6_a; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_perms_6_a <= r_10_3_entries_perms_6_a; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_perms_6_g <= l3_io_rresp_data_3_entries_perms_6_g; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_perms_6_g <= r_10_3_entries_perms_6_g; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_perms_6_u <= l3_io_rresp_data_3_entries_perms_6_u; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_perms_6_u <= r_10_3_entries_perms_6_u; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_perms_6_x <= l3_io_rresp_data_3_entries_perms_6_x; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_perms_6_x <= r_10_3_entries_perms_6_x; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_perms_6_w <= l3_io_rresp_data_3_entries_perms_6_w; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_perms_6_w <= r_10_3_entries_perms_6_w; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_perms_6_r <= l3_io_rresp_data_3_entries_perms_6_r; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_perms_6_r <= r_10_3_entries_perms_6_r; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_perms_7_d <= l3_io_rresp_data_3_entries_perms_7_d; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_perms_7_d <= r_10_3_entries_perms_7_d; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_perms_7_a <= l3_io_rresp_data_3_entries_perms_7_a; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_perms_7_a <= r_10_3_entries_perms_7_a; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_perms_7_g <= l3_io_rresp_data_3_entries_perms_7_g; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_perms_7_g <= r_10_3_entries_perms_7_g; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_perms_7_u <= l3_io_rresp_data_3_entries_perms_7_u; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_perms_7_u <= r_10_3_entries_perms_7_u; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_perms_7_x <= l3_io_rresp_data_3_entries_perms_7_x; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_perms_7_x <= r_10_3_entries_perms_7_x; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_perms_7_w <= l3_io_rresp_data_3_entries_perms_7_w; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_perms_7_w <= r_10_3_entries_perms_7_w; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_perms_7_r <= l3_io_rresp_data_3_entries_perms_7_r; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_perms_7_r <= r_10_3_entries_perms_7_r; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_entries_prefetch <= l3_io_rresp_data_3_entries_prefetch; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_entries_prefetch <= r_10_3_entries_prefetch; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_3_ecc <= l3_io_rresp_data_3_ecc; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_3_ecc <= r_10_3_ecc; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_tag <= l3_io_rresp_data_4_entries_tag; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_tag <= r_10_4_entries_tag; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_asid <= l3_io_rresp_data_4_entries_asid; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_asid <= r_10_4_entries_asid; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_ppns_0 <= l3_io_rresp_data_4_entries_ppns_0; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_ppns_0 <= r_10_4_entries_ppns_0; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_ppns_1 <= l3_io_rresp_data_4_entries_ppns_1; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_ppns_1 <= r_10_4_entries_ppns_1; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_ppns_2 <= l3_io_rresp_data_4_entries_ppns_2; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_ppns_2 <= r_10_4_entries_ppns_2; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_ppns_3 <= l3_io_rresp_data_4_entries_ppns_3; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_ppns_3 <= r_10_4_entries_ppns_3; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_ppns_4 <= l3_io_rresp_data_4_entries_ppns_4; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_ppns_4 <= r_10_4_entries_ppns_4; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_ppns_5 <= l3_io_rresp_data_4_entries_ppns_5; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_ppns_5 <= r_10_4_entries_ppns_5; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_ppns_6 <= l3_io_rresp_data_4_entries_ppns_6; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_ppns_6 <= r_10_4_entries_ppns_6; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_ppns_7 <= l3_io_rresp_data_4_entries_ppns_7; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_ppns_7 <= r_10_4_entries_ppns_7; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_vs_0 <= l3_io_rresp_data_4_entries_vs_0; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_vs_0 <= r_10_4_entries_vs_0; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_vs_1 <= l3_io_rresp_data_4_entries_vs_1; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_vs_1 <= r_10_4_entries_vs_1; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_vs_2 <= l3_io_rresp_data_4_entries_vs_2; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_vs_2 <= r_10_4_entries_vs_2; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_vs_3 <= l3_io_rresp_data_4_entries_vs_3; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_vs_3 <= r_10_4_entries_vs_3; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_vs_4 <= l3_io_rresp_data_4_entries_vs_4; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_vs_4 <= r_10_4_entries_vs_4; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_vs_5 <= l3_io_rresp_data_4_entries_vs_5; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_vs_5 <= r_10_4_entries_vs_5; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_vs_6 <= l3_io_rresp_data_4_entries_vs_6; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_vs_6 <= r_10_4_entries_vs_6; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_vs_7 <= l3_io_rresp_data_4_entries_vs_7; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_vs_7 <= r_10_4_entries_vs_7; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_perms_0_d <= l3_io_rresp_data_4_entries_perms_0_d; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_perms_0_d <= r_10_4_entries_perms_0_d; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_perms_0_a <= l3_io_rresp_data_4_entries_perms_0_a; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_perms_0_a <= r_10_4_entries_perms_0_a; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_perms_0_g <= l3_io_rresp_data_4_entries_perms_0_g; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_perms_0_g <= r_10_4_entries_perms_0_g; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_perms_0_u <= l3_io_rresp_data_4_entries_perms_0_u; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_perms_0_u <= r_10_4_entries_perms_0_u; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_perms_0_x <= l3_io_rresp_data_4_entries_perms_0_x; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_perms_0_x <= r_10_4_entries_perms_0_x; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_perms_0_w <= l3_io_rresp_data_4_entries_perms_0_w; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_perms_0_w <= r_10_4_entries_perms_0_w; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_perms_0_r <= l3_io_rresp_data_4_entries_perms_0_r; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_perms_0_r <= r_10_4_entries_perms_0_r; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_perms_1_d <= l3_io_rresp_data_4_entries_perms_1_d; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_perms_1_d <= r_10_4_entries_perms_1_d; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_perms_1_a <= l3_io_rresp_data_4_entries_perms_1_a; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_perms_1_a <= r_10_4_entries_perms_1_a; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_perms_1_g <= l3_io_rresp_data_4_entries_perms_1_g; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_perms_1_g <= r_10_4_entries_perms_1_g; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_perms_1_u <= l3_io_rresp_data_4_entries_perms_1_u; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_perms_1_u <= r_10_4_entries_perms_1_u; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_perms_1_x <= l3_io_rresp_data_4_entries_perms_1_x; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_perms_1_x <= r_10_4_entries_perms_1_x; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_perms_1_w <= l3_io_rresp_data_4_entries_perms_1_w; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_perms_1_w <= r_10_4_entries_perms_1_w; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_perms_1_r <= l3_io_rresp_data_4_entries_perms_1_r; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_perms_1_r <= r_10_4_entries_perms_1_r; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_perms_2_d <= l3_io_rresp_data_4_entries_perms_2_d; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_perms_2_d <= r_10_4_entries_perms_2_d; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_perms_2_a <= l3_io_rresp_data_4_entries_perms_2_a; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_perms_2_a <= r_10_4_entries_perms_2_a; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_perms_2_g <= l3_io_rresp_data_4_entries_perms_2_g; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_perms_2_g <= r_10_4_entries_perms_2_g; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_perms_2_u <= l3_io_rresp_data_4_entries_perms_2_u; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_perms_2_u <= r_10_4_entries_perms_2_u; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_perms_2_x <= l3_io_rresp_data_4_entries_perms_2_x; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_perms_2_x <= r_10_4_entries_perms_2_x; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_perms_2_w <= l3_io_rresp_data_4_entries_perms_2_w; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_perms_2_w <= r_10_4_entries_perms_2_w; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_perms_2_r <= l3_io_rresp_data_4_entries_perms_2_r; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_perms_2_r <= r_10_4_entries_perms_2_r; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_perms_3_d <= l3_io_rresp_data_4_entries_perms_3_d; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_perms_3_d <= r_10_4_entries_perms_3_d; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_perms_3_a <= l3_io_rresp_data_4_entries_perms_3_a; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_perms_3_a <= r_10_4_entries_perms_3_a; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_perms_3_g <= l3_io_rresp_data_4_entries_perms_3_g; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_perms_3_g <= r_10_4_entries_perms_3_g; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_perms_3_u <= l3_io_rresp_data_4_entries_perms_3_u; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_perms_3_u <= r_10_4_entries_perms_3_u; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_perms_3_x <= l3_io_rresp_data_4_entries_perms_3_x; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_perms_3_x <= r_10_4_entries_perms_3_x; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_perms_3_w <= l3_io_rresp_data_4_entries_perms_3_w; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_perms_3_w <= r_10_4_entries_perms_3_w; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_perms_3_r <= l3_io_rresp_data_4_entries_perms_3_r; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_perms_3_r <= r_10_4_entries_perms_3_r; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_perms_4_d <= l3_io_rresp_data_4_entries_perms_4_d; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_perms_4_d <= r_10_4_entries_perms_4_d; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_perms_4_a <= l3_io_rresp_data_4_entries_perms_4_a; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_perms_4_a <= r_10_4_entries_perms_4_a; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_perms_4_g <= l3_io_rresp_data_4_entries_perms_4_g; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_perms_4_g <= r_10_4_entries_perms_4_g; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_perms_4_u <= l3_io_rresp_data_4_entries_perms_4_u; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_perms_4_u <= r_10_4_entries_perms_4_u; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_perms_4_x <= l3_io_rresp_data_4_entries_perms_4_x; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_perms_4_x <= r_10_4_entries_perms_4_x; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_perms_4_w <= l3_io_rresp_data_4_entries_perms_4_w; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_perms_4_w <= r_10_4_entries_perms_4_w; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_perms_4_r <= l3_io_rresp_data_4_entries_perms_4_r; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_perms_4_r <= r_10_4_entries_perms_4_r; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_perms_5_d <= l3_io_rresp_data_4_entries_perms_5_d; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_perms_5_d <= r_10_4_entries_perms_5_d; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_perms_5_a <= l3_io_rresp_data_4_entries_perms_5_a; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_perms_5_a <= r_10_4_entries_perms_5_a; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_perms_5_g <= l3_io_rresp_data_4_entries_perms_5_g; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_perms_5_g <= r_10_4_entries_perms_5_g; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_perms_5_u <= l3_io_rresp_data_4_entries_perms_5_u; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_perms_5_u <= r_10_4_entries_perms_5_u; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_perms_5_x <= l3_io_rresp_data_4_entries_perms_5_x; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_perms_5_x <= r_10_4_entries_perms_5_x; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_perms_5_w <= l3_io_rresp_data_4_entries_perms_5_w; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_perms_5_w <= r_10_4_entries_perms_5_w; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_perms_5_r <= l3_io_rresp_data_4_entries_perms_5_r; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_perms_5_r <= r_10_4_entries_perms_5_r; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_perms_6_d <= l3_io_rresp_data_4_entries_perms_6_d; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_perms_6_d <= r_10_4_entries_perms_6_d; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_perms_6_a <= l3_io_rresp_data_4_entries_perms_6_a; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_perms_6_a <= r_10_4_entries_perms_6_a; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_perms_6_g <= l3_io_rresp_data_4_entries_perms_6_g; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_perms_6_g <= r_10_4_entries_perms_6_g; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_perms_6_u <= l3_io_rresp_data_4_entries_perms_6_u; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_perms_6_u <= r_10_4_entries_perms_6_u; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_perms_6_x <= l3_io_rresp_data_4_entries_perms_6_x; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_perms_6_x <= r_10_4_entries_perms_6_x; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_perms_6_w <= l3_io_rresp_data_4_entries_perms_6_w; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_perms_6_w <= r_10_4_entries_perms_6_w; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_perms_6_r <= l3_io_rresp_data_4_entries_perms_6_r; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_perms_6_r <= r_10_4_entries_perms_6_r; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_perms_7_d <= l3_io_rresp_data_4_entries_perms_7_d; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_perms_7_d <= r_10_4_entries_perms_7_d; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_perms_7_a <= l3_io_rresp_data_4_entries_perms_7_a; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_perms_7_a <= r_10_4_entries_perms_7_a; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_perms_7_g <= l3_io_rresp_data_4_entries_perms_7_g; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_perms_7_g <= r_10_4_entries_perms_7_g; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_perms_7_u <= l3_io_rresp_data_4_entries_perms_7_u; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_perms_7_u <= r_10_4_entries_perms_7_u; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_perms_7_x <= l3_io_rresp_data_4_entries_perms_7_x; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_perms_7_x <= r_10_4_entries_perms_7_x; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_perms_7_w <= l3_io_rresp_data_4_entries_perms_7_w; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_perms_7_w <= r_10_4_entries_perms_7_w; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_perms_7_r <= l3_io_rresp_data_4_entries_perms_7_r; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_perms_7_r <= r_10_4_entries_perms_7_r; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_entries_prefetch <= l3_io_rresp_data_4_entries_prefetch; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_entries_prefetch <= r_10_4_entries_prefetch; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_4_ecc <= l3_io_rresp_data_4_ecc; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_4_ecc <= r_10_4_ecc; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_tag <= l3_io_rresp_data_5_entries_tag; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_tag <= r_10_5_entries_tag; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_asid <= l3_io_rresp_data_5_entries_asid; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_asid <= r_10_5_entries_asid; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_ppns_0 <= l3_io_rresp_data_5_entries_ppns_0; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_ppns_0 <= r_10_5_entries_ppns_0; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_ppns_1 <= l3_io_rresp_data_5_entries_ppns_1; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_ppns_1 <= r_10_5_entries_ppns_1; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_ppns_2 <= l3_io_rresp_data_5_entries_ppns_2; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_ppns_2 <= r_10_5_entries_ppns_2; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_ppns_3 <= l3_io_rresp_data_5_entries_ppns_3; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_ppns_3 <= r_10_5_entries_ppns_3; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_ppns_4 <= l3_io_rresp_data_5_entries_ppns_4; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_ppns_4 <= r_10_5_entries_ppns_4; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_ppns_5 <= l3_io_rresp_data_5_entries_ppns_5; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_ppns_5 <= r_10_5_entries_ppns_5; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_ppns_6 <= l3_io_rresp_data_5_entries_ppns_6; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_ppns_6 <= r_10_5_entries_ppns_6; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_ppns_7 <= l3_io_rresp_data_5_entries_ppns_7; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_ppns_7 <= r_10_5_entries_ppns_7; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_vs_0 <= l3_io_rresp_data_5_entries_vs_0; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_vs_0 <= r_10_5_entries_vs_0; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_vs_1 <= l3_io_rresp_data_5_entries_vs_1; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_vs_1 <= r_10_5_entries_vs_1; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_vs_2 <= l3_io_rresp_data_5_entries_vs_2; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_vs_2 <= r_10_5_entries_vs_2; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_vs_3 <= l3_io_rresp_data_5_entries_vs_3; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_vs_3 <= r_10_5_entries_vs_3; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_vs_4 <= l3_io_rresp_data_5_entries_vs_4; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_vs_4 <= r_10_5_entries_vs_4; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_vs_5 <= l3_io_rresp_data_5_entries_vs_5; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_vs_5 <= r_10_5_entries_vs_5; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_vs_6 <= l3_io_rresp_data_5_entries_vs_6; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_vs_6 <= r_10_5_entries_vs_6; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_vs_7 <= l3_io_rresp_data_5_entries_vs_7; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_vs_7 <= r_10_5_entries_vs_7; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_perms_0_d <= l3_io_rresp_data_5_entries_perms_0_d; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_perms_0_d <= r_10_5_entries_perms_0_d; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_perms_0_a <= l3_io_rresp_data_5_entries_perms_0_a; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_perms_0_a <= r_10_5_entries_perms_0_a; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_perms_0_g <= l3_io_rresp_data_5_entries_perms_0_g; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_perms_0_g <= r_10_5_entries_perms_0_g; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_perms_0_u <= l3_io_rresp_data_5_entries_perms_0_u; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_perms_0_u <= r_10_5_entries_perms_0_u; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_perms_0_x <= l3_io_rresp_data_5_entries_perms_0_x; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_perms_0_x <= r_10_5_entries_perms_0_x; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_perms_0_w <= l3_io_rresp_data_5_entries_perms_0_w; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_perms_0_w <= r_10_5_entries_perms_0_w; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_perms_0_r <= l3_io_rresp_data_5_entries_perms_0_r; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_perms_0_r <= r_10_5_entries_perms_0_r; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_perms_1_d <= l3_io_rresp_data_5_entries_perms_1_d; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_perms_1_d <= r_10_5_entries_perms_1_d; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_perms_1_a <= l3_io_rresp_data_5_entries_perms_1_a; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_perms_1_a <= r_10_5_entries_perms_1_a; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_perms_1_g <= l3_io_rresp_data_5_entries_perms_1_g; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_perms_1_g <= r_10_5_entries_perms_1_g; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_perms_1_u <= l3_io_rresp_data_5_entries_perms_1_u; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_perms_1_u <= r_10_5_entries_perms_1_u; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_perms_1_x <= l3_io_rresp_data_5_entries_perms_1_x; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_perms_1_x <= r_10_5_entries_perms_1_x; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_perms_1_w <= l3_io_rresp_data_5_entries_perms_1_w; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_perms_1_w <= r_10_5_entries_perms_1_w; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_perms_1_r <= l3_io_rresp_data_5_entries_perms_1_r; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_perms_1_r <= r_10_5_entries_perms_1_r; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_perms_2_d <= l3_io_rresp_data_5_entries_perms_2_d; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_perms_2_d <= r_10_5_entries_perms_2_d; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_perms_2_a <= l3_io_rresp_data_5_entries_perms_2_a; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_perms_2_a <= r_10_5_entries_perms_2_a; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_perms_2_g <= l3_io_rresp_data_5_entries_perms_2_g; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_perms_2_g <= r_10_5_entries_perms_2_g; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_perms_2_u <= l3_io_rresp_data_5_entries_perms_2_u; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_perms_2_u <= r_10_5_entries_perms_2_u; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_perms_2_x <= l3_io_rresp_data_5_entries_perms_2_x; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_perms_2_x <= r_10_5_entries_perms_2_x; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_perms_2_w <= l3_io_rresp_data_5_entries_perms_2_w; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_perms_2_w <= r_10_5_entries_perms_2_w; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_perms_2_r <= l3_io_rresp_data_5_entries_perms_2_r; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_perms_2_r <= r_10_5_entries_perms_2_r; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_perms_3_d <= l3_io_rresp_data_5_entries_perms_3_d; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_perms_3_d <= r_10_5_entries_perms_3_d; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_perms_3_a <= l3_io_rresp_data_5_entries_perms_3_a; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_perms_3_a <= r_10_5_entries_perms_3_a; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_perms_3_g <= l3_io_rresp_data_5_entries_perms_3_g; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_perms_3_g <= r_10_5_entries_perms_3_g; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_perms_3_u <= l3_io_rresp_data_5_entries_perms_3_u; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_perms_3_u <= r_10_5_entries_perms_3_u; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_perms_3_x <= l3_io_rresp_data_5_entries_perms_3_x; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_perms_3_x <= r_10_5_entries_perms_3_x; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_perms_3_w <= l3_io_rresp_data_5_entries_perms_3_w; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_perms_3_w <= r_10_5_entries_perms_3_w; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_perms_3_r <= l3_io_rresp_data_5_entries_perms_3_r; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_perms_3_r <= r_10_5_entries_perms_3_r; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_perms_4_d <= l3_io_rresp_data_5_entries_perms_4_d; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_perms_4_d <= r_10_5_entries_perms_4_d; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_perms_4_a <= l3_io_rresp_data_5_entries_perms_4_a; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_perms_4_a <= r_10_5_entries_perms_4_a; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_perms_4_g <= l3_io_rresp_data_5_entries_perms_4_g; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_perms_4_g <= r_10_5_entries_perms_4_g; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_perms_4_u <= l3_io_rresp_data_5_entries_perms_4_u; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_perms_4_u <= r_10_5_entries_perms_4_u; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_perms_4_x <= l3_io_rresp_data_5_entries_perms_4_x; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_perms_4_x <= r_10_5_entries_perms_4_x; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_perms_4_w <= l3_io_rresp_data_5_entries_perms_4_w; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_perms_4_w <= r_10_5_entries_perms_4_w; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_perms_4_r <= l3_io_rresp_data_5_entries_perms_4_r; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_perms_4_r <= r_10_5_entries_perms_4_r; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_perms_5_d <= l3_io_rresp_data_5_entries_perms_5_d; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_perms_5_d <= r_10_5_entries_perms_5_d; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_perms_5_a <= l3_io_rresp_data_5_entries_perms_5_a; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_perms_5_a <= r_10_5_entries_perms_5_a; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_perms_5_g <= l3_io_rresp_data_5_entries_perms_5_g; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_perms_5_g <= r_10_5_entries_perms_5_g; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_perms_5_u <= l3_io_rresp_data_5_entries_perms_5_u; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_perms_5_u <= r_10_5_entries_perms_5_u; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_perms_5_x <= l3_io_rresp_data_5_entries_perms_5_x; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_perms_5_x <= r_10_5_entries_perms_5_x; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_perms_5_w <= l3_io_rresp_data_5_entries_perms_5_w; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_perms_5_w <= r_10_5_entries_perms_5_w; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_perms_5_r <= l3_io_rresp_data_5_entries_perms_5_r; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_perms_5_r <= r_10_5_entries_perms_5_r; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_perms_6_d <= l3_io_rresp_data_5_entries_perms_6_d; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_perms_6_d <= r_10_5_entries_perms_6_d; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_perms_6_a <= l3_io_rresp_data_5_entries_perms_6_a; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_perms_6_a <= r_10_5_entries_perms_6_a; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_perms_6_g <= l3_io_rresp_data_5_entries_perms_6_g; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_perms_6_g <= r_10_5_entries_perms_6_g; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_perms_6_u <= l3_io_rresp_data_5_entries_perms_6_u; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_perms_6_u <= r_10_5_entries_perms_6_u; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_perms_6_x <= l3_io_rresp_data_5_entries_perms_6_x; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_perms_6_x <= r_10_5_entries_perms_6_x; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_perms_6_w <= l3_io_rresp_data_5_entries_perms_6_w; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_perms_6_w <= r_10_5_entries_perms_6_w; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_perms_6_r <= l3_io_rresp_data_5_entries_perms_6_r; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_perms_6_r <= r_10_5_entries_perms_6_r; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_perms_7_d <= l3_io_rresp_data_5_entries_perms_7_d; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_perms_7_d <= r_10_5_entries_perms_7_d; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_perms_7_a <= l3_io_rresp_data_5_entries_perms_7_a; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_perms_7_a <= r_10_5_entries_perms_7_a; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_perms_7_g <= l3_io_rresp_data_5_entries_perms_7_g; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_perms_7_g <= r_10_5_entries_perms_7_g; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_perms_7_u <= l3_io_rresp_data_5_entries_perms_7_u; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_perms_7_u <= r_10_5_entries_perms_7_u; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_perms_7_x <= l3_io_rresp_data_5_entries_perms_7_x; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_perms_7_x <= r_10_5_entries_perms_7_x; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_perms_7_w <= l3_io_rresp_data_5_entries_perms_7_w; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_perms_7_w <= r_10_5_entries_perms_7_w; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_perms_7_r <= l3_io_rresp_data_5_entries_perms_7_r; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_perms_7_r <= r_10_5_entries_perms_7_r; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_entries_prefetch <= l3_io_rresp_data_5_entries_prefetch; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_entries_prefetch <= r_10_5_entries_prefetch; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_5_ecc <= l3_io_rresp_data_5_ecc; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_5_ecc <= r_10_5_ecc; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_tag <= l3_io_rresp_data_6_entries_tag; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_tag <= r_10_6_entries_tag; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_asid <= l3_io_rresp_data_6_entries_asid; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_asid <= r_10_6_entries_asid; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_ppns_0 <= l3_io_rresp_data_6_entries_ppns_0; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_ppns_0 <= r_10_6_entries_ppns_0; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_ppns_1 <= l3_io_rresp_data_6_entries_ppns_1; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_ppns_1 <= r_10_6_entries_ppns_1; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_ppns_2 <= l3_io_rresp_data_6_entries_ppns_2; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_ppns_2 <= r_10_6_entries_ppns_2; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_ppns_3 <= l3_io_rresp_data_6_entries_ppns_3; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_ppns_3 <= r_10_6_entries_ppns_3; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_ppns_4 <= l3_io_rresp_data_6_entries_ppns_4; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_ppns_4 <= r_10_6_entries_ppns_4; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_ppns_5 <= l3_io_rresp_data_6_entries_ppns_5; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_ppns_5 <= r_10_6_entries_ppns_5; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_ppns_6 <= l3_io_rresp_data_6_entries_ppns_6; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_ppns_6 <= r_10_6_entries_ppns_6; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_ppns_7 <= l3_io_rresp_data_6_entries_ppns_7; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_ppns_7 <= r_10_6_entries_ppns_7; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_vs_0 <= l3_io_rresp_data_6_entries_vs_0; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_vs_0 <= r_10_6_entries_vs_0; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_vs_1 <= l3_io_rresp_data_6_entries_vs_1; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_vs_1 <= r_10_6_entries_vs_1; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_vs_2 <= l3_io_rresp_data_6_entries_vs_2; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_vs_2 <= r_10_6_entries_vs_2; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_vs_3 <= l3_io_rresp_data_6_entries_vs_3; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_vs_3 <= r_10_6_entries_vs_3; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_vs_4 <= l3_io_rresp_data_6_entries_vs_4; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_vs_4 <= r_10_6_entries_vs_4; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_vs_5 <= l3_io_rresp_data_6_entries_vs_5; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_vs_5 <= r_10_6_entries_vs_5; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_vs_6 <= l3_io_rresp_data_6_entries_vs_6; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_vs_6 <= r_10_6_entries_vs_6; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_vs_7 <= l3_io_rresp_data_6_entries_vs_7; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_vs_7 <= r_10_6_entries_vs_7; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_perms_0_d <= l3_io_rresp_data_6_entries_perms_0_d; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_perms_0_d <= r_10_6_entries_perms_0_d; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_perms_0_a <= l3_io_rresp_data_6_entries_perms_0_a; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_perms_0_a <= r_10_6_entries_perms_0_a; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_perms_0_g <= l3_io_rresp_data_6_entries_perms_0_g; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_perms_0_g <= r_10_6_entries_perms_0_g; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_perms_0_u <= l3_io_rresp_data_6_entries_perms_0_u; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_perms_0_u <= r_10_6_entries_perms_0_u; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_perms_0_x <= l3_io_rresp_data_6_entries_perms_0_x; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_perms_0_x <= r_10_6_entries_perms_0_x; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_perms_0_w <= l3_io_rresp_data_6_entries_perms_0_w; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_perms_0_w <= r_10_6_entries_perms_0_w; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_perms_0_r <= l3_io_rresp_data_6_entries_perms_0_r; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_perms_0_r <= r_10_6_entries_perms_0_r; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_perms_1_d <= l3_io_rresp_data_6_entries_perms_1_d; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_perms_1_d <= r_10_6_entries_perms_1_d; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_perms_1_a <= l3_io_rresp_data_6_entries_perms_1_a; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_perms_1_a <= r_10_6_entries_perms_1_a; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_perms_1_g <= l3_io_rresp_data_6_entries_perms_1_g; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_perms_1_g <= r_10_6_entries_perms_1_g; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_perms_1_u <= l3_io_rresp_data_6_entries_perms_1_u; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_perms_1_u <= r_10_6_entries_perms_1_u; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_perms_1_x <= l3_io_rresp_data_6_entries_perms_1_x; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_perms_1_x <= r_10_6_entries_perms_1_x; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_perms_1_w <= l3_io_rresp_data_6_entries_perms_1_w; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_perms_1_w <= r_10_6_entries_perms_1_w; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_perms_1_r <= l3_io_rresp_data_6_entries_perms_1_r; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_perms_1_r <= r_10_6_entries_perms_1_r; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_perms_2_d <= l3_io_rresp_data_6_entries_perms_2_d; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_perms_2_d <= r_10_6_entries_perms_2_d; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_perms_2_a <= l3_io_rresp_data_6_entries_perms_2_a; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_perms_2_a <= r_10_6_entries_perms_2_a; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_perms_2_g <= l3_io_rresp_data_6_entries_perms_2_g; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_perms_2_g <= r_10_6_entries_perms_2_g; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_perms_2_u <= l3_io_rresp_data_6_entries_perms_2_u; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_perms_2_u <= r_10_6_entries_perms_2_u; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_perms_2_x <= l3_io_rresp_data_6_entries_perms_2_x; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_perms_2_x <= r_10_6_entries_perms_2_x; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_perms_2_w <= l3_io_rresp_data_6_entries_perms_2_w; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_perms_2_w <= r_10_6_entries_perms_2_w; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_perms_2_r <= l3_io_rresp_data_6_entries_perms_2_r; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_perms_2_r <= r_10_6_entries_perms_2_r; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_perms_3_d <= l3_io_rresp_data_6_entries_perms_3_d; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_perms_3_d <= r_10_6_entries_perms_3_d; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_perms_3_a <= l3_io_rresp_data_6_entries_perms_3_a; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_perms_3_a <= r_10_6_entries_perms_3_a; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_perms_3_g <= l3_io_rresp_data_6_entries_perms_3_g; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_perms_3_g <= r_10_6_entries_perms_3_g; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_perms_3_u <= l3_io_rresp_data_6_entries_perms_3_u; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_perms_3_u <= r_10_6_entries_perms_3_u; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_perms_3_x <= l3_io_rresp_data_6_entries_perms_3_x; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_perms_3_x <= r_10_6_entries_perms_3_x; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_perms_3_w <= l3_io_rresp_data_6_entries_perms_3_w; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_perms_3_w <= r_10_6_entries_perms_3_w; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_perms_3_r <= l3_io_rresp_data_6_entries_perms_3_r; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_perms_3_r <= r_10_6_entries_perms_3_r; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_perms_4_d <= l3_io_rresp_data_6_entries_perms_4_d; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_perms_4_d <= r_10_6_entries_perms_4_d; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_perms_4_a <= l3_io_rresp_data_6_entries_perms_4_a; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_perms_4_a <= r_10_6_entries_perms_4_a; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_perms_4_g <= l3_io_rresp_data_6_entries_perms_4_g; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_perms_4_g <= r_10_6_entries_perms_4_g; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_perms_4_u <= l3_io_rresp_data_6_entries_perms_4_u; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_perms_4_u <= r_10_6_entries_perms_4_u; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_perms_4_x <= l3_io_rresp_data_6_entries_perms_4_x; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_perms_4_x <= r_10_6_entries_perms_4_x; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_perms_4_w <= l3_io_rresp_data_6_entries_perms_4_w; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_perms_4_w <= r_10_6_entries_perms_4_w; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_perms_4_r <= l3_io_rresp_data_6_entries_perms_4_r; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_perms_4_r <= r_10_6_entries_perms_4_r; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_perms_5_d <= l3_io_rresp_data_6_entries_perms_5_d; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_perms_5_d <= r_10_6_entries_perms_5_d; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_perms_5_a <= l3_io_rresp_data_6_entries_perms_5_a; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_perms_5_a <= r_10_6_entries_perms_5_a; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_perms_5_g <= l3_io_rresp_data_6_entries_perms_5_g; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_perms_5_g <= r_10_6_entries_perms_5_g; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_perms_5_u <= l3_io_rresp_data_6_entries_perms_5_u; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_perms_5_u <= r_10_6_entries_perms_5_u; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_perms_5_x <= l3_io_rresp_data_6_entries_perms_5_x; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_perms_5_x <= r_10_6_entries_perms_5_x; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_perms_5_w <= l3_io_rresp_data_6_entries_perms_5_w; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_perms_5_w <= r_10_6_entries_perms_5_w; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_perms_5_r <= l3_io_rresp_data_6_entries_perms_5_r; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_perms_5_r <= r_10_6_entries_perms_5_r; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_perms_6_d <= l3_io_rresp_data_6_entries_perms_6_d; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_perms_6_d <= r_10_6_entries_perms_6_d; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_perms_6_a <= l3_io_rresp_data_6_entries_perms_6_a; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_perms_6_a <= r_10_6_entries_perms_6_a; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_perms_6_g <= l3_io_rresp_data_6_entries_perms_6_g; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_perms_6_g <= r_10_6_entries_perms_6_g; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_perms_6_u <= l3_io_rresp_data_6_entries_perms_6_u; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_perms_6_u <= r_10_6_entries_perms_6_u; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_perms_6_x <= l3_io_rresp_data_6_entries_perms_6_x; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_perms_6_x <= r_10_6_entries_perms_6_x; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_perms_6_w <= l3_io_rresp_data_6_entries_perms_6_w; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_perms_6_w <= r_10_6_entries_perms_6_w; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_perms_6_r <= l3_io_rresp_data_6_entries_perms_6_r; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_perms_6_r <= r_10_6_entries_perms_6_r; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_perms_7_d <= l3_io_rresp_data_6_entries_perms_7_d; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_perms_7_d <= r_10_6_entries_perms_7_d; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_perms_7_a <= l3_io_rresp_data_6_entries_perms_7_a; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_perms_7_a <= r_10_6_entries_perms_7_a; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_perms_7_g <= l3_io_rresp_data_6_entries_perms_7_g; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_perms_7_g <= r_10_6_entries_perms_7_g; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_perms_7_u <= l3_io_rresp_data_6_entries_perms_7_u; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_perms_7_u <= r_10_6_entries_perms_7_u; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_perms_7_x <= l3_io_rresp_data_6_entries_perms_7_x; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_perms_7_x <= r_10_6_entries_perms_7_x; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_perms_7_w <= l3_io_rresp_data_6_entries_perms_7_w; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_perms_7_w <= r_10_6_entries_perms_7_w; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_perms_7_r <= l3_io_rresp_data_6_entries_perms_7_r; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_perms_7_r <= r_10_6_entries_perms_7_r; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_entries_prefetch <= l3_io_rresp_data_6_entries_prefetch; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_entries_prefetch <= r_10_6_entries_prefetch; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_6_ecc <= l3_io_rresp_data_6_ecc; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_6_ecc <= r_10_6_ecc; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_tag <= l3_io_rresp_data_7_entries_tag; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_tag <= r_10_7_entries_tag; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_asid <= l3_io_rresp_data_7_entries_asid; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_asid <= r_10_7_entries_asid; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_ppns_0 <= l3_io_rresp_data_7_entries_ppns_0; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_ppns_0 <= r_10_7_entries_ppns_0; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_ppns_1 <= l3_io_rresp_data_7_entries_ppns_1; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_ppns_1 <= r_10_7_entries_ppns_1; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_ppns_2 <= l3_io_rresp_data_7_entries_ppns_2; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_ppns_2 <= r_10_7_entries_ppns_2; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_ppns_3 <= l3_io_rresp_data_7_entries_ppns_3; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_ppns_3 <= r_10_7_entries_ppns_3; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_ppns_4 <= l3_io_rresp_data_7_entries_ppns_4; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_ppns_4 <= r_10_7_entries_ppns_4; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_ppns_5 <= l3_io_rresp_data_7_entries_ppns_5; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_ppns_5 <= r_10_7_entries_ppns_5; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_ppns_6 <= l3_io_rresp_data_7_entries_ppns_6; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_ppns_6 <= r_10_7_entries_ppns_6; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_ppns_7 <= l3_io_rresp_data_7_entries_ppns_7; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_ppns_7 <= r_10_7_entries_ppns_7; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_vs_0 <= l3_io_rresp_data_7_entries_vs_0; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_vs_0 <= r_10_7_entries_vs_0; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_vs_1 <= l3_io_rresp_data_7_entries_vs_1; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_vs_1 <= r_10_7_entries_vs_1; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_vs_2 <= l3_io_rresp_data_7_entries_vs_2; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_vs_2 <= r_10_7_entries_vs_2; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_vs_3 <= l3_io_rresp_data_7_entries_vs_3; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_vs_3 <= r_10_7_entries_vs_3; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_vs_4 <= l3_io_rresp_data_7_entries_vs_4; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_vs_4 <= r_10_7_entries_vs_4; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_vs_5 <= l3_io_rresp_data_7_entries_vs_5; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_vs_5 <= r_10_7_entries_vs_5; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_vs_6 <= l3_io_rresp_data_7_entries_vs_6; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_vs_6 <= r_10_7_entries_vs_6; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_vs_7 <= l3_io_rresp_data_7_entries_vs_7; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_vs_7 <= r_10_7_entries_vs_7; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_perms_0_d <= l3_io_rresp_data_7_entries_perms_0_d; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_perms_0_d <= r_10_7_entries_perms_0_d; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_perms_0_a <= l3_io_rresp_data_7_entries_perms_0_a; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_perms_0_a <= r_10_7_entries_perms_0_a; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_perms_0_g <= l3_io_rresp_data_7_entries_perms_0_g; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_perms_0_g <= r_10_7_entries_perms_0_g; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_perms_0_u <= l3_io_rresp_data_7_entries_perms_0_u; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_perms_0_u <= r_10_7_entries_perms_0_u; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_perms_0_x <= l3_io_rresp_data_7_entries_perms_0_x; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_perms_0_x <= r_10_7_entries_perms_0_x; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_perms_0_w <= l3_io_rresp_data_7_entries_perms_0_w; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_perms_0_w <= r_10_7_entries_perms_0_w; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_perms_0_r <= l3_io_rresp_data_7_entries_perms_0_r; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_perms_0_r <= r_10_7_entries_perms_0_r; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_perms_1_d <= l3_io_rresp_data_7_entries_perms_1_d; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_perms_1_d <= r_10_7_entries_perms_1_d; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_perms_1_a <= l3_io_rresp_data_7_entries_perms_1_a; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_perms_1_a <= r_10_7_entries_perms_1_a; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_perms_1_g <= l3_io_rresp_data_7_entries_perms_1_g; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_perms_1_g <= r_10_7_entries_perms_1_g; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_perms_1_u <= l3_io_rresp_data_7_entries_perms_1_u; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_perms_1_u <= r_10_7_entries_perms_1_u; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_perms_1_x <= l3_io_rresp_data_7_entries_perms_1_x; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_perms_1_x <= r_10_7_entries_perms_1_x; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_perms_1_w <= l3_io_rresp_data_7_entries_perms_1_w; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_perms_1_w <= r_10_7_entries_perms_1_w; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_perms_1_r <= l3_io_rresp_data_7_entries_perms_1_r; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_perms_1_r <= r_10_7_entries_perms_1_r; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_perms_2_d <= l3_io_rresp_data_7_entries_perms_2_d; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_perms_2_d <= r_10_7_entries_perms_2_d; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_perms_2_a <= l3_io_rresp_data_7_entries_perms_2_a; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_perms_2_a <= r_10_7_entries_perms_2_a; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_perms_2_g <= l3_io_rresp_data_7_entries_perms_2_g; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_perms_2_g <= r_10_7_entries_perms_2_g; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_perms_2_u <= l3_io_rresp_data_7_entries_perms_2_u; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_perms_2_u <= r_10_7_entries_perms_2_u; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_perms_2_x <= l3_io_rresp_data_7_entries_perms_2_x; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_perms_2_x <= r_10_7_entries_perms_2_x; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_perms_2_w <= l3_io_rresp_data_7_entries_perms_2_w; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_perms_2_w <= r_10_7_entries_perms_2_w; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_perms_2_r <= l3_io_rresp_data_7_entries_perms_2_r; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_perms_2_r <= r_10_7_entries_perms_2_r; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_perms_3_d <= l3_io_rresp_data_7_entries_perms_3_d; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_perms_3_d <= r_10_7_entries_perms_3_d; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_perms_3_a <= l3_io_rresp_data_7_entries_perms_3_a; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_perms_3_a <= r_10_7_entries_perms_3_a; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_perms_3_g <= l3_io_rresp_data_7_entries_perms_3_g; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_perms_3_g <= r_10_7_entries_perms_3_g; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_perms_3_u <= l3_io_rresp_data_7_entries_perms_3_u; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_perms_3_u <= r_10_7_entries_perms_3_u; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_perms_3_x <= l3_io_rresp_data_7_entries_perms_3_x; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_perms_3_x <= r_10_7_entries_perms_3_x; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_perms_3_w <= l3_io_rresp_data_7_entries_perms_3_w; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_perms_3_w <= r_10_7_entries_perms_3_w; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_perms_3_r <= l3_io_rresp_data_7_entries_perms_3_r; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_perms_3_r <= r_10_7_entries_perms_3_r; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_perms_4_d <= l3_io_rresp_data_7_entries_perms_4_d; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_perms_4_d <= r_10_7_entries_perms_4_d; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_perms_4_a <= l3_io_rresp_data_7_entries_perms_4_a; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_perms_4_a <= r_10_7_entries_perms_4_a; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_perms_4_g <= l3_io_rresp_data_7_entries_perms_4_g; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_perms_4_g <= r_10_7_entries_perms_4_g; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_perms_4_u <= l3_io_rresp_data_7_entries_perms_4_u; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_perms_4_u <= r_10_7_entries_perms_4_u; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_perms_4_x <= l3_io_rresp_data_7_entries_perms_4_x; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_perms_4_x <= r_10_7_entries_perms_4_x; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_perms_4_w <= l3_io_rresp_data_7_entries_perms_4_w; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_perms_4_w <= r_10_7_entries_perms_4_w; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_perms_4_r <= l3_io_rresp_data_7_entries_perms_4_r; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_perms_4_r <= r_10_7_entries_perms_4_r; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_perms_5_d <= l3_io_rresp_data_7_entries_perms_5_d; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_perms_5_d <= r_10_7_entries_perms_5_d; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_perms_5_a <= l3_io_rresp_data_7_entries_perms_5_a; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_perms_5_a <= r_10_7_entries_perms_5_a; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_perms_5_g <= l3_io_rresp_data_7_entries_perms_5_g; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_perms_5_g <= r_10_7_entries_perms_5_g; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_perms_5_u <= l3_io_rresp_data_7_entries_perms_5_u; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_perms_5_u <= r_10_7_entries_perms_5_u; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_perms_5_x <= l3_io_rresp_data_7_entries_perms_5_x; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_perms_5_x <= r_10_7_entries_perms_5_x; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_perms_5_w <= l3_io_rresp_data_7_entries_perms_5_w; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_perms_5_w <= r_10_7_entries_perms_5_w; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_perms_5_r <= l3_io_rresp_data_7_entries_perms_5_r; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_perms_5_r <= r_10_7_entries_perms_5_r; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_perms_6_d <= l3_io_rresp_data_7_entries_perms_6_d; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_perms_6_d <= r_10_7_entries_perms_6_d; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_perms_6_a <= l3_io_rresp_data_7_entries_perms_6_a; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_perms_6_a <= r_10_7_entries_perms_6_a; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_perms_6_g <= l3_io_rresp_data_7_entries_perms_6_g; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_perms_6_g <= r_10_7_entries_perms_6_g; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_perms_6_u <= l3_io_rresp_data_7_entries_perms_6_u; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_perms_6_u <= r_10_7_entries_perms_6_u; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_perms_6_x <= l3_io_rresp_data_7_entries_perms_6_x; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_perms_6_x <= r_10_7_entries_perms_6_x; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_perms_6_w <= l3_io_rresp_data_7_entries_perms_6_w; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_perms_6_w <= r_10_7_entries_perms_6_w; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_perms_6_r <= l3_io_rresp_data_7_entries_perms_6_r; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_perms_6_r <= r_10_7_entries_perms_6_r; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_perms_7_d <= l3_io_rresp_data_7_entries_perms_7_d; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_perms_7_d <= r_10_7_entries_perms_7_d; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_perms_7_a <= l3_io_rresp_data_7_entries_perms_7_a; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_perms_7_a <= r_10_7_entries_perms_7_a; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_perms_7_g <= l3_io_rresp_data_7_entries_perms_7_g; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_perms_7_g <= r_10_7_entries_perms_7_g; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_perms_7_u <= l3_io_rresp_data_7_entries_perms_7_u; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_perms_7_u <= r_10_7_entries_perms_7_u; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_perms_7_x <= l3_io_rresp_data_7_entries_perms_7_x; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_perms_7_x <= r_10_7_entries_perms_7_x; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_perms_7_w <= l3_io_rresp_data_7_entries_perms_7_w; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_perms_7_w <= r_10_7_entries_perms_7_w; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_perms_7_r <= l3_io_rresp_data_7_entries_perms_7_r; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_perms_7_r <= r_10_7_entries_perms_7_r; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_entries_prefetch <= l3_io_rresp_data_7_entries_prefetch; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_entries_prefetch <= r_10_7_entries_prefetch; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (stageDelay_valid_1cycle) begin // @[Reg.scala 17:18]
        l3_ramDatas_7_ecc <= l3_io_rresp_data_7_ecc; // @[Reg.scala 17:22]
      end else begin
        l3_ramDatas_7_ecc <= r_10_7_ecc; // @[Reg.scala 16:16]
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      l3_hitVec_0 <= _T_158; // @[Reg.scala 17:22]
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      l3_hitVec_1 <= _T_163; // @[Reg.scala 17:22]
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      l3_hitVec_2 <= _T_168; // @[Reg.scala 17:22]
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      l3_hitVec_3 <= _T_173; // @[Reg.scala 17:22]
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      l3_hitVec_4 <= _T_178; // @[Reg.scala 17:22]
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      l3_hitVec_5 <= _T_183; // @[Reg.scala 17:22]
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      l3_hitVec_6 <= _T_188; // @[Reg.scala 17:22]
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      l3_hitVec_7 <= _T_193; // @[Reg.scala 17:22]
    end
    if (_stageDelay_valid_1cycle_T) begin // @[Reg.scala 17:18]
      r_13 <= sp_hitVecT_0; // @[Reg.scala 17:22]
    end
    if (_stageDelay_valid_1cycle_T) begin // @[Reg.scala 17:18]
      r_14 <= sp_hitVecT_1; // @[Reg.scala 17:22]
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      spHit <= _T_268; // @[Reg.scala 17:22]
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (r_13) begin // @[ParallelMux.scala 90:77]
        spHitData_ppn <= sp_0_ppn;
      end else begin
        spHitData_ppn <= sp_1_ppn;
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (r_13) begin // @[ParallelMux.scala 90:77]
        spHitData_perm_d <= sp_0_perm_d;
      end else begin
        spHitData_perm_d <= sp_1_perm_d;
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (r_13) begin // @[ParallelMux.scala 90:77]
        spHitData_perm_a <= sp_0_perm_a;
      end else begin
        spHitData_perm_a <= sp_1_perm_a;
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (r_13) begin // @[ParallelMux.scala 90:77]
        spHitData_perm_g <= sp_0_perm_g;
      end else begin
        spHitData_perm_g <= sp_1_perm_g;
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (r_13) begin // @[ParallelMux.scala 90:77]
        spHitData_perm_u <= sp_0_perm_u;
      end else begin
        spHitData_perm_u <= sp_1_perm_u;
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (r_13) begin // @[ParallelMux.scala 90:77]
        spHitData_perm_x <= sp_0_perm_x;
      end else begin
        spHitData_perm_x <= sp_1_perm_x;
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (r_13) begin // @[ParallelMux.scala 90:77]
        spHitData_perm_w <= sp_0_perm_w;
      end else begin
        spHitData_perm_w <= sp_1_perm_w;
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (r_13) begin // @[ParallelMux.scala 90:77]
        spHitData_perm_r <= sp_0_perm_r;
      end else begin
        spHitData_perm_r <= sp_1_perm_r;
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (r_13) begin // @[ParallelMux.scala 90:77]
        spHitData_level <= sp_0_level;
      end else begin
        spHitData_level <= sp_1_level;
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (r_13) begin // @[ParallelMux.scala 90:77]
        spPre <= sp_0_prefetch;
      end else begin
        spPre <= sp_1_prefetch;
      end
    end
    if (_stageCheck_valid_1cycle_T) begin // @[Reg.scala 17:18]
      if (r_13) begin // @[ParallelMux.scala 90:77]
        spValid <= sp_0_v;
      end else begin
        spValid <= sp_1_v;
      end
    end
    if (_stageResp_valid_1cycle_dup_0_T) begin // @[PageTableCache.scala 384:29]
      resp_res_l1_hit <= l1Hit; // @[PageTableCache.scala 384:40]
    end
    if (_stageResp_valid_1cycle_dup_0_T) begin // @[PageTableCache.scala 384:29]
      resp_res_l1_ppn <= l1HitPPN; // @[PageTableCache.scala 384:40]
    end
    if (_stageResp_valid_1cycle_dup_0_T) begin // @[PageTableCache.scala 384:29]
      resp_res_l2_hit <= check_res_l2_hit; // @[PageTableCache.scala 384:40]
    end
    if (_stageResp_valid_1cycle_dup_0_T) begin // @[PageTableCache.scala 384:29]
      if (3'h7 == data_1_req_info_vpn[11:9]) begin // @[PageTableCache.scala 49:14]
        if (l2_hitVec_0 | l2_hitVec_1) begin // @[ParallelMux.scala 90:77]
          if (l2_hitVec_0) begin // @[ParallelMux.scala 90:77]
            resp_res_l2_ppn <= l2_ramDatas_0_entries_ppns_7;
          end else begin
            resp_res_l2_ppn <= l2_ramDatas_1_entries_ppns_7;
          end
        end else if (l2_hitVec_2) begin // @[ParallelMux.scala 90:77]
          resp_res_l2_ppn <= l2_ramDatas_2_entries_ppns_7;
        end else begin
          resp_res_l2_ppn <= l2_ramDatas_3_entries_ppns_7;
        end
      end else if (3'h6 == data_1_req_info_vpn[11:9]) begin // @[PageTableCache.scala 49:14]
        if (l2_hitVec_0 | l2_hitVec_1) begin // @[ParallelMux.scala 90:77]
          resp_res_l2_ppn <= _T_114_entries_ppns_6;
        end else begin
          resp_res_l2_ppn <= _T_116_entries_ppns_6;
        end
      end else if (3'h5 == data_1_req_info_vpn[11:9]) begin // @[PageTableCache.scala 49:14]
        resp_res_l2_ppn <= _T_118_entries_ppns_5; // @[PageTableCache.scala 49:14]
      end else begin
        resp_res_l2_ppn <= _GEN_1541;
      end
    end
    if (_stageResp_valid_1cycle_dup_0_T) begin // @[PageTableCache.scala 384:29]
      resp_res_l2_ecc <= check_res_l2_ecc; // @[PageTableCache.scala 384:40]
    end
    if (_stageResp_valid_1cycle_dup_0_T) begin // @[PageTableCache.scala 384:29]
      resp_res_l3_hit <= check_res_l3_hit; // @[PageTableCache.scala 384:40]
    end
    if (_stageResp_valid_1cycle_dup_0_T) begin // @[PageTableCache.scala 384:29]
      if (l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3)) begin // @[ParallelMux.scala 90:77]
        if (l3_hitVec_0 | l3_hitVec_1) begin // @[ParallelMux.scala 90:77]
          if (l3_hitVec_0) begin // @[ParallelMux.scala 90:77]
            resp_res_l3_pre <= l3_ramDatas_0_entries_prefetch;
          end else begin
            resp_res_l3_pre <= l3_ramDatas_1_entries_prefetch;
          end
        end else if (l3_hitVec_2) begin // @[ParallelMux.scala 90:77]
          resp_res_l3_pre <= l3_ramDatas_2_entries_prefetch;
        end else begin
          resp_res_l3_pre <= l3_ramDatas_3_entries_prefetch;
        end
      end else if (l3_hitVec_4 | l3_hitVec_5) begin // @[ParallelMux.scala 90:77]
        if (l3_hitVec_4) begin // @[ParallelMux.scala 90:77]
          resp_res_l3_pre <= l3_ramDatas_4_entries_prefetch;
        end else begin
          resp_res_l3_pre <= l3_ramDatas_5_entries_prefetch;
        end
      end else if (l3_hitVec_6) begin // @[ParallelMux.scala 90:77]
        resp_res_l3_pre <= l3_ramDatas_6_entries_prefetch;
      end else begin
        resp_res_l3_pre <= l3_ramDatas_7_entries_prefetch;
      end
    end
    if (_stageResp_valid_1cycle_dup_0_T) begin // @[PageTableCache.scala 384:29]
      if (3'h7 == data_1_req_info_vpn[2:0]) begin // @[PageTableCache.scala 49:14]
        if (l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3)) begin // @[ParallelMux.scala 90:77]
          if (l3_hitVec_0 | l3_hitVec_1) begin // @[ParallelMux.scala 90:77]
            resp_res_l3_ppn <= _T_206_entries_ppns_7;
          end else begin
            resp_res_l3_ppn <= _T_208_entries_ppns_7;
          end
        end else if (l3_hitVec_4 | l3_hitVec_5) begin // @[ParallelMux.scala 90:77]
          resp_res_l3_ppn <= _T_212_entries_ppns_7;
        end else begin
          resp_res_l3_ppn <= _T_214_entries_ppns_7;
        end
      end else if (3'h6 == data_1_req_info_vpn[2:0]) begin // @[PageTableCache.scala 49:14]
        if (l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3)) begin // @[ParallelMux.scala 90:77]
          resp_res_l3_ppn <= _T_210_entries_ppns_6;
        end else begin
          resp_res_l3_ppn <= _T_216_entries_ppns_6;
        end
      end else if (3'h5 == data_1_req_info_vpn[2:0]) begin // @[PageTableCache.scala 49:14]
        resp_res_l3_ppn <= _T_218_entries_ppns_5; // @[PageTableCache.scala 49:14]
      end else begin
        resp_res_l3_ppn <= _GEN_1549;
      end
    end
    if (_stageResp_valid_1cycle_dup_0_T) begin // @[PageTableCache.scala 384:29]
      if (3'h7 == data_1_req_info_vpn[2:0]) begin // @[PageTableCache.scala 50:15]
        if (l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3)) begin // @[ParallelMux.scala 90:77]
          if (l3_hitVec_0 | l3_hitVec_1) begin // @[ParallelMux.scala 90:77]
            resp_res_l3_perm_d <= _T_206_entries_perms_7_d;
          end else begin
            resp_res_l3_perm_d <= _T_208_entries_perms_7_d;
          end
        end else if (l3_hitVec_4 | l3_hitVec_5) begin // @[ParallelMux.scala 90:77]
          resp_res_l3_perm_d <= _T_212_entries_perms_7_d;
        end else begin
          resp_res_l3_perm_d <= _T_214_entries_perms_7_d;
        end
      end else if (3'h6 == data_1_req_info_vpn[2:0]) begin // @[PageTableCache.scala 50:15]
        if (l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3)) begin // @[ParallelMux.scala 90:77]
          resp_res_l3_perm_d <= _T_210_entries_perms_6_d;
        end else begin
          resp_res_l3_perm_d <= _T_216_entries_perms_6_d;
        end
      end else if (3'h5 == data_1_req_info_vpn[2:0]) begin // @[PageTableCache.scala 50:15]
        resp_res_l3_perm_d <= _T_218_entries_perms_5_d; // @[PageTableCache.scala 50:15]
      end else begin
        resp_res_l3_perm_d <= _GEN_1557;
      end
    end
    if (_stageResp_valid_1cycle_dup_0_T) begin // @[PageTableCache.scala 384:29]
      if (3'h7 == data_1_req_info_vpn[2:0]) begin // @[PageTableCache.scala 50:15]
        if (l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3)) begin // @[ParallelMux.scala 90:77]
          if (l3_hitVec_0 | l3_hitVec_1) begin // @[ParallelMux.scala 90:77]
            resp_res_l3_perm_a <= _T_206_entries_perms_7_a;
          end else begin
            resp_res_l3_perm_a <= _T_208_entries_perms_7_a;
          end
        end else if (l3_hitVec_4 | l3_hitVec_5) begin // @[ParallelMux.scala 90:77]
          resp_res_l3_perm_a <= _T_212_entries_perms_7_a;
        end else begin
          resp_res_l3_perm_a <= _T_214_entries_perms_7_a;
        end
      end else if (3'h6 == data_1_req_info_vpn[2:0]) begin // @[PageTableCache.scala 50:15]
        if (l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3)) begin // @[ParallelMux.scala 90:77]
          resp_res_l3_perm_a <= _T_210_entries_perms_6_a;
        end else begin
          resp_res_l3_perm_a <= _T_216_entries_perms_6_a;
        end
      end else if (3'h5 == data_1_req_info_vpn[2:0]) begin // @[PageTableCache.scala 50:15]
        resp_res_l3_perm_a <= _T_218_entries_perms_5_a; // @[PageTableCache.scala 50:15]
      end else begin
        resp_res_l3_perm_a <= _GEN_1565;
      end
    end
    if (_stageResp_valid_1cycle_dup_0_T) begin // @[PageTableCache.scala 384:29]
      if (3'h7 == data_1_req_info_vpn[2:0]) begin // @[PageTableCache.scala 50:15]
        if (l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3)) begin // @[ParallelMux.scala 90:77]
          if (l3_hitVec_0 | l3_hitVec_1) begin // @[ParallelMux.scala 90:77]
            resp_res_l3_perm_g <= _T_206_entries_perms_7_g;
          end else begin
            resp_res_l3_perm_g <= _T_208_entries_perms_7_g;
          end
        end else if (l3_hitVec_4 | l3_hitVec_5) begin // @[ParallelMux.scala 90:77]
          resp_res_l3_perm_g <= _T_212_entries_perms_7_g;
        end else begin
          resp_res_l3_perm_g <= _T_214_entries_perms_7_g;
        end
      end else if (3'h6 == data_1_req_info_vpn[2:0]) begin // @[PageTableCache.scala 50:15]
        if (l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3)) begin // @[ParallelMux.scala 90:77]
          resp_res_l3_perm_g <= _T_210_entries_perms_6_g;
        end else begin
          resp_res_l3_perm_g <= _T_216_entries_perms_6_g;
        end
      end else if (3'h5 == data_1_req_info_vpn[2:0]) begin // @[PageTableCache.scala 50:15]
        resp_res_l3_perm_g <= _T_218_entries_perms_5_g; // @[PageTableCache.scala 50:15]
      end else begin
        resp_res_l3_perm_g <= _GEN_1573;
      end
    end
    if (_stageResp_valid_1cycle_dup_0_T) begin // @[PageTableCache.scala 384:29]
      if (3'h7 == data_1_req_info_vpn[2:0]) begin // @[PageTableCache.scala 50:15]
        if (l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3)) begin // @[ParallelMux.scala 90:77]
          if (l3_hitVec_0 | l3_hitVec_1) begin // @[ParallelMux.scala 90:77]
            resp_res_l3_perm_u <= _T_206_entries_perms_7_u;
          end else begin
            resp_res_l3_perm_u <= _T_208_entries_perms_7_u;
          end
        end else if (l3_hitVec_4 | l3_hitVec_5) begin // @[ParallelMux.scala 90:77]
          resp_res_l3_perm_u <= _T_212_entries_perms_7_u;
        end else begin
          resp_res_l3_perm_u <= _T_214_entries_perms_7_u;
        end
      end else if (3'h6 == data_1_req_info_vpn[2:0]) begin // @[PageTableCache.scala 50:15]
        if (l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3)) begin // @[ParallelMux.scala 90:77]
          resp_res_l3_perm_u <= _T_210_entries_perms_6_u;
        end else begin
          resp_res_l3_perm_u <= _T_216_entries_perms_6_u;
        end
      end else if (3'h5 == data_1_req_info_vpn[2:0]) begin // @[PageTableCache.scala 50:15]
        resp_res_l3_perm_u <= _T_218_entries_perms_5_u; // @[PageTableCache.scala 50:15]
      end else begin
        resp_res_l3_perm_u <= _GEN_1581;
      end
    end
    if (_stageResp_valid_1cycle_dup_0_T) begin // @[PageTableCache.scala 384:29]
      if (3'h7 == data_1_req_info_vpn[2:0]) begin // @[PageTableCache.scala 50:15]
        if (l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3)) begin // @[ParallelMux.scala 90:77]
          if (l3_hitVec_0 | l3_hitVec_1) begin // @[ParallelMux.scala 90:77]
            resp_res_l3_perm_x <= _T_206_entries_perms_7_x;
          end else begin
            resp_res_l3_perm_x <= _T_208_entries_perms_7_x;
          end
        end else if (l3_hitVec_4 | l3_hitVec_5) begin // @[ParallelMux.scala 90:77]
          resp_res_l3_perm_x <= _T_212_entries_perms_7_x;
        end else begin
          resp_res_l3_perm_x <= _T_214_entries_perms_7_x;
        end
      end else if (3'h6 == data_1_req_info_vpn[2:0]) begin // @[PageTableCache.scala 50:15]
        if (l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3)) begin // @[ParallelMux.scala 90:77]
          resp_res_l3_perm_x <= _T_210_entries_perms_6_x;
        end else begin
          resp_res_l3_perm_x <= _T_216_entries_perms_6_x;
        end
      end else if (3'h5 == data_1_req_info_vpn[2:0]) begin // @[PageTableCache.scala 50:15]
        resp_res_l3_perm_x <= _T_218_entries_perms_5_x; // @[PageTableCache.scala 50:15]
      end else begin
        resp_res_l3_perm_x <= _GEN_1589;
      end
    end
    if (_stageResp_valid_1cycle_dup_0_T) begin // @[PageTableCache.scala 384:29]
      if (3'h7 == data_1_req_info_vpn[2:0]) begin // @[PageTableCache.scala 50:15]
        if (l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3)) begin // @[ParallelMux.scala 90:77]
          if (l3_hitVec_0 | l3_hitVec_1) begin // @[ParallelMux.scala 90:77]
            resp_res_l3_perm_w <= _T_206_entries_perms_7_w;
          end else begin
            resp_res_l3_perm_w <= _T_208_entries_perms_7_w;
          end
        end else if (l3_hitVec_4 | l3_hitVec_5) begin // @[ParallelMux.scala 90:77]
          resp_res_l3_perm_w <= _T_212_entries_perms_7_w;
        end else begin
          resp_res_l3_perm_w <= _T_214_entries_perms_7_w;
        end
      end else if (3'h6 == data_1_req_info_vpn[2:0]) begin // @[PageTableCache.scala 50:15]
        if (l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3)) begin // @[ParallelMux.scala 90:77]
          resp_res_l3_perm_w <= _T_210_entries_perms_6_w;
        end else begin
          resp_res_l3_perm_w <= _T_216_entries_perms_6_w;
        end
      end else if (3'h5 == data_1_req_info_vpn[2:0]) begin // @[PageTableCache.scala 50:15]
        resp_res_l3_perm_w <= _T_218_entries_perms_5_w; // @[PageTableCache.scala 50:15]
      end else begin
        resp_res_l3_perm_w <= _GEN_1597;
      end
    end
    if (_stageResp_valid_1cycle_dup_0_T) begin // @[PageTableCache.scala 384:29]
      if (3'h7 == data_1_req_info_vpn[2:0]) begin // @[PageTableCache.scala 50:15]
        if (l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3)) begin // @[ParallelMux.scala 90:77]
          if (l3_hitVec_0 | l3_hitVec_1) begin // @[ParallelMux.scala 90:77]
            resp_res_l3_perm_r <= _T_206_entries_perms_7_r;
          end else begin
            resp_res_l3_perm_r <= _T_208_entries_perms_7_r;
          end
        end else if (l3_hitVec_4 | l3_hitVec_5) begin // @[ParallelMux.scala 90:77]
          resp_res_l3_perm_r <= _T_212_entries_perms_7_r;
        end else begin
          resp_res_l3_perm_r <= _T_214_entries_perms_7_r;
        end
      end else if (3'h6 == data_1_req_info_vpn[2:0]) begin // @[PageTableCache.scala 50:15]
        if (l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3)) begin // @[ParallelMux.scala 90:77]
          resp_res_l3_perm_r <= _T_210_entries_perms_6_r;
        end else begin
          resp_res_l3_perm_r <= _T_216_entries_perms_6_r;
        end
      end else if (3'h5 == data_1_req_info_vpn[2:0]) begin // @[PageTableCache.scala 50:15]
        resp_res_l3_perm_r <= _T_218_entries_perms_5_r; // @[PageTableCache.scala 50:15]
      end else begin
        resp_res_l3_perm_r <= _GEN_1605;
      end
    end
    if (_stageResp_valid_1cycle_dup_0_T) begin // @[PageTableCache.scala 384:29]
      resp_res_l3_ecc <= check_res_l3_ecc; // @[PageTableCache.scala 384:40]
    end
    if (_stageResp_valid_1cycle_dup_0_T) begin // @[PageTableCache.scala 384:29]
      if (3'h7 == data_1_req_info_vpn[2:0]) begin // @[PageTableCache.scala 53:12]
        if (l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3)) begin // @[ParallelMux.scala 90:77]
          if (l3_hitVec_0 | l3_hitVec_1) begin // @[ParallelMux.scala 90:77]
            resp_res_l3_v <= _T_206_entries_vs_7;
          end else begin
            resp_res_l3_v <= _T_208_entries_vs_7;
          end
        end else if (l3_hitVec_4 | l3_hitVec_5) begin // @[ParallelMux.scala 90:77]
          resp_res_l3_v <= _T_212_entries_vs_7;
        end else begin
          resp_res_l3_v <= _T_214_entries_vs_7;
        end
      end else if (3'h6 == data_1_req_info_vpn[2:0]) begin // @[PageTableCache.scala 53:12]
        if (l3_hitVec_0 | l3_hitVec_1 | (l3_hitVec_2 | l3_hitVec_3)) begin // @[ParallelMux.scala 90:77]
          resp_res_l3_v <= _T_210_entries_vs_6;
        end else begin
          resp_res_l3_v <= _T_216_entries_vs_6;
        end
      end else if (3'h5 == data_1_req_info_vpn[2:0]) begin // @[PageTableCache.scala 53:12]
        resp_res_l3_v <= _T_218_entries_vs_5; // @[PageTableCache.scala 53:12]
      end else begin
        resp_res_l3_v <= _GEN_1613;
      end
    end
    if (_stageResp_valid_1cycle_dup_0_T) begin // @[PageTableCache.scala 384:29]
      resp_res_sp_hit <= spHit; // @[PageTableCache.scala 384:40]
    end
    if (_stageResp_valid_1cycle_dup_0_T) begin // @[PageTableCache.scala 384:29]
      resp_res_sp_pre <= spPre; // @[PageTableCache.scala 384:40]
    end
    if (_stageResp_valid_1cycle_dup_0_T) begin // @[PageTableCache.scala 384:29]
      resp_res_sp_ppn <= spHitData_ppn; // @[PageTableCache.scala 384:40]
    end
    if (_stageResp_valid_1cycle_dup_0_T) begin // @[PageTableCache.scala 384:29]
      resp_res_sp_perm_d <= spHitData_perm_d; // @[PageTableCache.scala 384:40]
    end
    if (_stageResp_valid_1cycle_dup_0_T) begin // @[PageTableCache.scala 384:29]
      resp_res_sp_perm_a <= spHitData_perm_a; // @[PageTableCache.scala 384:40]
    end
    if (_stageResp_valid_1cycle_dup_0_T) begin // @[PageTableCache.scala 384:29]
      resp_res_sp_perm_g <= spHitData_perm_g; // @[PageTableCache.scala 384:40]
    end
    if (_stageResp_valid_1cycle_dup_0_T) begin // @[PageTableCache.scala 384:29]
      resp_res_sp_perm_u <= spHitData_perm_u; // @[PageTableCache.scala 384:40]
    end
    if (_stageResp_valid_1cycle_dup_0_T) begin // @[PageTableCache.scala 384:29]
      resp_res_sp_perm_x <= spHitData_perm_x; // @[PageTableCache.scala 384:40]
    end
    if (_stageResp_valid_1cycle_dup_0_T) begin // @[PageTableCache.scala 384:29]
      resp_res_sp_perm_w <= spHitData_perm_w; // @[PageTableCache.scala 384:40]
    end
    if (_stageResp_valid_1cycle_dup_0_T) begin // @[PageTableCache.scala 384:29]
      resp_res_sp_perm_r <= spHitData_perm_r; // @[PageTableCache.scala 384:40]
    end
    if (_stageResp_valid_1cycle_dup_0_T) begin // @[PageTableCache.scala 384:29]
      resp_res_sp_level <= spHitData_level; // @[PageTableCache.scala 384:40]
    end
    if (_stageResp_valid_1cycle_dup_0_T) begin // @[PageTableCache.scala 384:29]
      resp_res_sp_v <= spValid; // @[PageTableCache.scala 384:40]
    end
    io_perf_0_value_REG <= ~_base_valid_access_0_T & _base_valid_access_0_T_2; // @[PageTableCache.scala 673:69]
    io_perf_0_value_REG_1 <= io_perf_0_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_1_value_REG <= l1Hit; // @[PerfCounterUtils.scala 188:35]
    io_perf_1_value_REG_1 <= io_perf_1_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_2_value_REG <= _T_113 | _T_115; // @[ParallelMux.scala 36:53]
    io_perf_2_value_REG_1 <= io_perf_2_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_3_value_REG <= _T_209 | _T_215; // @[ParallelMux.scala 36:53]
    io_perf_3_value_REG_1 <= io_perf_3_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_4_value_REG <= spHit; // @[PerfCounterUtils.scala 188:35]
    io_perf_4_value_REG_1 <= io_perf_4_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_5_value_REG <= _T_217 | spHit; // @[PageTableCache.scala 769:33]
    io_perf_5_value_REG_1 <= io_perf_5_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_6_value_REG <= io_req_valid & _T_565; // @[PageTableCache.scala 770:41]
    io_perf_6_value_REG_1 <= io_perf_6_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_7_value_REG <= io_resp_valid & _T_567; // @[PageTableCache.scala 771:42]
    io_perf_7_value_REG_1 <= io_perf_7_value_REG; // @[PerfCounterUtils.scala 188:27]
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PipelineConnect.scala 112:20]
      valid <= 1'h0; // @[PipelineConnect.scala 112:28]
    end else if (flush) begin
      valid <= 1'h0;
    end else begin
      valid <= _GEN_13;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PipelineConnect.scala 112:20]
      valid_1 <= 1'h0; // @[PipelineConnect.scala 112:28]
    end else if (flush) begin
      valid_1 <= 1'h0;
    end else begin
      valid_1 <= _GEN_28;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PipelineConnect.scala 112:20]
      valid_2 <= 1'h0; // @[PipelineConnect.scala 112:28]
    end else if (flush) begin
      valid_2 <= 1'h0;
    end else begin
      valid_2 <= _GEN_43;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Hold.scala 57:18]
      stageDelay_valid_1cycle <= 1'h0; // @[Hold.scala 57:26]
    end else if (flush) begin
      stageDelay_valid_1cycle <= 1'h0;
    end else begin
      stageDelay_valid_1cycle <= _GEN_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Hold.scala 57:18]
      stageCheck_valid_1cycle <= 1'h0; // @[Hold.scala 57:26]
    end else if (flush) begin
      stageCheck_valid_1cycle <= 1'h0;
    end else begin
      stageCheck_valid_1cycle <= _GEN_4;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Hold.scala 57:18]
      stageResp_valid_1cycle_dup_0_valid <= 1'h0; // @[Hold.scala 57:26]
    end else if (flush) begin
      stageResp_valid_1cycle_dup_0_valid <= 1'h0;
    end else begin
      stageResp_valid_1cycle_dup_0_valid <= _GEN_7;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Hold.scala 57:18]
      stageResp_valid_1cycle_dup_1_valid <= 1'h0; // @[Hold.scala 57:26]
    end else if (flush) begin
      stageResp_valid_1cycle_dup_1_valid <= 1'h0;
    end else begin
      stageResp_valid_1cycle_dup_1_valid <= _GEN_10;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PageTableCache.scala 616:30]
      l1v <= 4'h0; // @[PageTableCache.scala 621:41 622:37 624:13 630:13]
    end else if (io_sfence_dup_0_valid) begin
      if (io_sfence_dup_0_bits_rs1) begin
        if (io_sfence_dup_0_bits_rs2) begin
          l1v <= 4'h0;
        end else begin
          l1v <= _l1v_T_3;
        end
      end else begin
        l1v <= _GEN_1728;
      end
    end else begin
      l1v <= _GEN_1728;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PageTableCache.scala 616:30]
      l2v <= 16'h0; // @[PageTableCache.scala 621:41 622:37 625:13 631:13]
    end else if (io_sfence_dup_0_valid) begin
      if (io_sfence_dup_0_bits_rs1) begin
        if (io_sfence_dup_0_bits_rs2) begin
          l2v <= 16'h0;
        end else begin
          l2v <= _l2v_T_3;
        end
      end else begin
        l2v <= _GEN_2533;
      end
    end else begin
      l2v <= _GEN_2533;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PageTableCache.scala 587:30]
      l3v <= 32'h0; // @[PageTableCache.scala 590:41 591:37 593:13 596:13 606:37 608:13 611:13]
    end else if (io_sfence_dup_3_valid) begin // @[PageTableCache.scala 579:21]
      if (io_sfence_dup_3_bits_rs1) begin // @[PageTableCache.scala 582:9]
        if (io_sfence_dup_3_bits_rs2) begin
          l3v <= 32'h0;
        end else begin
          l3v <= _l3v_T_3;
        end
      end else if (io_sfence_dup_3_bits_rs2) begin
        l3v <= _l3v_T_5;
      end else begin
        l3v <= _l3v_T_8;
      end
    end else if (l3eccFlush) begin // @[PageTableCache.scala 500:66]
      l3v <= _l3v_T_2; // @[PageTableCache.scala 520:9]
    end else if (~flush_dup_2 & io_refill_bits_levelOH_l3 & ~_T_377) begin // @[PageTableCache.scala 185:20]
      l3v <= _l3v_T;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PageTableCache.scala 616:30]
      spv <= 2'h0; // @[PageTableCache.scala 621:41 622:37 626:13 632:13 642:37 644:13 647:13]
    end else if (io_sfence_dup_0_valid) begin // @[PageTableCache.scala 540:129]
      if (io_sfence_dup_0_bits_rs1) begin // @[PageTableCache.scala 552:9]
        if (io_sfence_dup_0_bits_rs2) begin
          spv <= 2'h0;
        end else begin
          spv <= _spv_T_3;
        end
      end else if (io_sfence_dup_0_bits_rs2) begin
        spv <= _spv_T_14;
      end else begin
        spv <= _spv_T_26;
      end
    end else if (_T_296 & io_refill_bits_levelOH_sp & (_T_299 | _T_321) & _T_326) begin // @[PageTableCache.scala 204:20]
      spv <= _spv_T;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PageTableCache.scala 435:129]
      state_reg <= 3'h0; // @[Replacement.scala 172:15]
    end else if (~flush & io_refill_bits_levelOH_l1 & ~_T_299 & ~_T_321 & ~_T_325) begin // @[PageTableCache.scala 239:43]
      state_reg <= _state_reg_T_19; // @[Replacement.scala 172:15]
    end else if (_GEN_57 & stageDelay_valid_1cycle) begin // @[Replacement.scala 168:70]
      state_reg <= _state_reg_T_8;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PageTableCache.scala 462:129]
      state_vec__0 <= 3'h0; // @[Replacement.scala 308:{20,20}]
    end else if (~flush_dup_1 & io_refill_bits_levelOH_l2 & ~_T_336 & ~_T_358 & ~_T_362) begin
      if (2'h0 == l2_refillIdx) begin
        state_vec__0 <= _state_vec_T_40;
      end else begin
        state_vec__0 <= _GEN_272;
      end
    end else begin
      state_vec__0 <= _GEN_272;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PageTableCache.scala 462:129]
      state_vec__1 <= 3'h0; // @[Replacement.scala 308:{20,20}]
    end else if (~flush_dup_1 & io_refill_bits_levelOH_l2 & ~_T_336 & ~_T_358 & ~_T_362) begin
      if (2'h1 == l2_refillIdx) begin
        state_vec__1 <= _state_vec_T_40;
      end else begin
        state_vec__1 <= _GEN_273;
      end
    end else begin
      state_vec__1 <= _GEN_273;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PageTableCache.scala 462:129]
      state_vec__2 <= 3'h0; // @[Replacement.scala 308:{20,20}]
    end else if (~flush_dup_1 & io_refill_bits_levelOH_l2 & ~_T_336 & ~_T_358 & ~_T_362) begin
      if (2'h2 == l2_refillIdx) begin
        state_vec__2 <= _state_vec_T_40;
      end else begin
        state_vec__2 <= _GEN_274;
      end
    end else begin
      state_vec__2 <= _GEN_274;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PageTableCache.scala 462:129]
      state_vec__3 <= 3'h0; // @[Replacement.scala 308:{20,20}]
    end else if (~flush_dup_1 & io_refill_bits_levelOH_l2 & ~_T_336 & ~_T_358 & ~_T_362) begin
      if (2'h3 == l2_refillIdx) begin
        state_vec__3 <= _state_vec_T_40;
      end else begin
        state_vec__3 <= _GEN_275;
      end
    end else begin
      state_vec__3 <= _GEN_275;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PageTableCache.scala 500:66]
      state_vec_1_0 <= 7'h0; // @[Replacement.scala 308:{20,20}]
    end else if (~flush_dup_2 & io_refill_bits_levelOH_l3 & ~_T_377) begin
      if (2'h0 == l3_refillIdx) begin
        state_vec_1_0 <= _state_vec_T_63;
      end else begin
        state_vec_1_0 <= _GEN_1514;
      end
    end else begin
      state_vec_1_0 <= _GEN_1514;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PageTableCache.scala 500:66]
      state_vec_1_1 <= 7'h0; // @[Replacement.scala 308:{20,20}]
    end else if (~flush_dup_2 & io_refill_bits_levelOH_l3 & ~_T_377) begin
      if (2'h1 == l3_refillIdx) begin
        state_vec_1_1 <= _state_vec_T_63;
      end else begin
        state_vec_1_1 <= _GEN_1515;
      end
    end else begin
      state_vec_1_1 <= _GEN_1515;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PageTableCache.scala 500:66]
      state_vec_1_2 <= 7'h0; // @[Replacement.scala 308:{20,20}]
    end else if (~flush_dup_2 & io_refill_bits_levelOH_l3 & ~_T_377) begin
      if (2'h2 == l3_refillIdx) begin
        state_vec_1_2 <= _state_vec_T_63;
      end else begin
        state_vec_1_2 <= _GEN_1516;
      end
    end else begin
      state_vec_1_2 <= _GEN_1516;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PageTableCache.scala 500:66]
      state_vec_1_3 <= 7'h0; // @[Replacement.scala 308:{20,20}]
    end else if (~flush_dup_2 & io_refill_bits_levelOH_l3 & ~_T_377) begin
      if (2'h3 == l3_refillIdx) begin
        state_vec_1_3 <= _state_vec_T_63;
      end else begin
        state_vec_1_3 <= _GEN_1517;
      end
    end else begin
      state_vec_1_3 <= _GEN_1517;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PageTableCache.scala 540:129]
      state_reg_3 <= 1'h0; // @[Replacement.scala 172:15]
    end else if (_T_296 & io_refill_bits_levelOH_sp & (_T_299 | _T_321) & _T_326) begin // @[PageTableCache.scala 358:43]
      state_reg_3 <= _state_reg_T_21; // @[Replacement.scala 172:15]
    end else if (_T_268 & stageDelay_valid_1cycle) begin // @[Replacement.scala 168:70]
      state_reg_3 <= _state_reg_T_10;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Hold.scala 56:17]
      bypassed_0_valid <= 1'h0; // @[Hold.scala 56:25]
    end else begin
      bypassed_0_valid <= _stageResp_valid_1cycle_dup_0_T | _GEN_1669;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[MMUBundle.scala 798:20]
      bypassed_0_valid_1 <= 1'h0; // @[MMUBundle.scala 798:28]
    end else if (_bypassed_0_T_7) begin
      bypassed_0_valid_1 <= 1'h0;
    end else begin
      bypassed_0_valid_1 <= _GEN_1672;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Hold.scala 56:17]
      bypassed_1_valid <= 1'h0; // @[Hold.scala 56:25]
    end else begin
      bypassed_1_valid <= _stageResp_valid_1cycle_dup_0_T | _GEN_1675;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[MMUBundle.scala 798:20]
      bypassed_1_valid_1 <= 1'h0; // @[MMUBundle.scala 798:28]
    end else if (_bypassed_1_T_7) begin
      bypassed_1_valid_1 <= 1'h0;
    end else begin
      bypassed_1_valid_1 <= _GEN_1678;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Hold.scala 56:17]
      bypassed_2_valid <= 1'h0; // @[Hold.scala 56:25]
    end else begin
      bypassed_2_valid <= _stageResp_valid_1cycle_dup_0_T | _GEN_1681;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[MMUBundle.scala 798:20]
      bypassed_2_valid_1 <= 1'h0; // @[MMUBundle.scala 798:28]
    end else if (_bypassed_2_T_7) begin
      bypassed_2_valid_1 <= 1'h0;
    end else begin
      bypassed_2_valid_1 <= _GEN_1684;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  valid_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  valid_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  stageDelay_valid_1cycle = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  stageCheck_valid_1cycle = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  stageResp_valid_1cycle_dup_0_valid = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  stageResp_valid_1cycle_dup_1_valid = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  data_req_info_vpn = _RAND_7[26:0];
  _RAND_8 = {1{`RANDOM}};
  data_req_info_source = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  data_isFirst = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  bypassed_reg = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  bypassed_reg_1 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  bypassed_reg_2 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  data_1_req_info_vpn = _RAND_13[26:0];
  _RAND_14 = {1{`RANDOM}};
  data_1_req_info_source = _RAND_14[1:0];
  _RAND_15 = {1{`RANDOM}};
  data_1_isFirst = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  data_1_bypassed_0 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  data_1_bypassed_1 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  data_1_bypassed_2 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  bypassed_reg_3 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  bypassed_reg_4 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  bypassed_reg_5 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  data_2_req_info_vpn = _RAND_22[26:0];
  _RAND_23 = {1{`RANDOM}};
  data_2_req_info_source = _RAND_23[1:0];
  _RAND_24 = {1{`RANDOM}};
  data_2_isFirst = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  data_2_bypassed_0 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  data_2_bypassed_1 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  data_2_bypassed_2 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  l1_0_tag = _RAND_28[8:0];
  _RAND_29 = {1{`RANDOM}};
  l1_0_asid = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  l1_0_ppn = _RAND_30[23:0];
  _RAND_31 = {1{`RANDOM}};
  l1_1_tag = _RAND_31[8:0];
  _RAND_32 = {1{`RANDOM}};
  l1_1_asid = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  l1_1_ppn = _RAND_33[23:0];
  _RAND_34 = {1{`RANDOM}};
  l1_2_tag = _RAND_34[8:0];
  _RAND_35 = {1{`RANDOM}};
  l1_2_asid = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  l1_2_ppn = _RAND_36[23:0];
  _RAND_37 = {1{`RANDOM}};
  l1_3_tag = _RAND_37[8:0];
  _RAND_38 = {1{`RANDOM}};
  l1_3_asid = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  l1_3_ppn = _RAND_39[23:0];
  _RAND_40 = {1{`RANDOM}};
  l1v = _RAND_40[3:0];
  _RAND_41 = {1{`RANDOM}};
  l1g = _RAND_41[3:0];
  _RAND_42 = {1{`RANDOM}};
  l2v = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  l2g = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  l3v = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  l3g = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  sp_0_tag = _RAND_46[17:0];
  _RAND_47 = {1{`RANDOM}};
  sp_0_asid = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  sp_0_ppn = _RAND_48[23:0];
  _RAND_49 = {1{`RANDOM}};
  sp_0_perm_d = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  sp_0_perm_a = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  sp_0_perm_g = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  sp_0_perm_u = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  sp_0_perm_x = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  sp_0_perm_w = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  sp_0_perm_r = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  sp_0_level = _RAND_56[1:0];
  _RAND_57 = {1{`RANDOM}};
  sp_0_prefetch = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  sp_0_v = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  sp_1_tag = _RAND_59[17:0];
  _RAND_60 = {1{`RANDOM}};
  sp_1_asid = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  sp_1_ppn = _RAND_61[23:0];
  _RAND_62 = {1{`RANDOM}};
  sp_1_perm_d = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  sp_1_perm_a = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  sp_1_perm_g = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  sp_1_perm_u = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  sp_1_perm_x = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  sp_1_perm_w = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  sp_1_perm_r = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  sp_1_level = _RAND_69[1:0];
  _RAND_70 = {1{`RANDOM}};
  sp_1_prefetch = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  sp_1_v = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  spv = _RAND_72[1:0];
  _RAND_73 = {1{`RANDOM}};
  spg = _RAND_73[1:0];
  _RAND_74 = {1{`RANDOM}};
  state_reg = _RAND_74[2:0];
  _RAND_75 = {1{`RANDOM}};
  r = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  r_1 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  r_2 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  r_3 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  r_4 = _RAND_79[23:0];
  _RAND_80 = {1{`RANDOM}};
  r_6 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  l1Hit = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  l1HitPPN = _RAND_82[23:0];
  _RAND_83 = {1{`RANDOM}};
  state_vec__0 = _RAND_83[2:0];
  _RAND_84 = {1{`RANDOM}};
  state_vec__1 = _RAND_84[2:0];
  _RAND_85 = {1{`RANDOM}};
  state_vec__2 = _RAND_85[2:0];
  _RAND_86 = {1{`RANDOM}};
  state_vec__3 = _RAND_86[2:0];
  _RAND_87 = {1{`RANDOM}};
  r_7_0_entries_tag = _RAND_87[12:0];
  _RAND_88 = {1{`RANDOM}};
  r_7_0_entries_asid = _RAND_88[15:0];
  _RAND_89 = {1{`RANDOM}};
  r_7_0_entries_ppns_0 = _RAND_89[23:0];
  _RAND_90 = {1{`RANDOM}};
  r_7_0_entries_ppns_1 = _RAND_90[23:0];
  _RAND_91 = {1{`RANDOM}};
  r_7_0_entries_ppns_2 = _RAND_91[23:0];
  _RAND_92 = {1{`RANDOM}};
  r_7_0_entries_ppns_3 = _RAND_92[23:0];
  _RAND_93 = {1{`RANDOM}};
  r_7_0_entries_ppns_4 = _RAND_93[23:0];
  _RAND_94 = {1{`RANDOM}};
  r_7_0_entries_ppns_5 = _RAND_94[23:0];
  _RAND_95 = {1{`RANDOM}};
  r_7_0_entries_ppns_6 = _RAND_95[23:0];
  _RAND_96 = {1{`RANDOM}};
  r_7_0_entries_ppns_7 = _RAND_96[23:0];
  _RAND_97 = {1{`RANDOM}};
  r_7_0_entries_vs_0 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  r_7_0_entries_vs_1 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  r_7_0_entries_vs_2 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  r_7_0_entries_vs_3 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  r_7_0_entries_vs_4 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  r_7_0_entries_vs_5 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  r_7_0_entries_vs_6 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  r_7_0_entries_vs_7 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  r_7_0_entries_prefetch = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  r_7_0_ecc = _RAND_106[30:0];
  _RAND_107 = {1{`RANDOM}};
  r_7_1_entries_tag = _RAND_107[12:0];
  _RAND_108 = {1{`RANDOM}};
  r_7_1_entries_asid = _RAND_108[15:0];
  _RAND_109 = {1{`RANDOM}};
  r_7_1_entries_ppns_0 = _RAND_109[23:0];
  _RAND_110 = {1{`RANDOM}};
  r_7_1_entries_ppns_1 = _RAND_110[23:0];
  _RAND_111 = {1{`RANDOM}};
  r_7_1_entries_ppns_2 = _RAND_111[23:0];
  _RAND_112 = {1{`RANDOM}};
  r_7_1_entries_ppns_3 = _RAND_112[23:0];
  _RAND_113 = {1{`RANDOM}};
  r_7_1_entries_ppns_4 = _RAND_113[23:0];
  _RAND_114 = {1{`RANDOM}};
  r_7_1_entries_ppns_5 = _RAND_114[23:0];
  _RAND_115 = {1{`RANDOM}};
  r_7_1_entries_ppns_6 = _RAND_115[23:0];
  _RAND_116 = {1{`RANDOM}};
  r_7_1_entries_ppns_7 = _RAND_116[23:0];
  _RAND_117 = {1{`RANDOM}};
  r_7_1_entries_vs_0 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  r_7_1_entries_vs_1 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  r_7_1_entries_vs_2 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  r_7_1_entries_vs_3 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  r_7_1_entries_vs_4 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  r_7_1_entries_vs_5 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  r_7_1_entries_vs_6 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  r_7_1_entries_vs_7 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  r_7_1_entries_prefetch = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  r_7_1_ecc = _RAND_126[30:0];
  _RAND_127 = {1{`RANDOM}};
  r_7_2_entries_tag = _RAND_127[12:0];
  _RAND_128 = {1{`RANDOM}};
  r_7_2_entries_asid = _RAND_128[15:0];
  _RAND_129 = {1{`RANDOM}};
  r_7_2_entries_ppns_0 = _RAND_129[23:0];
  _RAND_130 = {1{`RANDOM}};
  r_7_2_entries_ppns_1 = _RAND_130[23:0];
  _RAND_131 = {1{`RANDOM}};
  r_7_2_entries_ppns_2 = _RAND_131[23:0];
  _RAND_132 = {1{`RANDOM}};
  r_7_2_entries_ppns_3 = _RAND_132[23:0];
  _RAND_133 = {1{`RANDOM}};
  r_7_2_entries_ppns_4 = _RAND_133[23:0];
  _RAND_134 = {1{`RANDOM}};
  r_7_2_entries_ppns_5 = _RAND_134[23:0];
  _RAND_135 = {1{`RANDOM}};
  r_7_2_entries_ppns_6 = _RAND_135[23:0];
  _RAND_136 = {1{`RANDOM}};
  r_7_2_entries_ppns_7 = _RAND_136[23:0];
  _RAND_137 = {1{`RANDOM}};
  r_7_2_entries_vs_0 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  r_7_2_entries_vs_1 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  r_7_2_entries_vs_2 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  r_7_2_entries_vs_3 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  r_7_2_entries_vs_4 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  r_7_2_entries_vs_5 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  r_7_2_entries_vs_6 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  r_7_2_entries_vs_7 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  r_7_2_entries_prefetch = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  r_7_2_ecc = _RAND_146[30:0];
  _RAND_147 = {1{`RANDOM}};
  r_7_3_entries_tag = _RAND_147[12:0];
  _RAND_148 = {1{`RANDOM}};
  r_7_3_entries_asid = _RAND_148[15:0];
  _RAND_149 = {1{`RANDOM}};
  r_7_3_entries_ppns_0 = _RAND_149[23:0];
  _RAND_150 = {1{`RANDOM}};
  r_7_3_entries_ppns_1 = _RAND_150[23:0];
  _RAND_151 = {1{`RANDOM}};
  r_7_3_entries_ppns_2 = _RAND_151[23:0];
  _RAND_152 = {1{`RANDOM}};
  r_7_3_entries_ppns_3 = _RAND_152[23:0];
  _RAND_153 = {1{`RANDOM}};
  r_7_3_entries_ppns_4 = _RAND_153[23:0];
  _RAND_154 = {1{`RANDOM}};
  r_7_3_entries_ppns_5 = _RAND_154[23:0];
  _RAND_155 = {1{`RANDOM}};
  r_7_3_entries_ppns_6 = _RAND_155[23:0];
  _RAND_156 = {1{`RANDOM}};
  r_7_3_entries_ppns_7 = _RAND_156[23:0];
  _RAND_157 = {1{`RANDOM}};
  r_7_3_entries_vs_0 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  r_7_3_entries_vs_1 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  r_7_3_entries_vs_2 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  r_7_3_entries_vs_3 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  r_7_3_entries_vs_4 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  r_7_3_entries_vs_5 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  r_7_3_entries_vs_6 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  r_7_3_entries_vs_7 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  r_7_3_entries_prefetch = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  r_7_3_ecc = _RAND_166[30:0];
  _RAND_167 = {1{`RANDOM}};
  r_8 = _RAND_167[3:0];
  _RAND_168 = {1{`RANDOM}};
  l2_ramDatas_0_entries_tag = _RAND_168[12:0];
  _RAND_169 = {1{`RANDOM}};
  l2_ramDatas_0_entries_asid = _RAND_169[15:0];
  _RAND_170 = {1{`RANDOM}};
  l2_ramDatas_0_entries_ppns_0 = _RAND_170[23:0];
  _RAND_171 = {1{`RANDOM}};
  l2_ramDatas_0_entries_ppns_1 = _RAND_171[23:0];
  _RAND_172 = {1{`RANDOM}};
  l2_ramDatas_0_entries_ppns_2 = _RAND_172[23:0];
  _RAND_173 = {1{`RANDOM}};
  l2_ramDatas_0_entries_ppns_3 = _RAND_173[23:0];
  _RAND_174 = {1{`RANDOM}};
  l2_ramDatas_0_entries_ppns_4 = _RAND_174[23:0];
  _RAND_175 = {1{`RANDOM}};
  l2_ramDatas_0_entries_ppns_5 = _RAND_175[23:0];
  _RAND_176 = {1{`RANDOM}};
  l2_ramDatas_0_entries_ppns_6 = _RAND_176[23:0];
  _RAND_177 = {1{`RANDOM}};
  l2_ramDatas_0_entries_ppns_7 = _RAND_177[23:0];
  _RAND_178 = {1{`RANDOM}};
  l2_ramDatas_0_entries_vs_0 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  l2_ramDatas_0_entries_vs_1 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  l2_ramDatas_0_entries_vs_2 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  l2_ramDatas_0_entries_vs_3 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  l2_ramDatas_0_entries_vs_4 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  l2_ramDatas_0_entries_vs_5 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  l2_ramDatas_0_entries_vs_6 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  l2_ramDatas_0_entries_vs_7 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  l2_ramDatas_0_entries_prefetch = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  l2_ramDatas_0_ecc = _RAND_187[30:0];
  _RAND_188 = {1{`RANDOM}};
  l2_ramDatas_1_entries_tag = _RAND_188[12:0];
  _RAND_189 = {1{`RANDOM}};
  l2_ramDatas_1_entries_asid = _RAND_189[15:0];
  _RAND_190 = {1{`RANDOM}};
  l2_ramDatas_1_entries_ppns_0 = _RAND_190[23:0];
  _RAND_191 = {1{`RANDOM}};
  l2_ramDatas_1_entries_ppns_1 = _RAND_191[23:0];
  _RAND_192 = {1{`RANDOM}};
  l2_ramDatas_1_entries_ppns_2 = _RAND_192[23:0];
  _RAND_193 = {1{`RANDOM}};
  l2_ramDatas_1_entries_ppns_3 = _RAND_193[23:0];
  _RAND_194 = {1{`RANDOM}};
  l2_ramDatas_1_entries_ppns_4 = _RAND_194[23:0];
  _RAND_195 = {1{`RANDOM}};
  l2_ramDatas_1_entries_ppns_5 = _RAND_195[23:0];
  _RAND_196 = {1{`RANDOM}};
  l2_ramDatas_1_entries_ppns_6 = _RAND_196[23:0];
  _RAND_197 = {1{`RANDOM}};
  l2_ramDatas_1_entries_ppns_7 = _RAND_197[23:0];
  _RAND_198 = {1{`RANDOM}};
  l2_ramDatas_1_entries_vs_0 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  l2_ramDatas_1_entries_vs_1 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  l2_ramDatas_1_entries_vs_2 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  l2_ramDatas_1_entries_vs_3 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  l2_ramDatas_1_entries_vs_4 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  l2_ramDatas_1_entries_vs_5 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  l2_ramDatas_1_entries_vs_6 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  l2_ramDatas_1_entries_vs_7 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  l2_ramDatas_1_entries_prefetch = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  l2_ramDatas_1_ecc = _RAND_207[30:0];
  _RAND_208 = {1{`RANDOM}};
  l2_ramDatas_2_entries_tag = _RAND_208[12:0];
  _RAND_209 = {1{`RANDOM}};
  l2_ramDatas_2_entries_asid = _RAND_209[15:0];
  _RAND_210 = {1{`RANDOM}};
  l2_ramDatas_2_entries_ppns_0 = _RAND_210[23:0];
  _RAND_211 = {1{`RANDOM}};
  l2_ramDatas_2_entries_ppns_1 = _RAND_211[23:0];
  _RAND_212 = {1{`RANDOM}};
  l2_ramDatas_2_entries_ppns_2 = _RAND_212[23:0];
  _RAND_213 = {1{`RANDOM}};
  l2_ramDatas_2_entries_ppns_3 = _RAND_213[23:0];
  _RAND_214 = {1{`RANDOM}};
  l2_ramDatas_2_entries_ppns_4 = _RAND_214[23:0];
  _RAND_215 = {1{`RANDOM}};
  l2_ramDatas_2_entries_ppns_5 = _RAND_215[23:0];
  _RAND_216 = {1{`RANDOM}};
  l2_ramDatas_2_entries_ppns_6 = _RAND_216[23:0];
  _RAND_217 = {1{`RANDOM}};
  l2_ramDatas_2_entries_ppns_7 = _RAND_217[23:0];
  _RAND_218 = {1{`RANDOM}};
  l2_ramDatas_2_entries_vs_0 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  l2_ramDatas_2_entries_vs_1 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  l2_ramDatas_2_entries_vs_2 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  l2_ramDatas_2_entries_vs_3 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  l2_ramDatas_2_entries_vs_4 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  l2_ramDatas_2_entries_vs_5 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  l2_ramDatas_2_entries_vs_6 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  l2_ramDatas_2_entries_vs_7 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  l2_ramDatas_2_entries_prefetch = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  l2_ramDatas_2_ecc = _RAND_227[30:0];
  _RAND_228 = {1{`RANDOM}};
  l2_ramDatas_3_entries_tag = _RAND_228[12:0];
  _RAND_229 = {1{`RANDOM}};
  l2_ramDatas_3_entries_asid = _RAND_229[15:0];
  _RAND_230 = {1{`RANDOM}};
  l2_ramDatas_3_entries_ppns_0 = _RAND_230[23:0];
  _RAND_231 = {1{`RANDOM}};
  l2_ramDatas_3_entries_ppns_1 = _RAND_231[23:0];
  _RAND_232 = {1{`RANDOM}};
  l2_ramDatas_3_entries_ppns_2 = _RAND_232[23:0];
  _RAND_233 = {1{`RANDOM}};
  l2_ramDatas_3_entries_ppns_3 = _RAND_233[23:0];
  _RAND_234 = {1{`RANDOM}};
  l2_ramDatas_3_entries_ppns_4 = _RAND_234[23:0];
  _RAND_235 = {1{`RANDOM}};
  l2_ramDatas_3_entries_ppns_5 = _RAND_235[23:0];
  _RAND_236 = {1{`RANDOM}};
  l2_ramDatas_3_entries_ppns_6 = _RAND_236[23:0];
  _RAND_237 = {1{`RANDOM}};
  l2_ramDatas_3_entries_ppns_7 = _RAND_237[23:0];
  _RAND_238 = {1{`RANDOM}};
  l2_ramDatas_3_entries_vs_0 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  l2_ramDatas_3_entries_vs_1 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  l2_ramDatas_3_entries_vs_2 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  l2_ramDatas_3_entries_vs_3 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  l2_ramDatas_3_entries_vs_4 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  l2_ramDatas_3_entries_vs_5 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  l2_ramDatas_3_entries_vs_6 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  l2_ramDatas_3_entries_vs_7 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  l2_ramDatas_3_entries_prefetch = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  l2_ramDatas_3_ecc = _RAND_247[30:0];
  _RAND_248 = {1{`RANDOM}};
  l2_hitVec_0 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  l2_hitVec_1 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  l2_hitVec_2 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  l2_hitVec_3 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  state_vec_1_0 = _RAND_252[6:0];
  _RAND_253 = {1{`RANDOM}};
  state_vec_1_1 = _RAND_253[6:0];
  _RAND_254 = {1{`RANDOM}};
  state_vec_1_2 = _RAND_254[6:0];
  _RAND_255 = {1{`RANDOM}};
  state_vec_1_3 = _RAND_255[6:0];
  _RAND_256 = {1{`RANDOM}};
  r_10_0_entries_tag = _RAND_256[21:0];
  _RAND_257 = {1{`RANDOM}};
  r_10_0_entries_asid = _RAND_257[15:0];
  _RAND_258 = {1{`RANDOM}};
  r_10_0_entries_ppns_0 = _RAND_258[23:0];
  _RAND_259 = {1{`RANDOM}};
  r_10_0_entries_ppns_1 = _RAND_259[23:0];
  _RAND_260 = {1{`RANDOM}};
  r_10_0_entries_ppns_2 = _RAND_260[23:0];
  _RAND_261 = {1{`RANDOM}};
  r_10_0_entries_ppns_3 = _RAND_261[23:0];
  _RAND_262 = {1{`RANDOM}};
  r_10_0_entries_ppns_4 = _RAND_262[23:0];
  _RAND_263 = {1{`RANDOM}};
  r_10_0_entries_ppns_5 = _RAND_263[23:0];
  _RAND_264 = {1{`RANDOM}};
  r_10_0_entries_ppns_6 = _RAND_264[23:0];
  _RAND_265 = {1{`RANDOM}};
  r_10_0_entries_ppns_7 = _RAND_265[23:0];
  _RAND_266 = {1{`RANDOM}};
  r_10_0_entries_vs_0 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  r_10_0_entries_vs_1 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  r_10_0_entries_vs_2 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  r_10_0_entries_vs_3 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  r_10_0_entries_vs_4 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  r_10_0_entries_vs_5 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  r_10_0_entries_vs_6 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  r_10_0_entries_vs_7 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  r_10_0_entries_perms_0_d = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  r_10_0_entries_perms_0_a = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  r_10_0_entries_perms_0_g = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  r_10_0_entries_perms_0_u = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  r_10_0_entries_perms_0_x = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  r_10_0_entries_perms_0_w = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  r_10_0_entries_perms_0_r = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  r_10_0_entries_perms_1_d = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  r_10_0_entries_perms_1_a = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  r_10_0_entries_perms_1_g = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  r_10_0_entries_perms_1_u = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  r_10_0_entries_perms_1_x = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  r_10_0_entries_perms_1_w = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  r_10_0_entries_perms_1_r = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  r_10_0_entries_perms_2_d = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  r_10_0_entries_perms_2_a = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  r_10_0_entries_perms_2_g = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  r_10_0_entries_perms_2_u = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  r_10_0_entries_perms_2_x = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  r_10_0_entries_perms_2_w = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  r_10_0_entries_perms_2_r = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  r_10_0_entries_perms_3_d = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  r_10_0_entries_perms_3_a = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  r_10_0_entries_perms_3_g = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  r_10_0_entries_perms_3_u = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  r_10_0_entries_perms_3_x = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  r_10_0_entries_perms_3_w = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  r_10_0_entries_perms_3_r = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  r_10_0_entries_perms_4_d = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  r_10_0_entries_perms_4_a = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  r_10_0_entries_perms_4_g = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  r_10_0_entries_perms_4_u = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  r_10_0_entries_perms_4_x = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  r_10_0_entries_perms_4_w = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  r_10_0_entries_perms_4_r = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  r_10_0_entries_perms_5_d = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  r_10_0_entries_perms_5_a = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  r_10_0_entries_perms_5_g = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  r_10_0_entries_perms_5_u = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  r_10_0_entries_perms_5_x = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  r_10_0_entries_perms_5_w = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  r_10_0_entries_perms_5_r = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  r_10_0_entries_perms_6_d = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  r_10_0_entries_perms_6_a = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  r_10_0_entries_perms_6_g = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  r_10_0_entries_perms_6_u = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  r_10_0_entries_perms_6_x = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  r_10_0_entries_perms_6_w = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  r_10_0_entries_perms_6_r = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  r_10_0_entries_perms_7_d = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  r_10_0_entries_perms_7_a = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  r_10_0_entries_perms_7_g = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  r_10_0_entries_perms_7_u = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  r_10_0_entries_perms_7_x = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  r_10_0_entries_perms_7_w = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  r_10_0_entries_perms_7_r = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  r_10_0_entries_prefetch = _RAND_330[0:0];
  _RAND_331 = {2{`RANDOM}};
  r_10_0_ecc = _RAND_331[38:0];
  _RAND_332 = {1{`RANDOM}};
  r_10_1_entries_tag = _RAND_332[21:0];
  _RAND_333 = {1{`RANDOM}};
  r_10_1_entries_asid = _RAND_333[15:0];
  _RAND_334 = {1{`RANDOM}};
  r_10_1_entries_ppns_0 = _RAND_334[23:0];
  _RAND_335 = {1{`RANDOM}};
  r_10_1_entries_ppns_1 = _RAND_335[23:0];
  _RAND_336 = {1{`RANDOM}};
  r_10_1_entries_ppns_2 = _RAND_336[23:0];
  _RAND_337 = {1{`RANDOM}};
  r_10_1_entries_ppns_3 = _RAND_337[23:0];
  _RAND_338 = {1{`RANDOM}};
  r_10_1_entries_ppns_4 = _RAND_338[23:0];
  _RAND_339 = {1{`RANDOM}};
  r_10_1_entries_ppns_5 = _RAND_339[23:0];
  _RAND_340 = {1{`RANDOM}};
  r_10_1_entries_ppns_6 = _RAND_340[23:0];
  _RAND_341 = {1{`RANDOM}};
  r_10_1_entries_ppns_7 = _RAND_341[23:0];
  _RAND_342 = {1{`RANDOM}};
  r_10_1_entries_vs_0 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  r_10_1_entries_vs_1 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  r_10_1_entries_vs_2 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  r_10_1_entries_vs_3 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  r_10_1_entries_vs_4 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  r_10_1_entries_vs_5 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  r_10_1_entries_vs_6 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  r_10_1_entries_vs_7 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  r_10_1_entries_perms_0_d = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  r_10_1_entries_perms_0_a = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  r_10_1_entries_perms_0_g = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  r_10_1_entries_perms_0_u = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  r_10_1_entries_perms_0_x = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  r_10_1_entries_perms_0_w = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  r_10_1_entries_perms_0_r = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  r_10_1_entries_perms_1_d = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  r_10_1_entries_perms_1_a = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  r_10_1_entries_perms_1_g = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  r_10_1_entries_perms_1_u = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  r_10_1_entries_perms_1_x = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  r_10_1_entries_perms_1_w = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  r_10_1_entries_perms_1_r = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  r_10_1_entries_perms_2_d = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  r_10_1_entries_perms_2_a = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  r_10_1_entries_perms_2_g = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  r_10_1_entries_perms_2_u = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  r_10_1_entries_perms_2_x = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  r_10_1_entries_perms_2_w = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  r_10_1_entries_perms_2_r = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  r_10_1_entries_perms_3_d = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  r_10_1_entries_perms_3_a = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  r_10_1_entries_perms_3_g = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  r_10_1_entries_perms_3_u = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  r_10_1_entries_perms_3_x = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  r_10_1_entries_perms_3_w = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  r_10_1_entries_perms_3_r = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  r_10_1_entries_perms_4_d = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  r_10_1_entries_perms_4_a = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  r_10_1_entries_perms_4_g = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  r_10_1_entries_perms_4_u = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  r_10_1_entries_perms_4_x = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  r_10_1_entries_perms_4_w = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  r_10_1_entries_perms_4_r = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  r_10_1_entries_perms_5_d = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  r_10_1_entries_perms_5_a = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  r_10_1_entries_perms_5_g = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  r_10_1_entries_perms_5_u = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  r_10_1_entries_perms_5_x = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  r_10_1_entries_perms_5_w = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  r_10_1_entries_perms_5_r = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  r_10_1_entries_perms_6_d = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  r_10_1_entries_perms_6_a = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  r_10_1_entries_perms_6_g = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  r_10_1_entries_perms_6_u = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  r_10_1_entries_perms_6_x = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  r_10_1_entries_perms_6_w = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  r_10_1_entries_perms_6_r = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  r_10_1_entries_perms_7_d = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  r_10_1_entries_perms_7_a = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  r_10_1_entries_perms_7_g = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  r_10_1_entries_perms_7_u = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  r_10_1_entries_perms_7_x = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  r_10_1_entries_perms_7_w = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  r_10_1_entries_perms_7_r = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  r_10_1_entries_prefetch = _RAND_406[0:0];
  _RAND_407 = {2{`RANDOM}};
  r_10_1_ecc = _RAND_407[38:0];
  _RAND_408 = {1{`RANDOM}};
  r_10_2_entries_tag = _RAND_408[21:0];
  _RAND_409 = {1{`RANDOM}};
  r_10_2_entries_asid = _RAND_409[15:0];
  _RAND_410 = {1{`RANDOM}};
  r_10_2_entries_ppns_0 = _RAND_410[23:0];
  _RAND_411 = {1{`RANDOM}};
  r_10_2_entries_ppns_1 = _RAND_411[23:0];
  _RAND_412 = {1{`RANDOM}};
  r_10_2_entries_ppns_2 = _RAND_412[23:0];
  _RAND_413 = {1{`RANDOM}};
  r_10_2_entries_ppns_3 = _RAND_413[23:0];
  _RAND_414 = {1{`RANDOM}};
  r_10_2_entries_ppns_4 = _RAND_414[23:0];
  _RAND_415 = {1{`RANDOM}};
  r_10_2_entries_ppns_5 = _RAND_415[23:0];
  _RAND_416 = {1{`RANDOM}};
  r_10_2_entries_ppns_6 = _RAND_416[23:0];
  _RAND_417 = {1{`RANDOM}};
  r_10_2_entries_ppns_7 = _RAND_417[23:0];
  _RAND_418 = {1{`RANDOM}};
  r_10_2_entries_vs_0 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  r_10_2_entries_vs_1 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  r_10_2_entries_vs_2 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  r_10_2_entries_vs_3 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  r_10_2_entries_vs_4 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  r_10_2_entries_vs_5 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  r_10_2_entries_vs_6 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  r_10_2_entries_vs_7 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  r_10_2_entries_perms_0_d = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  r_10_2_entries_perms_0_a = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  r_10_2_entries_perms_0_g = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  r_10_2_entries_perms_0_u = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  r_10_2_entries_perms_0_x = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  r_10_2_entries_perms_0_w = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  r_10_2_entries_perms_0_r = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  r_10_2_entries_perms_1_d = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  r_10_2_entries_perms_1_a = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  r_10_2_entries_perms_1_g = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  r_10_2_entries_perms_1_u = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  r_10_2_entries_perms_1_x = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  r_10_2_entries_perms_1_w = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  r_10_2_entries_perms_1_r = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  r_10_2_entries_perms_2_d = _RAND_440[0:0];
  _RAND_441 = {1{`RANDOM}};
  r_10_2_entries_perms_2_a = _RAND_441[0:0];
  _RAND_442 = {1{`RANDOM}};
  r_10_2_entries_perms_2_g = _RAND_442[0:0];
  _RAND_443 = {1{`RANDOM}};
  r_10_2_entries_perms_2_u = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  r_10_2_entries_perms_2_x = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  r_10_2_entries_perms_2_w = _RAND_445[0:0];
  _RAND_446 = {1{`RANDOM}};
  r_10_2_entries_perms_2_r = _RAND_446[0:0];
  _RAND_447 = {1{`RANDOM}};
  r_10_2_entries_perms_3_d = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  r_10_2_entries_perms_3_a = _RAND_448[0:0];
  _RAND_449 = {1{`RANDOM}};
  r_10_2_entries_perms_3_g = _RAND_449[0:0];
  _RAND_450 = {1{`RANDOM}};
  r_10_2_entries_perms_3_u = _RAND_450[0:0];
  _RAND_451 = {1{`RANDOM}};
  r_10_2_entries_perms_3_x = _RAND_451[0:0];
  _RAND_452 = {1{`RANDOM}};
  r_10_2_entries_perms_3_w = _RAND_452[0:0];
  _RAND_453 = {1{`RANDOM}};
  r_10_2_entries_perms_3_r = _RAND_453[0:0];
  _RAND_454 = {1{`RANDOM}};
  r_10_2_entries_perms_4_d = _RAND_454[0:0];
  _RAND_455 = {1{`RANDOM}};
  r_10_2_entries_perms_4_a = _RAND_455[0:0];
  _RAND_456 = {1{`RANDOM}};
  r_10_2_entries_perms_4_g = _RAND_456[0:0];
  _RAND_457 = {1{`RANDOM}};
  r_10_2_entries_perms_4_u = _RAND_457[0:0];
  _RAND_458 = {1{`RANDOM}};
  r_10_2_entries_perms_4_x = _RAND_458[0:0];
  _RAND_459 = {1{`RANDOM}};
  r_10_2_entries_perms_4_w = _RAND_459[0:0];
  _RAND_460 = {1{`RANDOM}};
  r_10_2_entries_perms_4_r = _RAND_460[0:0];
  _RAND_461 = {1{`RANDOM}};
  r_10_2_entries_perms_5_d = _RAND_461[0:0];
  _RAND_462 = {1{`RANDOM}};
  r_10_2_entries_perms_5_a = _RAND_462[0:0];
  _RAND_463 = {1{`RANDOM}};
  r_10_2_entries_perms_5_g = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  r_10_2_entries_perms_5_u = _RAND_464[0:0];
  _RAND_465 = {1{`RANDOM}};
  r_10_2_entries_perms_5_x = _RAND_465[0:0];
  _RAND_466 = {1{`RANDOM}};
  r_10_2_entries_perms_5_w = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  r_10_2_entries_perms_5_r = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  r_10_2_entries_perms_6_d = _RAND_468[0:0];
  _RAND_469 = {1{`RANDOM}};
  r_10_2_entries_perms_6_a = _RAND_469[0:0];
  _RAND_470 = {1{`RANDOM}};
  r_10_2_entries_perms_6_g = _RAND_470[0:0];
  _RAND_471 = {1{`RANDOM}};
  r_10_2_entries_perms_6_u = _RAND_471[0:0];
  _RAND_472 = {1{`RANDOM}};
  r_10_2_entries_perms_6_x = _RAND_472[0:0];
  _RAND_473 = {1{`RANDOM}};
  r_10_2_entries_perms_6_w = _RAND_473[0:0];
  _RAND_474 = {1{`RANDOM}};
  r_10_2_entries_perms_6_r = _RAND_474[0:0];
  _RAND_475 = {1{`RANDOM}};
  r_10_2_entries_perms_7_d = _RAND_475[0:0];
  _RAND_476 = {1{`RANDOM}};
  r_10_2_entries_perms_7_a = _RAND_476[0:0];
  _RAND_477 = {1{`RANDOM}};
  r_10_2_entries_perms_7_g = _RAND_477[0:0];
  _RAND_478 = {1{`RANDOM}};
  r_10_2_entries_perms_7_u = _RAND_478[0:0];
  _RAND_479 = {1{`RANDOM}};
  r_10_2_entries_perms_7_x = _RAND_479[0:0];
  _RAND_480 = {1{`RANDOM}};
  r_10_2_entries_perms_7_w = _RAND_480[0:0];
  _RAND_481 = {1{`RANDOM}};
  r_10_2_entries_perms_7_r = _RAND_481[0:0];
  _RAND_482 = {1{`RANDOM}};
  r_10_2_entries_prefetch = _RAND_482[0:0];
  _RAND_483 = {2{`RANDOM}};
  r_10_2_ecc = _RAND_483[38:0];
  _RAND_484 = {1{`RANDOM}};
  r_10_3_entries_tag = _RAND_484[21:0];
  _RAND_485 = {1{`RANDOM}};
  r_10_3_entries_asid = _RAND_485[15:0];
  _RAND_486 = {1{`RANDOM}};
  r_10_3_entries_ppns_0 = _RAND_486[23:0];
  _RAND_487 = {1{`RANDOM}};
  r_10_3_entries_ppns_1 = _RAND_487[23:0];
  _RAND_488 = {1{`RANDOM}};
  r_10_3_entries_ppns_2 = _RAND_488[23:0];
  _RAND_489 = {1{`RANDOM}};
  r_10_3_entries_ppns_3 = _RAND_489[23:0];
  _RAND_490 = {1{`RANDOM}};
  r_10_3_entries_ppns_4 = _RAND_490[23:0];
  _RAND_491 = {1{`RANDOM}};
  r_10_3_entries_ppns_5 = _RAND_491[23:0];
  _RAND_492 = {1{`RANDOM}};
  r_10_3_entries_ppns_6 = _RAND_492[23:0];
  _RAND_493 = {1{`RANDOM}};
  r_10_3_entries_ppns_7 = _RAND_493[23:0];
  _RAND_494 = {1{`RANDOM}};
  r_10_3_entries_vs_0 = _RAND_494[0:0];
  _RAND_495 = {1{`RANDOM}};
  r_10_3_entries_vs_1 = _RAND_495[0:0];
  _RAND_496 = {1{`RANDOM}};
  r_10_3_entries_vs_2 = _RAND_496[0:0];
  _RAND_497 = {1{`RANDOM}};
  r_10_3_entries_vs_3 = _RAND_497[0:0];
  _RAND_498 = {1{`RANDOM}};
  r_10_3_entries_vs_4 = _RAND_498[0:0];
  _RAND_499 = {1{`RANDOM}};
  r_10_3_entries_vs_5 = _RAND_499[0:0];
  _RAND_500 = {1{`RANDOM}};
  r_10_3_entries_vs_6 = _RAND_500[0:0];
  _RAND_501 = {1{`RANDOM}};
  r_10_3_entries_vs_7 = _RAND_501[0:0];
  _RAND_502 = {1{`RANDOM}};
  r_10_3_entries_perms_0_d = _RAND_502[0:0];
  _RAND_503 = {1{`RANDOM}};
  r_10_3_entries_perms_0_a = _RAND_503[0:0];
  _RAND_504 = {1{`RANDOM}};
  r_10_3_entries_perms_0_g = _RAND_504[0:0];
  _RAND_505 = {1{`RANDOM}};
  r_10_3_entries_perms_0_u = _RAND_505[0:0];
  _RAND_506 = {1{`RANDOM}};
  r_10_3_entries_perms_0_x = _RAND_506[0:0];
  _RAND_507 = {1{`RANDOM}};
  r_10_3_entries_perms_0_w = _RAND_507[0:0];
  _RAND_508 = {1{`RANDOM}};
  r_10_3_entries_perms_0_r = _RAND_508[0:0];
  _RAND_509 = {1{`RANDOM}};
  r_10_3_entries_perms_1_d = _RAND_509[0:0];
  _RAND_510 = {1{`RANDOM}};
  r_10_3_entries_perms_1_a = _RAND_510[0:0];
  _RAND_511 = {1{`RANDOM}};
  r_10_3_entries_perms_1_g = _RAND_511[0:0];
  _RAND_512 = {1{`RANDOM}};
  r_10_3_entries_perms_1_u = _RAND_512[0:0];
  _RAND_513 = {1{`RANDOM}};
  r_10_3_entries_perms_1_x = _RAND_513[0:0];
  _RAND_514 = {1{`RANDOM}};
  r_10_3_entries_perms_1_w = _RAND_514[0:0];
  _RAND_515 = {1{`RANDOM}};
  r_10_3_entries_perms_1_r = _RAND_515[0:0];
  _RAND_516 = {1{`RANDOM}};
  r_10_3_entries_perms_2_d = _RAND_516[0:0];
  _RAND_517 = {1{`RANDOM}};
  r_10_3_entries_perms_2_a = _RAND_517[0:0];
  _RAND_518 = {1{`RANDOM}};
  r_10_3_entries_perms_2_g = _RAND_518[0:0];
  _RAND_519 = {1{`RANDOM}};
  r_10_3_entries_perms_2_u = _RAND_519[0:0];
  _RAND_520 = {1{`RANDOM}};
  r_10_3_entries_perms_2_x = _RAND_520[0:0];
  _RAND_521 = {1{`RANDOM}};
  r_10_3_entries_perms_2_w = _RAND_521[0:0];
  _RAND_522 = {1{`RANDOM}};
  r_10_3_entries_perms_2_r = _RAND_522[0:0];
  _RAND_523 = {1{`RANDOM}};
  r_10_3_entries_perms_3_d = _RAND_523[0:0];
  _RAND_524 = {1{`RANDOM}};
  r_10_3_entries_perms_3_a = _RAND_524[0:0];
  _RAND_525 = {1{`RANDOM}};
  r_10_3_entries_perms_3_g = _RAND_525[0:0];
  _RAND_526 = {1{`RANDOM}};
  r_10_3_entries_perms_3_u = _RAND_526[0:0];
  _RAND_527 = {1{`RANDOM}};
  r_10_3_entries_perms_3_x = _RAND_527[0:0];
  _RAND_528 = {1{`RANDOM}};
  r_10_3_entries_perms_3_w = _RAND_528[0:0];
  _RAND_529 = {1{`RANDOM}};
  r_10_3_entries_perms_3_r = _RAND_529[0:0];
  _RAND_530 = {1{`RANDOM}};
  r_10_3_entries_perms_4_d = _RAND_530[0:0];
  _RAND_531 = {1{`RANDOM}};
  r_10_3_entries_perms_4_a = _RAND_531[0:0];
  _RAND_532 = {1{`RANDOM}};
  r_10_3_entries_perms_4_g = _RAND_532[0:0];
  _RAND_533 = {1{`RANDOM}};
  r_10_3_entries_perms_4_u = _RAND_533[0:0];
  _RAND_534 = {1{`RANDOM}};
  r_10_3_entries_perms_4_x = _RAND_534[0:0];
  _RAND_535 = {1{`RANDOM}};
  r_10_3_entries_perms_4_w = _RAND_535[0:0];
  _RAND_536 = {1{`RANDOM}};
  r_10_3_entries_perms_4_r = _RAND_536[0:0];
  _RAND_537 = {1{`RANDOM}};
  r_10_3_entries_perms_5_d = _RAND_537[0:0];
  _RAND_538 = {1{`RANDOM}};
  r_10_3_entries_perms_5_a = _RAND_538[0:0];
  _RAND_539 = {1{`RANDOM}};
  r_10_3_entries_perms_5_g = _RAND_539[0:0];
  _RAND_540 = {1{`RANDOM}};
  r_10_3_entries_perms_5_u = _RAND_540[0:0];
  _RAND_541 = {1{`RANDOM}};
  r_10_3_entries_perms_5_x = _RAND_541[0:0];
  _RAND_542 = {1{`RANDOM}};
  r_10_3_entries_perms_5_w = _RAND_542[0:0];
  _RAND_543 = {1{`RANDOM}};
  r_10_3_entries_perms_5_r = _RAND_543[0:0];
  _RAND_544 = {1{`RANDOM}};
  r_10_3_entries_perms_6_d = _RAND_544[0:0];
  _RAND_545 = {1{`RANDOM}};
  r_10_3_entries_perms_6_a = _RAND_545[0:0];
  _RAND_546 = {1{`RANDOM}};
  r_10_3_entries_perms_6_g = _RAND_546[0:0];
  _RAND_547 = {1{`RANDOM}};
  r_10_3_entries_perms_6_u = _RAND_547[0:0];
  _RAND_548 = {1{`RANDOM}};
  r_10_3_entries_perms_6_x = _RAND_548[0:0];
  _RAND_549 = {1{`RANDOM}};
  r_10_3_entries_perms_6_w = _RAND_549[0:0];
  _RAND_550 = {1{`RANDOM}};
  r_10_3_entries_perms_6_r = _RAND_550[0:0];
  _RAND_551 = {1{`RANDOM}};
  r_10_3_entries_perms_7_d = _RAND_551[0:0];
  _RAND_552 = {1{`RANDOM}};
  r_10_3_entries_perms_7_a = _RAND_552[0:0];
  _RAND_553 = {1{`RANDOM}};
  r_10_3_entries_perms_7_g = _RAND_553[0:0];
  _RAND_554 = {1{`RANDOM}};
  r_10_3_entries_perms_7_u = _RAND_554[0:0];
  _RAND_555 = {1{`RANDOM}};
  r_10_3_entries_perms_7_x = _RAND_555[0:0];
  _RAND_556 = {1{`RANDOM}};
  r_10_3_entries_perms_7_w = _RAND_556[0:0];
  _RAND_557 = {1{`RANDOM}};
  r_10_3_entries_perms_7_r = _RAND_557[0:0];
  _RAND_558 = {1{`RANDOM}};
  r_10_3_entries_prefetch = _RAND_558[0:0];
  _RAND_559 = {2{`RANDOM}};
  r_10_3_ecc = _RAND_559[38:0];
  _RAND_560 = {1{`RANDOM}};
  r_10_4_entries_tag = _RAND_560[21:0];
  _RAND_561 = {1{`RANDOM}};
  r_10_4_entries_asid = _RAND_561[15:0];
  _RAND_562 = {1{`RANDOM}};
  r_10_4_entries_ppns_0 = _RAND_562[23:0];
  _RAND_563 = {1{`RANDOM}};
  r_10_4_entries_ppns_1 = _RAND_563[23:0];
  _RAND_564 = {1{`RANDOM}};
  r_10_4_entries_ppns_2 = _RAND_564[23:0];
  _RAND_565 = {1{`RANDOM}};
  r_10_4_entries_ppns_3 = _RAND_565[23:0];
  _RAND_566 = {1{`RANDOM}};
  r_10_4_entries_ppns_4 = _RAND_566[23:0];
  _RAND_567 = {1{`RANDOM}};
  r_10_4_entries_ppns_5 = _RAND_567[23:0];
  _RAND_568 = {1{`RANDOM}};
  r_10_4_entries_ppns_6 = _RAND_568[23:0];
  _RAND_569 = {1{`RANDOM}};
  r_10_4_entries_ppns_7 = _RAND_569[23:0];
  _RAND_570 = {1{`RANDOM}};
  r_10_4_entries_vs_0 = _RAND_570[0:0];
  _RAND_571 = {1{`RANDOM}};
  r_10_4_entries_vs_1 = _RAND_571[0:0];
  _RAND_572 = {1{`RANDOM}};
  r_10_4_entries_vs_2 = _RAND_572[0:0];
  _RAND_573 = {1{`RANDOM}};
  r_10_4_entries_vs_3 = _RAND_573[0:0];
  _RAND_574 = {1{`RANDOM}};
  r_10_4_entries_vs_4 = _RAND_574[0:0];
  _RAND_575 = {1{`RANDOM}};
  r_10_4_entries_vs_5 = _RAND_575[0:0];
  _RAND_576 = {1{`RANDOM}};
  r_10_4_entries_vs_6 = _RAND_576[0:0];
  _RAND_577 = {1{`RANDOM}};
  r_10_4_entries_vs_7 = _RAND_577[0:0];
  _RAND_578 = {1{`RANDOM}};
  r_10_4_entries_perms_0_d = _RAND_578[0:0];
  _RAND_579 = {1{`RANDOM}};
  r_10_4_entries_perms_0_a = _RAND_579[0:0];
  _RAND_580 = {1{`RANDOM}};
  r_10_4_entries_perms_0_g = _RAND_580[0:0];
  _RAND_581 = {1{`RANDOM}};
  r_10_4_entries_perms_0_u = _RAND_581[0:0];
  _RAND_582 = {1{`RANDOM}};
  r_10_4_entries_perms_0_x = _RAND_582[0:0];
  _RAND_583 = {1{`RANDOM}};
  r_10_4_entries_perms_0_w = _RAND_583[0:0];
  _RAND_584 = {1{`RANDOM}};
  r_10_4_entries_perms_0_r = _RAND_584[0:0];
  _RAND_585 = {1{`RANDOM}};
  r_10_4_entries_perms_1_d = _RAND_585[0:0];
  _RAND_586 = {1{`RANDOM}};
  r_10_4_entries_perms_1_a = _RAND_586[0:0];
  _RAND_587 = {1{`RANDOM}};
  r_10_4_entries_perms_1_g = _RAND_587[0:0];
  _RAND_588 = {1{`RANDOM}};
  r_10_4_entries_perms_1_u = _RAND_588[0:0];
  _RAND_589 = {1{`RANDOM}};
  r_10_4_entries_perms_1_x = _RAND_589[0:0];
  _RAND_590 = {1{`RANDOM}};
  r_10_4_entries_perms_1_w = _RAND_590[0:0];
  _RAND_591 = {1{`RANDOM}};
  r_10_4_entries_perms_1_r = _RAND_591[0:0];
  _RAND_592 = {1{`RANDOM}};
  r_10_4_entries_perms_2_d = _RAND_592[0:0];
  _RAND_593 = {1{`RANDOM}};
  r_10_4_entries_perms_2_a = _RAND_593[0:0];
  _RAND_594 = {1{`RANDOM}};
  r_10_4_entries_perms_2_g = _RAND_594[0:0];
  _RAND_595 = {1{`RANDOM}};
  r_10_4_entries_perms_2_u = _RAND_595[0:0];
  _RAND_596 = {1{`RANDOM}};
  r_10_4_entries_perms_2_x = _RAND_596[0:0];
  _RAND_597 = {1{`RANDOM}};
  r_10_4_entries_perms_2_w = _RAND_597[0:0];
  _RAND_598 = {1{`RANDOM}};
  r_10_4_entries_perms_2_r = _RAND_598[0:0];
  _RAND_599 = {1{`RANDOM}};
  r_10_4_entries_perms_3_d = _RAND_599[0:0];
  _RAND_600 = {1{`RANDOM}};
  r_10_4_entries_perms_3_a = _RAND_600[0:0];
  _RAND_601 = {1{`RANDOM}};
  r_10_4_entries_perms_3_g = _RAND_601[0:0];
  _RAND_602 = {1{`RANDOM}};
  r_10_4_entries_perms_3_u = _RAND_602[0:0];
  _RAND_603 = {1{`RANDOM}};
  r_10_4_entries_perms_3_x = _RAND_603[0:0];
  _RAND_604 = {1{`RANDOM}};
  r_10_4_entries_perms_3_w = _RAND_604[0:0];
  _RAND_605 = {1{`RANDOM}};
  r_10_4_entries_perms_3_r = _RAND_605[0:0];
  _RAND_606 = {1{`RANDOM}};
  r_10_4_entries_perms_4_d = _RAND_606[0:0];
  _RAND_607 = {1{`RANDOM}};
  r_10_4_entries_perms_4_a = _RAND_607[0:0];
  _RAND_608 = {1{`RANDOM}};
  r_10_4_entries_perms_4_g = _RAND_608[0:0];
  _RAND_609 = {1{`RANDOM}};
  r_10_4_entries_perms_4_u = _RAND_609[0:0];
  _RAND_610 = {1{`RANDOM}};
  r_10_4_entries_perms_4_x = _RAND_610[0:0];
  _RAND_611 = {1{`RANDOM}};
  r_10_4_entries_perms_4_w = _RAND_611[0:0];
  _RAND_612 = {1{`RANDOM}};
  r_10_4_entries_perms_4_r = _RAND_612[0:0];
  _RAND_613 = {1{`RANDOM}};
  r_10_4_entries_perms_5_d = _RAND_613[0:0];
  _RAND_614 = {1{`RANDOM}};
  r_10_4_entries_perms_5_a = _RAND_614[0:0];
  _RAND_615 = {1{`RANDOM}};
  r_10_4_entries_perms_5_g = _RAND_615[0:0];
  _RAND_616 = {1{`RANDOM}};
  r_10_4_entries_perms_5_u = _RAND_616[0:0];
  _RAND_617 = {1{`RANDOM}};
  r_10_4_entries_perms_5_x = _RAND_617[0:0];
  _RAND_618 = {1{`RANDOM}};
  r_10_4_entries_perms_5_w = _RAND_618[0:0];
  _RAND_619 = {1{`RANDOM}};
  r_10_4_entries_perms_5_r = _RAND_619[0:0];
  _RAND_620 = {1{`RANDOM}};
  r_10_4_entries_perms_6_d = _RAND_620[0:0];
  _RAND_621 = {1{`RANDOM}};
  r_10_4_entries_perms_6_a = _RAND_621[0:0];
  _RAND_622 = {1{`RANDOM}};
  r_10_4_entries_perms_6_g = _RAND_622[0:0];
  _RAND_623 = {1{`RANDOM}};
  r_10_4_entries_perms_6_u = _RAND_623[0:0];
  _RAND_624 = {1{`RANDOM}};
  r_10_4_entries_perms_6_x = _RAND_624[0:0];
  _RAND_625 = {1{`RANDOM}};
  r_10_4_entries_perms_6_w = _RAND_625[0:0];
  _RAND_626 = {1{`RANDOM}};
  r_10_4_entries_perms_6_r = _RAND_626[0:0];
  _RAND_627 = {1{`RANDOM}};
  r_10_4_entries_perms_7_d = _RAND_627[0:0];
  _RAND_628 = {1{`RANDOM}};
  r_10_4_entries_perms_7_a = _RAND_628[0:0];
  _RAND_629 = {1{`RANDOM}};
  r_10_4_entries_perms_7_g = _RAND_629[0:0];
  _RAND_630 = {1{`RANDOM}};
  r_10_4_entries_perms_7_u = _RAND_630[0:0];
  _RAND_631 = {1{`RANDOM}};
  r_10_4_entries_perms_7_x = _RAND_631[0:0];
  _RAND_632 = {1{`RANDOM}};
  r_10_4_entries_perms_7_w = _RAND_632[0:0];
  _RAND_633 = {1{`RANDOM}};
  r_10_4_entries_perms_7_r = _RAND_633[0:0];
  _RAND_634 = {1{`RANDOM}};
  r_10_4_entries_prefetch = _RAND_634[0:0];
  _RAND_635 = {2{`RANDOM}};
  r_10_4_ecc = _RAND_635[38:0];
  _RAND_636 = {1{`RANDOM}};
  r_10_5_entries_tag = _RAND_636[21:0];
  _RAND_637 = {1{`RANDOM}};
  r_10_5_entries_asid = _RAND_637[15:0];
  _RAND_638 = {1{`RANDOM}};
  r_10_5_entries_ppns_0 = _RAND_638[23:0];
  _RAND_639 = {1{`RANDOM}};
  r_10_5_entries_ppns_1 = _RAND_639[23:0];
  _RAND_640 = {1{`RANDOM}};
  r_10_5_entries_ppns_2 = _RAND_640[23:0];
  _RAND_641 = {1{`RANDOM}};
  r_10_5_entries_ppns_3 = _RAND_641[23:0];
  _RAND_642 = {1{`RANDOM}};
  r_10_5_entries_ppns_4 = _RAND_642[23:0];
  _RAND_643 = {1{`RANDOM}};
  r_10_5_entries_ppns_5 = _RAND_643[23:0];
  _RAND_644 = {1{`RANDOM}};
  r_10_5_entries_ppns_6 = _RAND_644[23:0];
  _RAND_645 = {1{`RANDOM}};
  r_10_5_entries_ppns_7 = _RAND_645[23:0];
  _RAND_646 = {1{`RANDOM}};
  r_10_5_entries_vs_0 = _RAND_646[0:0];
  _RAND_647 = {1{`RANDOM}};
  r_10_5_entries_vs_1 = _RAND_647[0:0];
  _RAND_648 = {1{`RANDOM}};
  r_10_5_entries_vs_2 = _RAND_648[0:0];
  _RAND_649 = {1{`RANDOM}};
  r_10_5_entries_vs_3 = _RAND_649[0:0];
  _RAND_650 = {1{`RANDOM}};
  r_10_5_entries_vs_4 = _RAND_650[0:0];
  _RAND_651 = {1{`RANDOM}};
  r_10_5_entries_vs_5 = _RAND_651[0:0];
  _RAND_652 = {1{`RANDOM}};
  r_10_5_entries_vs_6 = _RAND_652[0:0];
  _RAND_653 = {1{`RANDOM}};
  r_10_5_entries_vs_7 = _RAND_653[0:0];
  _RAND_654 = {1{`RANDOM}};
  r_10_5_entries_perms_0_d = _RAND_654[0:0];
  _RAND_655 = {1{`RANDOM}};
  r_10_5_entries_perms_0_a = _RAND_655[0:0];
  _RAND_656 = {1{`RANDOM}};
  r_10_5_entries_perms_0_g = _RAND_656[0:0];
  _RAND_657 = {1{`RANDOM}};
  r_10_5_entries_perms_0_u = _RAND_657[0:0];
  _RAND_658 = {1{`RANDOM}};
  r_10_5_entries_perms_0_x = _RAND_658[0:0];
  _RAND_659 = {1{`RANDOM}};
  r_10_5_entries_perms_0_w = _RAND_659[0:0];
  _RAND_660 = {1{`RANDOM}};
  r_10_5_entries_perms_0_r = _RAND_660[0:0];
  _RAND_661 = {1{`RANDOM}};
  r_10_5_entries_perms_1_d = _RAND_661[0:0];
  _RAND_662 = {1{`RANDOM}};
  r_10_5_entries_perms_1_a = _RAND_662[0:0];
  _RAND_663 = {1{`RANDOM}};
  r_10_5_entries_perms_1_g = _RAND_663[0:0];
  _RAND_664 = {1{`RANDOM}};
  r_10_5_entries_perms_1_u = _RAND_664[0:0];
  _RAND_665 = {1{`RANDOM}};
  r_10_5_entries_perms_1_x = _RAND_665[0:0];
  _RAND_666 = {1{`RANDOM}};
  r_10_5_entries_perms_1_w = _RAND_666[0:0];
  _RAND_667 = {1{`RANDOM}};
  r_10_5_entries_perms_1_r = _RAND_667[0:0];
  _RAND_668 = {1{`RANDOM}};
  r_10_5_entries_perms_2_d = _RAND_668[0:0];
  _RAND_669 = {1{`RANDOM}};
  r_10_5_entries_perms_2_a = _RAND_669[0:0];
  _RAND_670 = {1{`RANDOM}};
  r_10_5_entries_perms_2_g = _RAND_670[0:0];
  _RAND_671 = {1{`RANDOM}};
  r_10_5_entries_perms_2_u = _RAND_671[0:0];
  _RAND_672 = {1{`RANDOM}};
  r_10_5_entries_perms_2_x = _RAND_672[0:0];
  _RAND_673 = {1{`RANDOM}};
  r_10_5_entries_perms_2_w = _RAND_673[0:0];
  _RAND_674 = {1{`RANDOM}};
  r_10_5_entries_perms_2_r = _RAND_674[0:0];
  _RAND_675 = {1{`RANDOM}};
  r_10_5_entries_perms_3_d = _RAND_675[0:0];
  _RAND_676 = {1{`RANDOM}};
  r_10_5_entries_perms_3_a = _RAND_676[0:0];
  _RAND_677 = {1{`RANDOM}};
  r_10_5_entries_perms_3_g = _RAND_677[0:0];
  _RAND_678 = {1{`RANDOM}};
  r_10_5_entries_perms_3_u = _RAND_678[0:0];
  _RAND_679 = {1{`RANDOM}};
  r_10_5_entries_perms_3_x = _RAND_679[0:0];
  _RAND_680 = {1{`RANDOM}};
  r_10_5_entries_perms_3_w = _RAND_680[0:0];
  _RAND_681 = {1{`RANDOM}};
  r_10_5_entries_perms_3_r = _RAND_681[0:0];
  _RAND_682 = {1{`RANDOM}};
  r_10_5_entries_perms_4_d = _RAND_682[0:0];
  _RAND_683 = {1{`RANDOM}};
  r_10_5_entries_perms_4_a = _RAND_683[0:0];
  _RAND_684 = {1{`RANDOM}};
  r_10_5_entries_perms_4_g = _RAND_684[0:0];
  _RAND_685 = {1{`RANDOM}};
  r_10_5_entries_perms_4_u = _RAND_685[0:0];
  _RAND_686 = {1{`RANDOM}};
  r_10_5_entries_perms_4_x = _RAND_686[0:0];
  _RAND_687 = {1{`RANDOM}};
  r_10_5_entries_perms_4_w = _RAND_687[0:0];
  _RAND_688 = {1{`RANDOM}};
  r_10_5_entries_perms_4_r = _RAND_688[0:0];
  _RAND_689 = {1{`RANDOM}};
  r_10_5_entries_perms_5_d = _RAND_689[0:0];
  _RAND_690 = {1{`RANDOM}};
  r_10_5_entries_perms_5_a = _RAND_690[0:0];
  _RAND_691 = {1{`RANDOM}};
  r_10_5_entries_perms_5_g = _RAND_691[0:0];
  _RAND_692 = {1{`RANDOM}};
  r_10_5_entries_perms_5_u = _RAND_692[0:0];
  _RAND_693 = {1{`RANDOM}};
  r_10_5_entries_perms_5_x = _RAND_693[0:0];
  _RAND_694 = {1{`RANDOM}};
  r_10_5_entries_perms_5_w = _RAND_694[0:0];
  _RAND_695 = {1{`RANDOM}};
  r_10_5_entries_perms_5_r = _RAND_695[0:0];
  _RAND_696 = {1{`RANDOM}};
  r_10_5_entries_perms_6_d = _RAND_696[0:0];
  _RAND_697 = {1{`RANDOM}};
  r_10_5_entries_perms_6_a = _RAND_697[0:0];
  _RAND_698 = {1{`RANDOM}};
  r_10_5_entries_perms_6_g = _RAND_698[0:0];
  _RAND_699 = {1{`RANDOM}};
  r_10_5_entries_perms_6_u = _RAND_699[0:0];
  _RAND_700 = {1{`RANDOM}};
  r_10_5_entries_perms_6_x = _RAND_700[0:0];
  _RAND_701 = {1{`RANDOM}};
  r_10_5_entries_perms_6_w = _RAND_701[0:0];
  _RAND_702 = {1{`RANDOM}};
  r_10_5_entries_perms_6_r = _RAND_702[0:0];
  _RAND_703 = {1{`RANDOM}};
  r_10_5_entries_perms_7_d = _RAND_703[0:0];
  _RAND_704 = {1{`RANDOM}};
  r_10_5_entries_perms_7_a = _RAND_704[0:0];
  _RAND_705 = {1{`RANDOM}};
  r_10_5_entries_perms_7_g = _RAND_705[0:0];
  _RAND_706 = {1{`RANDOM}};
  r_10_5_entries_perms_7_u = _RAND_706[0:0];
  _RAND_707 = {1{`RANDOM}};
  r_10_5_entries_perms_7_x = _RAND_707[0:0];
  _RAND_708 = {1{`RANDOM}};
  r_10_5_entries_perms_7_w = _RAND_708[0:0];
  _RAND_709 = {1{`RANDOM}};
  r_10_5_entries_perms_7_r = _RAND_709[0:0];
  _RAND_710 = {1{`RANDOM}};
  r_10_5_entries_prefetch = _RAND_710[0:0];
  _RAND_711 = {2{`RANDOM}};
  r_10_5_ecc = _RAND_711[38:0];
  _RAND_712 = {1{`RANDOM}};
  r_10_6_entries_tag = _RAND_712[21:0];
  _RAND_713 = {1{`RANDOM}};
  r_10_6_entries_asid = _RAND_713[15:0];
  _RAND_714 = {1{`RANDOM}};
  r_10_6_entries_ppns_0 = _RAND_714[23:0];
  _RAND_715 = {1{`RANDOM}};
  r_10_6_entries_ppns_1 = _RAND_715[23:0];
  _RAND_716 = {1{`RANDOM}};
  r_10_6_entries_ppns_2 = _RAND_716[23:0];
  _RAND_717 = {1{`RANDOM}};
  r_10_6_entries_ppns_3 = _RAND_717[23:0];
  _RAND_718 = {1{`RANDOM}};
  r_10_6_entries_ppns_4 = _RAND_718[23:0];
  _RAND_719 = {1{`RANDOM}};
  r_10_6_entries_ppns_5 = _RAND_719[23:0];
  _RAND_720 = {1{`RANDOM}};
  r_10_6_entries_ppns_6 = _RAND_720[23:0];
  _RAND_721 = {1{`RANDOM}};
  r_10_6_entries_ppns_7 = _RAND_721[23:0];
  _RAND_722 = {1{`RANDOM}};
  r_10_6_entries_vs_0 = _RAND_722[0:0];
  _RAND_723 = {1{`RANDOM}};
  r_10_6_entries_vs_1 = _RAND_723[0:0];
  _RAND_724 = {1{`RANDOM}};
  r_10_6_entries_vs_2 = _RAND_724[0:0];
  _RAND_725 = {1{`RANDOM}};
  r_10_6_entries_vs_3 = _RAND_725[0:0];
  _RAND_726 = {1{`RANDOM}};
  r_10_6_entries_vs_4 = _RAND_726[0:0];
  _RAND_727 = {1{`RANDOM}};
  r_10_6_entries_vs_5 = _RAND_727[0:0];
  _RAND_728 = {1{`RANDOM}};
  r_10_6_entries_vs_6 = _RAND_728[0:0];
  _RAND_729 = {1{`RANDOM}};
  r_10_6_entries_vs_7 = _RAND_729[0:0];
  _RAND_730 = {1{`RANDOM}};
  r_10_6_entries_perms_0_d = _RAND_730[0:0];
  _RAND_731 = {1{`RANDOM}};
  r_10_6_entries_perms_0_a = _RAND_731[0:0];
  _RAND_732 = {1{`RANDOM}};
  r_10_6_entries_perms_0_g = _RAND_732[0:0];
  _RAND_733 = {1{`RANDOM}};
  r_10_6_entries_perms_0_u = _RAND_733[0:0];
  _RAND_734 = {1{`RANDOM}};
  r_10_6_entries_perms_0_x = _RAND_734[0:0];
  _RAND_735 = {1{`RANDOM}};
  r_10_6_entries_perms_0_w = _RAND_735[0:0];
  _RAND_736 = {1{`RANDOM}};
  r_10_6_entries_perms_0_r = _RAND_736[0:0];
  _RAND_737 = {1{`RANDOM}};
  r_10_6_entries_perms_1_d = _RAND_737[0:0];
  _RAND_738 = {1{`RANDOM}};
  r_10_6_entries_perms_1_a = _RAND_738[0:0];
  _RAND_739 = {1{`RANDOM}};
  r_10_6_entries_perms_1_g = _RAND_739[0:0];
  _RAND_740 = {1{`RANDOM}};
  r_10_6_entries_perms_1_u = _RAND_740[0:0];
  _RAND_741 = {1{`RANDOM}};
  r_10_6_entries_perms_1_x = _RAND_741[0:0];
  _RAND_742 = {1{`RANDOM}};
  r_10_6_entries_perms_1_w = _RAND_742[0:0];
  _RAND_743 = {1{`RANDOM}};
  r_10_6_entries_perms_1_r = _RAND_743[0:0];
  _RAND_744 = {1{`RANDOM}};
  r_10_6_entries_perms_2_d = _RAND_744[0:0];
  _RAND_745 = {1{`RANDOM}};
  r_10_6_entries_perms_2_a = _RAND_745[0:0];
  _RAND_746 = {1{`RANDOM}};
  r_10_6_entries_perms_2_g = _RAND_746[0:0];
  _RAND_747 = {1{`RANDOM}};
  r_10_6_entries_perms_2_u = _RAND_747[0:0];
  _RAND_748 = {1{`RANDOM}};
  r_10_6_entries_perms_2_x = _RAND_748[0:0];
  _RAND_749 = {1{`RANDOM}};
  r_10_6_entries_perms_2_w = _RAND_749[0:0];
  _RAND_750 = {1{`RANDOM}};
  r_10_6_entries_perms_2_r = _RAND_750[0:0];
  _RAND_751 = {1{`RANDOM}};
  r_10_6_entries_perms_3_d = _RAND_751[0:0];
  _RAND_752 = {1{`RANDOM}};
  r_10_6_entries_perms_3_a = _RAND_752[0:0];
  _RAND_753 = {1{`RANDOM}};
  r_10_6_entries_perms_3_g = _RAND_753[0:0];
  _RAND_754 = {1{`RANDOM}};
  r_10_6_entries_perms_3_u = _RAND_754[0:0];
  _RAND_755 = {1{`RANDOM}};
  r_10_6_entries_perms_3_x = _RAND_755[0:0];
  _RAND_756 = {1{`RANDOM}};
  r_10_6_entries_perms_3_w = _RAND_756[0:0];
  _RAND_757 = {1{`RANDOM}};
  r_10_6_entries_perms_3_r = _RAND_757[0:0];
  _RAND_758 = {1{`RANDOM}};
  r_10_6_entries_perms_4_d = _RAND_758[0:0];
  _RAND_759 = {1{`RANDOM}};
  r_10_6_entries_perms_4_a = _RAND_759[0:0];
  _RAND_760 = {1{`RANDOM}};
  r_10_6_entries_perms_4_g = _RAND_760[0:0];
  _RAND_761 = {1{`RANDOM}};
  r_10_6_entries_perms_4_u = _RAND_761[0:0];
  _RAND_762 = {1{`RANDOM}};
  r_10_6_entries_perms_4_x = _RAND_762[0:0];
  _RAND_763 = {1{`RANDOM}};
  r_10_6_entries_perms_4_w = _RAND_763[0:0];
  _RAND_764 = {1{`RANDOM}};
  r_10_6_entries_perms_4_r = _RAND_764[0:0];
  _RAND_765 = {1{`RANDOM}};
  r_10_6_entries_perms_5_d = _RAND_765[0:0];
  _RAND_766 = {1{`RANDOM}};
  r_10_6_entries_perms_5_a = _RAND_766[0:0];
  _RAND_767 = {1{`RANDOM}};
  r_10_6_entries_perms_5_g = _RAND_767[0:0];
  _RAND_768 = {1{`RANDOM}};
  r_10_6_entries_perms_5_u = _RAND_768[0:0];
  _RAND_769 = {1{`RANDOM}};
  r_10_6_entries_perms_5_x = _RAND_769[0:0];
  _RAND_770 = {1{`RANDOM}};
  r_10_6_entries_perms_5_w = _RAND_770[0:0];
  _RAND_771 = {1{`RANDOM}};
  r_10_6_entries_perms_5_r = _RAND_771[0:0];
  _RAND_772 = {1{`RANDOM}};
  r_10_6_entries_perms_6_d = _RAND_772[0:0];
  _RAND_773 = {1{`RANDOM}};
  r_10_6_entries_perms_6_a = _RAND_773[0:0];
  _RAND_774 = {1{`RANDOM}};
  r_10_6_entries_perms_6_g = _RAND_774[0:0];
  _RAND_775 = {1{`RANDOM}};
  r_10_6_entries_perms_6_u = _RAND_775[0:0];
  _RAND_776 = {1{`RANDOM}};
  r_10_6_entries_perms_6_x = _RAND_776[0:0];
  _RAND_777 = {1{`RANDOM}};
  r_10_6_entries_perms_6_w = _RAND_777[0:0];
  _RAND_778 = {1{`RANDOM}};
  r_10_6_entries_perms_6_r = _RAND_778[0:0];
  _RAND_779 = {1{`RANDOM}};
  r_10_6_entries_perms_7_d = _RAND_779[0:0];
  _RAND_780 = {1{`RANDOM}};
  r_10_6_entries_perms_7_a = _RAND_780[0:0];
  _RAND_781 = {1{`RANDOM}};
  r_10_6_entries_perms_7_g = _RAND_781[0:0];
  _RAND_782 = {1{`RANDOM}};
  r_10_6_entries_perms_7_u = _RAND_782[0:0];
  _RAND_783 = {1{`RANDOM}};
  r_10_6_entries_perms_7_x = _RAND_783[0:0];
  _RAND_784 = {1{`RANDOM}};
  r_10_6_entries_perms_7_w = _RAND_784[0:0];
  _RAND_785 = {1{`RANDOM}};
  r_10_6_entries_perms_7_r = _RAND_785[0:0];
  _RAND_786 = {1{`RANDOM}};
  r_10_6_entries_prefetch = _RAND_786[0:0];
  _RAND_787 = {2{`RANDOM}};
  r_10_6_ecc = _RAND_787[38:0];
  _RAND_788 = {1{`RANDOM}};
  r_10_7_entries_tag = _RAND_788[21:0];
  _RAND_789 = {1{`RANDOM}};
  r_10_7_entries_asid = _RAND_789[15:0];
  _RAND_790 = {1{`RANDOM}};
  r_10_7_entries_ppns_0 = _RAND_790[23:0];
  _RAND_791 = {1{`RANDOM}};
  r_10_7_entries_ppns_1 = _RAND_791[23:0];
  _RAND_792 = {1{`RANDOM}};
  r_10_7_entries_ppns_2 = _RAND_792[23:0];
  _RAND_793 = {1{`RANDOM}};
  r_10_7_entries_ppns_3 = _RAND_793[23:0];
  _RAND_794 = {1{`RANDOM}};
  r_10_7_entries_ppns_4 = _RAND_794[23:0];
  _RAND_795 = {1{`RANDOM}};
  r_10_7_entries_ppns_5 = _RAND_795[23:0];
  _RAND_796 = {1{`RANDOM}};
  r_10_7_entries_ppns_6 = _RAND_796[23:0];
  _RAND_797 = {1{`RANDOM}};
  r_10_7_entries_ppns_7 = _RAND_797[23:0];
  _RAND_798 = {1{`RANDOM}};
  r_10_7_entries_vs_0 = _RAND_798[0:0];
  _RAND_799 = {1{`RANDOM}};
  r_10_7_entries_vs_1 = _RAND_799[0:0];
  _RAND_800 = {1{`RANDOM}};
  r_10_7_entries_vs_2 = _RAND_800[0:0];
  _RAND_801 = {1{`RANDOM}};
  r_10_7_entries_vs_3 = _RAND_801[0:0];
  _RAND_802 = {1{`RANDOM}};
  r_10_7_entries_vs_4 = _RAND_802[0:0];
  _RAND_803 = {1{`RANDOM}};
  r_10_7_entries_vs_5 = _RAND_803[0:0];
  _RAND_804 = {1{`RANDOM}};
  r_10_7_entries_vs_6 = _RAND_804[0:0];
  _RAND_805 = {1{`RANDOM}};
  r_10_7_entries_vs_7 = _RAND_805[0:0];
  _RAND_806 = {1{`RANDOM}};
  r_10_7_entries_perms_0_d = _RAND_806[0:0];
  _RAND_807 = {1{`RANDOM}};
  r_10_7_entries_perms_0_a = _RAND_807[0:0];
  _RAND_808 = {1{`RANDOM}};
  r_10_7_entries_perms_0_g = _RAND_808[0:0];
  _RAND_809 = {1{`RANDOM}};
  r_10_7_entries_perms_0_u = _RAND_809[0:0];
  _RAND_810 = {1{`RANDOM}};
  r_10_7_entries_perms_0_x = _RAND_810[0:0];
  _RAND_811 = {1{`RANDOM}};
  r_10_7_entries_perms_0_w = _RAND_811[0:0];
  _RAND_812 = {1{`RANDOM}};
  r_10_7_entries_perms_0_r = _RAND_812[0:0];
  _RAND_813 = {1{`RANDOM}};
  r_10_7_entries_perms_1_d = _RAND_813[0:0];
  _RAND_814 = {1{`RANDOM}};
  r_10_7_entries_perms_1_a = _RAND_814[0:0];
  _RAND_815 = {1{`RANDOM}};
  r_10_7_entries_perms_1_g = _RAND_815[0:0];
  _RAND_816 = {1{`RANDOM}};
  r_10_7_entries_perms_1_u = _RAND_816[0:0];
  _RAND_817 = {1{`RANDOM}};
  r_10_7_entries_perms_1_x = _RAND_817[0:0];
  _RAND_818 = {1{`RANDOM}};
  r_10_7_entries_perms_1_w = _RAND_818[0:0];
  _RAND_819 = {1{`RANDOM}};
  r_10_7_entries_perms_1_r = _RAND_819[0:0];
  _RAND_820 = {1{`RANDOM}};
  r_10_7_entries_perms_2_d = _RAND_820[0:0];
  _RAND_821 = {1{`RANDOM}};
  r_10_7_entries_perms_2_a = _RAND_821[0:0];
  _RAND_822 = {1{`RANDOM}};
  r_10_7_entries_perms_2_g = _RAND_822[0:0];
  _RAND_823 = {1{`RANDOM}};
  r_10_7_entries_perms_2_u = _RAND_823[0:0];
  _RAND_824 = {1{`RANDOM}};
  r_10_7_entries_perms_2_x = _RAND_824[0:0];
  _RAND_825 = {1{`RANDOM}};
  r_10_7_entries_perms_2_w = _RAND_825[0:0];
  _RAND_826 = {1{`RANDOM}};
  r_10_7_entries_perms_2_r = _RAND_826[0:0];
  _RAND_827 = {1{`RANDOM}};
  r_10_7_entries_perms_3_d = _RAND_827[0:0];
  _RAND_828 = {1{`RANDOM}};
  r_10_7_entries_perms_3_a = _RAND_828[0:0];
  _RAND_829 = {1{`RANDOM}};
  r_10_7_entries_perms_3_g = _RAND_829[0:0];
  _RAND_830 = {1{`RANDOM}};
  r_10_7_entries_perms_3_u = _RAND_830[0:0];
  _RAND_831 = {1{`RANDOM}};
  r_10_7_entries_perms_3_x = _RAND_831[0:0];
  _RAND_832 = {1{`RANDOM}};
  r_10_7_entries_perms_3_w = _RAND_832[0:0];
  _RAND_833 = {1{`RANDOM}};
  r_10_7_entries_perms_3_r = _RAND_833[0:0];
  _RAND_834 = {1{`RANDOM}};
  r_10_7_entries_perms_4_d = _RAND_834[0:0];
  _RAND_835 = {1{`RANDOM}};
  r_10_7_entries_perms_4_a = _RAND_835[0:0];
  _RAND_836 = {1{`RANDOM}};
  r_10_7_entries_perms_4_g = _RAND_836[0:0];
  _RAND_837 = {1{`RANDOM}};
  r_10_7_entries_perms_4_u = _RAND_837[0:0];
  _RAND_838 = {1{`RANDOM}};
  r_10_7_entries_perms_4_x = _RAND_838[0:0];
  _RAND_839 = {1{`RANDOM}};
  r_10_7_entries_perms_4_w = _RAND_839[0:0];
  _RAND_840 = {1{`RANDOM}};
  r_10_7_entries_perms_4_r = _RAND_840[0:0];
  _RAND_841 = {1{`RANDOM}};
  r_10_7_entries_perms_5_d = _RAND_841[0:0];
  _RAND_842 = {1{`RANDOM}};
  r_10_7_entries_perms_5_a = _RAND_842[0:0];
  _RAND_843 = {1{`RANDOM}};
  r_10_7_entries_perms_5_g = _RAND_843[0:0];
  _RAND_844 = {1{`RANDOM}};
  r_10_7_entries_perms_5_u = _RAND_844[0:0];
  _RAND_845 = {1{`RANDOM}};
  r_10_7_entries_perms_5_x = _RAND_845[0:0];
  _RAND_846 = {1{`RANDOM}};
  r_10_7_entries_perms_5_w = _RAND_846[0:0];
  _RAND_847 = {1{`RANDOM}};
  r_10_7_entries_perms_5_r = _RAND_847[0:0];
  _RAND_848 = {1{`RANDOM}};
  r_10_7_entries_perms_6_d = _RAND_848[0:0];
  _RAND_849 = {1{`RANDOM}};
  r_10_7_entries_perms_6_a = _RAND_849[0:0];
  _RAND_850 = {1{`RANDOM}};
  r_10_7_entries_perms_6_g = _RAND_850[0:0];
  _RAND_851 = {1{`RANDOM}};
  r_10_7_entries_perms_6_u = _RAND_851[0:0];
  _RAND_852 = {1{`RANDOM}};
  r_10_7_entries_perms_6_x = _RAND_852[0:0];
  _RAND_853 = {1{`RANDOM}};
  r_10_7_entries_perms_6_w = _RAND_853[0:0];
  _RAND_854 = {1{`RANDOM}};
  r_10_7_entries_perms_6_r = _RAND_854[0:0];
  _RAND_855 = {1{`RANDOM}};
  r_10_7_entries_perms_7_d = _RAND_855[0:0];
  _RAND_856 = {1{`RANDOM}};
  r_10_7_entries_perms_7_a = _RAND_856[0:0];
  _RAND_857 = {1{`RANDOM}};
  r_10_7_entries_perms_7_g = _RAND_857[0:0];
  _RAND_858 = {1{`RANDOM}};
  r_10_7_entries_perms_7_u = _RAND_858[0:0];
  _RAND_859 = {1{`RANDOM}};
  r_10_7_entries_perms_7_x = _RAND_859[0:0];
  _RAND_860 = {1{`RANDOM}};
  r_10_7_entries_perms_7_w = _RAND_860[0:0];
  _RAND_861 = {1{`RANDOM}};
  r_10_7_entries_perms_7_r = _RAND_861[0:0];
  _RAND_862 = {1{`RANDOM}};
  r_10_7_entries_prefetch = _RAND_862[0:0];
  _RAND_863 = {2{`RANDOM}};
  r_10_7_ecc = _RAND_863[38:0];
  _RAND_864 = {1{`RANDOM}};
  r_11 = _RAND_864[7:0];
  _RAND_865 = {1{`RANDOM}};
  l3_ramDatas_0_entries_tag = _RAND_865[21:0];
  _RAND_866 = {1{`RANDOM}};
  l3_ramDatas_0_entries_asid = _RAND_866[15:0];
  _RAND_867 = {1{`RANDOM}};
  l3_ramDatas_0_entries_ppns_0 = _RAND_867[23:0];
  _RAND_868 = {1{`RANDOM}};
  l3_ramDatas_0_entries_ppns_1 = _RAND_868[23:0];
  _RAND_869 = {1{`RANDOM}};
  l3_ramDatas_0_entries_ppns_2 = _RAND_869[23:0];
  _RAND_870 = {1{`RANDOM}};
  l3_ramDatas_0_entries_ppns_3 = _RAND_870[23:0];
  _RAND_871 = {1{`RANDOM}};
  l3_ramDatas_0_entries_ppns_4 = _RAND_871[23:0];
  _RAND_872 = {1{`RANDOM}};
  l3_ramDatas_0_entries_ppns_5 = _RAND_872[23:0];
  _RAND_873 = {1{`RANDOM}};
  l3_ramDatas_0_entries_ppns_6 = _RAND_873[23:0];
  _RAND_874 = {1{`RANDOM}};
  l3_ramDatas_0_entries_ppns_7 = _RAND_874[23:0];
  _RAND_875 = {1{`RANDOM}};
  l3_ramDatas_0_entries_vs_0 = _RAND_875[0:0];
  _RAND_876 = {1{`RANDOM}};
  l3_ramDatas_0_entries_vs_1 = _RAND_876[0:0];
  _RAND_877 = {1{`RANDOM}};
  l3_ramDatas_0_entries_vs_2 = _RAND_877[0:0];
  _RAND_878 = {1{`RANDOM}};
  l3_ramDatas_0_entries_vs_3 = _RAND_878[0:0];
  _RAND_879 = {1{`RANDOM}};
  l3_ramDatas_0_entries_vs_4 = _RAND_879[0:0];
  _RAND_880 = {1{`RANDOM}};
  l3_ramDatas_0_entries_vs_5 = _RAND_880[0:0];
  _RAND_881 = {1{`RANDOM}};
  l3_ramDatas_0_entries_vs_6 = _RAND_881[0:0];
  _RAND_882 = {1{`RANDOM}};
  l3_ramDatas_0_entries_vs_7 = _RAND_882[0:0];
  _RAND_883 = {1{`RANDOM}};
  l3_ramDatas_0_entries_perms_0_d = _RAND_883[0:0];
  _RAND_884 = {1{`RANDOM}};
  l3_ramDatas_0_entries_perms_0_a = _RAND_884[0:0];
  _RAND_885 = {1{`RANDOM}};
  l3_ramDatas_0_entries_perms_0_g = _RAND_885[0:0];
  _RAND_886 = {1{`RANDOM}};
  l3_ramDatas_0_entries_perms_0_u = _RAND_886[0:0];
  _RAND_887 = {1{`RANDOM}};
  l3_ramDatas_0_entries_perms_0_x = _RAND_887[0:0];
  _RAND_888 = {1{`RANDOM}};
  l3_ramDatas_0_entries_perms_0_w = _RAND_888[0:0];
  _RAND_889 = {1{`RANDOM}};
  l3_ramDatas_0_entries_perms_0_r = _RAND_889[0:0];
  _RAND_890 = {1{`RANDOM}};
  l3_ramDatas_0_entries_perms_1_d = _RAND_890[0:0];
  _RAND_891 = {1{`RANDOM}};
  l3_ramDatas_0_entries_perms_1_a = _RAND_891[0:0];
  _RAND_892 = {1{`RANDOM}};
  l3_ramDatas_0_entries_perms_1_g = _RAND_892[0:0];
  _RAND_893 = {1{`RANDOM}};
  l3_ramDatas_0_entries_perms_1_u = _RAND_893[0:0];
  _RAND_894 = {1{`RANDOM}};
  l3_ramDatas_0_entries_perms_1_x = _RAND_894[0:0];
  _RAND_895 = {1{`RANDOM}};
  l3_ramDatas_0_entries_perms_1_w = _RAND_895[0:0];
  _RAND_896 = {1{`RANDOM}};
  l3_ramDatas_0_entries_perms_1_r = _RAND_896[0:0];
  _RAND_897 = {1{`RANDOM}};
  l3_ramDatas_0_entries_perms_2_d = _RAND_897[0:0];
  _RAND_898 = {1{`RANDOM}};
  l3_ramDatas_0_entries_perms_2_a = _RAND_898[0:0];
  _RAND_899 = {1{`RANDOM}};
  l3_ramDatas_0_entries_perms_2_g = _RAND_899[0:0];
  _RAND_900 = {1{`RANDOM}};
  l3_ramDatas_0_entries_perms_2_u = _RAND_900[0:0];
  _RAND_901 = {1{`RANDOM}};
  l3_ramDatas_0_entries_perms_2_x = _RAND_901[0:0];
  _RAND_902 = {1{`RANDOM}};
  l3_ramDatas_0_entries_perms_2_w = _RAND_902[0:0];
  _RAND_903 = {1{`RANDOM}};
  l3_ramDatas_0_entries_perms_2_r = _RAND_903[0:0];
  _RAND_904 = {1{`RANDOM}};
  l3_ramDatas_0_entries_perms_3_d = _RAND_904[0:0];
  _RAND_905 = {1{`RANDOM}};
  l3_ramDatas_0_entries_perms_3_a = _RAND_905[0:0];
  _RAND_906 = {1{`RANDOM}};
  l3_ramDatas_0_entries_perms_3_g = _RAND_906[0:0];
  _RAND_907 = {1{`RANDOM}};
  l3_ramDatas_0_entries_perms_3_u = _RAND_907[0:0];
  _RAND_908 = {1{`RANDOM}};
  l3_ramDatas_0_entries_perms_3_x = _RAND_908[0:0];
  _RAND_909 = {1{`RANDOM}};
  l3_ramDatas_0_entries_perms_3_w = _RAND_909[0:0];
  _RAND_910 = {1{`RANDOM}};
  l3_ramDatas_0_entries_perms_3_r = _RAND_910[0:0];
  _RAND_911 = {1{`RANDOM}};
  l3_ramDatas_0_entries_perms_4_d = _RAND_911[0:0];
  _RAND_912 = {1{`RANDOM}};
  l3_ramDatas_0_entries_perms_4_a = _RAND_912[0:0];
  _RAND_913 = {1{`RANDOM}};
  l3_ramDatas_0_entries_perms_4_g = _RAND_913[0:0];
  _RAND_914 = {1{`RANDOM}};
  l3_ramDatas_0_entries_perms_4_u = _RAND_914[0:0];
  _RAND_915 = {1{`RANDOM}};
  l3_ramDatas_0_entries_perms_4_x = _RAND_915[0:0];
  _RAND_916 = {1{`RANDOM}};
  l3_ramDatas_0_entries_perms_4_w = _RAND_916[0:0];
  _RAND_917 = {1{`RANDOM}};
  l3_ramDatas_0_entries_perms_4_r = _RAND_917[0:0];
  _RAND_918 = {1{`RANDOM}};
  l3_ramDatas_0_entries_perms_5_d = _RAND_918[0:0];
  _RAND_919 = {1{`RANDOM}};
  l3_ramDatas_0_entries_perms_5_a = _RAND_919[0:0];
  _RAND_920 = {1{`RANDOM}};
  l3_ramDatas_0_entries_perms_5_g = _RAND_920[0:0];
  _RAND_921 = {1{`RANDOM}};
  l3_ramDatas_0_entries_perms_5_u = _RAND_921[0:0];
  _RAND_922 = {1{`RANDOM}};
  l3_ramDatas_0_entries_perms_5_x = _RAND_922[0:0];
  _RAND_923 = {1{`RANDOM}};
  l3_ramDatas_0_entries_perms_5_w = _RAND_923[0:0];
  _RAND_924 = {1{`RANDOM}};
  l3_ramDatas_0_entries_perms_5_r = _RAND_924[0:0];
  _RAND_925 = {1{`RANDOM}};
  l3_ramDatas_0_entries_perms_6_d = _RAND_925[0:0];
  _RAND_926 = {1{`RANDOM}};
  l3_ramDatas_0_entries_perms_6_a = _RAND_926[0:0];
  _RAND_927 = {1{`RANDOM}};
  l3_ramDatas_0_entries_perms_6_g = _RAND_927[0:0];
  _RAND_928 = {1{`RANDOM}};
  l3_ramDatas_0_entries_perms_6_u = _RAND_928[0:0];
  _RAND_929 = {1{`RANDOM}};
  l3_ramDatas_0_entries_perms_6_x = _RAND_929[0:0];
  _RAND_930 = {1{`RANDOM}};
  l3_ramDatas_0_entries_perms_6_w = _RAND_930[0:0];
  _RAND_931 = {1{`RANDOM}};
  l3_ramDatas_0_entries_perms_6_r = _RAND_931[0:0];
  _RAND_932 = {1{`RANDOM}};
  l3_ramDatas_0_entries_perms_7_d = _RAND_932[0:0];
  _RAND_933 = {1{`RANDOM}};
  l3_ramDatas_0_entries_perms_7_a = _RAND_933[0:0];
  _RAND_934 = {1{`RANDOM}};
  l3_ramDatas_0_entries_perms_7_g = _RAND_934[0:0];
  _RAND_935 = {1{`RANDOM}};
  l3_ramDatas_0_entries_perms_7_u = _RAND_935[0:0];
  _RAND_936 = {1{`RANDOM}};
  l3_ramDatas_0_entries_perms_7_x = _RAND_936[0:0];
  _RAND_937 = {1{`RANDOM}};
  l3_ramDatas_0_entries_perms_7_w = _RAND_937[0:0];
  _RAND_938 = {1{`RANDOM}};
  l3_ramDatas_0_entries_perms_7_r = _RAND_938[0:0];
  _RAND_939 = {1{`RANDOM}};
  l3_ramDatas_0_entries_prefetch = _RAND_939[0:0];
  _RAND_940 = {2{`RANDOM}};
  l3_ramDatas_0_ecc = _RAND_940[38:0];
  _RAND_941 = {1{`RANDOM}};
  l3_ramDatas_1_entries_tag = _RAND_941[21:0];
  _RAND_942 = {1{`RANDOM}};
  l3_ramDatas_1_entries_asid = _RAND_942[15:0];
  _RAND_943 = {1{`RANDOM}};
  l3_ramDatas_1_entries_ppns_0 = _RAND_943[23:0];
  _RAND_944 = {1{`RANDOM}};
  l3_ramDatas_1_entries_ppns_1 = _RAND_944[23:0];
  _RAND_945 = {1{`RANDOM}};
  l3_ramDatas_1_entries_ppns_2 = _RAND_945[23:0];
  _RAND_946 = {1{`RANDOM}};
  l3_ramDatas_1_entries_ppns_3 = _RAND_946[23:0];
  _RAND_947 = {1{`RANDOM}};
  l3_ramDatas_1_entries_ppns_4 = _RAND_947[23:0];
  _RAND_948 = {1{`RANDOM}};
  l3_ramDatas_1_entries_ppns_5 = _RAND_948[23:0];
  _RAND_949 = {1{`RANDOM}};
  l3_ramDatas_1_entries_ppns_6 = _RAND_949[23:0];
  _RAND_950 = {1{`RANDOM}};
  l3_ramDatas_1_entries_ppns_7 = _RAND_950[23:0];
  _RAND_951 = {1{`RANDOM}};
  l3_ramDatas_1_entries_vs_0 = _RAND_951[0:0];
  _RAND_952 = {1{`RANDOM}};
  l3_ramDatas_1_entries_vs_1 = _RAND_952[0:0];
  _RAND_953 = {1{`RANDOM}};
  l3_ramDatas_1_entries_vs_2 = _RAND_953[0:0];
  _RAND_954 = {1{`RANDOM}};
  l3_ramDatas_1_entries_vs_3 = _RAND_954[0:0];
  _RAND_955 = {1{`RANDOM}};
  l3_ramDatas_1_entries_vs_4 = _RAND_955[0:0];
  _RAND_956 = {1{`RANDOM}};
  l3_ramDatas_1_entries_vs_5 = _RAND_956[0:0];
  _RAND_957 = {1{`RANDOM}};
  l3_ramDatas_1_entries_vs_6 = _RAND_957[0:0];
  _RAND_958 = {1{`RANDOM}};
  l3_ramDatas_1_entries_vs_7 = _RAND_958[0:0];
  _RAND_959 = {1{`RANDOM}};
  l3_ramDatas_1_entries_perms_0_d = _RAND_959[0:0];
  _RAND_960 = {1{`RANDOM}};
  l3_ramDatas_1_entries_perms_0_a = _RAND_960[0:0];
  _RAND_961 = {1{`RANDOM}};
  l3_ramDatas_1_entries_perms_0_g = _RAND_961[0:0];
  _RAND_962 = {1{`RANDOM}};
  l3_ramDatas_1_entries_perms_0_u = _RAND_962[0:0];
  _RAND_963 = {1{`RANDOM}};
  l3_ramDatas_1_entries_perms_0_x = _RAND_963[0:0];
  _RAND_964 = {1{`RANDOM}};
  l3_ramDatas_1_entries_perms_0_w = _RAND_964[0:0];
  _RAND_965 = {1{`RANDOM}};
  l3_ramDatas_1_entries_perms_0_r = _RAND_965[0:0];
  _RAND_966 = {1{`RANDOM}};
  l3_ramDatas_1_entries_perms_1_d = _RAND_966[0:0];
  _RAND_967 = {1{`RANDOM}};
  l3_ramDatas_1_entries_perms_1_a = _RAND_967[0:0];
  _RAND_968 = {1{`RANDOM}};
  l3_ramDatas_1_entries_perms_1_g = _RAND_968[0:0];
  _RAND_969 = {1{`RANDOM}};
  l3_ramDatas_1_entries_perms_1_u = _RAND_969[0:0];
  _RAND_970 = {1{`RANDOM}};
  l3_ramDatas_1_entries_perms_1_x = _RAND_970[0:0];
  _RAND_971 = {1{`RANDOM}};
  l3_ramDatas_1_entries_perms_1_w = _RAND_971[0:0];
  _RAND_972 = {1{`RANDOM}};
  l3_ramDatas_1_entries_perms_1_r = _RAND_972[0:0];
  _RAND_973 = {1{`RANDOM}};
  l3_ramDatas_1_entries_perms_2_d = _RAND_973[0:0];
  _RAND_974 = {1{`RANDOM}};
  l3_ramDatas_1_entries_perms_2_a = _RAND_974[0:0];
  _RAND_975 = {1{`RANDOM}};
  l3_ramDatas_1_entries_perms_2_g = _RAND_975[0:0];
  _RAND_976 = {1{`RANDOM}};
  l3_ramDatas_1_entries_perms_2_u = _RAND_976[0:0];
  _RAND_977 = {1{`RANDOM}};
  l3_ramDatas_1_entries_perms_2_x = _RAND_977[0:0];
  _RAND_978 = {1{`RANDOM}};
  l3_ramDatas_1_entries_perms_2_w = _RAND_978[0:0];
  _RAND_979 = {1{`RANDOM}};
  l3_ramDatas_1_entries_perms_2_r = _RAND_979[0:0];
  _RAND_980 = {1{`RANDOM}};
  l3_ramDatas_1_entries_perms_3_d = _RAND_980[0:0];
  _RAND_981 = {1{`RANDOM}};
  l3_ramDatas_1_entries_perms_3_a = _RAND_981[0:0];
  _RAND_982 = {1{`RANDOM}};
  l3_ramDatas_1_entries_perms_3_g = _RAND_982[0:0];
  _RAND_983 = {1{`RANDOM}};
  l3_ramDatas_1_entries_perms_3_u = _RAND_983[0:0];
  _RAND_984 = {1{`RANDOM}};
  l3_ramDatas_1_entries_perms_3_x = _RAND_984[0:0];
  _RAND_985 = {1{`RANDOM}};
  l3_ramDatas_1_entries_perms_3_w = _RAND_985[0:0];
  _RAND_986 = {1{`RANDOM}};
  l3_ramDatas_1_entries_perms_3_r = _RAND_986[0:0];
  _RAND_987 = {1{`RANDOM}};
  l3_ramDatas_1_entries_perms_4_d = _RAND_987[0:0];
  _RAND_988 = {1{`RANDOM}};
  l3_ramDatas_1_entries_perms_4_a = _RAND_988[0:0];
  _RAND_989 = {1{`RANDOM}};
  l3_ramDatas_1_entries_perms_4_g = _RAND_989[0:0];
  _RAND_990 = {1{`RANDOM}};
  l3_ramDatas_1_entries_perms_4_u = _RAND_990[0:0];
  _RAND_991 = {1{`RANDOM}};
  l3_ramDatas_1_entries_perms_4_x = _RAND_991[0:0];
  _RAND_992 = {1{`RANDOM}};
  l3_ramDatas_1_entries_perms_4_w = _RAND_992[0:0];
  _RAND_993 = {1{`RANDOM}};
  l3_ramDatas_1_entries_perms_4_r = _RAND_993[0:0];
  _RAND_994 = {1{`RANDOM}};
  l3_ramDatas_1_entries_perms_5_d = _RAND_994[0:0];
  _RAND_995 = {1{`RANDOM}};
  l3_ramDatas_1_entries_perms_5_a = _RAND_995[0:0];
  _RAND_996 = {1{`RANDOM}};
  l3_ramDatas_1_entries_perms_5_g = _RAND_996[0:0];
  _RAND_997 = {1{`RANDOM}};
  l3_ramDatas_1_entries_perms_5_u = _RAND_997[0:0];
  _RAND_998 = {1{`RANDOM}};
  l3_ramDatas_1_entries_perms_5_x = _RAND_998[0:0];
  _RAND_999 = {1{`RANDOM}};
  l3_ramDatas_1_entries_perms_5_w = _RAND_999[0:0];
  _RAND_1000 = {1{`RANDOM}};
  l3_ramDatas_1_entries_perms_5_r = _RAND_1000[0:0];
  _RAND_1001 = {1{`RANDOM}};
  l3_ramDatas_1_entries_perms_6_d = _RAND_1001[0:0];
  _RAND_1002 = {1{`RANDOM}};
  l3_ramDatas_1_entries_perms_6_a = _RAND_1002[0:0];
  _RAND_1003 = {1{`RANDOM}};
  l3_ramDatas_1_entries_perms_6_g = _RAND_1003[0:0];
  _RAND_1004 = {1{`RANDOM}};
  l3_ramDatas_1_entries_perms_6_u = _RAND_1004[0:0];
  _RAND_1005 = {1{`RANDOM}};
  l3_ramDatas_1_entries_perms_6_x = _RAND_1005[0:0];
  _RAND_1006 = {1{`RANDOM}};
  l3_ramDatas_1_entries_perms_6_w = _RAND_1006[0:0];
  _RAND_1007 = {1{`RANDOM}};
  l3_ramDatas_1_entries_perms_6_r = _RAND_1007[0:0];
  _RAND_1008 = {1{`RANDOM}};
  l3_ramDatas_1_entries_perms_7_d = _RAND_1008[0:0];
  _RAND_1009 = {1{`RANDOM}};
  l3_ramDatas_1_entries_perms_7_a = _RAND_1009[0:0];
  _RAND_1010 = {1{`RANDOM}};
  l3_ramDatas_1_entries_perms_7_g = _RAND_1010[0:0];
  _RAND_1011 = {1{`RANDOM}};
  l3_ramDatas_1_entries_perms_7_u = _RAND_1011[0:0];
  _RAND_1012 = {1{`RANDOM}};
  l3_ramDatas_1_entries_perms_7_x = _RAND_1012[0:0];
  _RAND_1013 = {1{`RANDOM}};
  l3_ramDatas_1_entries_perms_7_w = _RAND_1013[0:0];
  _RAND_1014 = {1{`RANDOM}};
  l3_ramDatas_1_entries_perms_7_r = _RAND_1014[0:0];
  _RAND_1015 = {1{`RANDOM}};
  l3_ramDatas_1_entries_prefetch = _RAND_1015[0:0];
  _RAND_1016 = {2{`RANDOM}};
  l3_ramDatas_1_ecc = _RAND_1016[38:0];
  _RAND_1017 = {1{`RANDOM}};
  l3_ramDatas_2_entries_tag = _RAND_1017[21:0];
  _RAND_1018 = {1{`RANDOM}};
  l3_ramDatas_2_entries_asid = _RAND_1018[15:0];
  _RAND_1019 = {1{`RANDOM}};
  l3_ramDatas_2_entries_ppns_0 = _RAND_1019[23:0];
  _RAND_1020 = {1{`RANDOM}};
  l3_ramDatas_2_entries_ppns_1 = _RAND_1020[23:0];
  _RAND_1021 = {1{`RANDOM}};
  l3_ramDatas_2_entries_ppns_2 = _RAND_1021[23:0];
  _RAND_1022 = {1{`RANDOM}};
  l3_ramDatas_2_entries_ppns_3 = _RAND_1022[23:0];
  _RAND_1023 = {1{`RANDOM}};
  l3_ramDatas_2_entries_ppns_4 = _RAND_1023[23:0];
  _RAND_1024 = {1{`RANDOM}};
  l3_ramDatas_2_entries_ppns_5 = _RAND_1024[23:0];
  _RAND_1025 = {1{`RANDOM}};
  l3_ramDatas_2_entries_ppns_6 = _RAND_1025[23:0];
  _RAND_1026 = {1{`RANDOM}};
  l3_ramDatas_2_entries_ppns_7 = _RAND_1026[23:0];
  _RAND_1027 = {1{`RANDOM}};
  l3_ramDatas_2_entries_vs_0 = _RAND_1027[0:0];
  _RAND_1028 = {1{`RANDOM}};
  l3_ramDatas_2_entries_vs_1 = _RAND_1028[0:0];
  _RAND_1029 = {1{`RANDOM}};
  l3_ramDatas_2_entries_vs_2 = _RAND_1029[0:0];
  _RAND_1030 = {1{`RANDOM}};
  l3_ramDatas_2_entries_vs_3 = _RAND_1030[0:0];
  _RAND_1031 = {1{`RANDOM}};
  l3_ramDatas_2_entries_vs_4 = _RAND_1031[0:0];
  _RAND_1032 = {1{`RANDOM}};
  l3_ramDatas_2_entries_vs_5 = _RAND_1032[0:0];
  _RAND_1033 = {1{`RANDOM}};
  l3_ramDatas_2_entries_vs_6 = _RAND_1033[0:0];
  _RAND_1034 = {1{`RANDOM}};
  l3_ramDatas_2_entries_vs_7 = _RAND_1034[0:0];
  _RAND_1035 = {1{`RANDOM}};
  l3_ramDatas_2_entries_perms_0_d = _RAND_1035[0:0];
  _RAND_1036 = {1{`RANDOM}};
  l3_ramDatas_2_entries_perms_0_a = _RAND_1036[0:0];
  _RAND_1037 = {1{`RANDOM}};
  l3_ramDatas_2_entries_perms_0_g = _RAND_1037[0:0];
  _RAND_1038 = {1{`RANDOM}};
  l3_ramDatas_2_entries_perms_0_u = _RAND_1038[0:0];
  _RAND_1039 = {1{`RANDOM}};
  l3_ramDatas_2_entries_perms_0_x = _RAND_1039[0:0];
  _RAND_1040 = {1{`RANDOM}};
  l3_ramDatas_2_entries_perms_0_w = _RAND_1040[0:0];
  _RAND_1041 = {1{`RANDOM}};
  l3_ramDatas_2_entries_perms_0_r = _RAND_1041[0:0];
  _RAND_1042 = {1{`RANDOM}};
  l3_ramDatas_2_entries_perms_1_d = _RAND_1042[0:0];
  _RAND_1043 = {1{`RANDOM}};
  l3_ramDatas_2_entries_perms_1_a = _RAND_1043[0:0];
  _RAND_1044 = {1{`RANDOM}};
  l3_ramDatas_2_entries_perms_1_g = _RAND_1044[0:0];
  _RAND_1045 = {1{`RANDOM}};
  l3_ramDatas_2_entries_perms_1_u = _RAND_1045[0:0];
  _RAND_1046 = {1{`RANDOM}};
  l3_ramDatas_2_entries_perms_1_x = _RAND_1046[0:0];
  _RAND_1047 = {1{`RANDOM}};
  l3_ramDatas_2_entries_perms_1_w = _RAND_1047[0:0];
  _RAND_1048 = {1{`RANDOM}};
  l3_ramDatas_2_entries_perms_1_r = _RAND_1048[0:0];
  _RAND_1049 = {1{`RANDOM}};
  l3_ramDatas_2_entries_perms_2_d = _RAND_1049[0:0];
  _RAND_1050 = {1{`RANDOM}};
  l3_ramDatas_2_entries_perms_2_a = _RAND_1050[0:0];
  _RAND_1051 = {1{`RANDOM}};
  l3_ramDatas_2_entries_perms_2_g = _RAND_1051[0:0];
  _RAND_1052 = {1{`RANDOM}};
  l3_ramDatas_2_entries_perms_2_u = _RAND_1052[0:0];
  _RAND_1053 = {1{`RANDOM}};
  l3_ramDatas_2_entries_perms_2_x = _RAND_1053[0:0];
  _RAND_1054 = {1{`RANDOM}};
  l3_ramDatas_2_entries_perms_2_w = _RAND_1054[0:0];
  _RAND_1055 = {1{`RANDOM}};
  l3_ramDatas_2_entries_perms_2_r = _RAND_1055[0:0];
  _RAND_1056 = {1{`RANDOM}};
  l3_ramDatas_2_entries_perms_3_d = _RAND_1056[0:0];
  _RAND_1057 = {1{`RANDOM}};
  l3_ramDatas_2_entries_perms_3_a = _RAND_1057[0:0];
  _RAND_1058 = {1{`RANDOM}};
  l3_ramDatas_2_entries_perms_3_g = _RAND_1058[0:0];
  _RAND_1059 = {1{`RANDOM}};
  l3_ramDatas_2_entries_perms_3_u = _RAND_1059[0:0];
  _RAND_1060 = {1{`RANDOM}};
  l3_ramDatas_2_entries_perms_3_x = _RAND_1060[0:0];
  _RAND_1061 = {1{`RANDOM}};
  l3_ramDatas_2_entries_perms_3_w = _RAND_1061[0:0];
  _RAND_1062 = {1{`RANDOM}};
  l3_ramDatas_2_entries_perms_3_r = _RAND_1062[0:0];
  _RAND_1063 = {1{`RANDOM}};
  l3_ramDatas_2_entries_perms_4_d = _RAND_1063[0:0];
  _RAND_1064 = {1{`RANDOM}};
  l3_ramDatas_2_entries_perms_4_a = _RAND_1064[0:0];
  _RAND_1065 = {1{`RANDOM}};
  l3_ramDatas_2_entries_perms_4_g = _RAND_1065[0:0];
  _RAND_1066 = {1{`RANDOM}};
  l3_ramDatas_2_entries_perms_4_u = _RAND_1066[0:0];
  _RAND_1067 = {1{`RANDOM}};
  l3_ramDatas_2_entries_perms_4_x = _RAND_1067[0:0];
  _RAND_1068 = {1{`RANDOM}};
  l3_ramDatas_2_entries_perms_4_w = _RAND_1068[0:0];
  _RAND_1069 = {1{`RANDOM}};
  l3_ramDatas_2_entries_perms_4_r = _RAND_1069[0:0];
  _RAND_1070 = {1{`RANDOM}};
  l3_ramDatas_2_entries_perms_5_d = _RAND_1070[0:0];
  _RAND_1071 = {1{`RANDOM}};
  l3_ramDatas_2_entries_perms_5_a = _RAND_1071[0:0];
  _RAND_1072 = {1{`RANDOM}};
  l3_ramDatas_2_entries_perms_5_g = _RAND_1072[0:0];
  _RAND_1073 = {1{`RANDOM}};
  l3_ramDatas_2_entries_perms_5_u = _RAND_1073[0:0];
  _RAND_1074 = {1{`RANDOM}};
  l3_ramDatas_2_entries_perms_5_x = _RAND_1074[0:0];
  _RAND_1075 = {1{`RANDOM}};
  l3_ramDatas_2_entries_perms_5_w = _RAND_1075[0:0];
  _RAND_1076 = {1{`RANDOM}};
  l3_ramDatas_2_entries_perms_5_r = _RAND_1076[0:0];
  _RAND_1077 = {1{`RANDOM}};
  l3_ramDatas_2_entries_perms_6_d = _RAND_1077[0:0];
  _RAND_1078 = {1{`RANDOM}};
  l3_ramDatas_2_entries_perms_6_a = _RAND_1078[0:0];
  _RAND_1079 = {1{`RANDOM}};
  l3_ramDatas_2_entries_perms_6_g = _RAND_1079[0:0];
  _RAND_1080 = {1{`RANDOM}};
  l3_ramDatas_2_entries_perms_6_u = _RAND_1080[0:0];
  _RAND_1081 = {1{`RANDOM}};
  l3_ramDatas_2_entries_perms_6_x = _RAND_1081[0:0];
  _RAND_1082 = {1{`RANDOM}};
  l3_ramDatas_2_entries_perms_6_w = _RAND_1082[0:0];
  _RAND_1083 = {1{`RANDOM}};
  l3_ramDatas_2_entries_perms_6_r = _RAND_1083[0:0];
  _RAND_1084 = {1{`RANDOM}};
  l3_ramDatas_2_entries_perms_7_d = _RAND_1084[0:0];
  _RAND_1085 = {1{`RANDOM}};
  l3_ramDatas_2_entries_perms_7_a = _RAND_1085[0:0];
  _RAND_1086 = {1{`RANDOM}};
  l3_ramDatas_2_entries_perms_7_g = _RAND_1086[0:0];
  _RAND_1087 = {1{`RANDOM}};
  l3_ramDatas_2_entries_perms_7_u = _RAND_1087[0:0];
  _RAND_1088 = {1{`RANDOM}};
  l3_ramDatas_2_entries_perms_7_x = _RAND_1088[0:0];
  _RAND_1089 = {1{`RANDOM}};
  l3_ramDatas_2_entries_perms_7_w = _RAND_1089[0:0];
  _RAND_1090 = {1{`RANDOM}};
  l3_ramDatas_2_entries_perms_7_r = _RAND_1090[0:0];
  _RAND_1091 = {1{`RANDOM}};
  l3_ramDatas_2_entries_prefetch = _RAND_1091[0:0];
  _RAND_1092 = {2{`RANDOM}};
  l3_ramDatas_2_ecc = _RAND_1092[38:0];
  _RAND_1093 = {1{`RANDOM}};
  l3_ramDatas_3_entries_tag = _RAND_1093[21:0];
  _RAND_1094 = {1{`RANDOM}};
  l3_ramDatas_3_entries_asid = _RAND_1094[15:0];
  _RAND_1095 = {1{`RANDOM}};
  l3_ramDatas_3_entries_ppns_0 = _RAND_1095[23:0];
  _RAND_1096 = {1{`RANDOM}};
  l3_ramDatas_3_entries_ppns_1 = _RAND_1096[23:0];
  _RAND_1097 = {1{`RANDOM}};
  l3_ramDatas_3_entries_ppns_2 = _RAND_1097[23:0];
  _RAND_1098 = {1{`RANDOM}};
  l3_ramDatas_3_entries_ppns_3 = _RAND_1098[23:0];
  _RAND_1099 = {1{`RANDOM}};
  l3_ramDatas_3_entries_ppns_4 = _RAND_1099[23:0];
  _RAND_1100 = {1{`RANDOM}};
  l3_ramDatas_3_entries_ppns_5 = _RAND_1100[23:0];
  _RAND_1101 = {1{`RANDOM}};
  l3_ramDatas_3_entries_ppns_6 = _RAND_1101[23:0];
  _RAND_1102 = {1{`RANDOM}};
  l3_ramDatas_3_entries_ppns_7 = _RAND_1102[23:0];
  _RAND_1103 = {1{`RANDOM}};
  l3_ramDatas_3_entries_vs_0 = _RAND_1103[0:0];
  _RAND_1104 = {1{`RANDOM}};
  l3_ramDatas_3_entries_vs_1 = _RAND_1104[0:0];
  _RAND_1105 = {1{`RANDOM}};
  l3_ramDatas_3_entries_vs_2 = _RAND_1105[0:0];
  _RAND_1106 = {1{`RANDOM}};
  l3_ramDatas_3_entries_vs_3 = _RAND_1106[0:0];
  _RAND_1107 = {1{`RANDOM}};
  l3_ramDatas_3_entries_vs_4 = _RAND_1107[0:0];
  _RAND_1108 = {1{`RANDOM}};
  l3_ramDatas_3_entries_vs_5 = _RAND_1108[0:0];
  _RAND_1109 = {1{`RANDOM}};
  l3_ramDatas_3_entries_vs_6 = _RAND_1109[0:0];
  _RAND_1110 = {1{`RANDOM}};
  l3_ramDatas_3_entries_vs_7 = _RAND_1110[0:0];
  _RAND_1111 = {1{`RANDOM}};
  l3_ramDatas_3_entries_perms_0_d = _RAND_1111[0:0];
  _RAND_1112 = {1{`RANDOM}};
  l3_ramDatas_3_entries_perms_0_a = _RAND_1112[0:0];
  _RAND_1113 = {1{`RANDOM}};
  l3_ramDatas_3_entries_perms_0_g = _RAND_1113[0:0];
  _RAND_1114 = {1{`RANDOM}};
  l3_ramDatas_3_entries_perms_0_u = _RAND_1114[0:0];
  _RAND_1115 = {1{`RANDOM}};
  l3_ramDatas_3_entries_perms_0_x = _RAND_1115[0:0];
  _RAND_1116 = {1{`RANDOM}};
  l3_ramDatas_3_entries_perms_0_w = _RAND_1116[0:0];
  _RAND_1117 = {1{`RANDOM}};
  l3_ramDatas_3_entries_perms_0_r = _RAND_1117[0:0];
  _RAND_1118 = {1{`RANDOM}};
  l3_ramDatas_3_entries_perms_1_d = _RAND_1118[0:0];
  _RAND_1119 = {1{`RANDOM}};
  l3_ramDatas_3_entries_perms_1_a = _RAND_1119[0:0];
  _RAND_1120 = {1{`RANDOM}};
  l3_ramDatas_3_entries_perms_1_g = _RAND_1120[0:0];
  _RAND_1121 = {1{`RANDOM}};
  l3_ramDatas_3_entries_perms_1_u = _RAND_1121[0:0];
  _RAND_1122 = {1{`RANDOM}};
  l3_ramDatas_3_entries_perms_1_x = _RAND_1122[0:0];
  _RAND_1123 = {1{`RANDOM}};
  l3_ramDatas_3_entries_perms_1_w = _RAND_1123[0:0];
  _RAND_1124 = {1{`RANDOM}};
  l3_ramDatas_3_entries_perms_1_r = _RAND_1124[0:0];
  _RAND_1125 = {1{`RANDOM}};
  l3_ramDatas_3_entries_perms_2_d = _RAND_1125[0:0];
  _RAND_1126 = {1{`RANDOM}};
  l3_ramDatas_3_entries_perms_2_a = _RAND_1126[0:0];
  _RAND_1127 = {1{`RANDOM}};
  l3_ramDatas_3_entries_perms_2_g = _RAND_1127[0:0];
  _RAND_1128 = {1{`RANDOM}};
  l3_ramDatas_3_entries_perms_2_u = _RAND_1128[0:0];
  _RAND_1129 = {1{`RANDOM}};
  l3_ramDatas_3_entries_perms_2_x = _RAND_1129[0:0];
  _RAND_1130 = {1{`RANDOM}};
  l3_ramDatas_3_entries_perms_2_w = _RAND_1130[0:0];
  _RAND_1131 = {1{`RANDOM}};
  l3_ramDatas_3_entries_perms_2_r = _RAND_1131[0:0];
  _RAND_1132 = {1{`RANDOM}};
  l3_ramDatas_3_entries_perms_3_d = _RAND_1132[0:0];
  _RAND_1133 = {1{`RANDOM}};
  l3_ramDatas_3_entries_perms_3_a = _RAND_1133[0:0];
  _RAND_1134 = {1{`RANDOM}};
  l3_ramDatas_3_entries_perms_3_g = _RAND_1134[0:0];
  _RAND_1135 = {1{`RANDOM}};
  l3_ramDatas_3_entries_perms_3_u = _RAND_1135[0:0];
  _RAND_1136 = {1{`RANDOM}};
  l3_ramDatas_3_entries_perms_3_x = _RAND_1136[0:0];
  _RAND_1137 = {1{`RANDOM}};
  l3_ramDatas_3_entries_perms_3_w = _RAND_1137[0:0];
  _RAND_1138 = {1{`RANDOM}};
  l3_ramDatas_3_entries_perms_3_r = _RAND_1138[0:0];
  _RAND_1139 = {1{`RANDOM}};
  l3_ramDatas_3_entries_perms_4_d = _RAND_1139[0:0];
  _RAND_1140 = {1{`RANDOM}};
  l3_ramDatas_3_entries_perms_4_a = _RAND_1140[0:0];
  _RAND_1141 = {1{`RANDOM}};
  l3_ramDatas_3_entries_perms_4_g = _RAND_1141[0:0];
  _RAND_1142 = {1{`RANDOM}};
  l3_ramDatas_3_entries_perms_4_u = _RAND_1142[0:0];
  _RAND_1143 = {1{`RANDOM}};
  l3_ramDatas_3_entries_perms_4_x = _RAND_1143[0:0];
  _RAND_1144 = {1{`RANDOM}};
  l3_ramDatas_3_entries_perms_4_w = _RAND_1144[0:0];
  _RAND_1145 = {1{`RANDOM}};
  l3_ramDatas_3_entries_perms_4_r = _RAND_1145[0:0];
  _RAND_1146 = {1{`RANDOM}};
  l3_ramDatas_3_entries_perms_5_d = _RAND_1146[0:0];
  _RAND_1147 = {1{`RANDOM}};
  l3_ramDatas_3_entries_perms_5_a = _RAND_1147[0:0];
  _RAND_1148 = {1{`RANDOM}};
  l3_ramDatas_3_entries_perms_5_g = _RAND_1148[0:0];
  _RAND_1149 = {1{`RANDOM}};
  l3_ramDatas_3_entries_perms_5_u = _RAND_1149[0:0];
  _RAND_1150 = {1{`RANDOM}};
  l3_ramDatas_3_entries_perms_5_x = _RAND_1150[0:0];
  _RAND_1151 = {1{`RANDOM}};
  l3_ramDatas_3_entries_perms_5_w = _RAND_1151[0:0];
  _RAND_1152 = {1{`RANDOM}};
  l3_ramDatas_3_entries_perms_5_r = _RAND_1152[0:0];
  _RAND_1153 = {1{`RANDOM}};
  l3_ramDatas_3_entries_perms_6_d = _RAND_1153[0:0];
  _RAND_1154 = {1{`RANDOM}};
  l3_ramDatas_3_entries_perms_6_a = _RAND_1154[0:0];
  _RAND_1155 = {1{`RANDOM}};
  l3_ramDatas_3_entries_perms_6_g = _RAND_1155[0:0];
  _RAND_1156 = {1{`RANDOM}};
  l3_ramDatas_3_entries_perms_6_u = _RAND_1156[0:0];
  _RAND_1157 = {1{`RANDOM}};
  l3_ramDatas_3_entries_perms_6_x = _RAND_1157[0:0];
  _RAND_1158 = {1{`RANDOM}};
  l3_ramDatas_3_entries_perms_6_w = _RAND_1158[0:0];
  _RAND_1159 = {1{`RANDOM}};
  l3_ramDatas_3_entries_perms_6_r = _RAND_1159[0:0];
  _RAND_1160 = {1{`RANDOM}};
  l3_ramDatas_3_entries_perms_7_d = _RAND_1160[0:0];
  _RAND_1161 = {1{`RANDOM}};
  l3_ramDatas_3_entries_perms_7_a = _RAND_1161[0:0];
  _RAND_1162 = {1{`RANDOM}};
  l3_ramDatas_3_entries_perms_7_g = _RAND_1162[0:0];
  _RAND_1163 = {1{`RANDOM}};
  l3_ramDatas_3_entries_perms_7_u = _RAND_1163[0:0];
  _RAND_1164 = {1{`RANDOM}};
  l3_ramDatas_3_entries_perms_7_x = _RAND_1164[0:0];
  _RAND_1165 = {1{`RANDOM}};
  l3_ramDatas_3_entries_perms_7_w = _RAND_1165[0:0];
  _RAND_1166 = {1{`RANDOM}};
  l3_ramDatas_3_entries_perms_7_r = _RAND_1166[0:0];
  _RAND_1167 = {1{`RANDOM}};
  l3_ramDatas_3_entries_prefetch = _RAND_1167[0:0];
  _RAND_1168 = {2{`RANDOM}};
  l3_ramDatas_3_ecc = _RAND_1168[38:0];
  _RAND_1169 = {1{`RANDOM}};
  l3_ramDatas_4_entries_tag = _RAND_1169[21:0];
  _RAND_1170 = {1{`RANDOM}};
  l3_ramDatas_4_entries_asid = _RAND_1170[15:0];
  _RAND_1171 = {1{`RANDOM}};
  l3_ramDatas_4_entries_ppns_0 = _RAND_1171[23:0];
  _RAND_1172 = {1{`RANDOM}};
  l3_ramDatas_4_entries_ppns_1 = _RAND_1172[23:0];
  _RAND_1173 = {1{`RANDOM}};
  l3_ramDatas_4_entries_ppns_2 = _RAND_1173[23:0];
  _RAND_1174 = {1{`RANDOM}};
  l3_ramDatas_4_entries_ppns_3 = _RAND_1174[23:0];
  _RAND_1175 = {1{`RANDOM}};
  l3_ramDatas_4_entries_ppns_4 = _RAND_1175[23:0];
  _RAND_1176 = {1{`RANDOM}};
  l3_ramDatas_4_entries_ppns_5 = _RAND_1176[23:0];
  _RAND_1177 = {1{`RANDOM}};
  l3_ramDatas_4_entries_ppns_6 = _RAND_1177[23:0];
  _RAND_1178 = {1{`RANDOM}};
  l3_ramDatas_4_entries_ppns_7 = _RAND_1178[23:0];
  _RAND_1179 = {1{`RANDOM}};
  l3_ramDatas_4_entries_vs_0 = _RAND_1179[0:0];
  _RAND_1180 = {1{`RANDOM}};
  l3_ramDatas_4_entries_vs_1 = _RAND_1180[0:0];
  _RAND_1181 = {1{`RANDOM}};
  l3_ramDatas_4_entries_vs_2 = _RAND_1181[0:0];
  _RAND_1182 = {1{`RANDOM}};
  l3_ramDatas_4_entries_vs_3 = _RAND_1182[0:0];
  _RAND_1183 = {1{`RANDOM}};
  l3_ramDatas_4_entries_vs_4 = _RAND_1183[0:0];
  _RAND_1184 = {1{`RANDOM}};
  l3_ramDatas_4_entries_vs_5 = _RAND_1184[0:0];
  _RAND_1185 = {1{`RANDOM}};
  l3_ramDatas_4_entries_vs_6 = _RAND_1185[0:0];
  _RAND_1186 = {1{`RANDOM}};
  l3_ramDatas_4_entries_vs_7 = _RAND_1186[0:0];
  _RAND_1187 = {1{`RANDOM}};
  l3_ramDatas_4_entries_perms_0_d = _RAND_1187[0:0];
  _RAND_1188 = {1{`RANDOM}};
  l3_ramDatas_4_entries_perms_0_a = _RAND_1188[0:0];
  _RAND_1189 = {1{`RANDOM}};
  l3_ramDatas_4_entries_perms_0_g = _RAND_1189[0:0];
  _RAND_1190 = {1{`RANDOM}};
  l3_ramDatas_4_entries_perms_0_u = _RAND_1190[0:0];
  _RAND_1191 = {1{`RANDOM}};
  l3_ramDatas_4_entries_perms_0_x = _RAND_1191[0:0];
  _RAND_1192 = {1{`RANDOM}};
  l3_ramDatas_4_entries_perms_0_w = _RAND_1192[0:0];
  _RAND_1193 = {1{`RANDOM}};
  l3_ramDatas_4_entries_perms_0_r = _RAND_1193[0:0];
  _RAND_1194 = {1{`RANDOM}};
  l3_ramDatas_4_entries_perms_1_d = _RAND_1194[0:0];
  _RAND_1195 = {1{`RANDOM}};
  l3_ramDatas_4_entries_perms_1_a = _RAND_1195[0:0];
  _RAND_1196 = {1{`RANDOM}};
  l3_ramDatas_4_entries_perms_1_g = _RAND_1196[0:0];
  _RAND_1197 = {1{`RANDOM}};
  l3_ramDatas_4_entries_perms_1_u = _RAND_1197[0:0];
  _RAND_1198 = {1{`RANDOM}};
  l3_ramDatas_4_entries_perms_1_x = _RAND_1198[0:0];
  _RAND_1199 = {1{`RANDOM}};
  l3_ramDatas_4_entries_perms_1_w = _RAND_1199[0:0];
  _RAND_1200 = {1{`RANDOM}};
  l3_ramDatas_4_entries_perms_1_r = _RAND_1200[0:0];
  _RAND_1201 = {1{`RANDOM}};
  l3_ramDatas_4_entries_perms_2_d = _RAND_1201[0:0];
  _RAND_1202 = {1{`RANDOM}};
  l3_ramDatas_4_entries_perms_2_a = _RAND_1202[0:0];
  _RAND_1203 = {1{`RANDOM}};
  l3_ramDatas_4_entries_perms_2_g = _RAND_1203[0:0];
  _RAND_1204 = {1{`RANDOM}};
  l3_ramDatas_4_entries_perms_2_u = _RAND_1204[0:0];
  _RAND_1205 = {1{`RANDOM}};
  l3_ramDatas_4_entries_perms_2_x = _RAND_1205[0:0];
  _RAND_1206 = {1{`RANDOM}};
  l3_ramDatas_4_entries_perms_2_w = _RAND_1206[0:0];
  _RAND_1207 = {1{`RANDOM}};
  l3_ramDatas_4_entries_perms_2_r = _RAND_1207[0:0];
  _RAND_1208 = {1{`RANDOM}};
  l3_ramDatas_4_entries_perms_3_d = _RAND_1208[0:0];
  _RAND_1209 = {1{`RANDOM}};
  l3_ramDatas_4_entries_perms_3_a = _RAND_1209[0:0];
  _RAND_1210 = {1{`RANDOM}};
  l3_ramDatas_4_entries_perms_3_g = _RAND_1210[0:0];
  _RAND_1211 = {1{`RANDOM}};
  l3_ramDatas_4_entries_perms_3_u = _RAND_1211[0:0];
  _RAND_1212 = {1{`RANDOM}};
  l3_ramDatas_4_entries_perms_3_x = _RAND_1212[0:0];
  _RAND_1213 = {1{`RANDOM}};
  l3_ramDatas_4_entries_perms_3_w = _RAND_1213[0:0];
  _RAND_1214 = {1{`RANDOM}};
  l3_ramDatas_4_entries_perms_3_r = _RAND_1214[0:0];
  _RAND_1215 = {1{`RANDOM}};
  l3_ramDatas_4_entries_perms_4_d = _RAND_1215[0:0];
  _RAND_1216 = {1{`RANDOM}};
  l3_ramDatas_4_entries_perms_4_a = _RAND_1216[0:0];
  _RAND_1217 = {1{`RANDOM}};
  l3_ramDatas_4_entries_perms_4_g = _RAND_1217[0:0];
  _RAND_1218 = {1{`RANDOM}};
  l3_ramDatas_4_entries_perms_4_u = _RAND_1218[0:0];
  _RAND_1219 = {1{`RANDOM}};
  l3_ramDatas_4_entries_perms_4_x = _RAND_1219[0:0];
  _RAND_1220 = {1{`RANDOM}};
  l3_ramDatas_4_entries_perms_4_w = _RAND_1220[0:0];
  _RAND_1221 = {1{`RANDOM}};
  l3_ramDatas_4_entries_perms_4_r = _RAND_1221[0:0];
  _RAND_1222 = {1{`RANDOM}};
  l3_ramDatas_4_entries_perms_5_d = _RAND_1222[0:0];
  _RAND_1223 = {1{`RANDOM}};
  l3_ramDatas_4_entries_perms_5_a = _RAND_1223[0:0];
  _RAND_1224 = {1{`RANDOM}};
  l3_ramDatas_4_entries_perms_5_g = _RAND_1224[0:0];
  _RAND_1225 = {1{`RANDOM}};
  l3_ramDatas_4_entries_perms_5_u = _RAND_1225[0:0];
  _RAND_1226 = {1{`RANDOM}};
  l3_ramDatas_4_entries_perms_5_x = _RAND_1226[0:0];
  _RAND_1227 = {1{`RANDOM}};
  l3_ramDatas_4_entries_perms_5_w = _RAND_1227[0:0];
  _RAND_1228 = {1{`RANDOM}};
  l3_ramDatas_4_entries_perms_5_r = _RAND_1228[0:0];
  _RAND_1229 = {1{`RANDOM}};
  l3_ramDatas_4_entries_perms_6_d = _RAND_1229[0:0];
  _RAND_1230 = {1{`RANDOM}};
  l3_ramDatas_4_entries_perms_6_a = _RAND_1230[0:0];
  _RAND_1231 = {1{`RANDOM}};
  l3_ramDatas_4_entries_perms_6_g = _RAND_1231[0:0];
  _RAND_1232 = {1{`RANDOM}};
  l3_ramDatas_4_entries_perms_6_u = _RAND_1232[0:0];
  _RAND_1233 = {1{`RANDOM}};
  l3_ramDatas_4_entries_perms_6_x = _RAND_1233[0:0];
  _RAND_1234 = {1{`RANDOM}};
  l3_ramDatas_4_entries_perms_6_w = _RAND_1234[0:0];
  _RAND_1235 = {1{`RANDOM}};
  l3_ramDatas_4_entries_perms_6_r = _RAND_1235[0:0];
  _RAND_1236 = {1{`RANDOM}};
  l3_ramDatas_4_entries_perms_7_d = _RAND_1236[0:0];
  _RAND_1237 = {1{`RANDOM}};
  l3_ramDatas_4_entries_perms_7_a = _RAND_1237[0:0];
  _RAND_1238 = {1{`RANDOM}};
  l3_ramDatas_4_entries_perms_7_g = _RAND_1238[0:0];
  _RAND_1239 = {1{`RANDOM}};
  l3_ramDatas_4_entries_perms_7_u = _RAND_1239[0:0];
  _RAND_1240 = {1{`RANDOM}};
  l3_ramDatas_4_entries_perms_7_x = _RAND_1240[0:0];
  _RAND_1241 = {1{`RANDOM}};
  l3_ramDatas_4_entries_perms_7_w = _RAND_1241[0:0];
  _RAND_1242 = {1{`RANDOM}};
  l3_ramDatas_4_entries_perms_7_r = _RAND_1242[0:0];
  _RAND_1243 = {1{`RANDOM}};
  l3_ramDatas_4_entries_prefetch = _RAND_1243[0:0];
  _RAND_1244 = {2{`RANDOM}};
  l3_ramDatas_4_ecc = _RAND_1244[38:0];
  _RAND_1245 = {1{`RANDOM}};
  l3_ramDatas_5_entries_tag = _RAND_1245[21:0];
  _RAND_1246 = {1{`RANDOM}};
  l3_ramDatas_5_entries_asid = _RAND_1246[15:0];
  _RAND_1247 = {1{`RANDOM}};
  l3_ramDatas_5_entries_ppns_0 = _RAND_1247[23:0];
  _RAND_1248 = {1{`RANDOM}};
  l3_ramDatas_5_entries_ppns_1 = _RAND_1248[23:0];
  _RAND_1249 = {1{`RANDOM}};
  l3_ramDatas_5_entries_ppns_2 = _RAND_1249[23:0];
  _RAND_1250 = {1{`RANDOM}};
  l3_ramDatas_5_entries_ppns_3 = _RAND_1250[23:0];
  _RAND_1251 = {1{`RANDOM}};
  l3_ramDatas_5_entries_ppns_4 = _RAND_1251[23:0];
  _RAND_1252 = {1{`RANDOM}};
  l3_ramDatas_5_entries_ppns_5 = _RAND_1252[23:0];
  _RAND_1253 = {1{`RANDOM}};
  l3_ramDatas_5_entries_ppns_6 = _RAND_1253[23:0];
  _RAND_1254 = {1{`RANDOM}};
  l3_ramDatas_5_entries_ppns_7 = _RAND_1254[23:0];
  _RAND_1255 = {1{`RANDOM}};
  l3_ramDatas_5_entries_vs_0 = _RAND_1255[0:0];
  _RAND_1256 = {1{`RANDOM}};
  l3_ramDatas_5_entries_vs_1 = _RAND_1256[0:0];
  _RAND_1257 = {1{`RANDOM}};
  l3_ramDatas_5_entries_vs_2 = _RAND_1257[0:0];
  _RAND_1258 = {1{`RANDOM}};
  l3_ramDatas_5_entries_vs_3 = _RAND_1258[0:0];
  _RAND_1259 = {1{`RANDOM}};
  l3_ramDatas_5_entries_vs_4 = _RAND_1259[0:0];
  _RAND_1260 = {1{`RANDOM}};
  l3_ramDatas_5_entries_vs_5 = _RAND_1260[0:0];
  _RAND_1261 = {1{`RANDOM}};
  l3_ramDatas_5_entries_vs_6 = _RAND_1261[0:0];
  _RAND_1262 = {1{`RANDOM}};
  l3_ramDatas_5_entries_vs_7 = _RAND_1262[0:0];
  _RAND_1263 = {1{`RANDOM}};
  l3_ramDatas_5_entries_perms_0_d = _RAND_1263[0:0];
  _RAND_1264 = {1{`RANDOM}};
  l3_ramDatas_5_entries_perms_0_a = _RAND_1264[0:0];
  _RAND_1265 = {1{`RANDOM}};
  l3_ramDatas_5_entries_perms_0_g = _RAND_1265[0:0];
  _RAND_1266 = {1{`RANDOM}};
  l3_ramDatas_5_entries_perms_0_u = _RAND_1266[0:0];
  _RAND_1267 = {1{`RANDOM}};
  l3_ramDatas_5_entries_perms_0_x = _RAND_1267[0:0];
  _RAND_1268 = {1{`RANDOM}};
  l3_ramDatas_5_entries_perms_0_w = _RAND_1268[0:0];
  _RAND_1269 = {1{`RANDOM}};
  l3_ramDatas_5_entries_perms_0_r = _RAND_1269[0:0];
  _RAND_1270 = {1{`RANDOM}};
  l3_ramDatas_5_entries_perms_1_d = _RAND_1270[0:0];
  _RAND_1271 = {1{`RANDOM}};
  l3_ramDatas_5_entries_perms_1_a = _RAND_1271[0:0];
  _RAND_1272 = {1{`RANDOM}};
  l3_ramDatas_5_entries_perms_1_g = _RAND_1272[0:0];
  _RAND_1273 = {1{`RANDOM}};
  l3_ramDatas_5_entries_perms_1_u = _RAND_1273[0:0];
  _RAND_1274 = {1{`RANDOM}};
  l3_ramDatas_5_entries_perms_1_x = _RAND_1274[0:0];
  _RAND_1275 = {1{`RANDOM}};
  l3_ramDatas_5_entries_perms_1_w = _RAND_1275[0:0];
  _RAND_1276 = {1{`RANDOM}};
  l3_ramDatas_5_entries_perms_1_r = _RAND_1276[0:0];
  _RAND_1277 = {1{`RANDOM}};
  l3_ramDatas_5_entries_perms_2_d = _RAND_1277[0:0];
  _RAND_1278 = {1{`RANDOM}};
  l3_ramDatas_5_entries_perms_2_a = _RAND_1278[0:0];
  _RAND_1279 = {1{`RANDOM}};
  l3_ramDatas_5_entries_perms_2_g = _RAND_1279[0:0];
  _RAND_1280 = {1{`RANDOM}};
  l3_ramDatas_5_entries_perms_2_u = _RAND_1280[0:0];
  _RAND_1281 = {1{`RANDOM}};
  l3_ramDatas_5_entries_perms_2_x = _RAND_1281[0:0];
  _RAND_1282 = {1{`RANDOM}};
  l3_ramDatas_5_entries_perms_2_w = _RAND_1282[0:0];
  _RAND_1283 = {1{`RANDOM}};
  l3_ramDatas_5_entries_perms_2_r = _RAND_1283[0:0];
  _RAND_1284 = {1{`RANDOM}};
  l3_ramDatas_5_entries_perms_3_d = _RAND_1284[0:0];
  _RAND_1285 = {1{`RANDOM}};
  l3_ramDatas_5_entries_perms_3_a = _RAND_1285[0:0];
  _RAND_1286 = {1{`RANDOM}};
  l3_ramDatas_5_entries_perms_3_g = _RAND_1286[0:0];
  _RAND_1287 = {1{`RANDOM}};
  l3_ramDatas_5_entries_perms_3_u = _RAND_1287[0:0];
  _RAND_1288 = {1{`RANDOM}};
  l3_ramDatas_5_entries_perms_3_x = _RAND_1288[0:0];
  _RAND_1289 = {1{`RANDOM}};
  l3_ramDatas_5_entries_perms_3_w = _RAND_1289[0:0];
  _RAND_1290 = {1{`RANDOM}};
  l3_ramDatas_5_entries_perms_3_r = _RAND_1290[0:0];
  _RAND_1291 = {1{`RANDOM}};
  l3_ramDatas_5_entries_perms_4_d = _RAND_1291[0:0];
  _RAND_1292 = {1{`RANDOM}};
  l3_ramDatas_5_entries_perms_4_a = _RAND_1292[0:0];
  _RAND_1293 = {1{`RANDOM}};
  l3_ramDatas_5_entries_perms_4_g = _RAND_1293[0:0];
  _RAND_1294 = {1{`RANDOM}};
  l3_ramDatas_5_entries_perms_4_u = _RAND_1294[0:0];
  _RAND_1295 = {1{`RANDOM}};
  l3_ramDatas_5_entries_perms_4_x = _RAND_1295[0:0];
  _RAND_1296 = {1{`RANDOM}};
  l3_ramDatas_5_entries_perms_4_w = _RAND_1296[0:0];
  _RAND_1297 = {1{`RANDOM}};
  l3_ramDatas_5_entries_perms_4_r = _RAND_1297[0:0];
  _RAND_1298 = {1{`RANDOM}};
  l3_ramDatas_5_entries_perms_5_d = _RAND_1298[0:0];
  _RAND_1299 = {1{`RANDOM}};
  l3_ramDatas_5_entries_perms_5_a = _RAND_1299[0:0];
  _RAND_1300 = {1{`RANDOM}};
  l3_ramDatas_5_entries_perms_5_g = _RAND_1300[0:0];
  _RAND_1301 = {1{`RANDOM}};
  l3_ramDatas_5_entries_perms_5_u = _RAND_1301[0:0];
  _RAND_1302 = {1{`RANDOM}};
  l3_ramDatas_5_entries_perms_5_x = _RAND_1302[0:0];
  _RAND_1303 = {1{`RANDOM}};
  l3_ramDatas_5_entries_perms_5_w = _RAND_1303[0:0];
  _RAND_1304 = {1{`RANDOM}};
  l3_ramDatas_5_entries_perms_5_r = _RAND_1304[0:0];
  _RAND_1305 = {1{`RANDOM}};
  l3_ramDatas_5_entries_perms_6_d = _RAND_1305[0:0];
  _RAND_1306 = {1{`RANDOM}};
  l3_ramDatas_5_entries_perms_6_a = _RAND_1306[0:0];
  _RAND_1307 = {1{`RANDOM}};
  l3_ramDatas_5_entries_perms_6_g = _RAND_1307[0:0];
  _RAND_1308 = {1{`RANDOM}};
  l3_ramDatas_5_entries_perms_6_u = _RAND_1308[0:0];
  _RAND_1309 = {1{`RANDOM}};
  l3_ramDatas_5_entries_perms_6_x = _RAND_1309[0:0];
  _RAND_1310 = {1{`RANDOM}};
  l3_ramDatas_5_entries_perms_6_w = _RAND_1310[0:0];
  _RAND_1311 = {1{`RANDOM}};
  l3_ramDatas_5_entries_perms_6_r = _RAND_1311[0:0];
  _RAND_1312 = {1{`RANDOM}};
  l3_ramDatas_5_entries_perms_7_d = _RAND_1312[0:0];
  _RAND_1313 = {1{`RANDOM}};
  l3_ramDatas_5_entries_perms_7_a = _RAND_1313[0:0];
  _RAND_1314 = {1{`RANDOM}};
  l3_ramDatas_5_entries_perms_7_g = _RAND_1314[0:0];
  _RAND_1315 = {1{`RANDOM}};
  l3_ramDatas_5_entries_perms_7_u = _RAND_1315[0:0];
  _RAND_1316 = {1{`RANDOM}};
  l3_ramDatas_5_entries_perms_7_x = _RAND_1316[0:0];
  _RAND_1317 = {1{`RANDOM}};
  l3_ramDatas_5_entries_perms_7_w = _RAND_1317[0:0];
  _RAND_1318 = {1{`RANDOM}};
  l3_ramDatas_5_entries_perms_7_r = _RAND_1318[0:0];
  _RAND_1319 = {1{`RANDOM}};
  l3_ramDatas_5_entries_prefetch = _RAND_1319[0:0];
  _RAND_1320 = {2{`RANDOM}};
  l3_ramDatas_5_ecc = _RAND_1320[38:0];
  _RAND_1321 = {1{`RANDOM}};
  l3_ramDatas_6_entries_tag = _RAND_1321[21:0];
  _RAND_1322 = {1{`RANDOM}};
  l3_ramDatas_6_entries_asid = _RAND_1322[15:0];
  _RAND_1323 = {1{`RANDOM}};
  l3_ramDatas_6_entries_ppns_0 = _RAND_1323[23:0];
  _RAND_1324 = {1{`RANDOM}};
  l3_ramDatas_6_entries_ppns_1 = _RAND_1324[23:0];
  _RAND_1325 = {1{`RANDOM}};
  l3_ramDatas_6_entries_ppns_2 = _RAND_1325[23:0];
  _RAND_1326 = {1{`RANDOM}};
  l3_ramDatas_6_entries_ppns_3 = _RAND_1326[23:0];
  _RAND_1327 = {1{`RANDOM}};
  l3_ramDatas_6_entries_ppns_4 = _RAND_1327[23:0];
  _RAND_1328 = {1{`RANDOM}};
  l3_ramDatas_6_entries_ppns_5 = _RAND_1328[23:0];
  _RAND_1329 = {1{`RANDOM}};
  l3_ramDatas_6_entries_ppns_6 = _RAND_1329[23:0];
  _RAND_1330 = {1{`RANDOM}};
  l3_ramDatas_6_entries_ppns_7 = _RAND_1330[23:0];
  _RAND_1331 = {1{`RANDOM}};
  l3_ramDatas_6_entries_vs_0 = _RAND_1331[0:0];
  _RAND_1332 = {1{`RANDOM}};
  l3_ramDatas_6_entries_vs_1 = _RAND_1332[0:0];
  _RAND_1333 = {1{`RANDOM}};
  l3_ramDatas_6_entries_vs_2 = _RAND_1333[0:0];
  _RAND_1334 = {1{`RANDOM}};
  l3_ramDatas_6_entries_vs_3 = _RAND_1334[0:0];
  _RAND_1335 = {1{`RANDOM}};
  l3_ramDatas_6_entries_vs_4 = _RAND_1335[0:0];
  _RAND_1336 = {1{`RANDOM}};
  l3_ramDatas_6_entries_vs_5 = _RAND_1336[0:0];
  _RAND_1337 = {1{`RANDOM}};
  l3_ramDatas_6_entries_vs_6 = _RAND_1337[0:0];
  _RAND_1338 = {1{`RANDOM}};
  l3_ramDatas_6_entries_vs_7 = _RAND_1338[0:0];
  _RAND_1339 = {1{`RANDOM}};
  l3_ramDatas_6_entries_perms_0_d = _RAND_1339[0:0];
  _RAND_1340 = {1{`RANDOM}};
  l3_ramDatas_6_entries_perms_0_a = _RAND_1340[0:0];
  _RAND_1341 = {1{`RANDOM}};
  l3_ramDatas_6_entries_perms_0_g = _RAND_1341[0:0];
  _RAND_1342 = {1{`RANDOM}};
  l3_ramDatas_6_entries_perms_0_u = _RAND_1342[0:0];
  _RAND_1343 = {1{`RANDOM}};
  l3_ramDatas_6_entries_perms_0_x = _RAND_1343[0:0];
  _RAND_1344 = {1{`RANDOM}};
  l3_ramDatas_6_entries_perms_0_w = _RAND_1344[0:0];
  _RAND_1345 = {1{`RANDOM}};
  l3_ramDatas_6_entries_perms_0_r = _RAND_1345[0:0];
  _RAND_1346 = {1{`RANDOM}};
  l3_ramDatas_6_entries_perms_1_d = _RAND_1346[0:0];
  _RAND_1347 = {1{`RANDOM}};
  l3_ramDatas_6_entries_perms_1_a = _RAND_1347[0:0];
  _RAND_1348 = {1{`RANDOM}};
  l3_ramDatas_6_entries_perms_1_g = _RAND_1348[0:0];
  _RAND_1349 = {1{`RANDOM}};
  l3_ramDatas_6_entries_perms_1_u = _RAND_1349[0:0];
  _RAND_1350 = {1{`RANDOM}};
  l3_ramDatas_6_entries_perms_1_x = _RAND_1350[0:0];
  _RAND_1351 = {1{`RANDOM}};
  l3_ramDatas_6_entries_perms_1_w = _RAND_1351[0:0];
  _RAND_1352 = {1{`RANDOM}};
  l3_ramDatas_6_entries_perms_1_r = _RAND_1352[0:0];
  _RAND_1353 = {1{`RANDOM}};
  l3_ramDatas_6_entries_perms_2_d = _RAND_1353[0:0];
  _RAND_1354 = {1{`RANDOM}};
  l3_ramDatas_6_entries_perms_2_a = _RAND_1354[0:0];
  _RAND_1355 = {1{`RANDOM}};
  l3_ramDatas_6_entries_perms_2_g = _RAND_1355[0:0];
  _RAND_1356 = {1{`RANDOM}};
  l3_ramDatas_6_entries_perms_2_u = _RAND_1356[0:0];
  _RAND_1357 = {1{`RANDOM}};
  l3_ramDatas_6_entries_perms_2_x = _RAND_1357[0:0];
  _RAND_1358 = {1{`RANDOM}};
  l3_ramDatas_6_entries_perms_2_w = _RAND_1358[0:0];
  _RAND_1359 = {1{`RANDOM}};
  l3_ramDatas_6_entries_perms_2_r = _RAND_1359[0:0];
  _RAND_1360 = {1{`RANDOM}};
  l3_ramDatas_6_entries_perms_3_d = _RAND_1360[0:0];
  _RAND_1361 = {1{`RANDOM}};
  l3_ramDatas_6_entries_perms_3_a = _RAND_1361[0:0];
  _RAND_1362 = {1{`RANDOM}};
  l3_ramDatas_6_entries_perms_3_g = _RAND_1362[0:0];
  _RAND_1363 = {1{`RANDOM}};
  l3_ramDatas_6_entries_perms_3_u = _RAND_1363[0:0];
  _RAND_1364 = {1{`RANDOM}};
  l3_ramDatas_6_entries_perms_3_x = _RAND_1364[0:0];
  _RAND_1365 = {1{`RANDOM}};
  l3_ramDatas_6_entries_perms_3_w = _RAND_1365[0:0];
  _RAND_1366 = {1{`RANDOM}};
  l3_ramDatas_6_entries_perms_3_r = _RAND_1366[0:0];
  _RAND_1367 = {1{`RANDOM}};
  l3_ramDatas_6_entries_perms_4_d = _RAND_1367[0:0];
  _RAND_1368 = {1{`RANDOM}};
  l3_ramDatas_6_entries_perms_4_a = _RAND_1368[0:0];
  _RAND_1369 = {1{`RANDOM}};
  l3_ramDatas_6_entries_perms_4_g = _RAND_1369[0:0];
  _RAND_1370 = {1{`RANDOM}};
  l3_ramDatas_6_entries_perms_4_u = _RAND_1370[0:0];
  _RAND_1371 = {1{`RANDOM}};
  l3_ramDatas_6_entries_perms_4_x = _RAND_1371[0:0];
  _RAND_1372 = {1{`RANDOM}};
  l3_ramDatas_6_entries_perms_4_w = _RAND_1372[0:0];
  _RAND_1373 = {1{`RANDOM}};
  l3_ramDatas_6_entries_perms_4_r = _RAND_1373[0:0];
  _RAND_1374 = {1{`RANDOM}};
  l3_ramDatas_6_entries_perms_5_d = _RAND_1374[0:0];
  _RAND_1375 = {1{`RANDOM}};
  l3_ramDatas_6_entries_perms_5_a = _RAND_1375[0:0];
  _RAND_1376 = {1{`RANDOM}};
  l3_ramDatas_6_entries_perms_5_g = _RAND_1376[0:0];
  _RAND_1377 = {1{`RANDOM}};
  l3_ramDatas_6_entries_perms_5_u = _RAND_1377[0:0];
  _RAND_1378 = {1{`RANDOM}};
  l3_ramDatas_6_entries_perms_5_x = _RAND_1378[0:0];
  _RAND_1379 = {1{`RANDOM}};
  l3_ramDatas_6_entries_perms_5_w = _RAND_1379[0:0];
  _RAND_1380 = {1{`RANDOM}};
  l3_ramDatas_6_entries_perms_5_r = _RAND_1380[0:0];
  _RAND_1381 = {1{`RANDOM}};
  l3_ramDatas_6_entries_perms_6_d = _RAND_1381[0:0];
  _RAND_1382 = {1{`RANDOM}};
  l3_ramDatas_6_entries_perms_6_a = _RAND_1382[0:0];
  _RAND_1383 = {1{`RANDOM}};
  l3_ramDatas_6_entries_perms_6_g = _RAND_1383[0:0];
  _RAND_1384 = {1{`RANDOM}};
  l3_ramDatas_6_entries_perms_6_u = _RAND_1384[0:0];
  _RAND_1385 = {1{`RANDOM}};
  l3_ramDatas_6_entries_perms_6_x = _RAND_1385[0:0];
  _RAND_1386 = {1{`RANDOM}};
  l3_ramDatas_6_entries_perms_6_w = _RAND_1386[0:0];
  _RAND_1387 = {1{`RANDOM}};
  l3_ramDatas_6_entries_perms_6_r = _RAND_1387[0:0];
  _RAND_1388 = {1{`RANDOM}};
  l3_ramDatas_6_entries_perms_7_d = _RAND_1388[0:0];
  _RAND_1389 = {1{`RANDOM}};
  l3_ramDatas_6_entries_perms_7_a = _RAND_1389[0:0];
  _RAND_1390 = {1{`RANDOM}};
  l3_ramDatas_6_entries_perms_7_g = _RAND_1390[0:0];
  _RAND_1391 = {1{`RANDOM}};
  l3_ramDatas_6_entries_perms_7_u = _RAND_1391[0:0];
  _RAND_1392 = {1{`RANDOM}};
  l3_ramDatas_6_entries_perms_7_x = _RAND_1392[0:0];
  _RAND_1393 = {1{`RANDOM}};
  l3_ramDatas_6_entries_perms_7_w = _RAND_1393[0:0];
  _RAND_1394 = {1{`RANDOM}};
  l3_ramDatas_6_entries_perms_7_r = _RAND_1394[0:0];
  _RAND_1395 = {1{`RANDOM}};
  l3_ramDatas_6_entries_prefetch = _RAND_1395[0:0];
  _RAND_1396 = {2{`RANDOM}};
  l3_ramDatas_6_ecc = _RAND_1396[38:0];
  _RAND_1397 = {1{`RANDOM}};
  l3_ramDatas_7_entries_tag = _RAND_1397[21:0];
  _RAND_1398 = {1{`RANDOM}};
  l3_ramDatas_7_entries_asid = _RAND_1398[15:0];
  _RAND_1399 = {1{`RANDOM}};
  l3_ramDatas_7_entries_ppns_0 = _RAND_1399[23:0];
  _RAND_1400 = {1{`RANDOM}};
  l3_ramDatas_7_entries_ppns_1 = _RAND_1400[23:0];
  _RAND_1401 = {1{`RANDOM}};
  l3_ramDatas_7_entries_ppns_2 = _RAND_1401[23:0];
  _RAND_1402 = {1{`RANDOM}};
  l3_ramDatas_7_entries_ppns_3 = _RAND_1402[23:0];
  _RAND_1403 = {1{`RANDOM}};
  l3_ramDatas_7_entries_ppns_4 = _RAND_1403[23:0];
  _RAND_1404 = {1{`RANDOM}};
  l3_ramDatas_7_entries_ppns_5 = _RAND_1404[23:0];
  _RAND_1405 = {1{`RANDOM}};
  l3_ramDatas_7_entries_ppns_6 = _RAND_1405[23:0];
  _RAND_1406 = {1{`RANDOM}};
  l3_ramDatas_7_entries_ppns_7 = _RAND_1406[23:0];
  _RAND_1407 = {1{`RANDOM}};
  l3_ramDatas_7_entries_vs_0 = _RAND_1407[0:0];
  _RAND_1408 = {1{`RANDOM}};
  l3_ramDatas_7_entries_vs_1 = _RAND_1408[0:0];
  _RAND_1409 = {1{`RANDOM}};
  l3_ramDatas_7_entries_vs_2 = _RAND_1409[0:0];
  _RAND_1410 = {1{`RANDOM}};
  l3_ramDatas_7_entries_vs_3 = _RAND_1410[0:0];
  _RAND_1411 = {1{`RANDOM}};
  l3_ramDatas_7_entries_vs_4 = _RAND_1411[0:0];
  _RAND_1412 = {1{`RANDOM}};
  l3_ramDatas_7_entries_vs_5 = _RAND_1412[0:0];
  _RAND_1413 = {1{`RANDOM}};
  l3_ramDatas_7_entries_vs_6 = _RAND_1413[0:0];
  _RAND_1414 = {1{`RANDOM}};
  l3_ramDatas_7_entries_vs_7 = _RAND_1414[0:0];
  _RAND_1415 = {1{`RANDOM}};
  l3_ramDatas_7_entries_perms_0_d = _RAND_1415[0:0];
  _RAND_1416 = {1{`RANDOM}};
  l3_ramDatas_7_entries_perms_0_a = _RAND_1416[0:0];
  _RAND_1417 = {1{`RANDOM}};
  l3_ramDatas_7_entries_perms_0_g = _RAND_1417[0:0];
  _RAND_1418 = {1{`RANDOM}};
  l3_ramDatas_7_entries_perms_0_u = _RAND_1418[0:0];
  _RAND_1419 = {1{`RANDOM}};
  l3_ramDatas_7_entries_perms_0_x = _RAND_1419[0:0];
  _RAND_1420 = {1{`RANDOM}};
  l3_ramDatas_7_entries_perms_0_w = _RAND_1420[0:0];
  _RAND_1421 = {1{`RANDOM}};
  l3_ramDatas_7_entries_perms_0_r = _RAND_1421[0:0];
  _RAND_1422 = {1{`RANDOM}};
  l3_ramDatas_7_entries_perms_1_d = _RAND_1422[0:0];
  _RAND_1423 = {1{`RANDOM}};
  l3_ramDatas_7_entries_perms_1_a = _RAND_1423[0:0];
  _RAND_1424 = {1{`RANDOM}};
  l3_ramDatas_7_entries_perms_1_g = _RAND_1424[0:0];
  _RAND_1425 = {1{`RANDOM}};
  l3_ramDatas_7_entries_perms_1_u = _RAND_1425[0:0];
  _RAND_1426 = {1{`RANDOM}};
  l3_ramDatas_7_entries_perms_1_x = _RAND_1426[0:0];
  _RAND_1427 = {1{`RANDOM}};
  l3_ramDatas_7_entries_perms_1_w = _RAND_1427[0:0];
  _RAND_1428 = {1{`RANDOM}};
  l3_ramDatas_7_entries_perms_1_r = _RAND_1428[0:0];
  _RAND_1429 = {1{`RANDOM}};
  l3_ramDatas_7_entries_perms_2_d = _RAND_1429[0:0];
  _RAND_1430 = {1{`RANDOM}};
  l3_ramDatas_7_entries_perms_2_a = _RAND_1430[0:0];
  _RAND_1431 = {1{`RANDOM}};
  l3_ramDatas_7_entries_perms_2_g = _RAND_1431[0:0];
  _RAND_1432 = {1{`RANDOM}};
  l3_ramDatas_7_entries_perms_2_u = _RAND_1432[0:0];
  _RAND_1433 = {1{`RANDOM}};
  l3_ramDatas_7_entries_perms_2_x = _RAND_1433[0:0];
  _RAND_1434 = {1{`RANDOM}};
  l3_ramDatas_7_entries_perms_2_w = _RAND_1434[0:0];
  _RAND_1435 = {1{`RANDOM}};
  l3_ramDatas_7_entries_perms_2_r = _RAND_1435[0:0];
  _RAND_1436 = {1{`RANDOM}};
  l3_ramDatas_7_entries_perms_3_d = _RAND_1436[0:0];
  _RAND_1437 = {1{`RANDOM}};
  l3_ramDatas_7_entries_perms_3_a = _RAND_1437[0:0];
  _RAND_1438 = {1{`RANDOM}};
  l3_ramDatas_7_entries_perms_3_g = _RAND_1438[0:0];
  _RAND_1439 = {1{`RANDOM}};
  l3_ramDatas_7_entries_perms_3_u = _RAND_1439[0:0];
  _RAND_1440 = {1{`RANDOM}};
  l3_ramDatas_7_entries_perms_3_x = _RAND_1440[0:0];
  _RAND_1441 = {1{`RANDOM}};
  l3_ramDatas_7_entries_perms_3_w = _RAND_1441[0:0];
  _RAND_1442 = {1{`RANDOM}};
  l3_ramDatas_7_entries_perms_3_r = _RAND_1442[0:0];
  _RAND_1443 = {1{`RANDOM}};
  l3_ramDatas_7_entries_perms_4_d = _RAND_1443[0:0];
  _RAND_1444 = {1{`RANDOM}};
  l3_ramDatas_7_entries_perms_4_a = _RAND_1444[0:0];
  _RAND_1445 = {1{`RANDOM}};
  l3_ramDatas_7_entries_perms_4_g = _RAND_1445[0:0];
  _RAND_1446 = {1{`RANDOM}};
  l3_ramDatas_7_entries_perms_4_u = _RAND_1446[0:0];
  _RAND_1447 = {1{`RANDOM}};
  l3_ramDatas_7_entries_perms_4_x = _RAND_1447[0:0];
  _RAND_1448 = {1{`RANDOM}};
  l3_ramDatas_7_entries_perms_4_w = _RAND_1448[0:0];
  _RAND_1449 = {1{`RANDOM}};
  l3_ramDatas_7_entries_perms_4_r = _RAND_1449[0:0];
  _RAND_1450 = {1{`RANDOM}};
  l3_ramDatas_7_entries_perms_5_d = _RAND_1450[0:0];
  _RAND_1451 = {1{`RANDOM}};
  l3_ramDatas_7_entries_perms_5_a = _RAND_1451[0:0];
  _RAND_1452 = {1{`RANDOM}};
  l3_ramDatas_7_entries_perms_5_g = _RAND_1452[0:0];
  _RAND_1453 = {1{`RANDOM}};
  l3_ramDatas_7_entries_perms_5_u = _RAND_1453[0:0];
  _RAND_1454 = {1{`RANDOM}};
  l3_ramDatas_7_entries_perms_5_x = _RAND_1454[0:0];
  _RAND_1455 = {1{`RANDOM}};
  l3_ramDatas_7_entries_perms_5_w = _RAND_1455[0:0];
  _RAND_1456 = {1{`RANDOM}};
  l3_ramDatas_7_entries_perms_5_r = _RAND_1456[0:0];
  _RAND_1457 = {1{`RANDOM}};
  l3_ramDatas_7_entries_perms_6_d = _RAND_1457[0:0];
  _RAND_1458 = {1{`RANDOM}};
  l3_ramDatas_7_entries_perms_6_a = _RAND_1458[0:0];
  _RAND_1459 = {1{`RANDOM}};
  l3_ramDatas_7_entries_perms_6_g = _RAND_1459[0:0];
  _RAND_1460 = {1{`RANDOM}};
  l3_ramDatas_7_entries_perms_6_u = _RAND_1460[0:0];
  _RAND_1461 = {1{`RANDOM}};
  l3_ramDatas_7_entries_perms_6_x = _RAND_1461[0:0];
  _RAND_1462 = {1{`RANDOM}};
  l3_ramDatas_7_entries_perms_6_w = _RAND_1462[0:0];
  _RAND_1463 = {1{`RANDOM}};
  l3_ramDatas_7_entries_perms_6_r = _RAND_1463[0:0];
  _RAND_1464 = {1{`RANDOM}};
  l3_ramDatas_7_entries_perms_7_d = _RAND_1464[0:0];
  _RAND_1465 = {1{`RANDOM}};
  l3_ramDatas_7_entries_perms_7_a = _RAND_1465[0:0];
  _RAND_1466 = {1{`RANDOM}};
  l3_ramDatas_7_entries_perms_7_g = _RAND_1466[0:0];
  _RAND_1467 = {1{`RANDOM}};
  l3_ramDatas_7_entries_perms_7_u = _RAND_1467[0:0];
  _RAND_1468 = {1{`RANDOM}};
  l3_ramDatas_7_entries_perms_7_x = _RAND_1468[0:0];
  _RAND_1469 = {1{`RANDOM}};
  l3_ramDatas_7_entries_perms_7_w = _RAND_1469[0:0];
  _RAND_1470 = {1{`RANDOM}};
  l3_ramDatas_7_entries_perms_7_r = _RAND_1470[0:0];
  _RAND_1471 = {1{`RANDOM}};
  l3_ramDatas_7_entries_prefetch = _RAND_1471[0:0];
  _RAND_1472 = {2{`RANDOM}};
  l3_ramDatas_7_ecc = _RAND_1472[38:0];
  _RAND_1473 = {1{`RANDOM}};
  l3_hitVec_0 = _RAND_1473[0:0];
  _RAND_1474 = {1{`RANDOM}};
  l3_hitVec_1 = _RAND_1474[0:0];
  _RAND_1475 = {1{`RANDOM}};
  l3_hitVec_2 = _RAND_1475[0:0];
  _RAND_1476 = {1{`RANDOM}};
  l3_hitVec_3 = _RAND_1476[0:0];
  _RAND_1477 = {1{`RANDOM}};
  l3_hitVec_4 = _RAND_1477[0:0];
  _RAND_1478 = {1{`RANDOM}};
  l3_hitVec_5 = _RAND_1478[0:0];
  _RAND_1479 = {1{`RANDOM}};
  l3_hitVec_6 = _RAND_1479[0:0];
  _RAND_1480 = {1{`RANDOM}};
  l3_hitVec_7 = _RAND_1480[0:0];
  _RAND_1481 = {1{`RANDOM}};
  state_reg_3 = _RAND_1481[0:0];
  _RAND_1482 = {1{`RANDOM}};
  r_13 = _RAND_1482[0:0];
  _RAND_1483 = {1{`RANDOM}};
  r_14 = _RAND_1483[0:0];
  _RAND_1484 = {1{`RANDOM}};
  spHit = _RAND_1484[0:0];
  _RAND_1485 = {1{`RANDOM}};
  spHitData_ppn = _RAND_1485[23:0];
  _RAND_1486 = {1{`RANDOM}};
  spHitData_perm_d = _RAND_1486[0:0];
  _RAND_1487 = {1{`RANDOM}};
  spHitData_perm_a = _RAND_1487[0:0];
  _RAND_1488 = {1{`RANDOM}};
  spHitData_perm_g = _RAND_1488[0:0];
  _RAND_1489 = {1{`RANDOM}};
  spHitData_perm_u = _RAND_1489[0:0];
  _RAND_1490 = {1{`RANDOM}};
  spHitData_perm_x = _RAND_1490[0:0];
  _RAND_1491 = {1{`RANDOM}};
  spHitData_perm_w = _RAND_1491[0:0];
  _RAND_1492 = {1{`RANDOM}};
  spHitData_perm_r = _RAND_1492[0:0];
  _RAND_1493 = {1{`RANDOM}};
  spHitData_level = _RAND_1493[1:0];
  _RAND_1494 = {1{`RANDOM}};
  spPre = _RAND_1494[0:0];
  _RAND_1495 = {1{`RANDOM}};
  spValid = _RAND_1495[0:0];
  _RAND_1496 = {1{`RANDOM}};
  resp_res_l1_hit = _RAND_1496[0:0];
  _RAND_1497 = {1{`RANDOM}};
  resp_res_l1_ppn = _RAND_1497[23:0];
  _RAND_1498 = {1{`RANDOM}};
  resp_res_l2_hit = _RAND_1498[0:0];
  _RAND_1499 = {1{`RANDOM}};
  resp_res_l2_ppn = _RAND_1499[23:0];
  _RAND_1500 = {1{`RANDOM}};
  resp_res_l2_ecc = _RAND_1500[0:0];
  _RAND_1501 = {1{`RANDOM}};
  resp_res_l3_hit = _RAND_1501[0:0];
  _RAND_1502 = {1{`RANDOM}};
  resp_res_l3_pre = _RAND_1502[0:0];
  _RAND_1503 = {1{`RANDOM}};
  resp_res_l3_ppn = _RAND_1503[23:0];
  _RAND_1504 = {1{`RANDOM}};
  resp_res_l3_perm_d = _RAND_1504[0:0];
  _RAND_1505 = {1{`RANDOM}};
  resp_res_l3_perm_a = _RAND_1505[0:0];
  _RAND_1506 = {1{`RANDOM}};
  resp_res_l3_perm_g = _RAND_1506[0:0];
  _RAND_1507 = {1{`RANDOM}};
  resp_res_l3_perm_u = _RAND_1507[0:0];
  _RAND_1508 = {1{`RANDOM}};
  resp_res_l3_perm_x = _RAND_1508[0:0];
  _RAND_1509 = {1{`RANDOM}};
  resp_res_l3_perm_w = _RAND_1509[0:0];
  _RAND_1510 = {1{`RANDOM}};
  resp_res_l3_perm_r = _RAND_1510[0:0];
  _RAND_1511 = {1{`RANDOM}};
  resp_res_l3_ecc = _RAND_1511[0:0];
  _RAND_1512 = {1{`RANDOM}};
  resp_res_l3_v = _RAND_1512[0:0];
  _RAND_1513 = {1{`RANDOM}};
  resp_res_sp_hit = _RAND_1513[0:0];
  _RAND_1514 = {1{`RANDOM}};
  resp_res_sp_pre = _RAND_1514[0:0];
  _RAND_1515 = {1{`RANDOM}};
  resp_res_sp_ppn = _RAND_1515[23:0];
  _RAND_1516 = {1{`RANDOM}};
  resp_res_sp_perm_d = _RAND_1516[0:0];
  _RAND_1517 = {1{`RANDOM}};
  resp_res_sp_perm_a = _RAND_1517[0:0];
  _RAND_1518 = {1{`RANDOM}};
  resp_res_sp_perm_g = _RAND_1518[0:0];
  _RAND_1519 = {1{`RANDOM}};
  resp_res_sp_perm_u = _RAND_1519[0:0];
  _RAND_1520 = {1{`RANDOM}};
  resp_res_sp_perm_x = _RAND_1520[0:0];
  _RAND_1521 = {1{`RANDOM}};
  resp_res_sp_perm_w = _RAND_1521[0:0];
  _RAND_1522 = {1{`RANDOM}};
  resp_res_sp_perm_r = _RAND_1522[0:0];
  _RAND_1523 = {1{`RANDOM}};
  resp_res_sp_level = _RAND_1523[1:0];
  _RAND_1524 = {1{`RANDOM}};
  resp_res_sp_v = _RAND_1524[0:0];
  _RAND_1525 = {1{`RANDOM}};
  bypassed_0_valid = _RAND_1525[0:0];
  _RAND_1526 = {1{`RANDOM}};
  bypassed_0_valid_1 = _RAND_1526[0:0];
  _RAND_1527 = {1{`RANDOM}};
  bypassed_1_valid = _RAND_1527[0:0];
  _RAND_1528 = {1{`RANDOM}};
  bypassed_1_valid_1 = _RAND_1528[0:0];
  _RAND_1529 = {1{`RANDOM}};
  bypassed_2_valid = _RAND_1529[0:0];
  _RAND_1530 = {1{`RANDOM}};
  bypassed_2_valid_1 = _RAND_1530[0:0];
  _RAND_1531 = {1{`RANDOM}};
  io_perf_0_value_REG = _RAND_1531[0:0];
  _RAND_1532 = {1{`RANDOM}};
  io_perf_0_value_REG_1 = _RAND_1532[0:0];
  _RAND_1533 = {1{`RANDOM}};
  io_perf_1_value_REG = _RAND_1533[0:0];
  _RAND_1534 = {1{`RANDOM}};
  io_perf_1_value_REG_1 = _RAND_1534[0:0];
  _RAND_1535 = {1{`RANDOM}};
  io_perf_2_value_REG = _RAND_1535[0:0];
  _RAND_1536 = {1{`RANDOM}};
  io_perf_2_value_REG_1 = _RAND_1536[0:0];
  _RAND_1537 = {1{`RANDOM}};
  io_perf_3_value_REG = _RAND_1537[0:0];
  _RAND_1538 = {1{`RANDOM}};
  io_perf_3_value_REG_1 = _RAND_1538[0:0];
  _RAND_1539 = {1{`RANDOM}};
  io_perf_4_value_REG = _RAND_1539[0:0];
  _RAND_1540 = {1{`RANDOM}};
  io_perf_4_value_REG_1 = _RAND_1540[0:0];
  _RAND_1541 = {1{`RANDOM}};
  io_perf_5_value_REG = _RAND_1541[0:0];
  _RAND_1542 = {1{`RANDOM}};
  io_perf_5_value_REG_1 = _RAND_1542[0:0];
  _RAND_1543 = {1{`RANDOM}};
  io_perf_6_value_REG = _RAND_1543[0:0];
  _RAND_1544 = {1{`RANDOM}};
  io_perf_6_value_REG_1 = _RAND_1544[0:0];
  _RAND_1545 = {1{`RANDOM}};
  io_perf_7_value_REG = _RAND_1545[0:0];
  _RAND_1546 = {1{`RANDOM}};
  io_perf_7_value_REG_1 = _RAND_1546[0:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    valid = 1'h0;
  end
  if (reset) begin
    valid_1 = 1'h0;
  end
  if (reset) begin
    valid_2 = 1'h0;
  end
  if (reset) begin
    stageDelay_valid_1cycle = 1'h0;
  end
  if (reset) begin
    stageCheck_valid_1cycle = 1'h0;
  end
  if (reset) begin
    stageResp_valid_1cycle_dup_0_valid = 1'h0;
  end
  if (reset) begin
    stageResp_valid_1cycle_dup_1_valid = 1'h0;
  end
  if (reset) begin
    l1v = 4'h0;
  end
  if (reset) begin
    l2v = 16'h0;
  end
  if (reset) begin
    l3v = 32'h0;
  end
  if (reset) begin
    spv = 2'h0;
  end
  if (reset) begin
    state_reg = 3'h0;
  end
  if (reset) begin
    state_vec__0 = 3'h0;
  end
  if (reset) begin
    state_vec__1 = 3'h0;
  end
  if (reset) begin
    state_vec__2 = 3'h0;
  end
  if (reset) begin
    state_vec__3 = 3'h0;
  end
  if (reset) begin
    state_vec_1_0 = 7'h0;
  end
  if (reset) begin
    state_vec_1_1 = 7'h0;
  end
  if (reset) begin
    state_vec_1_2 = 7'h0;
  end
  if (reset) begin
    state_vec_1_3 = 7'h0;
  end
  if (reset) begin
    state_reg_3 = 1'h0;
  end
  if (reset) begin
    bypassed_0_valid = 1'h0;
  end
  if (reset) begin
    bypassed_0_valid_1 = 1'h0;
  end
  if (reset) begin
    bypassed_1_valid = 1'h0;
  end
  if (reset) begin
    bypassed_1_valid_1 = 1'h0;
  end
  if (reset) begin
    bypassed_2_valid = 1'h0;
  end
  if (reset) begin
    bypassed_2_valid_1 = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule

