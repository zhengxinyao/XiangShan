module ReservationStation_1(
  input         clock,
  input         reset,
  input         io_redirect_valid,
  input         io_redirect_bits_robIdx_flag,
  input  [4:0]  io_redirect_bits_robIdx_value,
  input         io_redirect_bits_level,
  output        io_fromDispatch_0_ready,
  input         io_fromDispatch_0_valid,
  input  [1:0]  io_fromDispatch_0_bits_ctrl_srcType_0,
  input  [1:0]  io_fromDispatch_0_bits_ctrl_srcType_1,
  input  [3:0]  io_fromDispatch_0_bits_ctrl_fuType,
  input  [6:0]  io_fromDispatch_0_bits_ctrl_fuOpType,
  input         io_fromDispatch_0_bits_ctrl_rfWen,
  input         io_fromDispatch_0_bits_ctrl_fpWen,
  input  [19:0] io_fromDispatch_0_bits_ctrl_imm,
  input         io_fromDispatch_0_bits_srcState_0,
  input         io_fromDispatch_0_bits_srcState_1,
  input  [5:0]  io_fromDispatch_0_bits_psrc_0,
  input  [5:0]  io_fromDispatch_0_bits_psrc_1,
  input  [5:0]  io_fromDispatch_0_bits_pdest,
  input         io_fromDispatch_0_bits_robIdx_flag,
  input  [4:0]  io_fromDispatch_0_bits_robIdx_value,
  output        io_fromDispatch_1_ready,
  input         io_fromDispatch_1_valid,
  input  [1:0]  io_fromDispatch_1_bits_ctrl_srcType_0,
  input  [1:0]  io_fromDispatch_1_bits_ctrl_srcType_1,
  input  [3:0]  io_fromDispatch_1_bits_ctrl_fuType,
  input  [6:0]  io_fromDispatch_1_bits_ctrl_fuOpType,
  input         io_fromDispatch_1_bits_ctrl_rfWen,
  input         io_fromDispatch_1_bits_ctrl_fpWen,
  input  [19:0] io_fromDispatch_1_bits_ctrl_imm,
  input         io_fromDispatch_1_bits_srcState_0,
  input         io_fromDispatch_1_bits_srcState_1,
  input  [5:0]  io_fromDispatch_1_bits_psrc_0,
  input  [5:0]  io_fromDispatch_1_bits_psrc_1,
  input  [5:0]  io_fromDispatch_1_bits_pdest,
  input         io_fromDispatch_1_bits_robIdx_flag,
  input  [4:0]  io_fromDispatch_1_bits_robIdx_value,
  input  [63:0] io_srcRegValue_0_0,
  input  [63:0] io_srcRegValue_0_1,
  input  [63:0] io_srcRegValue_1_0,
  input  [63:0] io_srcRegValue_1_1,
  input         io_deq_0_ready,
  output        io_deq_0_valid,
  output [3:0]  io_deq_0_bits_uop_ctrl_fuType,
  output [6:0]  io_deq_0_bits_uop_ctrl_fuOpType,
  output        io_deq_0_bits_uop_ctrl_rfWen,
  output        io_deq_0_bits_uop_ctrl_fpWen,
  output [5:0]  io_deq_0_bits_uop_pdest,
  output        io_deq_0_bits_uop_robIdx_flag,
  output [4:0]  io_deq_0_bits_uop_robIdx_value,
  output [63:0] io_deq_0_bits_src_0,
  output [63:0] io_deq_0_bits_src_1,
  input         io_fastUopsIn_0_valid,
  input         io_fastUopsIn_0_bits_ctrl_rfWen,
  input  [5:0]  io_fastUopsIn_0_bits_pdest,
  input  [63:0] io_fastDatas_0,
  input         io_slowPorts_0_valid,
  input         io_slowPorts_0_bits_uop_ctrl_rfWen,
  input  [5:0]  io_slowPorts_0_bits_uop_pdest,
  input  [63:0] io_slowPorts_0_bits_data,
  input         io_slowPorts_1_valid,
  input         io_slowPorts_1_bits_uop_ctrl_rfWen,
  input  [5:0]  io_slowPorts_1_bits_uop_pdest,
  input  [63:0] io_slowPorts_1_bits_data,
  input         io_slowPorts_2_valid,
  input         io_slowPorts_2_bits_uop_ctrl_rfWen,
  input  [5:0]  io_slowPorts_2_bits_uop_pdest,
  input  [63:0] io_slowPorts_2_bits_data,
  input         io_slowPorts_3_valid,
  input         io_slowPorts_3_bits_uop_ctrl_rfWen,
  input  [5:0]  io_slowPorts_3_bits_uop_pdest,
  input  [63:0] io_slowPorts_3_bits_data,
  input         io_slowPorts_4_valid,
  input         io_slowPorts_4_bits_uop_ctrl_rfWen,
  input  [5:0]  io_slowPorts_4_bits_uop_pdest,
  input  [63:0] io_slowPorts_4_bits_data,
  output        io_fastWakeup_0_valid,
  output        io_fastWakeup_0_bits_ctrl_rfWen,
  output [5:0]  io_fastWakeup_0_bits_pdest,
  output [5:0]  io_perf_0_value
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [63:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [63:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [63:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [63:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [63:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
`endif // RANDOMIZE_REG_INIT
  wire  statusArray_clock; // @[ReservationStation.scala 261:27]
  wire  statusArray_reset; // @[ReservationStation.scala 261:27]
  wire  statusArray_io_redirect_valid; // @[ReservationStation.scala 261:27]
  wire  statusArray_io_redirect_bits_robIdx_flag; // @[ReservationStation.scala 261:27]
  wire [4:0] statusArray_io_redirect_bits_robIdx_value; // @[ReservationStation.scala 261:27]
  wire  statusArray_io_redirect_bits_level; // @[ReservationStation.scala 261:27]
  wire [7:0] statusArray_io_isValid; // @[ReservationStation.scala 261:27]
  wire [7:0] statusArray_io_isValidNext; // @[ReservationStation.scala 261:27]
  wire [7:0] statusArray_io_canIssue; // @[ReservationStation.scala 261:27]
  wire [7:0] statusArray_io_flushed; // @[ReservationStation.scala 261:27]
  wire  statusArray_io_update_0_enable; // @[ReservationStation.scala 261:27]
  wire [7:0] statusArray_io_update_0_addr; // @[ReservationStation.scala 261:27]
  wire  statusArray_io_update_0_data_srcState_0; // @[ReservationStation.scala 261:27]
  wire  statusArray_io_update_0_data_srcState_1; // @[ReservationStation.scala 261:27]
  wire [5:0] statusArray_io_update_0_data_psrc_0; // @[ReservationStation.scala 261:27]
  wire [5:0] statusArray_io_update_0_data_psrc_1; // @[ReservationStation.scala 261:27]
  wire [1:0] statusArray_io_update_0_data_srcType_0; // @[ReservationStation.scala 261:27]
  wire [1:0] statusArray_io_update_0_data_srcType_1; // @[ReservationStation.scala 261:27]
  wire  statusArray_io_update_0_data_robIdx_flag; // @[ReservationStation.scala 261:27]
  wire [4:0] statusArray_io_update_0_data_robIdx_value; // @[ReservationStation.scala 261:27]
  wire  statusArray_io_update_1_enable; // @[ReservationStation.scala 261:27]
  wire [7:0] statusArray_io_update_1_addr; // @[ReservationStation.scala 261:27]
  wire  statusArray_io_update_1_data_srcState_0; // @[ReservationStation.scala 261:27]
  wire  statusArray_io_update_1_data_srcState_1; // @[ReservationStation.scala 261:27]
  wire [5:0] statusArray_io_update_1_data_psrc_0; // @[ReservationStation.scala 261:27]
  wire [5:0] statusArray_io_update_1_data_psrc_1; // @[ReservationStation.scala 261:27]
  wire [1:0] statusArray_io_update_1_data_srcType_0; // @[ReservationStation.scala 261:27]
  wire [1:0] statusArray_io_update_1_data_srcType_1; // @[ReservationStation.scala 261:27]
  wire  statusArray_io_update_1_data_robIdx_flag; // @[ReservationStation.scala 261:27]
  wire [4:0] statusArray_io_update_1_data_robIdx_value; // @[ReservationStation.scala 261:27]
  wire  statusArray_io_wakeup_0_valid; // @[ReservationStation.scala 261:27]
  wire  statusArray_io_wakeup_0_bits_ctrl_rfWen; // @[ReservationStation.scala 261:27]
  wire [5:0] statusArray_io_wakeup_0_bits_pdest; // @[ReservationStation.scala 261:27]
  wire  statusArray_io_wakeup_1_valid; // @[ReservationStation.scala 261:27]
  wire  statusArray_io_wakeup_1_bits_ctrl_rfWen; // @[ReservationStation.scala 261:27]
  wire [5:0] statusArray_io_wakeup_1_bits_pdest; // @[ReservationStation.scala 261:27]
  wire  statusArray_io_wakeup_2_valid; // @[ReservationStation.scala 261:27]
  wire  statusArray_io_wakeup_2_bits_ctrl_rfWen; // @[ReservationStation.scala 261:27]
  wire [5:0] statusArray_io_wakeup_2_bits_pdest; // @[ReservationStation.scala 261:27]
  wire  statusArray_io_wakeup_3_valid; // @[ReservationStation.scala 261:27]
  wire  statusArray_io_wakeup_3_bits_ctrl_rfWen; // @[ReservationStation.scala 261:27]
  wire [5:0] statusArray_io_wakeup_3_bits_pdest; // @[ReservationStation.scala 261:27]
  wire  statusArray_io_wakeup_4_valid; // @[ReservationStation.scala 261:27]
  wire  statusArray_io_wakeup_4_bits_ctrl_rfWen; // @[ReservationStation.scala 261:27]
  wire [5:0] statusArray_io_wakeup_4_bits_pdest; // @[ReservationStation.scala 261:27]
  wire  statusArray_io_wakeup_5_valid; // @[ReservationStation.scala 261:27]
  wire  statusArray_io_wakeup_5_bits_ctrl_rfWen; // @[ReservationStation.scala 261:27]
  wire [5:0] statusArray_io_wakeup_5_bits_pdest; // @[ReservationStation.scala 261:27]
  wire [5:0] statusArray_io_wakeupMatch_0_0; // @[ReservationStation.scala 261:27]
  wire [5:0] statusArray_io_wakeupMatch_0_1; // @[ReservationStation.scala 261:27]
  wire [5:0] statusArray_io_wakeupMatch_1_0; // @[ReservationStation.scala 261:27]
  wire [5:0] statusArray_io_wakeupMatch_1_1; // @[ReservationStation.scala 261:27]
  wire [5:0] statusArray_io_wakeupMatch_2_0; // @[ReservationStation.scala 261:27]
  wire [5:0] statusArray_io_wakeupMatch_2_1; // @[ReservationStation.scala 261:27]
  wire [5:0] statusArray_io_wakeupMatch_3_0; // @[ReservationStation.scala 261:27]
  wire [5:0] statusArray_io_wakeupMatch_3_1; // @[ReservationStation.scala 261:27]
  wire [5:0] statusArray_io_wakeupMatch_4_0; // @[ReservationStation.scala 261:27]
  wire [5:0] statusArray_io_wakeupMatch_4_1; // @[ReservationStation.scala 261:27]
  wire [5:0] statusArray_io_wakeupMatch_5_0; // @[ReservationStation.scala 261:27]
  wire [5:0] statusArray_io_wakeupMatch_5_1; // @[ReservationStation.scala 261:27]
  wire [5:0] statusArray_io_wakeupMatch_6_0; // @[ReservationStation.scala 261:27]
  wire [5:0] statusArray_io_wakeupMatch_6_1; // @[ReservationStation.scala 261:27]
  wire [5:0] statusArray_io_wakeupMatch_7_0; // @[ReservationStation.scala 261:27]
  wire [5:0] statusArray_io_wakeupMatch_7_1; // @[ReservationStation.scala 261:27]
  wire  statusArray_io_deqResp_0_valid; // @[ReservationStation.scala 261:27]
  wire [7:0] statusArray_io_deqResp_0_bits_rsMask; // @[ReservationStation.scala 261:27]
  wire  statusArray_io_deqResp_0_bits_success; // @[ReservationStation.scala 261:27]
  wire  statusArray_io_deqResp_1_valid; // @[ReservationStation.scala 261:27]
  wire [7:0] statusArray_io_deqResp_1_bits_rsMask; // @[ReservationStation.scala 261:27]
  wire  statusArray_io_deqResp_1_bits_success; // @[ReservationStation.scala 261:27]
  wire  statusArray_io_deqResp_2_valid; // @[ReservationStation.scala 261:27]
  wire [7:0] statusArray_io_deqResp_2_bits_rsMask; // @[ReservationStation.scala 261:27]
  wire  statusArray_io_deqResp_2_bits_success; // @[ReservationStation.scala 261:27]
  wire [7:0] select_io_validVec; // @[ReservationStation.scala 262:22]
  wire [7:0] select_io_allocate_0_bits; // @[ReservationStation.scala 262:22]
  wire [7:0] select_io_allocate_1_bits; // @[ReservationStation.scala 262:22]
  wire [7:0] select_io_request; // @[ReservationStation.scala 262:22]
  wire  select_io_grant_0_valid; // @[ReservationStation.scala 262:22]
  wire [7:0] select_io_grant_0_bits; // @[ReservationStation.scala 262:22]
  wire  dataArray_clock; // @[ReservationStation.scala 263:25]
  wire [7:0] dataArray_io_read_0_addr; // @[ReservationStation.scala 263:25]
  wire [63:0] dataArray_io_read_0_data_0; // @[ReservationStation.scala 263:25]
  wire [63:0] dataArray_io_read_0_data_1; // @[ReservationStation.scala 263:25]
  wire [7:0] dataArray_io_read_1_addr; // @[ReservationStation.scala 263:25]
  wire [63:0] dataArray_io_read_1_data_0; // @[ReservationStation.scala 263:25]
  wire [63:0] dataArray_io_read_1_data_1; // @[ReservationStation.scala 263:25]
  wire  dataArray_io_write_0_enable; // @[ReservationStation.scala 263:25]
  wire  dataArray_io_write_0_mask_0; // @[ReservationStation.scala 263:25]
  wire  dataArray_io_write_0_mask_1; // @[ReservationStation.scala 263:25]
  wire [7:0] dataArray_io_write_0_addr; // @[ReservationStation.scala 263:25]
  wire [63:0] dataArray_io_write_0_data_0; // @[ReservationStation.scala 263:25]
  wire [63:0] dataArray_io_write_0_data_1; // @[ReservationStation.scala 263:25]
  wire  dataArray_io_write_1_enable; // @[ReservationStation.scala 263:25]
  wire  dataArray_io_write_1_mask_0; // @[ReservationStation.scala 263:25]
  wire  dataArray_io_write_1_mask_1; // @[ReservationStation.scala 263:25]
  wire [7:0] dataArray_io_write_1_addr; // @[ReservationStation.scala 263:25]
  wire [63:0] dataArray_io_write_1_data_0; // @[ReservationStation.scala 263:25]
  wire [63:0] dataArray_io_write_1_data_1; // @[ReservationStation.scala 263:25]
  wire  dataArray_io_multiWrite_0_enable; // @[ReservationStation.scala 263:25]
  wire [7:0] dataArray_io_multiWrite_0_addr_0; // @[ReservationStation.scala 263:25]
  wire [7:0] dataArray_io_multiWrite_0_addr_1; // @[ReservationStation.scala 263:25]
  wire [63:0] dataArray_io_multiWrite_0_data; // @[ReservationStation.scala 263:25]
  wire  dataArray_io_multiWrite_1_enable; // @[ReservationStation.scala 263:25]
  wire [7:0] dataArray_io_multiWrite_1_addr_0; // @[ReservationStation.scala 263:25]
  wire [7:0] dataArray_io_multiWrite_1_addr_1; // @[ReservationStation.scala 263:25]
  wire [63:0] dataArray_io_multiWrite_1_data; // @[ReservationStation.scala 263:25]
  wire  dataArray_io_multiWrite_2_enable; // @[ReservationStation.scala 263:25]
  wire [7:0] dataArray_io_multiWrite_2_addr_0; // @[ReservationStation.scala 263:25]
  wire [7:0] dataArray_io_multiWrite_2_addr_1; // @[ReservationStation.scala 263:25]
  wire [63:0] dataArray_io_multiWrite_2_data; // @[ReservationStation.scala 263:25]
  wire  dataArray_io_multiWrite_3_enable; // @[ReservationStation.scala 263:25]
  wire [7:0] dataArray_io_multiWrite_3_addr_0; // @[ReservationStation.scala 263:25]
  wire [7:0] dataArray_io_multiWrite_3_addr_1; // @[ReservationStation.scala 263:25]
  wire [63:0] dataArray_io_multiWrite_3_data; // @[ReservationStation.scala 263:25]
  wire  dataArray_io_multiWrite_4_enable; // @[ReservationStation.scala 263:25]
  wire [7:0] dataArray_io_multiWrite_4_addr_0; // @[ReservationStation.scala 263:25]
  wire [7:0] dataArray_io_multiWrite_4_addr_1; // @[ReservationStation.scala 263:25]
  wire [63:0] dataArray_io_multiWrite_4_data; // @[ReservationStation.scala 263:25]
  wire  payloadArray_clock; // @[ReservationStation.scala 264:28]
  wire [7:0] payloadArray_io_read_0_addr; // @[ReservationStation.scala 264:28]
  wire [3:0] payloadArray_io_read_0_data_ctrl_fuType; // @[ReservationStation.scala 264:28]
  wire [6:0] payloadArray_io_read_0_data_ctrl_fuOpType; // @[ReservationStation.scala 264:28]
  wire  payloadArray_io_read_0_data_ctrl_rfWen; // @[ReservationStation.scala 264:28]
  wire  payloadArray_io_read_0_data_ctrl_fpWen; // @[ReservationStation.scala 264:28]
  wire [5:0] payloadArray_io_read_0_data_pdest; // @[ReservationStation.scala 264:28]
  wire  payloadArray_io_read_0_data_robIdx_flag; // @[ReservationStation.scala 264:28]
  wire [4:0] payloadArray_io_read_0_data_robIdx_value; // @[ReservationStation.scala 264:28]
  wire [7:0] payloadArray_io_read_1_addr; // @[ReservationStation.scala 264:28]
  wire [3:0] payloadArray_io_read_1_data_ctrl_fuType; // @[ReservationStation.scala 264:28]
  wire [6:0] payloadArray_io_read_1_data_ctrl_fuOpType; // @[ReservationStation.scala 264:28]
  wire  payloadArray_io_read_1_data_ctrl_rfWen; // @[ReservationStation.scala 264:28]
  wire  payloadArray_io_read_1_data_ctrl_fpWen; // @[ReservationStation.scala 264:28]
  wire [5:0] payloadArray_io_read_1_data_pdest; // @[ReservationStation.scala 264:28]
  wire  payloadArray_io_read_1_data_robIdx_flag; // @[ReservationStation.scala 264:28]
  wire [4:0] payloadArray_io_read_1_data_robIdx_value; // @[ReservationStation.scala 264:28]
  wire  payloadArray_io_write_0_enable; // @[ReservationStation.scala 264:28]
  wire [7:0] payloadArray_io_write_0_addr; // @[ReservationStation.scala 264:28]
  wire [3:0] payloadArray_io_write_0_data_ctrl_fuType; // @[ReservationStation.scala 264:28]
  wire [6:0] payloadArray_io_write_0_data_ctrl_fuOpType; // @[ReservationStation.scala 264:28]
  wire  payloadArray_io_write_0_data_ctrl_rfWen; // @[ReservationStation.scala 264:28]
  wire  payloadArray_io_write_0_data_ctrl_fpWen; // @[ReservationStation.scala 264:28]
  wire [5:0] payloadArray_io_write_0_data_pdest; // @[ReservationStation.scala 264:28]
  wire  payloadArray_io_write_0_data_robIdx_flag; // @[ReservationStation.scala 264:28]
  wire [4:0] payloadArray_io_write_0_data_robIdx_value; // @[ReservationStation.scala 264:28]
  wire  payloadArray_io_write_1_enable; // @[ReservationStation.scala 264:28]
  wire [7:0] payloadArray_io_write_1_addr; // @[ReservationStation.scala 264:28]
  wire [3:0] payloadArray_io_write_1_data_ctrl_fuType; // @[ReservationStation.scala 264:28]
  wire [6:0] payloadArray_io_write_1_data_ctrl_fuOpType; // @[ReservationStation.scala 264:28]
  wire  payloadArray_io_write_1_data_ctrl_rfWen; // @[ReservationStation.scala 264:28]
  wire  payloadArray_io_write_1_data_ctrl_fpWen; // @[ReservationStation.scala 264:28]
  wire [5:0] payloadArray_io_write_1_data_pdest; // @[ReservationStation.scala 264:28]
  wire  payloadArray_io_write_1_data_robIdx_flag; // @[ReservationStation.scala 264:28]
  wire [4:0] payloadArray_io_write_1_data_robIdx_value; // @[ReservationStation.scala 264:28]
  wire  s1_oldestSel_age_clock; // @[SelectPolicy.scala 174:21]
  wire  s1_oldestSel_age_reset; // @[SelectPolicy.scala 174:21]
  wire [7:0] s1_oldestSel_age_io_enq_0; // @[SelectPolicy.scala 174:21]
  wire [7:0] s1_oldestSel_age_io_enq_1; // @[SelectPolicy.scala 174:21]
  wire [7:0] s1_oldestSel_age_io_deq; // @[SelectPolicy.scala 174:21]
  wire [7:0] s1_oldestSel_age_io_out; // @[SelectPolicy.scala 174:21]
  wire  oldestSelection_io_oldest_valid; // @[ReservationStation.scala 499:33]
  wire  oldestSelection_io_isOverrided_0; // @[ReservationStation.scala 499:33]
  wire  wakeupQueue_clock; // @[ReservationStation.scala 564:31]
  wire  wakeupQueue_reset; // @[ReservationStation.scala 564:31]
  wire  wakeupQueue_io_in_valid; // @[ReservationStation.scala 564:31]
  wire  wakeupQueue_io_in_bits_ctrl_rfWen; // @[ReservationStation.scala 564:31]
  wire [5:0] wakeupQueue_io_in_bits_pdest; // @[ReservationStation.scala 564:31]
  wire  wakeupQueue_io_in_bits_robIdx_flag; // @[ReservationStation.scala 564:31]
  wire [4:0] wakeupQueue_io_in_bits_robIdx_value; // @[ReservationStation.scala 564:31]
  wire  wakeupQueue_io_out_valid; // @[ReservationStation.scala 564:31]
  wire  wakeupQueue_io_out_bits_ctrl_rfWen; // @[ReservationStation.scala 564:31]
  wire [5:0] wakeupQueue_io_out_bits_pdest; // @[ReservationStation.scala 564:31]
  wire  wakeupQueue_io_redirect_valid; // @[ReservationStation.scala 564:31]
  wire  wakeupQueue_io_redirect_bits_robIdx_flag; // @[ReservationStation.scala 564:31]
  wire [4:0] wakeupQueue_io_redirect_bits_robIdx_value; // @[ReservationStation.scala 564:31]
  wire  wakeupQueue_io_redirect_bits_level; // @[ReservationStation.scala 564:31]
  wire [1:0] immExt_io_uop_ctrl_srcType_1; // @[DataArray.scala 159:36]
  wire [19:0] immExt_io_uop_ctrl_imm; // @[DataArray.scala 159:36]
  wire [63:0] immExt_io_data_in_0; // @[DataArray.scala 159:36]
  wire [63:0] immExt_io_data_in_1; // @[DataArray.scala 159:36]
  wire [63:0] immExt_io_data_out_0; // @[DataArray.scala 159:36]
  wire [63:0] immExt_io_data_out_1; // @[DataArray.scala 159:36]
  wire [1:0] immExt_1_io_uop_ctrl_srcType_1; // @[DataArray.scala 159:36]
  wire [19:0] immExt_1_io_uop_ctrl_imm; // @[DataArray.scala 159:36]
  wire [63:0] immExt_1_io_data_in_0; // @[DataArray.scala 159:36]
  wire [63:0] immExt_1_io_data_in_1; // @[DataArray.scala 159:36]
  wire [63:0] immExt_1_io_data_out_0; // @[DataArray.scala 159:36]
  wire [63:0] immExt_1_io_data_out_1; // @[DataArray.scala 159:36]
  wire  dataSelect_io_doOverride_0; // @[ReservationStation.scala 691:26]
  wire [63:0] dataSelect_io_readData_0_0; // @[ReservationStation.scala 691:26]
  wire [63:0] dataSelect_io_readData_0_1; // @[ReservationStation.scala 691:26]
  wire [63:0] dataSelect_io_readData_1_0; // @[ReservationStation.scala 691:26]
  wire [63:0] dataSelect_io_readData_1_1; // @[ReservationStation.scala 691:26]
  wire [4:0] dataSelect_io_fromSlowPorts_0_0; // @[ReservationStation.scala 691:26]
  wire [4:0] dataSelect_io_fromSlowPorts_0_1; // @[ReservationStation.scala 691:26]
  wire [4:0] dataSelect_io_fromSlowPorts_1_0; // @[ReservationStation.scala 691:26]
  wire [4:0] dataSelect_io_fromSlowPorts_1_1; // @[ReservationStation.scala 691:26]
  wire [4:0] dataSelect_io_fromSlowPorts_2_0; // @[ReservationStation.scala 691:26]
  wire [4:0] dataSelect_io_fromSlowPorts_2_1; // @[ReservationStation.scala 691:26]
  wire [63:0] dataSelect_io_slowData_0; // @[ReservationStation.scala 691:26]
  wire [63:0] dataSelect_io_slowData_1; // @[ReservationStation.scala 691:26]
  wire [63:0] dataSelect_io_slowData_2; // @[ReservationStation.scala 691:26]
  wire [63:0] dataSelect_io_slowData_3; // @[ReservationStation.scala 691:26]
  wire [63:0] dataSelect_io_slowData_4; // @[ReservationStation.scala 691:26]
  wire  dataSelect_io_enqBypass_0_0; // @[ReservationStation.scala 691:26]
  wire [63:0] dataSelect_io_enqData_0_0_bits; // @[ReservationStation.scala 691:26]
  wire [63:0] dataSelect_io_enqData_0_1_bits; // @[ReservationStation.scala 691:26]
  wire [63:0] dataSelect_io_deqData_0_0; // @[ReservationStation.scala 691:26]
  wire [63:0] dataSelect_io_deqData_0_1; // @[ReservationStation.scala 691:26]
  wire  bypassNetwork_clock; // @[BypassNetwork.scala 111:13]
  wire  bypassNetwork_io_hold; // @[BypassNetwork.scala 111:13]
  wire [63:0] bypassNetwork_io_source_0; // @[BypassNetwork.scala 111:13]
  wire [63:0] bypassNetwork_io_source_1; // @[BypassNetwork.scala 111:13]
  wire [63:0] bypassNetwork_io_target_0; // @[BypassNetwork.scala 111:13]
  wire [63:0] bypassNetwork_io_target_1; // @[BypassNetwork.scala 111:13]
  wire  bypassNetwork_io_bypass_0_valid_0; // @[BypassNetwork.scala 111:13]
  wire  bypassNetwork_io_bypass_0_valid_1; // @[BypassNetwork.scala 111:13]
  wire [63:0] bypassNetwork_io_bypass_0_data; // @[BypassNetwork.scala 111:13]
  wire [7:0] s0_allocatePtrOH_0 = select_io_allocate_0_bits; // @[ReservationStation.scala 273:{33,33}]
  wire [7:0] s0_allocatePtrOH_1 = select_io_allocate_1_bits; // @[ReservationStation.scala 273:{33,33}]
  reg [7:0] validAfterAllocate; // @[ReservationStation.scala 282:35]
  wire  _s0_doEnqueue_0_T = io_fromDispatch_0_ready & io_fromDispatch_0_valid; // @[Decoupled.scala 50:35]
  wire  _s0_doEnqueue_0_T_1 = ~io_redirect_valid; // @[ReservationStation.scala 336:51]
  wire  s0_doEnqueue_0 = _s0_doEnqueue_0_T & ~io_redirect_valid; // @[ReservationStation.scala 336:48]
  wire [7:0] validUpdateByAllocate_xs_0 = s0_doEnqueue_0 ? s0_allocatePtrOH_0 : 8'h0; // @[ParallelMux.scala 64:44]
  wire  _s0_doEnqueue_1_T = io_fromDispatch_1_ready & io_fromDispatch_1_valid; // @[Decoupled.scala 50:35]
  wire  s0_doEnqueue_1 = _s0_doEnqueue_1_T & ~io_redirect_valid; // @[ReservationStation.scala 336:48]
  wire [7:0] validUpdateByAllocate_xs_1 = s0_doEnqueue_1 ? s0_allocatePtrOH_1 : 8'h0; // @[ParallelMux.scala 64:44]
  wire [7:0] validUpdateByAllocate = validUpdateByAllocate_xs_0 | validUpdateByAllocate_xs_1; // @[ParallelMux.scala 36:53]
  wire  _numEmptyEntries_T_8 = ~statusArray_io_isValid[0]; // @[ReservationStation.scala 311:76]
  wire  _numEmptyEntries_T_9 = ~statusArray_io_isValid[1]; // @[ReservationStation.scala 311:76]
  wire  _numEmptyEntries_T_10 = ~statusArray_io_isValid[2]; // @[ReservationStation.scala 311:76]
  wire  _numEmptyEntries_T_11 = ~statusArray_io_isValid[3]; // @[ReservationStation.scala 311:76]
  wire  _numEmptyEntries_T_12 = ~statusArray_io_isValid[4]; // @[ReservationStation.scala 311:76]
  wire  _numEmptyEntries_T_13 = ~statusArray_io_isValid[5]; // @[ReservationStation.scala 311:76]
  wire  _numEmptyEntries_T_14 = ~statusArray_io_isValid[6]; // @[ReservationStation.scala 311:76]
  wire  _numEmptyEntries_T_15 = ~statusArray_io_isValid[7]; // @[ReservationStation.scala 311:76]
  wire [1:0] _numEmptyEntries_T_16 = _numEmptyEntries_T_8 + _numEmptyEntries_T_9; // @[Bitwise.scala 48:55]
  wire [1:0] _numEmptyEntries_T_18 = _numEmptyEntries_T_10 + _numEmptyEntries_T_11; // @[Bitwise.scala 48:55]
  wire [2:0] _numEmptyEntries_T_20 = _numEmptyEntries_T_16 + _numEmptyEntries_T_18; // @[Bitwise.scala 48:55]
  wire [1:0] _numEmptyEntries_T_22 = _numEmptyEntries_T_12 + _numEmptyEntries_T_13; // @[Bitwise.scala 48:55]
  wire [1:0] _numEmptyEntries_T_24 = _numEmptyEntries_T_14 + _numEmptyEntries_T_15; // @[Bitwise.scala 48:55]
  wire [2:0] _numEmptyEntries_T_26 = _numEmptyEntries_T_22 + _numEmptyEntries_T_24; // @[Bitwise.scala 48:55]
  wire [3:0] numEmptyEntries = _numEmptyEntries_T_20 + _numEmptyEntries_T_26; // @[Bitwise.scala 48:55]
  wire [1:0] numAllocateS1 = statusArray_io_update_0_enable + statusArray_io_update_1_enable; // @[Bitwise.scala 48:55]
  wire [3:0] _GEN_771 = {{2'd0}, numAllocateS1}; // @[ReservationStation.scala 313:47]
  wire [3:0] realNumEmptyAfterS1 = numEmptyEntries - _GEN_771; // @[ReservationStation.scala 313:47]
  wire [1:0] highBits = realNumEmptyAfterS1[3:2]; // @[ReservationStation.scala 315:41]
  wire [2:0] numEmptyAfterS1 = |highBits ? 3'h4 : {{1'd0}, realNumEmptyAfterS1[1:0]}; // @[ReservationStation.scala 316:27]
  wire  _numDeq_T = statusArray_io_deqResp_0_valid & statusArray_io_deqResp_0_bits_success; // @[ReservationStation.scala 317:81]
  wire  _numDeq_T_1 = statusArray_io_deqResp_1_valid & statusArray_io_deqResp_1_bits_success; // @[ReservationStation.scala 317:81]
  wire  _numDeq_T_2 = statusArray_io_deqResp_2_valid & statusArray_io_deqResp_2_bits_success; // @[ReservationStation.scala 317:81]
  wire [1:0] _numDeq_T_3 = _numDeq_T_1 + _numDeq_T_2; // @[Bitwise.scala 48:55]
  wire [1:0] _GEN_772 = {{1'd0}, _numDeq_T}; // @[Bitwise.scala 48:55]
  wire [2:0] _numDeq_T_5 = _GEN_772 + _numDeq_T_3; // @[Bitwise.scala 48:55]
  wire [1:0] numDeq = _numDeq_T_5[1:0]; // @[Bitwise.scala 48:55]
  reg [2:0] emptyThisCycle; // @[ReservationStation.scala 318:29]
  wire [2:0] _GEN_773 = {{1'd0}, numDeq}; // @[ReservationStation.scala 319:39]
  wire [1:0] numAllocateS0 = s0_doEnqueue_0 + s0_doEnqueue_1; // @[Bitwise.scala 48:55]
  reg [1:0] allocateThisCycle; // @[ReservationStation.scala 322:34]
  wire [2:0] _allocateThisCycle_T = {{1'd0}, numAllocateS0}; // @[ReservationStation.scala 323:42]
  wire [2:0] _GEN_774 = {{1'd0}, allocateThisCycle}; // @[ReservationStation.scala 324:42]
  reg [1:0] allocateThisCycle_1; // @[ReservationStation.scala 322:34]
  wire [2:0] _allocateThisCycle_T_1 = numAllocateS0 + 2'h1; // @[ReservationStation.scala 323:42]
  wire [2:0] _GEN_775 = {{1'd0}, allocateThisCycle_1}; // @[ReservationStation.scala 324:42]
  wire  pdestMatch = io_slowPorts_0_bits_uop_pdest == io_fromDispatch_0_bits_psrc_0; // @[Bundle.scala 262:30]
  wire  stateCond = pdestMatch & io_slowPorts_0_bits_uop_ctrl_rfWen; // @[Bundle.scala 268:34]
  wire  rfDataMatch = io_slowPorts_0_bits_uop_ctrl_rfWen & io_fromDispatch_0_bits_psrc_0 != 6'h0; // @[Bundle.scala 270:58]
  wire  _dataCond_T = io_fromDispatch_0_bits_ctrl_srcType_0 == 2'h0; // @[package.scala 37:39]
  wire  dataCond = pdestMatch & (rfDataMatch & _dataCond_T); // @[Bundle.scala 271:33]
  wire  pdestMatch_1 = io_slowPorts_0_bits_uop_pdest == io_fromDispatch_0_bits_psrc_1; // @[Bundle.scala 262:30]
  wire  stateCond_1 = pdestMatch_1 & io_slowPorts_0_bits_uop_ctrl_rfWen; // @[Bundle.scala 268:34]
  wire  rfDataMatch_1 = io_slowPorts_0_bits_uop_ctrl_rfWen & io_fromDispatch_0_bits_psrc_1 != 6'h0; // @[Bundle.scala 270:58]
  wire  _dataCond_T_5 = io_fromDispatch_0_bits_ctrl_srcType_1 == 2'h0; // @[package.scala 37:39]
  wire  dataCond_1 = pdestMatch_1 & (rfDataMatch_1 & _dataCond_T_5); // @[Bundle.scala 271:33]
  wire  pdestMatch_3 = io_slowPorts_1_bits_uop_pdest == io_fromDispatch_0_bits_psrc_0; // @[Bundle.scala 262:30]
  wire  stateCond_3 = pdestMatch_3 & io_slowPorts_1_bits_uop_ctrl_rfWen; // @[Bundle.scala 268:34]
  wire  rfDataMatch_3 = io_slowPorts_1_bits_uop_ctrl_rfWen & io_fromDispatch_0_bits_psrc_0 != 6'h0; // @[Bundle.scala 270:58]
  wire  dataCond_3 = pdestMatch_3 & (rfDataMatch_3 & _dataCond_T); // @[Bundle.scala 271:33]
  wire  pdestMatch_4 = io_slowPorts_1_bits_uop_pdest == io_fromDispatch_0_bits_psrc_1; // @[Bundle.scala 262:30]
  wire  stateCond_4 = pdestMatch_4 & io_slowPorts_1_bits_uop_ctrl_rfWen; // @[Bundle.scala 268:34]
  wire  rfDataMatch_4 = io_slowPorts_1_bits_uop_ctrl_rfWen & io_fromDispatch_0_bits_psrc_1 != 6'h0; // @[Bundle.scala 270:58]
  wire  dataCond_4 = pdestMatch_4 & (rfDataMatch_4 & _dataCond_T_5); // @[Bundle.scala 271:33]
  wire  pdestMatch_6 = io_slowPorts_2_bits_uop_pdest == io_fromDispatch_0_bits_psrc_0; // @[Bundle.scala 262:30]
  wire  stateCond_6 = pdestMatch_6 & io_slowPorts_2_bits_uop_ctrl_rfWen; // @[Bundle.scala 268:34]
  wire  rfDataMatch_6 = io_slowPorts_2_bits_uop_ctrl_rfWen & io_fromDispatch_0_bits_psrc_0 != 6'h0; // @[Bundle.scala 270:58]
  wire  dataCond_6 = pdestMatch_6 & (rfDataMatch_6 & _dataCond_T); // @[Bundle.scala 271:33]
  wire  pdestMatch_7 = io_slowPorts_2_bits_uop_pdest == io_fromDispatch_0_bits_psrc_1; // @[Bundle.scala 262:30]
  wire  stateCond_7 = pdestMatch_7 & io_slowPorts_2_bits_uop_ctrl_rfWen; // @[Bundle.scala 268:34]
  wire  rfDataMatch_7 = io_slowPorts_2_bits_uop_ctrl_rfWen & io_fromDispatch_0_bits_psrc_1 != 6'h0; // @[Bundle.scala 270:58]
  wire  dataCond_7 = pdestMatch_7 & (rfDataMatch_7 & _dataCond_T_5); // @[Bundle.scala 271:33]
  wire  pdestMatch_9 = io_slowPorts_3_bits_uop_pdest == io_fromDispatch_0_bits_psrc_0; // @[Bundle.scala 262:30]
  wire  stateCond_9 = pdestMatch_9 & io_slowPorts_3_bits_uop_ctrl_rfWen; // @[Bundle.scala 268:34]
  wire  rfDataMatch_9 = io_slowPorts_3_bits_uop_ctrl_rfWen & io_fromDispatch_0_bits_psrc_0 != 6'h0; // @[Bundle.scala 270:58]
  wire  dataCond_9 = pdestMatch_9 & (rfDataMatch_9 & _dataCond_T); // @[Bundle.scala 271:33]
  wire  pdestMatch_10 = io_slowPorts_3_bits_uop_pdest == io_fromDispatch_0_bits_psrc_1; // @[Bundle.scala 262:30]
  wire  stateCond_10 = pdestMatch_10 & io_slowPorts_3_bits_uop_ctrl_rfWen; // @[Bundle.scala 268:34]
  wire  rfDataMatch_10 = io_slowPorts_3_bits_uop_ctrl_rfWen & io_fromDispatch_0_bits_psrc_1 != 6'h0; // @[Bundle.scala 270:58]
  wire  dataCond_10 = pdestMatch_10 & (rfDataMatch_10 & _dataCond_T_5); // @[Bundle.scala 271:33]
  wire  pdestMatch_12 = io_slowPorts_4_bits_uop_pdest == io_fromDispatch_0_bits_psrc_0; // @[Bundle.scala 262:30]
  wire  stateCond_12 = pdestMatch_12 & io_slowPorts_4_bits_uop_ctrl_rfWen; // @[Bundle.scala 268:34]
  wire  rfDataMatch_12 = io_slowPorts_4_bits_uop_ctrl_rfWen & io_fromDispatch_0_bits_psrc_0 != 6'h0; // @[Bundle.scala 270:58]
  wire  dataCond_12 = pdestMatch_12 & (rfDataMatch_12 & _dataCond_T); // @[Bundle.scala 271:33]
  wire  pdestMatch_13 = io_slowPorts_4_bits_uop_pdest == io_fromDispatch_0_bits_psrc_1; // @[Bundle.scala 262:30]
  wire  stateCond_13 = pdestMatch_13 & io_slowPorts_4_bits_uop_ctrl_rfWen; // @[Bundle.scala 268:34]
  wire  rfDataMatch_13 = io_slowPorts_4_bits_uop_ctrl_rfWen & io_fromDispatch_0_bits_psrc_1 != 6'h0; // @[Bundle.scala 270:58]
  wire  dataCond_13 = pdestMatch_13 & (rfDataMatch_13 & _dataCond_T_5); // @[Bundle.scala 271:33]
  wire  pdestMatch_15 = io_fastUopsIn_0_bits_pdest == io_fromDispatch_0_bits_psrc_0; // @[Bundle.scala 262:30]
  wire  rfDataMatch_15 = io_fastUopsIn_0_bits_ctrl_rfWen & io_fromDispatch_0_bits_psrc_0 != 6'h0; // @[Bundle.scala 270:58]
  wire  dataCond_15 = pdestMatch_15 & (rfDataMatch_15 & _dataCond_T); // @[Bundle.scala 271:33]
  wire  pdestMatch_16 = io_fastUopsIn_0_bits_pdest == io_fromDispatch_0_bits_psrc_1; // @[Bundle.scala 262:30]
  wire  rfDataMatch_16 = io_fastUopsIn_0_bits_ctrl_rfWen & io_fromDispatch_0_bits_psrc_1 != 6'h0; // @[Bundle.scala 270:58]
  wire  dataCond_16 = pdestMatch_16 & (rfDataMatch_16 & _dataCond_T_5); // @[Bundle.scala 271:33]
  wire  _s0_enqWakeup_0_0_T = io_slowPorts_0_valid & stateCond; // @[ReservationStation.scala 341:90]
  wire  _s0_enqWakeup_0_0_T_1 = io_slowPorts_1_valid & stateCond_3; // @[ReservationStation.scala 341:90]
  wire  _s0_enqWakeup_0_0_T_2 = io_slowPorts_2_valid & stateCond_6; // @[ReservationStation.scala 341:90]
  wire  _s0_enqWakeup_0_0_T_3 = io_slowPorts_3_valid & stateCond_9; // @[ReservationStation.scala 341:90]
  wire  _s0_enqWakeup_0_0_T_4 = io_slowPorts_4_valid & stateCond_12; // @[ReservationStation.scala 341:90]
  wire [1:0] s0_enqWakeup_0_0_lo = {_s0_enqWakeup_0_0_T_1,_s0_enqWakeup_0_0_T}; // @[ReservationStation.scala 341:100]
  wire [2:0] s0_enqWakeup_0_0_hi = {_s0_enqWakeup_0_0_T_4,_s0_enqWakeup_0_0_T_3,_s0_enqWakeup_0_0_T_2}; // @[ReservationStation.scala 341:100]
  wire  _s0_enqDataCapture_0_0_T = io_slowPorts_0_valid & dataCond; // @[ReservationStation.scala 342:94]
  wire  _s0_enqDataCapture_0_0_T_1 = io_slowPorts_1_valid & dataCond_3; // @[ReservationStation.scala 342:94]
  wire  _s0_enqDataCapture_0_0_T_2 = io_slowPorts_2_valid & dataCond_6; // @[ReservationStation.scala 342:94]
  wire  _s0_enqDataCapture_0_0_T_3 = io_slowPorts_3_valid & dataCond_9; // @[ReservationStation.scala 342:94]
  wire  _s0_enqDataCapture_0_0_T_4 = io_slowPorts_4_valid & dataCond_12; // @[ReservationStation.scala 342:94]
  wire [1:0] s0_enqDataCapture_0_0_lo = {_s0_enqDataCapture_0_0_T_1,_s0_enqDataCapture_0_0_T}; // @[ReservationStation.scala 342:104]
  wire [2:0] s0_enqDataCapture_0_0_hi = {_s0_enqDataCapture_0_0_T_4,_s0_enqDataCapture_0_0_T_3,
    _s0_enqDataCapture_0_0_T_2}; // @[ReservationStation.scala 342:104]
  wire  _s0_enqWakeup_0_1_T = io_slowPorts_0_valid & stateCond_1; // @[ReservationStation.scala 341:90]
  wire  _s0_enqWakeup_0_1_T_1 = io_slowPorts_1_valid & stateCond_4; // @[ReservationStation.scala 341:90]
  wire  _s0_enqWakeup_0_1_T_2 = io_slowPorts_2_valid & stateCond_7; // @[ReservationStation.scala 341:90]
  wire  _s0_enqWakeup_0_1_T_3 = io_slowPorts_3_valid & stateCond_10; // @[ReservationStation.scala 341:90]
  wire  _s0_enqWakeup_0_1_T_4 = io_slowPorts_4_valid & stateCond_13; // @[ReservationStation.scala 341:90]
  wire [1:0] s0_enqWakeup_0_1_lo = {_s0_enqWakeup_0_1_T_1,_s0_enqWakeup_0_1_T}; // @[ReservationStation.scala 341:100]
  wire [2:0] s0_enqWakeup_0_1_hi = {_s0_enqWakeup_0_1_T_4,_s0_enqWakeup_0_1_T_3,_s0_enqWakeup_0_1_T_2}; // @[ReservationStation.scala 341:100]
  wire  _s0_enqDataCapture_0_1_T = io_slowPorts_0_valid & dataCond_1; // @[ReservationStation.scala 342:94]
  wire  _s0_enqDataCapture_0_1_T_1 = io_slowPorts_1_valid & dataCond_4; // @[ReservationStation.scala 342:94]
  wire  _s0_enqDataCapture_0_1_T_2 = io_slowPorts_2_valid & dataCond_7; // @[ReservationStation.scala 342:94]
  wire  _s0_enqDataCapture_0_1_T_3 = io_slowPorts_3_valid & dataCond_10; // @[ReservationStation.scala 342:94]
  wire  _s0_enqDataCapture_0_1_T_4 = io_slowPorts_4_valid & dataCond_13; // @[ReservationStation.scala 342:94]
  wire [1:0] s0_enqDataCapture_0_1_lo = {_s0_enqDataCapture_0_1_T_1,_s0_enqDataCapture_0_1_T}; // @[ReservationStation.scala 342:104]
  wire [2:0] s0_enqDataCapture_0_1_hi = {_s0_enqDataCapture_0_1_T_4,_s0_enqDataCapture_0_1_T_3,
    _s0_enqDataCapture_0_1_T_2}; // @[ReservationStation.scala 342:104]
  wire  pdestMatch_18 = io_slowPorts_0_bits_uop_pdest == io_fromDispatch_1_bits_psrc_0; // @[Bundle.scala 262:30]
  wire  stateCond_18 = pdestMatch_18 & io_slowPorts_0_bits_uop_ctrl_rfWen; // @[Bundle.scala 268:34]
  wire  rfDataMatch_18 = io_slowPorts_0_bits_uop_ctrl_rfWen & io_fromDispatch_1_bits_psrc_0 != 6'h0; // @[Bundle.scala 270:58]
  wire  _dataCond_T_90 = io_fromDispatch_1_bits_ctrl_srcType_0 == 2'h0; // @[package.scala 37:39]
  wire  dataCond_18 = pdestMatch_18 & (rfDataMatch_18 & _dataCond_T_90); // @[Bundle.scala 271:33]
  wire  pdestMatch_19 = io_slowPorts_0_bits_uop_pdest == io_fromDispatch_1_bits_psrc_1; // @[Bundle.scala 262:30]
  wire  stateCond_19 = pdestMatch_19 & io_slowPorts_0_bits_uop_ctrl_rfWen; // @[Bundle.scala 268:34]
  wire  rfDataMatch_19 = io_slowPorts_0_bits_uop_ctrl_rfWen & io_fromDispatch_1_bits_psrc_1 != 6'h0; // @[Bundle.scala 270:58]
  wire  _dataCond_T_95 = io_fromDispatch_1_bits_ctrl_srcType_1 == 2'h0; // @[package.scala 37:39]
  wire  dataCond_19 = pdestMatch_19 & (rfDataMatch_19 & _dataCond_T_95); // @[Bundle.scala 271:33]
  wire  pdestMatch_21 = io_slowPorts_1_bits_uop_pdest == io_fromDispatch_1_bits_psrc_0; // @[Bundle.scala 262:30]
  wire  stateCond_21 = pdestMatch_21 & io_slowPorts_1_bits_uop_ctrl_rfWen; // @[Bundle.scala 268:34]
  wire  rfDataMatch_21 = io_slowPorts_1_bits_uop_ctrl_rfWen & io_fromDispatch_1_bits_psrc_0 != 6'h0; // @[Bundle.scala 270:58]
  wire  dataCond_21 = pdestMatch_21 & (rfDataMatch_21 & _dataCond_T_90); // @[Bundle.scala 271:33]
  wire  pdestMatch_22 = io_slowPorts_1_bits_uop_pdest == io_fromDispatch_1_bits_psrc_1; // @[Bundle.scala 262:30]
  wire  stateCond_22 = pdestMatch_22 & io_slowPorts_1_bits_uop_ctrl_rfWen; // @[Bundle.scala 268:34]
  wire  rfDataMatch_22 = io_slowPorts_1_bits_uop_ctrl_rfWen & io_fromDispatch_1_bits_psrc_1 != 6'h0; // @[Bundle.scala 270:58]
  wire  dataCond_22 = pdestMatch_22 & (rfDataMatch_22 & _dataCond_T_95); // @[Bundle.scala 271:33]
  wire  pdestMatch_24 = io_slowPorts_2_bits_uop_pdest == io_fromDispatch_1_bits_psrc_0; // @[Bundle.scala 262:30]
  wire  stateCond_24 = pdestMatch_24 & io_slowPorts_2_bits_uop_ctrl_rfWen; // @[Bundle.scala 268:34]
  wire  rfDataMatch_24 = io_slowPorts_2_bits_uop_ctrl_rfWen & io_fromDispatch_1_bits_psrc_0 != 6'h0; // @[Bundle.scala 270:58]
  wire  dataCond_24 = pdestMatch_24 & (rfDataMatch_24 & _dataCond_T_90); // @[Bundle.scala 271:33]
  wire  pdestMatch_25 = io_slowPorts_2_bits_uop_pdest == io_fromDispatch_1_bits_psrc_1; // @[Bundle.scala 262:30]
  wire  stateCond_25 = pdestMatch_25 & io_slowPorts_2_bits_uop_ctrl_rfWen; // @[Bundle.scala 268:34]
  wire  rfDataMatch_25 = io_slowPorts_2_bits_uop_ctrl_rfWen & io_fromDispatch_1_bits_psrc_1 != 6'h0; // @[Bundle.scala 270:58]
  wire  dataCond_25 = pdestMatch_25 & (rfDataMatch_25 & _dataCond_T_95); // @[Bundle.scala 271:33]
  wire  pdestMatch_27 = io_slowPorts_3_bits_uop_pdest == io_fromDispatch_1_bits_psrc_0; // @[Bundle.scala 262:30]
  wire  stateCond_27 = pdestMatch_27 & io_slowPorts_3_bits_uop_ctrl_rfWen; // @[Bundle.scala 268:34]
  wire  rfDataMatch_27 = io_slowPorts_3_bits_uop_ctrl_rfWen & io_fromDispatch_1_bits_psrc_0 != 6'h0; // @[Bundle.scala 270:58]
  wire  dataCond_27 = pdestMatch_27 & (rfDataMatch_27 & _dataCond_T_90); // @[Bundle.scala 271:33]
  wire  pdestMatch_28 = io_slowPorts_3_bits_uop_pdest == io_fromDispatch_1_bits_psrc_1; // @[Bundle.scala 262:30]
  wire  stateCond_28 = pdestMatch_28 & io_slowPorts_3_bits_uop_ctrl_rfWen; // @[Bundle.scala 268:34]
  wire  rfDataMatch_28 = io_slowPorts_3_bits_uop_ctrl_rfWen & io_fromDispatch_1_bits_psrc_1 != 6'h0; // @[Bundle.scala 270:58]
  wire  dataCond_28 = pdestMatch_28 & (rfDataMatch_28 & _dataCond_T_95); // @[Bundle.scala 271:33]
  wire  pdestMatch_30 = io_slowPorts_4_bits_uop_pdest == io_fromDispatch_1_bits_psrc_0; // @[Bundle.scala 262:30]
  wire  stateCond_30 = pdestMatch_30 & io_slowPorts_4_bits_uop_ctrl_rfWen; // @[Bundle.scala 268:34]
  wire  rfDataMatch_30 = io_slowPorts_4_bits_uop_ctrl_rfWen & io_fromDispatch_1_bits_psrc_0 != 6'h0; // @[Bundle.scala 270:58]
  wire  dataCond_30 = pdestMatch_30 & (rfDataMatch_30 & _dataCond_T_90); // @[Bundle.scala 271:33]
  wire  pdestMatch_31 = io_slowPorts_4_bits_uop_pdest == io_fromDispatch_1_bits_psrc_1; // @[Bundle.scala 262:30]
  wire  stateCond_31 = pdestMatch_31 & io_slowPorts_4_bits_uop_ctrl_rfWen; // @[Bundle.scala 268:34]
  wire  rfDataMatch_31 = io_slowPorts_4_bits_uop_ctrl_rfWen & io_fromDispatch_1_bits_psrc_1 != 6'h0; // @[Bundle.scala 270:58]
  wire  dataCond_31 = pdestMatch_31 & (rfDataMatch_31 & _dataCond_T_95); // @[Bundle.scala 271:33]
  wire  pdestMatch_33 = io_fastUopsIn_0_bits_pdest == io_fromDispatch_1_bits_psrc_0; // @[Bundle.scala 262:30]
  wire  rfDataMatch_33 = io_fastUopsIn_0_bits_ctrl_rfWen & io_fromDispatch_1_bits_psrc_0 != 6'h0; // @[Bundle.scala 270:58]
  wire  dataCond_33 = pdestMatch_33 & (rfDataMatch_33 & _dataCond_T_90); // @[Bundle.scala 271:33]
  wire  pdestMatch_34 = io_fastUopsIn_0_bits_pdest == io_fromDispatch_1_bits_psrc_1; // @[Bundle.scala 262:30]
  wire  rfDataMatch_34 = io_fastUopsIn_0_bits_ctrl_rfWen & io_fromDispatch_1_bits_psrc_1 != 6'h0; // @[Bundle.scala 270:58]
  wire  dataCond_34 = pdestMatch_34 & (rfDataMatch_34 & _dataCond_T_95); // @[Bundle.scala 271:33]
  wire  _s0_enqWakeup_1_0_T = io_slowPorts_0_valid & stateCond_18; // @[ReservationStation.scala 341:90]
  wire  _s0_enqWakeup_1_0_T_1 = io_slowPorts_1_valid & stateCond_21; // @[ReservationStation.scala 341:90]
  wire  _s0_enqWakeup_1_0_T_2 = io_slowPorts_2_valid & stateCond_24; // @[ReservationStation.scala 341:90]
  wire  _s0_enqWakeup_1_0_T_3 = io_slowPorts_3_valid & stateCond_27; // @[ReservationStation.scala 341:90]
  wire  _s0_enqWakeup_1_0_T_4 = io_slowPorts_4_valid & stateCond_30; // @[ReservationStation.scala 341:90]
  wire [1:0] s0_enqWakeup_1_0_lo = {_s0_enqWakeup_1_0_T_1,_s0_enqWakeup_1_0_T}; // @[ReservationStation.scala 341:100]
  wire [2:0] s0_enqWakeup_1_0_hi = {_s0_enqWakeup_1_0_T_4,_s0_enqWakeup_1_0_T_3,_s0_enqWakeup_1_0_T_2}; // @[ReservationStation.scala 341:100]
  wire  _s0_enqDataCapture_1_0_T = io_slowPorts_0_valid & dataCond_18; // @[ReservationStation.scala 342:94]
  wire  _s0_enqDataCapture_1_0_T_1 = io_slowPorts_1_valid & dataCond_21; // @[ReservationStation.scala 342:94]
  wire  _s0_enqDataCapture_1_0_T_2 = io_slowPorts_2_valid & dataCond_24; // @[ReservationStation.scala 342:94]
  wire  _s0_enqDataCapture_1_0_T_3 = io_slowPorts_3_valid & dataCond_27; // @[ReservationStation.scala 342:94]
  wire  _s0_enqDataCapture_1_0_T_4 = io_slowPorts_4_valid & dataCond_30; // @[ReservationStation.scala 342:94]
  wire [1:0] s0_enqDataCapture_1_0_lo = {_s0_enqDataCapture_1_0_T_1,_s0_enqDataCapture_1_0_T}; // @[ReservationStation.scala 342:104]
  wire [2:0] s0_enqDataCapture_1_0_hi = {_s0_enqDataCapture_1_0_T_4,_s0_enqDataCapture_1_0_T_3,
    _s0_enqDataCapture_1_0_T_2}; // @[ReservationStation.scala 342:104]
  wire  _s0_enqWakeup_1_1_T = io_slowPorts_0_valid & stateCond_19; // @[ReservationStation.scala 341:90]
  wire  _s0_enqWakeup_1_1_T_1 = io_slowPorts_1_valid & stateCond_22; // @[ReservationStation.scala 341:90]
  wire  _s0_enqWakeup_1_1_T_2 = io_slowPorts_2_valid & stateCond_25; // @[ReservationStation.scala 341:90]
  wire  _s0_enqWakeup_1_1_T_3 = io_slowPorts_3_valid & stateCond_28; // @[ReservationStation.scala 341:90]
  wire  _s0_enqWakeup_1_1_T_4 = io_slowPorts_4_valid & stateCond_31; // @[ReservationStation.scala 341:90]
  wire [1:0] s0_enqWakeup_1_1_lo = {_s0_enqWakeup_1_1_T_1,_s0_enqWakeup_1_1_T}; // @[ReservationStation.scala 341:100]
  wire [2:0] s0_enqWakeup_1_1_hi = {_s0_enqWakeup_1_1_T_4,_s0_enqWakeup_1_1_T_3,_s0_enqWakeup_1_1_T_2}; // @[ReservationStation.scala 341:100]
  wire  _s0_enqDataCapture_1_1_T = io_slowPorts_0_valid & dataCond_19; // @[ReservationStation.scala 342:94]
  wire  _s0_enqDataCapture_1_1_T_1 = io_slowPorts_1_valid & dataCond_22; // @[ReservationStation.scala 342:94]
  wire  _s0_enqDataCapture_1_1_T_2 = io_slowPorts_2_valid & dataCond_25; // @[ReservationStation.scala 342:94]
  wire  _s0_enqDataCapture_1_1_T_3 = io_slowPorts_3_valid & dataCond_28; // @[ReservationStation.scala 342:94]
  wire  _s0_enqDataCapture_1_1_T_4 = io_slowPorts_4_valid & dataCond_31; // @[ReservationStation.scala 342:94]
  wire [1:0] s0_enqDataCapture_1_1_lo = {_s0_enqDataCapture_1_1_T_1,_s0_enqDataCapture_1_1_T}; // @[ReservationStation.scala 342:104]
  wire [2:0] s0_enqDataCapture_1_1_hi = {_s0_enqDataCapture_1_1_T_4,_s0_enqDataCapture_1_1_T_3,
    _s0_enqDataCapture_1_1_T_2}; // @[ReservationStation.scala 342:104]
  reg [7:0] enqVec_REG; // @[ReservationStation.scala 361:86]
  reg [7:0] enqVec_REG_1; // @[ReservationStation.scala 361:86]
  wire [7:0] _s1_oldestSel_out_valid_T = statusArray_io_canIssue & s1_oldestSel_age_io_out; // @[SelectPolicy.scala 178:28]
  reg  s1_dispatchUops_dup_0_0_valid; // @[ReservationStation.scala 391:32]
  reg [1:0] s1_dispatchUops_dup_0_0_bits_ctrl_srcType_0; // @[ReservationStation.scala 391:32]
  reg [1:0] s1_dispatchUops_dup_0_0_bits_ctrl_srcType_1; // @[ReservationStation.scala 391:32]
  reg [3:0] s1_dispatchUops_dup_0_0_bits_ctrl_fuType; // @[ReservationStation.scala 391:32]
  reg [6:0] s1_dispatchUops_dup_0_0_bits_ctrl_fuOpType; // @[ReservationStation.scala 391:32]
  reg  s1_dispatchUops_dup_0_0_bits_ctrl_rfWen; // @[ReservationStation.scala 391:32]
  reg  s1_dispatchUops_dup_0_0_bits_ctrl_fpWen; // @[ReservationStation.scala 391:32]
  reg  s1_dispatchUops_dup_0_0_bits_srcState_0; // @[ReservationStation.scala 391:32]
  reg  s1_dispatchUops_dup_0_0_bits_srcState_1; // @[ReservationStation.scala 391:32]
  reg [5:0] s1_dispatchUops_dup_0_0_bits_psrc_0; // @[ReservationStation.scala 391:32]
  reg [5:0] s1_dispatchUops_dup_0_0_bits_psrc_1; // @[ReservationStation.scala 391:32]
  reg [5:0] s1_dispatchUops_dup_0_0_bits_pdest; // @[ReservationStation.scala 391:32]
  reg  s1_dispatchUops_dup_0_0_bits_robIdx_flag; // @[ReservationStation.scala 391:32]
  reg [4:0] s1_dispatchUops_dup_0_0_bits_robIdx_value; // @[ReservationStation.scala 391:32]
  reg  s1_dispatchUops_dup_0_1_valid; // @[ReservationStation.scala 391:32]
  reg [1:0] s1_dispatchUops_dup_0_1_bits_ctrl_srcType_0; // @[ReservationStation.scala 391:32]
  reg [1:0] s1_dispatchUops_dup_0_1_bits_ctrl_srcType_1; // @[ReservationStation.scala 391:32]
  reg  s1_dispatchUops_dup_0_1_bits_srcState_0; // @[ReservationStation.scala 391:32]
  reg  s1_dispatchUops_dup_0_1_bits_srcState_1; // @[ReservationStation.scala 391:32]
  reg [5:0] s1_dispatchUops_dup_0_1_bits_psrc_0; // @[ReservationStation.scala 391:32]
  reg [5:0] s1_dispatchUops_dup_0_1_bits_psrc_1; // @[ReservationStation.scala 391:32]
  reg  s1_dispatchUops_dup_0_1_bits_robIdx_flag; // @[ReservationStation.scala 391:32]
  reg [4:0] s1_dispatchUops_dup_0_1_bits_robIdx_value; // @[ReservationStation.scala 391:32]
  reg  s1_dispatchUops_dup_1_0_valid; // @[ReservationStation.scala 391:32]
  reg [3:0] s1_dispatchUops_dup_1_0_bits_ctrl_fuType; // @[ReservationStation.scala 391:32]
  reg [6:0] s1_dispatchUops_dup_1_0_bits_ctrl_fuOpType; // @[ReservationStation.scala 391:32]
  reg  s1_dispatchUops_dup_1_0_bits_ctrl_rfWen; // @[ReservationStation.scala 391:32]
  reg  s1_dispatchUops_dup_1_0_bits_ctrl_fpWen; // @[ReservationStation.scala 391:32]
  reg [5:0] s1_dispatchUops_dup_1_0_bits_pdest; // @[ReservationStation.scala 391:32]
  reg  s1_dispatchUops_dup_1_0_bits_robIdx_flag; // @[ReservationStation.scala 391:32]
  reg [4:0] s1_dispatchUops_dup_1_0_bits_robIdx_value; // @[ReservationStation.scala 391:32]
  reg  s1_dispatchUops_dup_1_1_valid; // @[ReservationStation.scala 391:32]
  reg [3:0] s1_dispatchUops_dup_1_1_bits_ctrl_fuType; // @[ReservationStation.scala 391:32]
  reg [6:0] s1_dispatchUops_dup_1_1_bits_ctrl_fuOpType; // @[ReservationStation.scala 391:32]
  reg  s1_dispatchUops_dup_1_1_bits_ctrl_rfWen; // @[ReservationStation.scala 391:32]
  reg  s1_dispatchUops_dup_1_1_bits_ctrl_fpWen; // @[ReservationStation.scala 391:32]
  reg [5:0] s1_dispatchUops_dup_1_1_bits_pdest; // @[ReservationStation.scala 391:32]
  reg  s1_dispatchUops_dup_1_1_bits_robIdx_flag; // @[ReservationStation.scala 391:32]
  reg [4:0] s1_dispatchUops_dup_1_1_bits_robIdx_value; // @[ReservationStation.scala 391:32]
  reg  s1_dispatchUops_dup_2_0_valid; // @[ReservationStation.scala 391:32]
  reg [1:0] s1_dispatchUops_dup_2_0_bits_ctrl_srcType_0; // @[ReservationStation.scala 391:32]
  reg [1:0] s1_dispatchUops_dup_2_0_bits_ctrl_srcType_1; // @[ReservationStation.scala 391:32]
  reg [19:0] s1_dispatchUops_dup_2_0_bits_ctrl_imm; // @[ReservationStation.scala 391:32]
  reg  s1_dispatchUops_dup_2_0_bits_srcState_0; // @[ReservationStation.scala 391:32]
  reg  s1_dispatchUops_dup_2_0_bits_srcState_1; // @[ReservationStation.scala 391:32]
  reg  s1_dispatchUops_dup_2_1_valid; // @[ReservationStation.scala 391:32]
  reg [1:0] s1_dispatchUops_dup_2_1_bits_ctrl_srcType_0; // @[ReservationStation.scala 391:32]
  reg [1:0] s1_dispatchUops_dup_2_1_bits_ctrl_srcType_1; // @[ReservationStation.scala 391:32]
  reg [19:0] s1_dispatchUops_dup_2_1_bits_ctrl_imm; // @[ReservationStation.scala 391:32]
  reg  s1_dispatchUops_dup_2_1_bits_srcState_0; // @[ReservationStation.scala 391:32]
  reg  s1_dispatchUops_dup_2_1_bits_srcState_1; // @[ReservationStation.scala 391:32]
  reg [7:0] s1_allocatePtrOH_dup_0_0; // @[ReservationStation.scala 393:37]
  reg [7:0] s1_allocatePtrOH_dup_0_1; // @[ReservationStation.scala 393:37]
  reg [7:0] s1_allocatePtrOH_dup_1_0; // @[ReservationStation.scala 393:37]
  reg [7:0] s1_allocatePtrOH_dup_1_1; // @[ReservationStation.scala 393:37]
  reg [7:0] s1_allocatePtrOH_dup_2_0; // @[ReservationStation.scala 393:37]
  reg [7:0] s1_allocatePtrOH_dup_2_1; // @[ReservationStation.scala 393:37]
  reg [4:0] s1_enqWakeup_0_0; // @[ReservationStation.scala 395:29]
  reg [4:0] s1_enqWakeup_0_1; // @[ReservationStation.scala 395:29]
  reg [4:0] s1_enqWakeup_1_0; // @[ReservationStation.scala 395:29]
  reg [4:0] s1_enqWakeup_1_1; // @[ReservationStation.scala 395:29]
  reg [4:0] s1_enqDataCapture_0_0; // @[ReservationStation.scala 396:34]
  reg [4:0] s1_enqDataCapture_0_1; // @[ReservationStation.scala 396:34]
  reg [4:0] s1_enqDataCapture_1_0; // @[ReservationStation.scala 396:34]
  reg [4:0] s1_enqDataCapture_1_1; // @[ReservationStation.scala 396:34]
  reg  s1_fastWakeup_0_0_0; // @[ReservationStation.scala 397:30]
  reg  s1_fastWakeup_0_1_0; // @[ReservationStation.scala 397:30]
  reg  s1_fastWakeup_1_0_0; // @[ReservationStation.scala 397:30]
  reg  s1_fastWakeup_1_1_0; // @[ReservationStation.scala 397:30]
  wire  s1_issue_oldest_0 = oldestSelection_io_isOverrided_0; // @[ReservationStation.scala 402:29 504:21]
  wire [7:0] s1_in_oldestPtrOH_bits = s1_oldestSel_age_io_out; // @[SelectPolicy.scala 177:19 179:14]
  wire  _s1_issuePtrOH_0_valid_T = s1_issue_oldest_0 | select_io_grant_0_valid; // @[ReservationStation.scala 514:50]
  wire  _canBypass_WIRE_1 = statusArray_io_update_0_data_srcState_1; // @[StatusArray.scala 61:{13,13}]
  wire  _canBypass_WIRE_0 = statusArray_io_update_0_data_srcState_0; // @[StatusArray.scala 61:{13,13}]
  wire [1:0] _canBypass_T = {_canBypass_WIRE_1,_canBypass_WIRE_0}; // @[StatusArray.scala 61:31]
  wire  _canBypass_T_1 = &_canBypass_T; // @[StatusArray.scala 61:38]
  wire  canBypass = s1_dispatchUops_dup_0_0_valid & _canBypass_T_1; // @[ReservationStation.scala 511:55]
  wire  s1_issuePtrOH_0_valid = s1_issue_oldest_0 | select_io_grant_0_valid | canBypass; // @[ReservationStation.scala 514:77]
  wire  _statusArray_io_update_0_data_srcState_0_T_2 = s1_dispatchUops_dup_0_0_bits_ctrl_srcType_0[0] |
    s1_dispatchUops_dup_0_0_bits_srcState_0; // @[Bundle.scala 245:81]
  wire  _statusArray_io_update_0_data_srcState_0_T_5 = s1_dispatchUops_dup_0_0_bits_ctrl_srcType_1[0] |
    s1_dispatchUops_dup_0_0_bits_srcState_1; // @[Bundle.scala 245:81]
  wire  _statusArray_io_update_1_data_srcState_0_T_2 = s1_dispatchUops_dup_0_1_bits_ctrl_srcType_0[0] |
    s1_dispatchUops_dup_0_1_bits_srcState_0; // @[Bundle.scala 245:81]
  wire  _statusArray_io_update_1_data_srcState_0_T_5 = s1_dispatchUops_dup_0_1_bits_ctrl_srcType_1[0] |
    s1_dispatchUops_dup_0_1_bits_srcState_1; // @[Bundle.scala 245:81]
  wire  _s1_issue_dispatch_0_T = ~s1_issue_oldest_0; // @[ReservationStation.scala 512:42]
  wire  s1_issue_dispatch_0 = canBypass & ~s1_issue_oldest_0 & ~select_io_grant_0_valid; // @[ReservationStation.scala 512:62]
  reg  valid; // @[PipelineConnect.scala 108:24]
  wire  s2_deq_0_ready = ~valid | io_deq_0_ready; // @[ReservationStation.scala 747:41]
  wire  _statusArray_io_issueGranted_2_valid_T_1 = select_io_grant_0_valid & _s1_issue_dispatch_0_T; // @[ReservationStation.scala 484:49]
  wire  statusArray_io_issueGranted_3_valid_xs_0 = s1_issue_oldest_0 & s2_deq_0_ready; // @[ParallelMux.scala 64:44]
  wire [3:0] _s1_out_0_bits_uop_T_ctrl_fuType = select_io_grant_0_valid ? payloadArray_io_read_0_data_ctrl_fuType :
    s1_dispatchUops_dup_0_0_bits_ctrl_fuType; // @[ReservationStation.scala 519:10]
  wire  _s1_out_0_bits_uop_T_ctrl_rfWen = select_io_grant_0_valid ? payloadArray_io_read_0_data_ctrl_rfWen :
    s1_dispatchUops_dup_0_0_bits_ctrl_rfWen; // @[ReservationStation.scala 519:10]
  wire [5:0] _s1_out_0_bits_uop_T_pdest = select_io_grant_0_valid ? payloadArray_io_read_0_data_pdest :
    s1_dispatchUops_dup_0_0_bits_pdest; // @[ReservationStation.scala 519:10]
  wire  _s1_out_0_bits_uop_T_robIdx_flag = select_io_grant_0_valid ? payloadArray_io_read_0_data_robIdx_flag :
    s1_dispatchUops_dup_0_0_bits_robIdx_flag; // @[ReservationStation.scala 519:10]
  wire [4:0] _s1_out_0_bits_uop_T_robIdx_value = select_io_grant_0_valid ? payloadArray_io_read_0_data_robIdx_value :
    s1_dispatchUops_dup_0_0_bits_robIdx_value; // @[ReservationStation.scala 519:10]
  wire [3:0] s1_out_0_bits_uop_ctrl_fuType = s1_issue_oldest_0 ? payloadArray_io_read_1_data_ctrl_fuType :
    _s1_out_0_bits_uop_T_ctrl_fuType; // @[ReservationStation.scala 518:30]
  wire  s1_out_0_bits_uop_robIdx_flag = s1_issue_oldest_0 ? payloadArray_io_read_1_data_robIdx_flag :
    _s1_out_0_bits_uop_T_robIdx_flag; // @[ReservationStation.scala 518:30]
  wire [4:0] s1_out_0_bits_uop_robIdx_value = s1_issue_oldest_0 ? payloadArray_io_read_1_data_robIdx_value :
    _s1_out_0_bits_uop_T_robIdx_value; // @[ReservationStation.scala 518:30]
  wire [5:0] _s1_out_0_valid_flushItself_T_1 = {s1_out_0_bits_uop_robIdx_flag,s1_out_0_bits_uop_robIdx_value}; // @[CircularQueuePtr.scala 61:50]
  wire [5:0] _s1_out_0_valid_flushItself_T_2 = {io_redirect_bits_robIdx_flag,io_redirect_bits_robIdx_value}; // @[CircularQueuePtr.scala 61:70]
  wire  _s1_out_0_valid_flushItself_T_3 = _s1_out_0_valid_flushItself_T_1 == _s1_out_0_valid_flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  s1_out_0_valid_flushItself = io_redirect_bits_level & _s1_out_0_valid_flushItself_T_3; // @[Rob.scala 122:51]
  wire  s1_out_0_valid_differentFlag = s1_out_0_bits_uop_robIdx_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  s1_out_0_valid_compare = s1_out_0_bits_uop_robIdx_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _s1_out_0_valid_T = s1_out_0_valid_differentFlag ^ s1_out_0_valid_compare; // @[CircularQueuePtr.scala 88:19]
  wire  _s1_out_0_valid_T_2 = io_redirect_valid & (s1_out_0_valid_flushItself | _s1_out_0_valid_T); // @[Rob.scala 123:20]
  wire  s1_out_0_valid = s1_issuePtrOH_0_valid & ~_s1_out_0_valid_T_2; // @[ReservationStation.scala 532:47]
  wire  fuCheck = s1_out_0_bits_uop_ctrl_fuType == 4'h4; // @[ReservationStation.scala 565:70]
  wire  _T_18 = ~s2_deq_0_ready; // @[ReservationStation.scala 572:81]
  reg [4:0] slowWakeupMatchVec_0_0; // @[ReservationStation.scala 626:31]
  reg [4:0] slowWakeupMatchVec_0_1; // @[ReservationStation.scala 626:31]
  reg [4:0] slowWakeupMatchVec_1_0; // @[ReservationStation.scala 626:31]
  reg [4:0] slowWakeupMatchVec_1_1; // @[ReservationStation.scala 626:31]
  reg [4:0] slowWakeupMatchVec_2_0; // @[ReservationStation.scala 626:31]
  reg [4:0] slowWakeupMatchVec_2_1; // @[ReservationStation.scala 626:31]
  reg [4:0] slowWakeupMatchVec_3_0; // @[ReservationStation.scala 626:31]
  reg [4:0] slowWakeupMatchVec_3_1; // @[ReservationStation.scala 626:31]
  reg [4:0] slowWakeupMatchVec_4_0; // @[ReservationStation.scala 626:31]
  reg [4:0] slowWakeupMatchVec_4_1; // @[ReservationStation.scala 626:31]
  reg [4:0] slowWakeupMatchVec_5_0; // @[ReservationStation.scala 626:31]
  reg [4:0] slowWakeupMatchVec_5_1; // @[ReservationStation.scala 626:31]
  reg [4:0] slowWakeupMatchVec_6_0; // @[ReservationStation.scala 626:31]
  reg [4:0] slowWakeupMatchVec_6_1; // @[ReservationStation.scala 626:31]
  reg [4:0] slowWakeupMatchVec_7_0; // @[ReservationStation.scala 626:31]
  reg [4:0] slowWakeupMatchVec_7_1; // @[ReservationStation.scala 626:31]
  reg  dataArray_io_multiWrite_0_enable_REG; // @[ReservationStation.scala 633:24]
  wire  allocateValid_0 = s1_enqDataCapture_0_0[0] & s1_dispatchUops_dup_2_0_valid; // @[ReservationStation.scala 635:93]
  wire  allocateValid_1 = s1_enqDataCapture_1_0[0] & s1_dispatchUops_dup_2_1_valid; // @[ReservationStation.scala 635:93]
  wire [7:0] allocateDataCapture_xs_0 = allocateValid_0 ? s1_allocatePtrOH_dup_2_0 : 8'h0; // @[ParallelMux.scala 64:44]
  wire [7:0] allocateDataCapture_xs_1 = allocateValid_1 ? s1_allocatePtrOH_dup_2_1 : 8'h0; // @[ParallelMux.scala 64:44]
  wire [7:0] allocateDataCapture = allocateDataCapture_xs_0 | allocateDataCapture_xs_1; // @[ParallelMux.scala 36:53]
  wire [7:0] _dataArray_io_multiWrite_0_addr_0_T_8 = {slowWakeupMatchVec_7_0[0],slowWakeupMatchVec_6_0[0],
    slowWakeupMatchVec_5_0[0],slowWakeupMatchVec_4_0[0],slowWakeupMatchVec_3_0[0],slowWakeupMatchVec_2_0[0],
    slowWakeupMatchVec_1_0[0],slowWakeupMatchVec_0_0[0]}; // @[ReservationStation.scala 637:61]
  wire  allocateValid_0_1 = s1_enqDataCapture_0_1[0] & s1_dispatchUops_dup_2_0_valid; // @[ReservationStation.scala 635:93]
  wire  allocateValid_1_1 = s1_enqDataCapture_1_1[0] & s1_dispatchUops_dup_2_1_valid; // @[ReservationStation.scala 635:93]
  wire [7:0] allocateDataCapture_xs_0_1 = allocateValid_0_1 ? s1_allocatePtrOH_dup_2_0 : 8'h0; // @[ParallelMux.scala 64:44]
  wire [7:0] allocateDataCapture_xs_1_1 = allocateValid_1_1 ? s1_allocatePtrOH_dup_2_1 : 8'h0; // @[ParallelMux.scala 64:44]
  wire [7:0] allocateDataCapture_1 = allocateDataCapture_xs_0_1 | allocateDataCapture_xs_1_1; // @[ParallelMux.scala 36:53]
  wire [7:0] _dataArray_io_multiWrite_0_addr_1_T_8 = {slowWakeupMatchVec_7_1[0],slowWakeupMatchVec_6_1[0],
    slowWakeupMatchVec_5_1[0],slowWakeupMatchVec_4_1[0],slowWakeupMatchVec_3_1[0],slowWakeupMatchVec_2_1[0],
    slowWakeupMatchVec_1_1[0],slowWakeupMatchVec_0_1[0]}; // @[ReservationStation.scala 637:61]
  reg [63:0] dataArray_io_multiWrite_0_data_r; // @[Reg.scala 16:16]
  reg  dataArray_io_multiWrite_1_enable_REG; // @[ReservationStation.scala 633:24]
  wire  allocateValid_0_2 = s1_enqDataCapture_0_0[1] & s1_dispatchUops_dup_2_0_valid; // @[ReservationStation.scala 635:93]
  wire  allocateValid_1_2 = s1_enqDataCapture_1_0[1] & s1_dispatchUops_dup_2_1_valid; // @[ReservationStation.scala 635:93]
  wire [7:0] allocateDataCapture_xs_0_2 = allocateValid_0_2 ? s1_allocatePtrOH_dup_2_0 : 8'h0; // @[ParallelMux.scala 64:44]
  wire [7:0] allocateDataCapture_xs_1_2 = allocateValid_1_2 ? s1_allocatePtrOH_dup_2_1 : 8'h0; // @[ParallelMux.scala 64:44]
  wire [7:0] allocateDataCapture_2 = allocateDataCapture_xs_0_2 | allocateDataCapture_xs_1_2; // @[ParallelMux.scala 36:53]
  wire [7:0] _dataArray_io_multiWrite_1_addr_0_T_8 = {slowWakeupMatchVec_7_0[1],slowWakeupMatchVec_6_0[1],
    slowWakeupMatchVec_5_0[1],slowWakeupMatchVec_4_0[1],slowWakeupMatchVec_3_0[1],slowWakeupMatchVec_2_0[1],
    slowWakeupMatchVec_1_0[1],slowWakeupMatchVec_0_0[1]}; // @[ReservationStation.scala 637:61]
  wire  allocateValid_0_3 = s1_enqDataCapture_0_1[1] & s1_dispatchUops_dup_2_0_valid; // @[ReservationStation.scala 635:93]
  wire  allocateValid_1_3 = s1_enqDataCapture_1_1[1] & s1_dispatchUops_dup_2_1_valid; // @[ReservationStation.scala 635:93]
  wire [7:0] allocateDataCapture_xs_0_3 = allocateValid_0_3 ? s1_allocatePtrOH_dup_2_0 : 8'h0; // @[ParallelMux.scala 64:44]
  wire [7:0] allocateDataCapture_xs_1_3 = allocateValid_1_3 ? s1_allocatePtrOH_dup_2_1 : 8'h0; // @[ParallelMux.scala 64:44]
  wire [7:0] allocateDataCapture_3 = allocateDataCapture_xs_0_3 | allocateDataCapture_xs_1_3; // @[ParallelMux.scala 36:53]
  wire [7:0] _dataArray_io_multiWrite_1_addr_1_T_8 = {slowWakeupMatchVec_7_1[1],slowWakeupMatchVec_6_1[1],
    slowWakeupMatchVec_5_1[1],slowWakeupMatchVec_4_1[1],slowWakeupMatchVec_3_1[1],slowWakeupMatchVec_2_1[1],
    slowWakeupMatchVec_1_1[1],slowWakeupMatchVec_0_1[1]}; // @[ReservationStation.scala 637:61]
  reg [63:0] dataArray_io_multiWrite_1_data_r; // @[Reg.scala 16:16]
  reg  dataArray_io_multiWrite_2_enable_REG; // @[ReservationStation.scala 633:24]
  wire  allocateValid_0_4 = s1_enqDataCapture_0_0[2] & s1_dispatchUops_dup_2_0_valid; // @[ReservationStation.scala 635:93]
  wire  allocateValid_1_4 = s1_enqDataCapture_1_0[2] & s1_dispatchUops_dup_2_1_valid; // @[ReservationStation.scala 635:93]
  wire [7:0] allocateDataCapture_xs_0_4 = allocateValid_0_4 ? s1_allocatePtrOH_dup_2_0 : 8'h0; // @[ParallelMux.scala 64:44]
  wire [7:0] allocateDataCapture_xs_1_4 = allocateValid_1_4 ? s1_allocatePtrOH_dup_2_1 : 8'h0; // @[ParallelMux.scala 64:44]
  wire [7:0] allocateDataCapture_4 = allocateDataCapture_xs_0_4 | allocateDataCapture_xs_1_4; // @[ParallelMux.scala 36:53]
  wire [7:0] _dataArray_io_multiWrite_2_addr_0_T_8 = {slowWakeupMatchVec_7_0[2],slowWakeupMatchVec_6_0[2],
    slowWakeupMatchVec_5_0[2],slowWakeupMatchVec_4_0[2],slowWakeupMatchVec_3_0[2],slowWakeupMatchVec_2_0[2],
    slowWakeupMatchVec_1_0[2],slowWakeupMatchVec_0_0[2]}; // @[ReservationStation.scala 637:61]
  wire  allocateValid_0_5 = s1_enqDataCapture_0_1[2] & s1_dispatchUops_dup_2_0_valid; // @[ReservationStation.scala 635:93]
  wire  allocateValid_1_5 = s1_enqDataCapture_1_1[2] & s1_dispatchUops_dup_2_1_valid; // @[ReservationStation.scala 635:93]
  wire [7:0] allocateDataCapture_xs_0_5 = allocateValid_0_5 ? s1_allocatePtrOH_dup_2_0 : 8'h0; // @[ParallelMux.scala 64:44]
  wire [7:0] allocateDataCapture_xs_1_5 = allocateValid_1_5 ? s1_allocatePtrOH_dup_2_1 : 8'h0; // @[ParallelMux.scala 64:44]
  wire [7:0] allocateDataCapture_5 = allocateDataCapture_xs_0_5 | allocateDataCapture_xs_1_5; // @[ParallelMux.scala 36:53]
  wire [7:0] _dataArray_io_multiWrite_2_addr_1_T_8 = {slowWakeupMatchVec_7_1[2],slowWakeupMatchVec_6_1[2],
    slowWakeupMatchVec_5_1[2],slowWakeupMatchVec_4_1[2],slowWakeupMatchVec_3_1[2],slowWakeupMatchVec_2_1[2],
    slowWakeupMatchVec_1_1[2],slowWakeupMatchVec_0_1[2]}; // @[ReservationStation.scala 637:61]
  reg [63:0] dataArray_io_multiWrite_2_data_r; // @[Reg.scala 16:16]
  reg  dataArray_io_multiWrite_3_enable_REG; // @[ReservationStation.scala 633:24]
  wire  allocateValid_0_6 = s1_enqDataCapture_0_0[3] & s1_dispatchUops_dup_2_0_valid; // @[ReservationStation.scala 635:93]
  wire  allocateValid_1_6 = s1_enqDataCapture_1_0[3] & s1_dispatchUops_dup_2_1_valid; // @[ReservationStation.scala 635:93]
  wire [7:0] allocateDataCapture_xs_0_6 = allocateValid_0_6 ? s1_allocatePtrOH_dup_2_0 : 8'h0; // @[ParallelMux.scala 64:44]
  wire [7:0] allocateDataCapture_xs_1_6 = allocateValid_1_6 ? s1_allocatePtrOH_dup_2_1 : 8'h0; // @[ParallelMux.scala 64:44]
  wire [7:0] allocateDataCapture_6 = allocateDataCapture_xs_0_6 | allocateDataCapture_xs_1_6; // @[ParallelMux.scala 36:53]
  wire [7:0] _dataArray_io_multiWrite_3_addr_0_T_8 = {slowWakeupMatchVec_7_0[3],slowWakeupMatchVec_6_0[3],
    slowWakeupMatchVec_5_0[3],slowWakeupMatchVec_4_0[3],slowWakeupMatchVec_3_0[3],slowWakeupMatchVec_2_0[3],
    slowWakeupMatchVec_1_0[3],slowWakeupMatchVec_0_0[3]}; // @[ReservationStation.scala 637:61]
  wire  allocateValid_0_7 = s1_enqDataCapture_0_1[3] & s1_dispatchUops_dup_2_0_valid; // @[ReservationStation.scala 635:93]
  wire  allocateValid_1_7 = s1_enqDataCapture_1_1[3] & s1_dispatchUops_dup_2_1_valid; // @[ReservationStation.scala 635:93]
  wire [7:0] allocateDataCapture_xs_0_7 = allocateValid_0_7 ? s1_allocatePtrOH_dup_2_0 : 8'h0; // @[ParallelMux.scala 64:44]
  wire [7:0] allocateDataCapture_xs_1_7 = allocateValid_1_7 ? s1_allocatePtrOH_dup_2_1 : 8'h0; // @[ParallelMux.scala 64:44]
  wire [7:0] allocateDataCapture_7 = allocateDataCapture_xs_0_7 | allocateDataCapture_xs_1_7; // @[ParallelMux.scala 36:53]
  wire [7:0] _dataArray_io_multiWrite_3_addr_1_T_8 = {slowWakeupMatchVec_7_1[3],slowWakeupMatchVec_6_1[3],
    slowWakeupMatchVec_5_1[3],slowWakeupMatchVec_4_1[3],slowWakeupMatchVec_3_1[3],slowWakeupMatchVec_2_1[3],
    slowWakeupMatchVec_1_1[3],slowWakeupMatchVec_0_1[3]}; // @[ReservationStation.scala 637:61]
  reg [63:0] dataArray_io_multiWrite_3_data_r; // @[Reg.scala 16:16]
  reg  dataArray_io_multiWrite_4_enable_REG; // @[ReservationStation.scala 633:24]
  wire  allocateValid_0_8 = s1_enqDataCapture_0_0[4] & s1_dispatchUops_dup_2_0_valid; // @[ReservationStation.scala 635:93]
  wire  allocateValid_1_8 = s1_enqDataCapture_1_0[4] & s1_dispatchUops_dup_2_1_valid; // @[ReservationStation.scala 635:93]
  wire [7:0] allocateDataCapture_xs_0_8 = allocateValid_0_8 ? s1_allocatePtrOH_dup_2_0 : 8'h0; // @[ParallelMux.scala 64:44]
  wire [7:0] allocateDataCapture_xs_1_8 = allocateValid_1_8 ? s1_allocatePtrOH_dup_2_1 : 8'h0; // @[ParallelMux.scala 64:44]
  wire [7:0] allocateDataCapture_8 = allocateDataCapture_xs_0_8 | allocateDataCapture_xs_1_8; // @[ParallelMux.scala 36:53]
  wire [7:0] _dataArray_io_multiWrite_4_addr_0_T_8 = {slowWakeupMatchVec_7_0[4],slowWakeupMatchVec_6_0[4],
    slowWakeupMatchVec_5_0[4],slowWakeupMatchVec_4_0[4],slowWakeupMatchVec_3_0[4],slowWakeupMatchVec_2_0[4],
    slowWakeupMatchVec_1_0[4],slowWakeupMatchVec_0_0[4]}; // @[ReservationStation.scala 637:61]
  wire  allocateValid_0_9 = s1_enqDataCapture_0_1[4] & s1_dispatchUops_dup_2_0_valid; // @[ReservationStation.scala 635:93]
  wire  allocateValid_1_9 = s1_enqDataCapture_1_1[4] & s1_dispatchUops_dup_2_1_valid; // @[ReservationStation.scala 635:93]
  wire [7:0] allocateDataCapture_xs_0_9 = allocateValid_0_9 ? s1_allocatePtrOH_dup_2_0 : 8'h0; // @[ParallelMux.scala 64:44]
  wire [7:0] allocateDataCapture_xs_1_9 = allocateValid_1_9 ? s1_allocatePtrOH_dup_2_1 : 8'h0; // @[ParallelMux.scala 64:44]
  wire [7:0] allocateDataCapture_9 = allocateDataCapture_xs_0_9 | allocateDataCapture_xs_1_9; // @[ParallelMux.scala 36:53]
  wire [7:0] _dataArray_io_multiWrite_4_addr_1_T_8 = {slowWakeupMatchVec_7_1[4],slowWakeupMatchVec_6_1[4],
    slowWakeupMatchVec_5_1[4],slowWakeupMatchVec_4_1[4],slowWakeupMatchVec_3_1[4],slowWakeupMatchVec_2_1[4],
    slowWakeupMatchVec_1_1[4],slowWakeupMatchVec_0_1[4]}; // @[ReservationStation.scala 637:61]
  reg [63:0] dataArray_io_multiWrite_4_data_r; // @[Reg.scala 16:16]
  wire [7:0] _dataSelect_io_fromSlowPorts_0_0_T = dataArray_io_read_0_addr & dataArray_io_multiWrite_0_addr_0; // @[ReservationStation.scala 697:77]
  wire  _dataSelect_io_fromSlowPorts_0_0_T_2 = dataArray_io_multiWrite_0_enable & |_dataSelect_io_fromSlowPorts_0_0_T; // @[ReservationStation.scala 697:68]
  wire [7:0] _dataSelect_io_fromSlowPorts_0_0_T_3 = dataArray_io_read_0_addr & dataArray_io_multiWrite_1_addr_0; // @[ReservationStation.scala 697:77]
  wire  _dataSelect_io_fromSlowPorts_0_0_T_5 = dataArray_io_multiWrite_1_enable & |_dataSelect_io_fromSlowPorts_0_0_T_3; // @[ReservationStation.scala 697:68]
  wire [7:0] _dataSelect_io_fromSlowPorts_0_0_T_6 = dataArray_io_read_0_addr & dataArray_io_multiWrite_2_addr_0; // @[ReservationStation.scala 697:77]
  wire  _dataSelect_io_fromSlowPorts_0_0_T_8 = dataArray_io_multiWrite_2_enable & |_dataSelect_io_fromSlowPorts_0_0_T_6; // @[ReservationStation.scala 697:68]
  wire [7:0] _dataSelect_io_fromSlowPorts_0_0_T_9 = dataArray_io_read_0_addr & dataArray_io_multiWrite_3_addr_0; // @[ReservationStation.scala 697:77]
  wire  _dataSelect_io_fromSlowPorts_0_0_T_11 = dataArray_io_multiWrite_3_enable & |_dataSelect_io_fromSlowPorts_0_0_T_9
    ; // @[ReservationStation.scala 697:68]
  wire [7:0] _dataSelect_io_fromSlowPorts_0_0_T_12 = dataArray_io_read_0_addr & dataArray_io_multiWrite_4_addr_0; // @[ReservationStation.scala 697:77]
  wire  _dataSelect_io_fromSlowPorts_0_0_T_14 = dataArray_io_multiWrite_4_enable & |
    _dataSelect_io_fromSlowPorts_0_0_T_12; // @[ReservationStation.scala 697:68]
  wire [1:0] dataSelect_io_fromSlowPorts_0_0_lo = {_dataSelect_io_fromSlowPorts_0_0_T_5,
    _dataSelect_io_fromSlowPorts_0_0_T_2}; // @[ReservationStation.scala 697:103]
  wire [2:0] dataSelect_io_fromSlowPorts_0_0_hi = {_dataSelect_io_fromSlowPorts_0_0_T_14,
    _dataSelect_io_fromSlowPorts_0_0_T_11,_dataSelect_io_fromSlowPorts_0_0_T_8}; // @[ReservationStation.scala 697:103]
  wire [7:0] _dataSelect_io_fromSlowPorts_0_1_T = dataArray_io_read_0_addr & dataArray_io_multiWrite_0_addr_1; // @[ReservationStation.scala 697:77]
  wire  _dataSelect_io_fromSlowPorts_0_1_T_2 = dataArray_io_multiWrite_0_enable & |_dataSelect_io_fromSlowPorts_0_1_T; // @[ReservationStation.scala 697:68]
  wire [7:0] _dataSelect_io_fromSlowPorts_0_1_T_3 = dataArray_io_read_0_addr & dataArray_io_multiWrite_1_addr_1; // @[ReservationStation.scala 697:77]
  wire  _dataSelect_io_fromSlowPorts_0_1_T_5 = dataArray_io_multiWrite_1_enable & |_dataSelect_io_fromSlowPorts_0_1_T_3; // @[ReservationStation.scala 697:68]
  wire [7:0] _dataSelect_io_fromSlowPorts_0_1_T_6 = dataArray_io_read_0_addr & dataArray_io_multiWrite_2_addr_1; // @[ReservationStation.scala 697:77]
  wire  _dataSelect_io_fromSlowPorts_0_1_T_8 = dataArray_io_multiWrite_2_enable & |_dataSelect_io_fromSlowPorts_0_1_T_6; // @[ReservationStation.scala 697:68]
  wire [7:0] _dataSelect_io_fromSlowPorts_0_1_T_9 = dataArray_io_read_0_addr & dataArray_io_multiWrite_3_addr_1; // @[ReservationStation.scala 697:77]
  wire  _dataSelect_io_fromSlowPorts_0_1_T_11 = dataArray_io_multiWrite_3_enable & |_dataSelect_io_fromSlowPorts_0_1_T_9
    ; // @[ReservationStation.scala 697:68]
  wire [7:0] _dataSelect_io_fromSlowPorts_0_1_T_12 = dataArray_io_read_0_addr & dataArray_io_multiWrite_4_addr_1; // @[ReservationStation.scala 697:77]
  wire  _dataSelect_io_fromSlowPorts_0_1_T_14 = dataArray_io_multiWrite_4_enable & |
    _dataSelect_io_fromSlowPorts_0_1_T_12; // @[ReservationStation.scala 697:68]
  wire [1:0] dataSelect_io_fromSlowPorts_0_1_lo = {_dataSelect_io_fromSlowPorts_0_1_T_5,
    _dataSelect_io_fromSlowPorts_0_1_T_2}; // @[ReservationStation.scala 697:103]
  wire [2:0] dataSelect_io_fromSlowPorts_0_1_hi = {_dataSelect_io_fromSlowPorts_0_1_T_14,
    _dataSelect_io_fromSlowPorts_0_1_T_11,_dataSelect_io_fromSlowPorts_0_1_T_8}; // @[ReservationStation.scala 697:103]
  wire [7:0] _dataSelect_io_fromSlowPorts_1_0_T = dataArray_io_read_1_addr & dataArray_io_multiWrite_0_addr_0; // @[ReservationStation.scala 697:77]
  wire  _dataSelect_io_fromSlowPorts_1_0_T_2 = dataArray_io_multiWrite_0_enable & |_dataSelect_io_fromSlowPorts_1_0_T; // @[ReservationStation.scala 697:68]
  wire [7:0] _dataSelect_io_fromSlowPorts_1_0_T_3 = dataArray_io_read_1_addr & dataArray_io_multiWrite_1_addr_0; // @[ReservationStation.scala 697:77]
  wire  _dataSelect_io_fromSlowPorts_1_0_T_5 = dataArray_io_multiWrite_1_enable & |_dataSelect_io_fromSlowPorts_1_0_T_3; // @[ReservationStation.scala 697:68]
  wire [7:0] _dataSelect_io_fromSlowPorts_1_0_T_6 = dataArray_io_read_1_addr & dataArray_io_multiWrite_2_addr_0; // @[ReservationStation.scala 697:77]
  wire  _dataSelect_io_fromSlowPorts_1_0_T_8 = dataArray_io_multiWrite_2_enable & |_dataSelect_io_fromSlowPorts_1_0_T_6; // @[ReservationStation.scala 697:68]
  wire [7:0] _dataSelect_io_fromSlowPorts_1_0_T_9 = dataArray_io_read_1_addr & dataArray_io_multiWrite_3_addr_0; // @[ReservationStation.scala 697:77]
  wire  _dataSelect_io_fromSlowPorts_1_0_T_11 = dataArray_io_multiWrite_3_enable & |_dataSelect_io_fromSlowPorts_1_0_T_9
    ; // @[ReservationStation.scala 697:68]
  wire [7:0] _dataSelect_io_fromSlowPorts_1_0_T_12 = dataArray_io_read_1_addr & dataArray_io_multiWrite_4_addr_0; // @[ReservationStation.scala 697:77]
  wire  _dataSelect_io_fromSlowPorts_1_0_T_14 = dataArray_io_multiWrite_4_enable & |
    _dataSelect_io_fromSlowPorts_1_0_T_12; // @[ReservationStation.scala 697:68]
  wire [1:0] dataSelect_io_fromSlowPorts_1_0_lo = {_dataSelect_io_fromSlowPorts_1_0_T_5,
    _dataSelect_io_fromSlowPorts_1_0_T_2}; // @[ReservationStation.scala 697:103]
  wire [2:0] dataSelect_io_fromSlowPorts_1_0_hi = {_dataSelect_io_fromSlowPorts_1_0_T_14,
    _dataSelect_io_fromSlowPorts_1_0_T_11,_dataSelect_io_fromSlowPorts_1_0_T_8}; // @[ReservationStation.scala 697:103]
  wire [7:0] _dataSelect_io_fromSlowPorts_1_1_T = dataArray_io_read_1_addr & dataArray_io_multiWrite_0_addr_1; // @[ReservationStation.scala 697:77]
  wire  _dataSelect_io_fromSlowPorts_1_1_T_2 = dataArray_io_multiWrite_0_enable & |_dataSelect_io_fromSlowPorts_1_1_T; // @[ReservationStation.scala 697:68]
  wire [7:0] _dataSelect_io_fromSlowPorts_1_1_T_3 = dataArray_io_read_1_addr & dataArray_io_multiWrite_1_addr_1; // @[ReservationStation.scala 697:77]
  wire  _dataSelect_io_fromSlowPorts_1_1_T_5 = dataArray_io_multiWrite_1_enable & |_dataSelect_io_fromSlowPorts_1_1_T_3; // @[ReservationStation.scala 697:68]
  wire [7:0] _dataSelect_io_fromSlowPorts_1_1_T_6 = dataArray_io_read_1_addr & dataArray_io_multiWrite_2_addr_1; // @[ReservationStation.scala 697:77]
  wire  _dataSelect_io_fromSlowPorts_1_1_T_8 = dataArray_io_multiWrite_2_enable & |_dataSelect_io_fromSlowPorts_1_1_T_6; // @[ReservationStation.scala 697:68]
  wire [7:0] _dataSelect_io_fromSlowPorts_1_1_T_9 = dataArray_io_read_1_addr & dataArray_io_multiWrite_3_addr_1; // @[ReservationStation.scala 697:77]
  wire  _dataSelect_io_fromSlowPorts_1_1_T_11 = dataArray_io_multiWrite_3_enable & |_dataSelect_io_fromSlowPorts_1_1_T_9
    ; // @[ReservationStation.scala 697:68]
  wire [7:0] _dataSelect_io_fromSlowPorts_1_1_T_12 = dataArray_io_read_1_addr & dataArray_io_multiWrite_4_addr_1; // @[ReservationStation.scala 697:77]
  wire  _dataSelect_io_fromSlowPorts_1_1_T_14 = dataArray_io_multiWrite_4_enable & |
    _dataSelect_io_fromSlowPorts_1_1_T_12; // @[ReservationStation.scala 697:68]
  wire [1:0] dataSelect_io_fromSlowPorts_1_1_lo = {_dataSelect_io_fromSlowPorts_1_1_T_5,
    _dataSelect_io_fromSlowPorts_1_1_T_2}; // @[ReservationStation.scala 697:103]
  wire [2:0] dataSelect_io_fromSlowPorts_1_1_hi = {_dataSelect_io_fromSlowPorts_1_1_T_14,
    _dataSelect_io_fromSlowPorts_1_1_T_11,_dataSelect_io_fromSlowPorts_1_1_T_8}; // @[ReservationStation.scala 697:103]
  wire [7:0] _dataSelect_io_fromSlowPorts_2_0_T = dataArray_io_write_0_addr & dataArray_io_multiWrite_0_addr_0; // @[ReservationStation.scala 697:77]
  wire  _dataSelect_io_fromSlowPorts_2_0_T_2 = dataArray_io_multiWrite_0_enable & |_dataSelect_io_fromSlowPorts_2_0_T; // @[ReservationStation.scala 697:68]
  wire [7:0] _dataSelect_io_fromSlowPorts_2_0_T_3 = dataArray_io_write_0_addr & dataArray_io_multiWrite_1_addr_0; // @[ReservationStation.scala 697:77]
  wire  _dataSelect_io_fromSlowPorts_2_0_T_5 = dataArray_io_multiWrite_1_enable & |_dataSelect_io_fromSlowPorts_2_0_T_3; // @[ReservationStation.scala 697:68]
  wire [7:0] _dataSelect_io_fromSlowPorts_2_0_T_6 = dataArray_io_write_0_addr & dataArray_io_multiWrite_2_addr_0; // @[ReservationStation.scala 697:77]
  wire  _dataSelect_io_fromSlowPorts_2_0_T_8 = dataArray_io_multiWrite_2_enable & |_dataSelect_io_fromSlowPorts_2_0_T_6; // @[ReservationStation.scala 697:68]
  wire [7:0] _dataSelect_io_fromSlowPorts_2_0_T_9 = dataArray_io_write_0_addr & dataArray_io_multiWrite_3_addr_0; // @[ReservationStation.scala 697:77]
  wire  _dataSelect_io_fromSlowPorts_2_0_T_11 = dataArray_io_multiWrite_3_enable & |_dataSelect_io_fromSlowPorts_2_0_T_9
    ; // @[ReservationStation.scala 697:68]
  wire [7:0] _dataSelect_io_fromSlowPorts_2_0_T_12 = dataArray_io_write_0_addr & dataArray_io_multiWrite_4_addr_0; // @[ReservationStation.scala 697:77]
  wire  _dataSelect_io_fromSlowPorts_2_0_T_14 = dataArray_io_multiWrite_4_enable & |
    _dataSelect_io_fromSlowPorts_2_0_T_12; // @[ReservationStation.scala 697:68]
  wire [1:0] dataSelect_io_fromSlowPorts_2_0_lo = {_dataSelect_io_fromSlowPorts_2_0_T_5,
    _dataSelect_io_fromSlowPorts_2_0_T_2}; // @[ReservationStation.scala 697:103]
  wire [2:0] dataSelect_io_fromSlowPorts_2_0_hi = {_dataSelect_io_fromSlowPorts_2_0_T_14,
    _dataSelect_io_fromSlowPorts_2_0_T_11,_dataSelect_io_fromSlowPorts_2_0_T_8}; // @[ReservationStation.scala 697:103]
  wire [7:0] _dataSelect_io_fromSlowPorts_2_1_T = dataArray_io_write_0_addr & dataArray_io_multiWrite_0_addr_1; // @[ReservationStation.scala 697:77]
  wire  _dataSelect_io_fromSlowPorts_2_1_T_2 = dataArray_io_multiWrite_0_enable & |_dataSelect_io_fromSlowPorts_2_1_T; // @[ReservationStation.scala 697:68]
  wire [7:0] _dataSelect_io_fromSlowPorts_2_1_T_3 = dataArray_io_write_0_addr & dataArray_io_multiWrite_1_addr_1; // @[ReservationStation.scala 697:77]
  wire  _dataSelect_io_fromSlowPorts_2_1_T_5 = dataArray_io_multiWrite_1_enable & |_dataSelect_io_fromSlowPorts_2_1_T_3; // @[ReservationStation.scala 697:68]
  wire [7:0] _dataSelect_io_fromSlowPorts_2_1_T_6 = dataArray_io_write_0_addr & dataArray_io_multiWrite_2_addr_1; // @[ReservationStation.scala 697:77]
  wire  _dataSelect_io_fromSlowPorts_2_1_T_8 = dataArray_io_multiWrite_2_enable & |_dataSelect_io_fromSlowPorts_2_1_T_6; // @[ReservationStation.scala 697:68]
  wire [7:0] _dataSelect_io_fromSlowPorts_2_1_T_9 = dataArray_io_write_0_addr & dataArray_io_multiWrite_3_addr_1; // @[ReservationStation.scala 697:77]
  wire  _dataSelect_io_fromSlowPorts_2_1_T_11 = dataArray_io_multiWrite_3_enable & |_dataSelect_io_fromSlowPorts_2_1_T_9
    ; // @[ReservationStation.scala 697:68]
  wire [7:0] _dataSelect_io_fromSlowPorts_2_1_T_12 = dataArray_io_write_0_addr & dataArray_io_multiWrite_4_addr_1; // @[ReservationStation.scala 697:77]
  wire  _dataSelect_io_fromSlowPorts_2_1_T_14 = dataArray_io_multiWrite_4_enable & |
    _dataSelect_io_fromSlowPorts_2_1_T_12; // @[ReservationStation.scala 697:68]
  wire [1:0] dataSelect_io_fromSlowPorts_2_1_lo = {_dataSelect_io_fromSlowPorts_2_1_T_5,
    _dataSelect_io_fromSlowPorts_2_1_T_2}; // @[ReservationStation.scala 697:103]
  wire [2:0] dataSelect_io_fromSlowPorts_2_1_hi = {_dataSelect_io_fromSlowPorts_2_1_T_14,
    _dataSelect_io_fromSlowPorts_2_1_T_11,_dataSelect_io_fromSlowPorts_2_1_T_8}; // @[ReservationStation.scala 697:103]
  reg  fastWakeupMatch_0_0_0; // @[ReservationStation.scala 718:28]
  reg  fastWakeupMatch_0_1_0; // @[ReservationStation.scala 718:28]
  reg  fastWakeupMatch_1_0_0; // @[ReservationStation.scala 718:28]
  reg  fastWakeupMatch_1_1_0; // @[ReservationStation.scala 718:28]
  reg  fastWakeupMatch_2_0_0; // @[ReservationStation.scala 718:28]
  reg  fastWakeupMatch_2_1_0; // @[ReservationStation.scala 718:28]
  reg  fastWakeupMatch_3_0_0; // @[ReservationStation.scala 718:28]
  reg  fastWakeupMatch_3_1_0; // @[ReservationStation.scala 718:28]
  reg  fastWakeupMatch_4_0_0; // @[ReservationStation.scala 718:28]
  reg  fastWakeupMatch_4_1_0; // @[ReservationStation.scala 718:28]
  reg  fastWakeupMatch_5_0_0; // @[ReservationStation.scala 718:28]
  reg  fastWakeupMatch_5_1_0; // @[ReservationStation.scala 718:28]
  reg  fastWakeupMatch_6_0_0; // @[ReservationStation.scala 718:28]
  reg  fastWakeupMatch_6_1_0; // @[ReservationStation.scala 718:28]
  reg  fastWakeupMatch_7_0_0; // @[ReservationStation.scala 718:28]
  reg  fastWakeupMatch_7_1_0; // @[ReservationStation.scala 718:28]
  wire  s1_out_fire_0 = s1_out_0_valid & s2_deq_0_ready; // @[ReservationStation.scala 728:60]
  reg  data_uop_robIdx_flag; // @[Reg.scala 16:16]
  reg [4:0] data_uop_robIdx_value; // @[Reg.scala 16:16]
  wire [5:0] _flushItself_T_1 = {data_uop_robIdx_flag,data_uop_robIdx_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_3 = _flushItself_T_1 == _s1_out_0_valid_flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself = io_redirect_bits_level & _flushItself_T_3; // @[Rob.scala 122:51]
  wire  differentFlag = data_uop_robIdx_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare = data_uop_robIdx_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_134 = differentFlag ^ compare; // @[CircularQueuePtr.scala 88:19]
  wire  _T_136 = io_redirect_valid & (flushItself | _T_134); // @[Rob.scala 123:20]
  wire  _T_137 = s2_deq_0_ready | _T_136; // @[ReservationStation.scala 736:59]
  wire  _GEN_657 = _T_137 ? 1'h0 : valid; // @[PipelineConnect.scala 108:24 110:{25,33}]
  reg [3:0] data_uop_ctrl_fuType; // @[Reg.scala 16:16]
  reg [6:0] data_uop_ctrl_fuOpType; // @[Reg.scala 16:16]
  reg  data_uop_ctrl_rfWen; // @[Reg.scala 16:16]
  reg  data_uop_ctrl_fpWen; // @[Reg.scala 16:16]
  reg [5:0] data_uop_pdest; // @[Reg.scala 16:16]
  wire [7:0] normalIssuePtrOH = s1_issue_oldest_0 ? s1_in_oldestPtrOH_bits : select_io_grant_0_bits; // @[ReservationStation.scala 756:33]
  wire  normalFastWakeupMatch_0_0 = normalIssuePtrOH[0] & fastWakeupMatch_0_0_0 | normalIssuePtrOH[1] &
    fastWakeupMatch_1_0_0 | normalIssuePtrOH[2] & fastWakeupMatch_2_0_0 | normalIssuePtrOH[3] & fastWakeupMatch_3_0_0 |
    normalIssuePtrOH[4] & fastWakeupMatch_4_0_0 | normalIssuePtrOH[5] & fastWakeupMatch_5_0_0 | normalIssuePtrOH[6] &
    fastWakeupMatch_6_0_0 | normalIssuePtrOH[7] & fastWakeupMatch_7_0_0; // @[Mux.scala 27:73]
  wire  normalFastWakeupMatch_1_0 = normalIssuePtrOH[0] & fastWakeupMatch_0_1_0 | normalIssuePtrOH[1] &
    fastWakeupMatch_1_1_0 | normalIssuePtrOH[2] & fastWakeupMatch_2_1_0 | normalIssuePtrOH[3] & fastWakeupMatch_3_1_0 |
    normalIssuePtrOH[4] & fastWakeupMatch_4_1_0 | normalIssuePtrOH[5] & fastWakeupMatch_5_1_0 | normalIssuePtrOH[6] &
    fastWakeupMatch_6_1_0 | normalIssuePtrOH[7] & fastWakeupMatch_7_1_0; // @[Mux.scala 27:73]
  reg  io_perf_0_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg  io_perf_0_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  StatusArray_1 statusArray ( // @[ReservationStation.scala 261:27]
    .clock(statusArray_clock),
    .reset(statusArray_reset),
    .io_redirect_valid(statusArray_io_redirect_valid),
    .io_redirect_bits_robIdx_flag(statusArray_io_redirect_bits_robIdx_flag),
    .io_redirect_bits_robIdx_value(statusArray_io_redirect_bits_robIdx_value),
    .io_redirect_bits_level(statusArray_io_redirect_bits_level),
    .io_isValid(statusArray_io_isValid),
    .io_isValidNext(statusArray_io_isValidNext),
    .io_canIssue(statusArray_io_canIssue),
    .io_flushed(statusArray_io_flushed),
    .io_update_0_enable(statusArray_io_update_0_enable),
    .io_update_0_addr(statusArray_io_update_0_addr),
    .io_update_0_data_srcState_0(statusArray_io_update_0_data_srcState_0),
    .io_update_0_data_srcState_1(statusArray_io_update_0_data_srcState_1),
    .io_update_0_data_psrc_0(statusArray_io_update_0_data_psrc_0),
    .io_update_0_data_psrc_1(statusArray_io_update_0_data_psrc_1),
    .io_update_0_data_srcType_0(statusArray_io_update_0_data_srcType_0),
    .io_update_0_data_srcType_1(statusArray_io_update_0_data_srcType_1),
    .io_update_0_data_robIdx_flag(statusArray_io_update_0_data_robIdx_flag),
    .io_update_0_data_robIdx_value(statusArray_io_update_0_data_robIdx_value),
    .io_update_1_enable(statusArray_io_update_1_enable),
    .io_update_1_addr(statusArray_io_update_1_addr),
    .io_update_1_data_srcState_0(statusArray_io_update_1_data_srcState_0),
    .io_update_1_data_srcState_1(statusArray_io_update_1_data_srcState_1),
    .io_update_1_data_psrc_0(statusArray_io_update_1_data_psrc_0),
    .io_update_1_data_psrc_1(statusArray_io_update_1_data_psrc_1),
    .io_update_1_data_srcType_0(statusArray_io_update_1_data_srcType_0),
    .io_update_1_data_srcType_1(statusArray_io_update_1_data_srcType_1),
    .io_update_1_data_robIdx_flag(statusArray_io_update_1_data_robIdx_flag),
    .io_update_1_data_robIdx_value(statusArray_io_update_1_data_robIdx_value),
    .io_wakeup_0_valid(statusArray_io_wakeup_0_valid),
    .io_wakeup_0_bits_ctrl_rfWen(statusArray_io_wakeup_0_bits_ctrl_rfWen),
    .io_wakeup_0_bits_pdest(statusArray_io_wakeup_0_bits_pdest),
    .io_wakeup_1_valid(statusArray_io_wakeup_1_valid),
    .io_wakeup_1_bits_ctrl_rfWen(statusArray_io_wakeup_1_bits_ctrl_rfWen),
    .io_wakeup_1_bits_pdest(statusArray_io_wakeup_1_bits_pdest),
    .io_wakeup_2_valid(statusArray_io_wakeup_2_valid),
    .io_wakeup_2_bits_ctrl_rfWen(statusArray_io_wakeup_2_bits_ctrl_rfWen),
    .io_wakeup_2_bits_pdest(statusArray_io_wakeup_2_bits_pdest),
    .io_wakeup_3_valid(statusArray_io_wakeup_3_valid),
    .io_wakeup_3_bits_ctrl_rfWen(statusArray_io_wakeup_3_bits_ctrl_rfWen),
    .io_wakeup_3_bits_pdest(statusArray_io_wakeup_3_bits_pdest),
    .io_wakeup_4_valid(statusArray_io_wakeup_4_valid),
    .io_wakeup_4_bits_ctrl_rfWen(statusArray_io_wakeup_4_bits_ctrl_rfWen),
    .io_wakeup_4_bits_pdest(statusArray_io_wakeup_4_bits_pdest),
    .io_wakeup_5_valid(statusArray_io_wakeup_5_valid),
    .io_wakeup_5_bits_ctrl_rfWen(statusArray_io_wakeup_5_bits_ctrl_rfWen),
    .io_wakeup_5_bits_pdest(statusArray_io_wakeup_5_bits_pdest),
    .io_wakeupMatch_0_0(statusArray_io_wakeupMatch_0_0),
    .io_wakeupMatch_0_1(statusArray_io_wakeupMatch_0_1),
    .io_wakeupMatch_1_0(statusArray_io_wakeupMatch_1_0),
    .io_wakeupMatch_1_1(statusArray_io_wakeupMatch_1_1),
    .io_wakeupMatch_2_0(statusArray_io_wakeupMatch_2_0),
    .io_wakeupMatch_2_1(statusArray_io_wakeupMatch_2_1),
    .io_wakeupMatch_3_0(statusArray_io_wakeupMatch_3_0),
    .io_wakeupMatch_3_1(statusArray_io_wakeupMatch_3_1),
    .io_wakeupMatch_4_0(statusArray_io_wakeupMatch_4_0),
    .io_wakeupMatch_4_1(statusArray_io_wakeupMatch_4_1),
    .io_wakeupMatch_5_0(statusArray_io_wakeupMatch_5_0),
    .io_wakeupMatch_5_1(statusArray_io_wakeupMatch_5_1),
    .io_wakeupMatch_6_0(statusArray_io_wakeupMatch_6_0),
    .io_wakeupMatch_6_1(statusArray_io_wakeupMatch_6_1),
    .io_wakeupMatch_7_0(statusArray_io_wakeupMatch_7_0),
    .io_wakeupMatch_7_1(statusArray_io_wakeupMatch_7_1),
    .io_deqResp_0_valid(statusArray_io_deqResp_0_valid),
    .io_deqResp_0_bits_rsMask(statusArray_io_deqResp_0_bits_rsMask),
    .io_deqResp_0_bits_success(statusArray_io_deqResp_0_bits_success),
    .io_deqResp_1_valid(statusArray_io_deqResp_1_valid),
    .io_deqResp_1_bits_rsMask(statusArray_io_deqResp_1_bits_rsMask),
    .io_deqResp_1_bits_success(statusArray_io_deqResp_1_bits_success),
    .io_deqResp_2_valid(statusArray_io_deqResp_2_valid),
    .io_deqResp_2_bits_rsMask(statusArray_io_deqResp_2_bits_rsMask),
    .io_deqResp_2_bits_success(statusArray_io_deqResp_2_bits_success)
  );
  SelectPolicy_1 select ( // @[ReservationStation.scala 262:22]
    .io_validVec(select_io_validVec),
    .io_allocate_0_bits(select_io_allocate_0_bits),
    .io_allocate_1_bits(select_io_allocate_1_bits),
    .io_request(select_io_request),
    .io_grant_0_valid(select_io_grant_0_valid),
    .io_grant_0_bits(select_io_grant_0_bits)
  );
  DataArray_1 dataArray ( // @[ReservationStation.scala 263:25]
    .clock(dataArray_clock),
    .io_read_0_addr(dataArray_io_read_0_addr),
    .io_read_0_data_0(dataArray_io_read_0_data_0),
    .io_read_0_data_1(dataArray_io_read_0_data_1),
    .io_read_1_addr(dataArray_io_read_1_addr),
    .io_read_1_data_0(dataArray_io_read_1_data_0),
    .io_read_1_data_1(dataArray_io_read_1_data_1),
    .io_write_0_enable(dataArray_io_write_0_enable),
    .io_write_0_mask_0(dataArray_io_write_0_mask_0),
    .io_write_0_mask_1(dataArray_io_write_0_mask_1),
    .io_write_0_addr(dataArray_io_write_0_addr),
    .io_write_0_data_0(dataArray_io_write_0_data_0),
    .io_write_0_data_1(dataArray_io_write_0_data_1),
    .io_write_1_enable(dataArray_io_write_1_enable),
    .io_write_1_mask_0(dataArray_io_write_1_mask_0),
    .io_write_1_mask_1(dataArray_io_write_1_mask_1),
    .io_write_1_addr(dataArray_io_write_1_addr),
    .io_write_1_data_0(dataArray_io_write_1_data_0),
    .io_write_1_data_1(dataArray_io_write_1_data_1),
    .io_multiWrite_0_enable(dataArray_io_multiWrite_0_enable),
    .io_multiWrite_0_addr_0(dataArray_io_multiWrite_0_addr_0),
    .io_multiWrite_0_addr_1(dataArray_io_multiWrite_0_addr_1),
    .io_multiWrite_0_data(dataArray_io_multiWrite_0_data),
    .io_multiWrite_1_enable(dataArray_io_multiWrite_1_enable),
    .io_multiWrite_1_addr_0(dataArray_io_multiWrite_1_addr_0),
    .io_multiWrite_1_addr_1(dataArray_io_multiWrite_1_addr_1),
    .io_multiWrite_1_data(dataArray_io_multiWrite_1_data),
    .io_multiWrite_2_enable(dataArray_io_multiWrite_2_enable),
    .io_multiWrite_2_addr_0(dataArray_io_multiWrite_2_addr_0),
    .io_multiWrite_2_addr_1(dataArray_io_multiWrite_2_addr_1),
    .io_multiWrite_2_data(dataArray_io_multiWrite_2_data),
    .io_multiWrite_3_enable(dataArray_io_multiWrite_3_enable),
    .io_multiWrite_3_addr_0(dataArray_io_multiWrite_3_addr_0),
    .io_multiWrite_3_addr_1(dataArray_io_multiWrite_3_addr_1),
    .io_multiWrite_3_data(dataArray_io_multiWrite_3_data),
    .io_multiWrite_4_enable(dataArray_io_multiWrite_4_enable),
    .io_multiWrite_4_addr_0(dataArray_io_multiWrite_4_addr_0),
    .io_multiWrite_4_addr_1(dataArray_io_multiWrite_4_addr_1),
    .io_multiWrite_4_data(dataArray_io_multiWrite_4_data)
  );
  PayloadArray_1 payloadArray ( // @[ReservationStation.scala 264:28]
    .clock(payloadArray_clock),
    .io_read_0_addr(payloadArray_io_read_0_addr),
    .io_read_0_data_ctrl_fuType(payloadArray_io_read_0_data_ctrl_fuType),
    .io_read_0_data_ctrl_fuOpType(payloadArray_io_read_0_data_ctrl_fuOpType),
    .io_read_0_data_ctrl_rfWen(payloadArray_io_read_0_data_ctrl_rfWen),
    .io_read_0_data_ctrl_fpWen(payloadArray_io_read_0_data_ctrl_fpWen),
    .io_read_0_data_pdest(payloadArray_io_read_0_data_pdest),
    .io_read_0_data_robIdx_flag(payloadArray_io_read_0_data_robIdx_flag),
    .io_read_0_data_robIdx_value(payloadArray_io_read_0_data_robIdx_value),
    .io_read_1_addr(payloadArray_io_read_1_addr),
    .io_read_1_data_ctrl_fuType(payloadArray_io_read_1_data_ctrl_fuType),
    .io_read_1_data_ctrl_fuOpType(payloadArray_io_read_1_data_ctrl_fuOpType),
    .io_read_1_data_ctrl_rfWen(payloadArray_io_read_1_data_ctrl_rfWen),
    .io_read_1_data_ctrl_fpWen(payloadArray_io_read_1_data_ctrl_fpWen),
    .io_read_1_data_pdest(payloadArray_io_read_1_data_pdest),
    .io_read_1_data_robIdx_flag(payloadArray_io_read_1_data_robIdx_flag),
    .io_read_1_data_robIdx_value(payloadArray_io_read_1_data_robIdx_value),
    .io_write_0_enable(payloadArray_io_write_0_enable),
    .io_write_0_addr(payloadArray_io_write_0_addr),
    .io_write_0_data_ctrl_fuType(payloadArray_io_write_0_data_ctrl_fuType),
    .io_write_0_data_ctrl_fuOpType(payloadArray_io_write_0_data_ctrl_fuOpType),
    .io_write_0_data_ctrl_rfWen(payloadArray_io_write_0_data_ctrl_rfWen),
    .io_write_0_data_ctrl_fpWen(payloadArray_io_write_0_data_ctrl_fpWen),
    .io_write_0_data_pdest(payloadArray_io_write_0_data_pdest),
    .io_write_0_data_robIdx_flag(payloadArray_io_write_0_data_robIdx_flag),
    .io_write_0_data_robIdx_value(payloadArray_io_write_0_data_robIdx_value),
    .io_write_1_enable(payloadArray_io_write_1_enable),
    .io_write_1_addr(payloadArray_io_write_1_addr),
    .io_write_1_data_ctrl_fuType(payloadArray_io_write_1_data_ctrl_fuType),
    .io_write_1_data_ctrl_fuOpType(payloadArray_io_write_1_data_ctrl_fuOpType),
    .io_write_1_data_ctrl_rfWen(payloadArray_io_write_1_data_ctrl_rfWen),
    .io_write_1_data_ctrl_fpWen(payloadArray_io_write_1_data_ctrl_fpWen),
    .io_write_1_data_pdest(payloadArray_io_write_1_data_pdest),
    .io_write_1_data_robIdx_flag(payloadArray_io_write_1_data_robIdx_flag),
    .io_write_1_data_robIdx_value(payloadArray_io_write_1_data_robIdx_value)
  );
  AgeDetector_1 s1_oldestSel_age ( // @[SelectPolicy.scala 174:21]
    .clock(s1_oldestSel_age_clock),
    .reset(s1_oldestSel_age_reset),
    .io_enq_0(s1_oldestSel_age_io_enq_0),
    .io_enq_1(s1_oldestSel_age_io_enq_1),
    .io_deq(s1_oldestSel_age_io_deq),
    .io_out(s1_oldestSel_age_io_out)
  );
  OldestSelection_1 oldestSelection ( // @[ReservationStation.scala 499:33]
    .io_oldest_valid(oldestSelection_io_oldest_valid),
    .io_isOverrided_0(oldestSelection_io_isOverrided_0)
  );
  WakeupQueue_2 wakeupQueue ( // @[ReservationStation.scala 564:31]
    .clock(wakeupQueue_clock),
    .reset(wakeupQueue_reset),
    .io_in_valid(wakeupQueue_io_in_valid),
    .io_in_bits_ctrl_rfWen(wakeupQueue_io_in_bits_ctrl_rfWen),
    .io_in_bits_pdest(wakeupQueue_io_in_bits_pdest),
    .io_in_bits_robIdx_flag(wakeupQueue_io_in_bits_robIdx_flag),
    .io_in_bits_robIdx_value(wakeupQueue_io_in_bits_robIdx_value),
    .io_out_valid(wakeupQueue_io_out_valid),
    .io_out_bits_ctrl_rfWen(wakeupQueue_io_out_bits_ctrl_rfWen),
    .io_out_bits_pdest(wakeupQueue_io_out_bits_pdest),
    .io_redirect_valid(wakeupQueue_io_redirect_valid),
    .io_redirect_bits_robIdx_flag(wakeupQueue_io_redirect_bits_robIdx_flag),
    .io_redirect_bits_robIdx_value(wakeupQueue_io_redirect_bits_robIdx_value),
    .io_redirect_bits_level(wakeupQueue_io_redirect_bits_level)
  );
  MduImmExtractor immExt ( // @[DataArray.scala 159:36]
    .io_uop_ctrl_srcType_1(immExt_io_uop_ctrl_srcType_1),
    .io_uop_ctrl_imm(immExt_io_uop_ctrl_imm),
    .io_data_in_0(immExt_io_data_in_0),
    .io_data_in_1(immExt_io_data_in_1),
    .io_data_out_0(immExt_io_data_out_0),
    .io_data_out_1(immExt_io_data_out_1)
  );
  MduImmExtractor immExt_1 ( // @[DataArray.scala 159:36]
    .io_uop_ctrl_srcType_1(immExt_1_io_uop_ctrl_srcType_1),
    .io_uop_ctrl_imm(immExt_1_io_uop_ctrl_imm),
    .io_data_in_0(immExt_1_io_data_in_0),
    .io_data_in_1(immExt_1_io_data_in_1),
    .io_data_out_0(immExt_1_io_data_out_0),
    .io_data_out_1(immExt_1_io_data_out_1)
  );
  DataSelect_1 dataSelect ( // @[ReservationStation.scala 691:26]
    .io_doOverride_0(dataSelect_io_doOverride_0),
    .io_readData_0_0(dataSelect_io_readData_0_0),
    .io_readData_0_1(dataSelect_io_readData_0_1),
    .io_readData_1_0(dataSelect_io_readData_1_0),
    .io_readData_1_1(dataSelect_io_readData_1_1),
    .io_fromSlowPorts_0_0(dataSelect_io_fromSlowPorts_0_0),
    .io_fromSlowPorts_0_1(dataSelect_io_fromSlowPorts_0_1),
    .io_fromSlowPorts_1_0(dataSelect_io_fromSlowPorts_1_0),
    .io_fromSlowPorts_1_1(dataSelect_io_fromSlowPorts_1_1),
    .io_fromSlowPorts_2_0(dataSelect_io_fromSlowPorts_2_0),
    .io_fromSlowPorts_2_1(dataSelect_io_fromSlowPorts_2_1),
    .io_slowData_0(dataSelect_io_slowData_0),
    .io_slowData_1(dataSelect_io_slowData_1),
    .io_slowData_2(dataSelect_io_slowData_2),
    .io_slowData_3(dataSelect_io_slowData_3),
    .io_slowData_4(dataSelect_io_slowData_4),
    .io_enqBypass_0_0(dataSelect_io_enqBypass_0_0),
    .io_enqData_0_0_bits(dataSelect_io_enqData_0_0_bits),
    .io_enqData_0_1_bits(dataSelect_io_enqData_0_1_bits),
    .io_deqData_0_0(dataSelect_io_deqData_0_0),
    .io_deqData_0_1(dataSelect_io_deqData_0_1)
  );
  BypassNetworkLeft_2 bypassNetwork ( // @[BypassNetwork.scala 111:13]
    .clock(bypassNetwork_clock),
    .io_hold(bypassNetwork_io_hold),
    .io_source_0(bypassNetwork_io_source_0),
    .io_source_1(bypassNetwork_io_source_1),
    .io_target_0(bypassNetwork_io_target_0),
    .io_target_1(bypassNetwork_io_target_1),
    .io_bypass_0_valid_0(bypassNetwork_io_bypass_0_valid_0),
    .io_bypass_0_valid_1(bypassNetwork_io_bypass_0_valid_1),
    .io_bypass_0_data(bypassNetwork_io_bypass_0_data)
  );
  assign io_fromDispatch_0_ready = emptyThisCycle > _GEN_774; // @[ReservationStation.scala 324:42]
  assign io_fromDispatch_1_ready = emptyThisCycle > _GEN_775; // @[ReservationStation.scala 324:42]
  assign io_deq_0_valid = valid; // @[PipelineConnect.scala 117:17 ReservationStation.scala 266:20]
  assign io_deq_0_bits_uop_ctrl_fuType = data_uop_ctrl_fuType; // @[PipelineConnect.scala 116:16 ReservationStation.scala 266:20]
  assign io_deq_0_bits_uop_ctrl_fuOpType = data_uop_ctrl_fuOpType; // @[PipelineConnect.scala 116:16 ReservationStation.scala 266:20]
  assign io_deq_0_bits_uop_ctrl_rfWen = data_uop_ctrl_rfWen; // @[PipelineConnect.scala 116:16 ReservationStation.scala 266:20]
  assign io_deq_0_bits_uop_ctrl_fpWen = data_uop_ctrl_fpWen; // @[PipelineConnect.scala 116:16 ReservationStation.scala 266:20]
  assign io_deq_0_bits_uop_pdest = data_uop_pdest; // @[PipelineConnect.scala 116:16 ReservationStation.scala 266:20]
  assign io_deq_0_bits_uop_robIdx_flag = data_uop_robIdx_flag; // @[PipelineConnect.scala 116:16 ReservationStation.scala 266:20]
  assign io_deq_0_bits_uop_robIdx_value = data_uop_robIdx_value; // @[PipelineConnect.scala 116:16 ReservationStation.scala 266:20]
  assign io_deq_0_bits_src_0 = bypassNetwork_io_target_0; // @[ReservationStation.scala 266:20 772:31]
  assign io_deq_0_bits_src_1 = bypassNetwork_io_target_1; // @[ReservationStation.scala 266:20 772:31]
  assign io_fastWakeup_0_valid = wakeupQueue_io_out_valid; // @[ReservationStation.scala 571:28]
  assign io_fastWakeup_0_bits_ctrl_rfWen = wakeupQueue_io_out_bits_ctrl_rfWen; // @[ReservationStation.scala 571:28]
  assign io_fastWakeup_0_bits_pdest = wakeupQueue_io_out_bits_pdest; // @[ReservationStation.scala 571:28]
  assign io_perf_0_value = {{5'd0}, io_perf_0_value_REG_1}; // @[PerfCounterUtils.scala 188:17]
  assign statusArray_clock = clock;
  assign statusArray_reset = reset;
  assign statusArray_io_redirect_valid = io_redirect_valid; // @[ReservationStation.scala 437:27]
  assign statusArray_io_redirect_bits_robIdx_flag = io_redirect_bits_robIdx_flag; // @[ReservationStation.scala 437:27]
  assign statusArray_io_redirect_bits_robIdx_value = io_redirect_bits_robIdx_value; // @[ReservationStation.scala 437:27]
  assign statusArray_io_redirect_bits_level = io_redirect_bits_level; // @[ReservationStation.scala 437:27]
  assign statusArray_io_update_0_enable = s1_dispatchUops_dup_0_0_valid; // @[ReservationStation.scala 445:25]
  assign statusArray_io_update_0_addr = s1_allocatePtrOH_dup_0_0; // @[ReservationStation.scala 446:23]
  assign statusArray_io_update_0_data_srcState_0 = _statusArray_io_update_0_data_srcState_0_T_2 | |s1_enqWakeup_0_0 | |
    s1_fastWakeup_0_0_0; // @[ReservationStation.scala 452:96]
  assign statusArray_io_update_0_data_srcState_1 = _statusArray_io_update_0_data_srcState_0_T_5 | |s1_enqWakeup_0_1 | |
    s1_fastWakeup_0_1_0; // @[ReservationStation.scala 452:96]
  assign statusArray_io_update_0_data_psrc_0 = s1_dispatchUops_dup_0_0_bits_psrc_0; // @[ReservationStation.scala 455:28]
  assign statusArray_io_update_0_data_psrc_1 = s1_dispatchUops_dup_0_0_bits_psrc_1; // @[ReservationStation.scala 455:28]
  assign statusArray_io_update_0_data_srcType_0 = s1_dispatchUops_dup_0_0_bits_ctrl_srcType_0; // @[ReservationStation.scala 456:31]
  assign statusArray_io_update_0_data_srcType_1 = s1_dispatchUops_dup_0_0_bits_ctrl_srcType_1; // @[ReservationStation.scala 456:31]
  assign statusArray_io_update_0_data_robIdx_flag = s1_dispatchUops_dup_0_0_bits_robIdx_flag; // @[ReservationStation.scala 457:30]
  assign statusArray_io_update_0_data_robIdx_value = s1_dispatchUops_dup_0_0_bits_robIdx_value; // @[ReservationStation.scala 457:30]
  assign statusArray_io_update_1_enable = s1_dispatchUops_dup_0_1_valid; // @[ReservationStation.scala 445:25]
  assign statusArray_io_update_1_addr = s1_allocatePtrOH_dup_0_1; // @[ReservationStation.scala 446:23]
  assign statusArray_io_update_1_data_srcState_0 = _statusArray_io_update_1_data_srcState_0_T_2 | |s1_enqWakeup_1_0 | |
    s1_fastWakeup_1_0_0; // @[ReservationStation.scala 452:96]
  assign statusArray_io_update_1_data_srcState_1 = _statusArray_io_update_1_data_srcState_0_T_5 | |s1_enqWakeup_1_1 | |
    s1_fastWakeup_1_1_0; // @[ReservationStation.scala 452:96]
  assign statusArray_io_update_1_data_psrc_0 = s1_dispatchUops_dup_0_1_bits_psrc_0; // @[ReservationStation.scala 455:28]
  assign statusArray_io_update_1_data_psrc_1 = s1_dispatchUops_dup_0_1_bits_psrc_1; // @[ReservationStation.scala 455:28]
  assign statusArray_io_update_1_data_srcType_0 = s1_dispatchUops_dup_0_1_bits_ctrl_srcType_0; // @[ReservationStation.scala 456:31]
  assign statusArray_io_update_1_data_srcType_1 = s1_dispatchUops_dup_0_1_bits_ctrl_srcType_1; // @[ReservationStation.scala 456:31]
  assign statusArray_io_update_1_data_robIdx_flag = s1_dispatchUops_dup_0_1_bits_robIdx_flag; // @[ReservationStation.scala 457:30]
  assign statusArray_io_update_1_data_robIdx_value = s1_dispatchUops_dup_0_1_bits_robIdx_value; // @[ReservationStation.scala 457:30]
  assign statusArray_io_wakeup_0_valid = io_fastUopsIn_0_valid; // @[ReservationStation.scala 352:18]
  assign statusArray_io_wakeup_0_bits_ctrl_rfWen = io_fastUopsIn_0_bits_ctrl_rfWen; // @[ReservationStation.scala 353:17]
  assign statusArray_io_wakeup_0_bits_pdest = io_fastUopsIn_0_bits_pdest; // @[ReservationStation.scala 353:17]
  assign statusArray_io_wakeup_1_valid = io_slowPorts_0_valid; // @[ReservationStation.scala 352:18]
  assign statusArray_io_wakeup_1_bits_ctrl_rfWen = io_slowPorts_0_bits_uop_ctrl_rfWen; // @[ReservationStation.scala 353:17]
  assign statusArray_io_wakeup_1_bits_pdest = io_slowPorts_0_bits_uop_pdest; // @[ReservationStation.scala 353:17]
  assign statusArray_io_wakeup_2_valid = io_slowPorts_1_valid; // @[ReservationStation.scala 352:18]
  assign statusArray_io_wakeup_2_bits_ctrl_rfWen = io_slowPorts_1_bits_uop_ctrl_rfWen; // @[ReservationStation.scala 353:17]
  assign statusArray_io_wakeup_2_bits_pdest = io_slowPorts_1_bits_uop_pdest; // @[ReservationStation.scala 353:17]
  assign statusArray_io_wakeup_3_valid = io_slowPorts_2_valid; // @[ReservationStation.scala 352:18]
  assign statusArray_io_wakeup_3_bits_ctrl_rfWen = io_slowPorts_2_bits_uop_ctrl_rfWen; // @[ReservationStation.scala 353:17]
  assign statusArray_io_wakeup_3_bits_pdest = io_slowPorts_2_bits_uop_pdest; // @[ReservationStation.scala 353:17]
  assign statusArray_io_wakeup_4_valid = io_slowPorts_3_valid; // @[ReservationStation.scala 352:18]
  assign statusArray_io_wakeup_4_bits_ctrl_rfWen = io_slowPorts_3_bits_uop_ctrl_rfWen; // @[ReservationStation.scala 353:17]
  assign statusArray_io_wakeup_4_bits_pdest = io_slowPorts_3_bits_uop_pdest; // @[ReservationStation.scala 353:17]
  assign statusArray_io_wakeup_5_valid = io_slowPorts_4_valid; // @[ReservationStation.scala 352:18]
  assign statusArray_io_wakeup_5_bits_ctrl_rfWen = io_slowPorts_4_bits_uop_ctrl_rfWen; // @[ReservationStation.scala 353:17]
  assign statusArray_io_wakeup_5_bits_pdest = io_slowPorts_4_bits_uop_pdest; // @[ReservationStation.scala 353:17]
  assign statusArray_io_deqResp_0_valid = _statusArray_io_issueGranted_2_valid_T_1 & s2_deq_0_ready; // @[ReservationStation.scala 550:91]
  assign statusArray_io_deqResp_0_bits_rsMask = select_io_grant_0_bits; // @[ReservationStation.scala 551:47]
  assign statusArray_io_deqResp_0_bits_success = ~valid | io_deq_0_ready; // @[ReservationStation.scala 747:41]
  assign statusArray_io_deqResp_1_valid = s1_issue_dispatch_0 & s2_deq_0_ready; // @[ReservationStation.scala 556:67]
  assign statusArray_io_deqResp_1_bits_rsMask = s1_allocatePtrOH_dup_0_0; // @[ReservationStation.scala 557:49]
  assign statusArray_io_deqResp_1_bits_success = ~valid | io_deq_0_ready; // @[ReservationStation.scala 747:41]
  assign statusArray_io_deqResp_2_valid = |s1_issue_oldest_0 & statusArray_io_issueGranted_3_valid_xs_0; // @[ReservationStation.scala 577:69]
  assign statusArray_io_deqResp_2_bits_rsMask = s1_oldestSel_age_io_out; // @[SelectPolicy.scala 177:19 179:14]
  assign statusArray_io_deqResp_2_bits_success = s1_issue_oldest_0 & s2_deq_0_ready; // @[ParallelMux.scala 64:44]
  assign select_io_validVec = validAfterAllocate; // @[ReservationStation.scala 285:22]
  assign select_io_request = statusArray_io_canIssue; // @[ReservationStation.scala 358:21]
  assign dataArray_clock = clock;
  assign dataArray_io_read_0_addr = select_io_grant_0_bits; // @[ReservationStation.scala 376:31]
  assign dataArray_io_read_1_addr = s1_oldestSel_age_io_out; // @[SelectPolicy.scala 177:19 179:14]
  assign dataArray_io_write_0_enable = s1_dispatchUops_dup_2_0_valid; // @[ReservationStation.scala 603:34]
  assign dataArray_io_write_0_mask_0 = s1_dispatchUops_dup_2_0_bits_ctrl_srcType_0[0] |
    s1_dispatchUops_dup_2_0_bits_srcState_0; // @[Bundle.scala 245:81]
  assign dataArray_io_write_0_mask_1 = s1_dispatchUops_dup_2_0_bits_ctrl_srcType_1[0] |
    s1_dispatchUops_dup_2_0_bits_srcState_1; // @[Bundle.scala 245:81]
  assign dataArray_io_write_0_addr = s1_allocatePtrOH_dup_2_0; // @[ReservationStation.scala 605:32]
  assign dataArray_io_write_0_data_0 = immExt_io_data_out_0; // @[ReservationStation.scala 589:29 593:12]
  assign dataArray_io_write_0_data_1 = immExt_io_data_out_1; // @[ReservationStation.scala 589:29 593:12]
  assign dataArray_io_write_1_enable = s1_dispatchUops_dup_2_1_valid; // @[ReservationStation.scala 603:34]
  assign dataArray_io_write_1_mask_0 = s1_dispatchUops_dup_2_1_bits_ctrl_srcType_0[0] |
    s1_dispatchUops_dup_2_1_bits_srcState_0; // @[Bundle.scala 245:81]
  assign dataArray_io_write_1_mask_1 = s1_dispatchUops_dup_2_1_bits_ctrl_srcType_1[0] |
    s1_dispatchUops_dup_2_1_bits_srcState_1; // @[Bundle.scala 245:81]
  assign dataArray_io_write_1_addr = s1_allocatePtrOH_dup_2_1; // @[ReservationStation.scala 605:32]
  assign dataArray_io_write_1_data_0 = immExt_1_io_data_out_0; // @[ReservationStation.scala 589:29 593:12]
  assign dataArray_io_write_1_data_1 = immExt_1_io_data_out_1; // @[ReservationStation.scala 589:29 593:12]
  assign dataArray_io_multiWrite_0_enable = dataArray_io_multiWrite_0_enable_REG; // @[ReservationStation.scala 633:14]
  assign dataArray_io_multiWrite_0_addr_0 = _dataArray_io_multiWrite_0_addr_0_T_8 | allocateDataCapture; // @[ReservationStation.scala 637:68]
  assign dataArray_io_multiWrite_0_addr_1 = _dataArray_io_multiWrite_0_addr_1_T_8 | allocateDataCapture_1; // @[ReservationStation.scala 637:68]
  assign dataArray_io_multiWrite_0_data = dataArray_io_multiWrite_0_data_r; // @[ReservationStation.scala 639:12]
  assign dataArray_io_multiWrite_1_enable = dataArray_io_multiWrite_1_enable_REG; // @[ReservationStation.scala 633:14]
  assign dataArray_io_multiWrite_1_addr_0 = _dataArray_io_multiWrite_1_addr_0_T_8 | allocateDataCapture_2; // @[ReservationStation.scala 637:68]
  assign dataArray_io_multiWrite_1_addr_1 = _dataArray_io_multiWrite_1_addr_1_T_8 | allocateDataCapture_3; // @[ReservationStation.scala 637:68]
  assign dataArray_io_multiWrite_1_data = dataArray_io_multiWrite_1_data_r; // @[ReservationStation.scala 639:12]
  assign dataArray_io_multiWrite_2_enable = dataArray_io_multiWrite_2_enable_REG; // @[ReservationStation.scala 633:14]
  assign dataArray_io_multiWrite_2_addr_0 = _dataArray_io_multiWrite_2_addr_0_T_8 | allocateDataCapture_4; // @[ReservationStation.scala 637:68]
  assign dataArray_io_multiWrite_2_addr_1 = _dataArray_io_multiWrite_2_addr_1_T_8 | allocateDataCapture_5; // @[ReservationStation.scala 637:68]
  assign dataArray_io_multiWrite_2_data = dataArray_io_multiWrite_2_data_r; // @[ReservationStation.scala 639:12]
  assign dataArray_io_multiWrite_3_enable = dataArray_io_multiWrite_3_enable_REG; // @[ReservationStation.scala 633:14]
  assign dataArray_io_multiWrite_3_addr_0 = _dataArray_io_multiWrite_3_addr_0_T_8 | allocateDataCapture_6; // @[ReservationStation.scala 637:68]
  assign dataArray_io_multiWrite_3_addr_1 = _dataArray_io_multiWrite_3_addr_1_T_8 | allocateDataCapture_7; // @[ReservationStation.scala 637:68]
  assign dataArray_io_multiWrite_3_data = dataArray_io_multiWrite_3_data_r; // @[ReservationStation.scala 639:12]
  assign dataArray_io_multiWrite_4_enable = dataArray_io_multiWrite_4_enable_REG; // @[ReservationStation.scala 633:14]
  assign dataArray_io_multiWrite_4_addr_0 = _dataArray_io_multiWrite_4_addr_0_T_8 | allocateDataCapture_8; // @[ReservationStation.scala 637:68]
  assign dataArray_io_multiWrite_4_addr_1 = _dataArray_io_multiWrite_4_addr_1_T_8 | allocateDataCapture_9; // @[ReservationStation.scala 637:68]
  assign dataArray_io_multiWrite_4_data = dataArray_io_multiWrite_4_data_r; // @[ReservationStation.scala 639:12]
  assign payloadArray_clock = clock;
  assign payloadArray_io_read_0_addr = select_io_grant_0_bits; // @[ReservationStation.scala 368:34]
  assign payloadArray_io_read_1_addr = s1_oldestSel_age_io_out; // @[SelectPolicy.scala 177:19 179:14]
  assign payloadArray_io_write_0_enable = s1_dispatchUops_dup_1_0_valid; // @[ReservationStation.scala 471:25]
  assign payloadArray_io_write_0_addr = s1_allocatePtrOH_dup_1_0; // @[ReservationStation.scala 472:23]
  assign payloadArray_io_write_0_data_ctrl_fuType = s1_dispatchUops_dup_1_0_bits_ctrl_fuType; // @[ReservationStation.scala 473:23]
  assign payloadArray_io_write_0_data_ctrl_fuOpType = s1_dispatchUops_dup_1_0_bits_ctrl_fuOpType; // @[ReservationStation.scala 473:23]
  assign payloadArray_io_write_0_data_ctrl_rfWen = s1_dispatchUops_dup_1_0_bits_ctrl_rfWen; // @[ReservationStation.scala 473:23]
  assign payloadArray_io_write_0_data_ctrl_fpWen = s1_dispatchUops_dup_1_0_bits_ctrl_fpWen; // @[ReservationStation.scala 473:23]
  assign payloadArray_io_write_0_data_pdest = s1_dispatchUops_dup_1_0_bits_pdest; // @[ReservationStation.scala 473:23]
  assign payloadArray_io_write_0_data_robIdx_flag = s1_dispatchUops_dup_1_0_bits_robIdx_flag; // @[ReservationStation.scala 473:23]
  assign payloadArray_io_write_0_data_robIdx_value = s1_dispatchUops_dup_1_0_bits_robIdx_value; // @[ReservationStation.scala 473:23]
  assign payloadArray_io_write_1_enable = s1_dispatchUops_dup_1_1_valid; // @[ReservationStation.scala 471:25]
  assign payloadArray_io_write_1_addr = s1_allocatePtrOH_dup_1_1; // @[ReservationStation.scala 472:23]
  assign payloadArray_io_write_1_data_ctrl_fuType = s1_dispatchUops_dup_1_1_bits_ctrl_fuType; // @[ReservationStation.scala 473:23]
  assign payloadArray_io_write_1_data_ctrl_fuOpType = s1_dispatchUops_dup_1_1_bits_ctrl_fuOpType; // @[ReservationStation.scala 473:23]
  assign payloadArray_io_write_1_data_ctrl_rfWen = s1_dispatchUops_dup_1_1_bits_ctrl_rfWen; // @[ReservationStation.scala 473:23]
  assign payloadArray_io_write_1_data_ctrl_fpWen = s1_dispatchUops_dup_1_1_bits_ctrl_fpWen; // @[ReservationStation.scala 473:23]
  assign payloadArray_io_write_1_data_pdest = s1_dispatchUops_dup_1_1_bits_pdest; // @[ReservationStation.scala 473:23]
  assign payloadArray_io_write_1_data_robIdx_flag = s1_dispatchUops_dup_1_1_bits_robIdx_flag; // @[ReservationStation.scala 473:23]
  assign payloadArray_io_write_1_data_robIdx_value = s1_dispatchUops_dup_1_1_bits_robIdx_value; // @[ReservationStation.scala 473:23]
  assign s1_oldestSel_age_clock = clock;
  assign s1_oldestSel_age_reset = reset;
  assign s1_oldestSel_age_io_enq_0 = enqVec_REG; // @[ReservationStation.scala 361:{23,23}]
  assign s1_oldestSel_age_io_enq_1 = enqVec_REG_1; // @[ReservationStation.scala 361:{23,23}]
  assign s1_oldestSel_age_io_deq = statusArray_io_flushed; // @[SelectPolicy.scala 176:16]
  assign oldestSelection_io_oldest_valid = |_s1_oldestSel_out_valid_T; // @[SelectPolicy.scala 178:42]
  assign wakeupQueue_clock = clock;
  assign wakeupQueue_reset = reset;
  assign wakeupQueue_io_in_valid = s1_issuePtrOH_0_valid & s2_deq_0_ready & fuCheck; // @[ReservationStation.scala 567:76]
  assign wakeupQueue_io_in_bits_ctrl_rfWen = s1_issue_oldest_0 ? payloadArray_io_read_1_data_ctrl_rfWen :
    _s1_out_0_bits_uop_T_ctrl_rfWen; // @[ReservationStation.scala 518:30]
  assign wakeupQueue_io_in_bits_pdest = s1_issue_oldest_0 ? payloadArray_io_read_1_data_pdest :
    _s1_out_0_bits_uop_T_pdest; // @[ReservationStation.scala 518:30]
  assign wakeupQueue_io_in_bits_robIdx_flag = s1_issue_oldest_0 ? payloadArray_io_read_1_data_robIdx_flag :
    _s1_out_0_bits_uop_T_robIdx_flag; // @[ReservationStation.scala 518:30]
  assign wakeupQueue_io_in_bits_robIdx_value = s1_issue_oldest_0 ? payloadArray_io_read_1_data_robIdx_value :
    _s1_out_0_bits_uop_T_robIdx_value; // @[ReservationStation.scala 518:30]
  assign wakeupQueue_io_redirect_valid = io_redirect_valid; // @[ReservationStation.scala 570:31]
  assign wakeupQueue_io_redirect_bits_robIdx_flag = io_redirect_bits_robIdx_flag; // @[ReservationStation.scala 570:31]
  assign wakeupQueue_io_redirect_bits_robIdx_value = io_redirect_bits_robIdx_value; // @[ReservationStation.scala 570:31]
  assign wakeupQueue_io_redirect_bits_level = io_redirect_bits_level; // @[ReservationStation.scala 570:31]
  assign immExt_io_uop_ctrl_srcType_1 = s1_dispatchUops_dup_2_0_bits_ctrl_srcType_1; // @[DataArray.scala 162:19]
  assign immExt_io_uop_ctrl_imm = s1_dispatchUops_dup_2_0_bits_ctrl_imm; // @[DataArray.scala 162:19]
  assign immExt_io_data_in_0 = io_srcRegValue_0_0; // @[DataArray.scala 163:23]
  assign immExt_io_data_in_1 = io_srcRegValue_0_1; // @[DataArray.scala 163:23]
  assign immExt_1_io_uop_ctrl_srcType_1 = s1_dispatchUops_dup_2_1_bits_ctrl_srcType_1; // @[DataArray.scala 162:19]
  assign immExt_1_io_uop_ctrl_imm = s1_dispatchUops_dup_2_1_bits_ctrl_imm; // @[DataArray.scala 162:19]
  assign immExt_1_io_data_in_0 = io_srcRegValue_1_0; // @[DataArray.scala 163:23]
  assign immExt_1_io_data_in_1 = io_srcRegValue_1_1; // @[DataArray.scala 163:23]
  assign dataSelect_io_doOverride_0 = oldestSelection_io_isOverrided_0; // @[ReservationStation.scala 402:29 504:21]
  assign dataSelect_io_readData_0_0 = dataArray_io_read_0_data_0; // @[ReservationStation.scala 693:26]
  assign dataSelect_io_readData_0_1 = dataArray_io_read_0_data_1; // @[ReservationStation.scala 693:26]
  assign dataSelect_io_readData_1_0 = dataArray_io_read_1_data_0; // @[ReservationStation.scala 693:26]
  assign dataSelect_io_readData_1_1 = dataArray_io_read_1_data_1; // @[ReservationStation.scala 693:26]
  assign dataSelect_io_fromSlowPorts_0_0 = {dataSelect_io_fromSlowPorts_0_0_hi,dataSelect_io_fromSlowPorts_0_0_lo}; // @[ReservationStation.scala 697:103]
  assign dataSelect_io_fromSlowPorts_0_1 = {dataSelect_io_fromSlowPorts_0_1_hi,dataSelect_io_fromSlowPorts_0_1_lo}; // @[ReservationStation.scala 697:103]
  assign dataSelect_io_fromSlowPorts_1_0 = {dataSelect_io_fromSlowPorts_1_0_hi,dataSelect_io_fromSlowPorts_1_0_lo}; // @[ReservationStation.scala 697:103]
  assign dataSelect_io_fromSlowPorts_1_1 = {dataSelect_io_fromSlowPorts_1_1_hi,dataSelect_io_fromSlowPorts_1_1_lo}; // @[ReservationStation.scala 697:103]
  assign dataSelect_io_fromSlowPorts_2_0 = {dataSelect_io_fromSlowPorts_2_0_hi,dataSelect_io_fromSlowPorts_2_0_lo}; // @[ReservationStation.scala 697:103]
  assign dataSelect_io_fromSlowPorts_2_1 = {dataSelect_io_fromSlowPorts_2_1_hi,dataSelect_io_fromSlowPorts_2_1_lo}; // @[ReservationStation.scala 697:103]
  assign dataSelect_io_slowData_0 = dataArray_io_multiWrite_0_data; // @[ReservationStation.scala 700:26]
  assign dataSelect_io_slowData_1 = dataArray_io_multiWrite_1_data; // @[ReservationStation.scala 700:26]
  assign dataSelect_io_slowData_2 = dataArray_io_multiWrite_2_data; // @[ReservationStation.scala 700:26]
  assign dataSelect_io_slowData_3 = dataArray_io_multiWrite_3_data; // @[ReservationStation.scala 700:26]
  assign dataSelect_io_slowData_4 = dataArray_io_multiWrite_4_data; // @[ReservationStation.scala 700:26]
  assign dataSelect_io_enqBypass_0_0 = canBypass & ~s1_issue_oldest_0 & ~select_io_grant_0_valid; // @[ReservationStation.scala 512:62]
  assign dataSelect_io_enqData_0_0_bits = immExt_io_data_out_0; // @[ReservationStation.scala 589:29 593:12]
  assign dataSelect_io_enqData_0_1_bits = immExt_io_data_out_1; // @[ReservationStation.scala 589:29 593:12]
  assign bypassNetwork_clock = clock;
  assign bypassNetwork_io_hold = _T_18 | ~s1_out_0_valid; // @[ReservationStation.scala 766:49]
  assign bypassNetwork_io_source_0 = dataSelect_io_deqData_0_0; // @[ReservationStation.scala 404:20 710:29]
  assign bypassNetwork_io_source_1 = dataSelect_io_deqData_0_1; // @[ReservationStation.scala 404:20 710:29]
  assign bypassNetwork_io_bypass_0_valid_0 = _s1_issuePtrOH_0_valid_T ? normalFastWakeupMatch_0_0 : s1_fastWakeup_0_0_0; // @[ReservationStation.scala 761:40]
  assign bypassNetwork_io_bypass_0_valid_1 = _s1_issuePtrOH_0_valid_T ? normalFastWakeupMatch_1_0 : s1_fastWakeup_0_1_0; // @[ReservationStation.scala 761:40]
  assign bypassNetwork_io_bypass_0_data = io_fastDatas_0; // @[ReservationStation.scala 770:17]
  always @(posedge clock) begin
    emptyThisCycle <= numEmptyAfterS1 + _GEN_773; // @[ReservationStation.scala 319:39]
    allocateThisCycle <= _allocateThisCycle_T[1:0]; // @[ReservationStation.scala 323:25]
    allocateThisCycle_1 <= _allocateThisCycle_T_1[1:0]; // @[ReservationStation.scala 323:25]
    if (s0_doEnqueue_0) begin // @[ReservationStation.scala 361:90]
      enqVec_REG <= s0_allocatePtrOH_0;
    end else begin
      enqVec_REG <= 8'h0;
    end
    if (s0_doEnqueue_1) begin // @[ReservationStation.scala 361:90]
      enqVec_REG_1 <= s0_allocatePtrOH_1;
    end else begin
      enqVec_REG_1 <= 8'h0;
    end
    s1_dispatchUops_dup_0_0_valid <= _s0_doEnqueue_0_T & _s0_doEnqueue_0_T_1; // @[ReservationStation.scala 416:28]
    if (s0_doEnqueue_0) begin // @[ReservationStation.scala 418:21]
      s1_dispatchUops_dup_0_0_bits_ctrl_srcType_0 <= io_fromDispatch_0_bits_ctrl_srcType_0; // @[ReservationStation.scala 419:16]
    end
    if (s0_doEnqueue_0) begin // @[ReservationStation.scala 418:21]
      s1_dispatchUops_dup_0_0_bits_ctrl_srcType_1 <= io_fromDispatch_0_bits_ctrl_srcType_1; // @[ReservationStation.scala 419:16]
    end
    if (s0_doEnqueue_0) begin // @[ReservationStation.scala 418:21]
      s1_dispatchUops_dup_0_0_bits_ctrl_fuType <= io_fromDispatch_0_bits_ctrl_fuType; // @[ReservationStation.scala 419:16]
    end
    if (s0_doEnqueue_0) begin // @[ReservationStation.scala 418:21]
      s1_dispatchUops_dup_0_0_bits_ctrl_fuOpType <= io_fromDispatch_0_bits_ctrl_fuOpType; // @[ReservationStation.scala 419:16]
    end
    if (s0_doEnqueue_0) begin // @[ReservationStation.scala 418:21]
      s1_dispatchUops_dup_0_0_bits_ctrl_rfWen <= io_fromDispatch_0_bits_ctrl_rfWen; // @[ReservationStation.scala 419:16]
    end
    if (s0_doEnqueue_0) begin // @[ReservationStation.scala 418:21]
      s1_dispatchUops_dup_0_0_bits_ctrl_fpWen <= io_fromDispatch_0_bits_ctrl_fpWen; // @[ReservationStation.scala 419:16]
    end
    if (s0_doEnqueue_0) begin // @[ReservationStation.scala 418:21]
      s1_dispatchUops_dup_0_0_bits_srcState_0 <= io_fromDispatch_0_bits_srcState_0; // @[ReservationStation.scala 419:16]
    end
    if (s0_doEnqueue_0) begin // @[ReservationStation.scala 418:21]
      s1_dispatchUops_dup_0_0_bits_srcState_1 <= io_fromDispatch_0_bits_srcState_1; // @[ReservationStation.scala 419:16]
    end
    if (s0_doEnqueue_0) begin // @[ReservationStation.scala 418:21]
      s1_dispatchUops_dup_0_0_bits_psrc_0 <= io_fromDispatch_0_bits_psrc_0; // @[ReservationStation.scala 419:16]
    end
    if (s0_doEnqueue_0) begin // @[ReservationStation.scala 418:21]
      s1_dispatchUops_dup_0_0_bits_psrc_1 <= io_fromDispatch_0_bits_psrc_1; // @[ReservationStation.scala 419:16]
    end
    if (s0_doEnqueue_0) begin // @[ReservationStation.scala 418:21]
      s1_dispatchUops_dup_0_0_bits_pdest <= io_fromDispatch_0_bits_pdest; // @[ReservationStation.scala 419:16]
    end
    if (s0_doEnqueue_0) begin // @[ReservationStation.scala 418:21]
      s1_dispatchUops_dup_0_0_bits_robIdx_flag <= io_fromDispatch_0_bits_robIdx_flag; // @[ReservationStation.scala 419:16]
    end
    if (s0_doEnqueue_0) begin // @[ReservationStation.scala 418:21]
      s1_dispatchUops_dup_0_0_bits_robIdx_value <= io_fromDispatch_0_bits_robIdx_value; // @[ReservationStation.scala 419:16]
    end
    s1_dispatchUops_dup_0_1_valid <= _s0_doEnqueue_1_T & _s0_doEnqueue_0_T_1; // @[ReservationStation.scala 416:28]
    if (s0_doEnqueue_1) begin // @[ReservationStation.scala 418:21]
      s1_dispatchUops_dup_0_1_bits_ctrl_srcType_0 <= io_fromDispatch_1_bits_ctrl_srcType_0; // @[ReservationStation.scala 419:16]
    end
    if (s0_doEnqueue_1) begin // @[ReservationStation.scala 418:21]
      s1_dispatchUops_dup_0_1_bits_ctrl_srcType_1 <= io_fromDispatch_1_bits_ctrl_srcType_1; // @[ReservationStation.scala 419:16]
    end
    if (s0_doEnqueue_1) begin // @[ReservationStation.scala 418:21]
      s1_dispatchUops_dup_0_1_bits_srcState_0 <= io_fromDispatch_1_bits_srcState_0; // @[ReservationStation.scala 419:16]
    end
    if (s0_doEnqueue_1) begin // @[ReservationStation.scala 418:21]
      s1_dispatchUops_dup_0_1_bits_srcState_1 <= io_fromDispatch_1_bits_srcState_1; // @[ReservationStation.scala 419:16]
    end
    if (s0_doEnqueue_1) begin // @[ReservationStation.scala 418:21]
      s1_dispatchUops_dup_0_1_bits_psrc_0 <= io_fromDispatch_1_bits_psrc_0; // @[ReservationStation.scala 419:16]
    end
    if (s0_doEnqueue_1) begin // @[ReservationStation.scala 418:21]
      s1_dispatchUops_dup_0_1_bits_psrc_1 <= io_fromDispatch_1_bits_psrc_1; // @[ReservationStation.scala 419:16]
    end
    if (s0_doEnqueue_1) begin // @[ReservationStation.scala 418:21]
      s1_dispatchUops_dup_0_1_bits_robIdx_flag <= io_fromDispatch_1_bits_robIdx_flag; // @[ReservationStation.scala 419:16]
    end
    if (s0_doEnqueue_1) begin // @[ReservationStation.scala 418:21]
      s1_dispatchUops_dup_0_1_bits_robIdx_value <= io_fromDispatch_1_bits_robIdx_value; // @[ReservationStation.scala 419:16]
    end
    s1_dispatchUops_dup_1_0_valid <= _s0_doEnqueue_0_T & _s0_doEnqueue_0_T_1; // @[ReservationStation.scala 416:28]
    if (s0_doEnqueue_0) begin // @[ReservationStation.scala 418:21]
      s1_dispatchUops_dup_1_0_bits_ctrl_fuType <= io_fromDispatch_0_bits_ctrl_fuType; // @[ReservationStation.scala 419:16]
    end
    if (s0_doEnqueue_0) begin // @[ReservationStation.scala 418:21]
      s1_dispatchUops_dup_1_0_bits_ctrl_fuOpType <= io_fromDispatch_0_bits_ctrl_fuOpType; // @[ReservationStation.scala 419:16]
    end
    if (s0_doEnqueue_0) begin // @[ReservationStation.scala 418:21]
      s1_dispatchUops_dup_1_0_bits_ctrl_rfWen <= io_fromDispatch_0_bits_ctrl_rfWen; // @[ReservationStation.scala 419:16]
    end
    if (s0_doEnqueue_0) begin // @[ReservationStation.scala 418:21]
      s1_dispatchUops_dup_1_0_bits_ctrl_fpWen <= io_fromDispatch_0_bits_ctrl_fpWen; // @[ReservationStation.scala 419:16]
    end
    if (s0_doEnqueue_0) begin // @[ReservationStation.scala 418:21]
      s1_dispatchUops_dup_1_0_bits_pdest <= io_fromDispatch_0_bits_pdest; // @[ReservationStation.scala 419:16]
    end
    if (s0_doEnqueue_0) begin // @[ReservationStation.scala 418:21]
      s1_dispatchUops_dup_1_0_bits_robIdx_flag <= io_fromDispatch_0_bits_robIdx_flag; // @[ReservationStation.scala 419:16]
    end
    if (s0_doEnqueue_0) begin // @[ReservationStation.scala 418:21]
      s1_dispatchUops_dup_1_0_bits_robIdx_value <= io_fromDispatch_0_bits_robIdx_value; // @[ReservationStation.scala 419:16]
    end
    s1_dispatchUops_dup_1_1_valid <= _s0_doEnqueue_1_T & _s0_doEnqueue_0_T_1; // @[ReservationStation.scala 416:28]
    if (s0_doEnqueue_1) begin // @[ReservationStation.scala 418:21]
      s1_dispatchUops_dup_1_1_bits_ctrl_fuType <= io_fromDispatch_1_bits_ctrl_fuType; // @[ReservationStation.scala 419:16]
    end
    if (s0_doEnqueue_1) begin // @[ReservationStation.scala 418:21]
      s1_dispatchUops_dup_1_1_bits_ctrl_fuOpType <= io_fromDispatch_1_bits_ctrl_fuOpType; // @[ReservationStation.scala 419:16]
    end
    if (s0_doEnqueue_1) begin // @[ReservationStation.scala 418:21]
      s1_dispatchUops_dup_1_1_bits_ctrl_rfWen <= io_fromDispatch_1_bits_ctrl_rfWen; // @[ReservationStation.scala 419:16]
    end
    if (s0_doEnqueue_1) begin // @[ReservationStation.scala 418:21]
      s1_dispatchUops_dup_1_1_bits_ctrl_fpWen <= io_fromDispatch_1_bits_ctrl_fpWen; // @[ReservationStation.scala 419:16]
    end
    if (s0_doEnqueue_1) begin // @[ReservationStation.scala 418:21]
      s1_dispatchUops_dup_1_1_bits_pdest <= io_fromDispatch_1_bits_pdest; // @[ReservationStation.scala 419:16]
    end
    if (s0_doEnqueue_1) begin // @[ReservationStation.scala 418:21]
      s1_dispatchUops_dup_1_1_bits_robIdx_flag <= io_fromDispatch_1_bits_robIdx_flag; // @[ReservationStation.scala 419:16]
    end
    if (s0_doEnqueue_1) begin // @[ReservationStation.scala 418:21]
      s1_dispatchUops_dup_1_1_bits_robIdx_value <= io_fromDispatch_1_bits_robIdx_value; // @[ReservationStation.scala 419:16]
    end
    s1_dispatchUops_dup_2_0_valid <= _s0_doEnqueue_0_T & _s0_doEnqueue_0_T_1; // @[ReservationStation.scala 416:28]
    if (s0_doEnqueue_0) begin // @[ReservationStation.scala 418:21]
      s1_dispatchUops_dup_2_0_bits_ctrl_srcType_0 <= io_fromDispatch_0_bits_ctrl_srcType_0; // @[ReservationStation.scala 419:16]
    end
    if (s0_doEnqueue_0) begin // @[ReservationStation.scala 418:21]
      s1_dispatchUops_dup_2_0_bits_ctrl_srcType_1 <= io_fromDispatch_0_bits_ctrl_srcType_1; // @[ReservationStation.scala 419:16]
    end
    if (s0_doEnqueue_0) begin // @[ReservationStation.scala 418:21]
      s1_dispatchUops_dup_2_0_bits_ctrl_imm <= io_fromDispatch_0_bits_ctrl_imm; // @[ReservationStation.scala 419:16]
    end
    if (s0_doEnqueue_0) begin // @[ReservationStation.scala 418:21]
      s1_dispatchUops_dup_2_0_bits_srcState_0 <= io_fromDispatch_0_bits_srcState_0; // @[ReservationStation.scala 419:16]
    end
    if (s0_doEnqueue_0) begin // @[ReservationStation.scala 418:21]
      s1_dispatchUops_dup_2_0_bits_srcState_1 <= io_fromDispatch_0_bits_srcState_1; // @[ReservationStation.scala 419:16]
    end
    s1_dispatchUops_dup_2_1_valid <= _s0_doEnqueue_1_T & _s0_doEnqueue_0_T_1; // @[ReservationStation.scala 416:28]
    if (s0_doEnqueue_1) begin // @[ReservationStation.scala 418:21]
      s1_dispatchUops_dup_2_1_bits_ctrl_srcType_0 <= io_fromDispatch_1_bits_ctrl_srcType_0; // @[ReservationStation.scala 419:16]
    end
    if (s0_doEnqueue_1) begin // @[ReservationStation.scala 418:21]
      s1_dispatchUops_dup_2_1_bits_ctrl_srcType_1 <= io_fromDispatch_1_bits_ctrl_srcType_1; // @[ReservationStation.scala 419:16]
    end
    if (s0_doEnqueue_1) begin // @[ReservationStation.scala 418:21]
      s1_dispatchUops_dup_2_1_bits_ctrl_imm <= io_fromDispatch_1_bits_ctrl_imm; // @[ReservationStation.scala 419:16]
    end
    if (s0_doEnqueue_1) begin // @[ReservationStation.scala 418:21]
      s1_dispatchUops_dup_2_1_bits_srcState_0 <= io_fromDispatch_1_bits_srcState_0; // @[ReservationStation.scala 419:16]
    end
    if (s0_doEnqueue_1) begin // @[ReservationStation.scala 418:21]
      s1_dispatchUops_dup_2_1_bits_srcState_1 <= io_fromDispatch_1_bits_srcState_1; // @[ReservationStation.scala 419:16]
    end
    s1_allocatePtrOH_dup_0_0 <= select_io_allocate_0_bits; // @[ReservationStation.scala 273:{33,33}]
    s1_allocatePtrOH_dup_0_1 <= select_io_allocate_1_bits; // @[ReservationStation.scala 273:{33,33}]
    s1_allocatePtrOH_dup_1_0 <= select_io_allocate_0_bits; // @[ReservationStation.scala 273:{33,33}]
    s1_allocatePtrOH_dup_1_1 <= select_io_allocate_1_bits; // @[ReservationStation.scala 273:{33,33}]
    s1_allocatePtrOH_dup_2_0 <= select_io_allocate_0_bits; // @[ReservationStation.scala 273:{33,33}]
    s1_allocatePtrOH_dup_2_1 <= select_io_allocate_1_bits; // @[ReservationStation.scala 273:{33,33}]
    s1_enqWakeup_0_0 <= {s0_enqWakeup_0_0_hi,s0_enqWakeup_0_0_lo}; // @[ReservationStation.scala 341:100]
    s1_enqWakeup_0_1 <= {s0_enqWakeup_0_1_hi,s0_enqWakeup_0_1_lo}; // @[ReservationStation.scala 341:100]
    s1_enqWakeup_1_0 <= {s0_enqWakeup_1_0_hi,s0_enqWakeup_1_0_lo}; // @[ReservationStation.scala 341:100]
    s1_enqWakeup_1_1 <= {s0_enqWakeup_1_1_hi,s0_enqWakeup_1_1_lo}; // @[ReservationStation.scala 341:100]
    s1_enqDataCapture_0_0 <= {s0_enqDataCapture_0_0_hi,s0_enqDataCapture_0_0_lo}; // @[ReservationStation.scala 342:104]
    s1_enqDataCapture_0_1 <= {s0_enqDataCapture_0_1_hi,s0_enqDataCapture_0_1_lo}; // @[ReservationStation.scala 342:104]
    s1_enqDataCapture_1_0 <= {s0_enqDataCapture_1_0_hi,s0_enqDataCapture_1_0_lo}; // @[ReservationStation.scala 342:104]
    s1_enqDataCapture_1_1 <= {s0_enqDataCapture_1_1_hi,s0_enqDataCapture_1_1_lo}; // @[ReservationStation.scala 342:104]
    s1_fastWakeup_0_0_0 <= io_fastUopsIn_0_valid & dataCond_15; // @[ReservationStation.scala 344:83]
    s1_fastWakeup_0_1_0 <= io_fastUopsIn_0_valid & dataCond_16; // @[ReservationStation.scala 344:83]
    s1_fastWakeup_1_0_0 <= io_fastUopsIn_0_valid & dataCond_33; // @[ReservationStation.scala 344:83]
    s1_fastWakeup_1_1_0 <= io_fastUopsIn_0_valid & dataCond_34; // @[ReservationStation.scala 344:83]
    slowWakeupMatchVec_0_0 <= statusArray_io_wakeupMatch_0_0[5:1]; // @[ReservationStation.scala 629:67]
    slowWakeupMatchVec_0_1 <= statusArray_io_wakeupMatch_0_1[5:1]; // @[ReservationStation.scala 629:67]
    slowWakeupMatchVec_1_0 <= statusArray_io_wakeupMatch_1_0[5:1]; // @[ReservationStation.scala 629:67]
    slowWakeupMatchVec_1_1 <= statusArray_io_wakeupMatch_1_1[5:1]; // @[ReservationStation.scala 629:67]
    slowWakeupMatchVec_2_0 <= statusArray_io_wakeupMatch_2_0[5:1]; // @[ReservationStation.scala 629:67]
    slowWakeupMatchVec_2_1 <= statusArray_io_wakeupMatch_2_1[5:1]; // @[ReservationStation.scala 629:67]
    slowWakeupMatchVec_3_0 <= statusArray_io_wakeupMatch_3_0[5:1]; // @[ReservationStation.scala 629:67]
    slowWakeupMatchVec_3_1 <= statusArray_io_wakeupMatch_3_1[5:1]; // @[ReservationStation.scala 629:67]
    slowWakeupMatchVec_4_0 <= statusArray_io_wakeupMatch_4_0[5:1]; // @[ReservationStation.scala 629:67]
    slowWakeupMatchVec_4_1 <= statusArray_io_wakeupMatch_4_1[5:1]; // @[ReservationStation.scala 629:67]
    slowWakeupMatchVec_5_0 <= statusArray_io_wakeupMatch_5_0[5:1]; // @[ReservationStation.scala 629:67]
    slowWakeupMatchVec_5_1 <= statusArray_io_wakeupMatch_5_1[5:1]; // @[ReservationStation.scala 629:67]
    slowWakeupMatchVec_6_0 <= statusArray_io_wakeupMatch_6_0[5:1]; // @[ReservationStation.scala 629:67]
    slowWakeupMatchVec_6_1 <= statusArray_io_wakeupMatch_6_1[5:1]; // @[ReservationStation.scala 629:67]
    slowWakeupMatchVec_7_0 <= statusArray_io_wakeupMatch_7_0[5:1]; // @[ReservationStation.scala 629:67]
    slowWakeupMatchVec_7_1 <= statusArray_io_wakeupMatch_7_1[5:1]; // @[ReservationStation.scala 629:67]
    dataArray_io_multiWrite_0_enable_REG <= io_slowPorts_0_valid; // @[ReservationStation.scala 633:24]
    if (io_slowPorts_0_valid) begin // @[Reg.scala 17:18]
      dataArray_io_multiWrite_0_data_r <= io_slowPorts_0_bits_data; // @[Reg.scala 17:22]
    end
    dataArray_io_multiWrite_1_enable_REG <= io_slowPorts_1_valid; // @[ReservationStation.scala 633:24]
    if (io_slowPorts_1_valid) begin // @[Reg.scala 17:18]
      dataArray_io_multiWrite_1_data_r <= io_slowPorts_1_bits_data; // @[Reg.scala 17:22]
    end
    dataArray_io_multiWrite_2_enable_REG <= io_slowPorts_2_valid; // @[ReservationStation.scala 633:24]
    if (io_slowPorts_2_valid) begin // @[Reg.scala 17:18]
      dataArray_io_multiWrite_2_data_r <= io_slowPorts_2_bits_data; // @[Reg.scala 17:22]
    end
    dataArray_io_multiWrite_3_enable_REG <= io_slowPorts_3_valid; // @[ReservationStation.scala 633:24]
    if (io_slowPorts_3_valid) begin // @[Reg.scala 17:18]
      dataArray_io_multiWrite_3_data_r <= io_slowPorts_3_bits_data; // @[Reg.scala 17:22]
    end
    dataArray_io_multiWrite_4_enable_REG <= io_slowPorts_4_valid; // @[ReservationStation.scala 633:24]
    if (io_slowPorts_4_valid) begin // @[Reg.scala 17:18]
      dataArray_io_multiWrite_4_data_r <= io_slowPorts_4_bits_data; // @[Reg.scala 17:22]
    end
    fastWakeupMatch_0_0_0 <= statusArray_io_wakeupMatch_0_0[0]; // @[ReservationStation.scala 721:65]
    fastWakeupMatch_0_1_0 <= statusArray_io_wakeupMatch_0_1[0]; // @[ReservationStation.scala 721:65]
    fastWakeupMatch_1_0_0 <= statusArray_io_wakeupMatch_1_0[0]; // @[ReservationStation.scala 721:65]
    fastWakeupMatch_1_1_0 <= statusArray_io_wakeupMatch_1_1[0]; // @[ReservationStation.scala 721:65]
    fastWakeupMatch_2_0_0 <= statusArray_io_wakeupMatch_2_0[0]; // @[ReservationStation.scala 721:65]
    fastWakeupMatch_2_1_0 <= statusArray_io_wakeupMatch_2_1[0]; // @[ReservationStation.scala 721:65]
    fastWakeupMatch_3_0_0 <= statusArray_io_wakeupMatch_3_0[0]; // @[ReservationStation.scala 721:65]
    fastWakeupMatch_3_1_0 <= statusArray_io_wakeupMatch_3_1[0]; // @[ReservationStation.scala 721:65]
    fastWakeupMatch_4_0_0 <= statusArray_io_wakeupMatch_4_0[0]; // @[ReservationStation.scala 721:65]
    fastWakeupMatch_4_1_0 <= statusArray_io_wakeupMatch_4_1[0]; // @[ReservationStation.scala 721:65]
    fastWakeupMatch_5_0_0 <= statusArray_io_wakeupMatch_5_0[0]; // @[ReservationStation.scala 721:65]
    fastWakeupMatch_5_1_0 <= statusArray_io_wakeupMatch_5_1[0]; // @[ReservationStation.scala 721:65]
    fastWakeupMatch_6_0_0 <= statusArray_io_wakeupMatch_6_0[0]; // @[ReservationStation.scala 721:65]
    fastWakeupMatch_6_1_0 <= statusArray_io_wakeupMatch_6_1[0]; // @[ReservationStation.scala 721:65]
    fastWakeupMatch_7_0_0 <= statusArray_io_wakeupMatch_7_0[0]; // @[ReservationStation.scala 721:65]
    fastWakeupMatch_7_1_0 <= statusArray_io_wakeupMatch_7_1[0]; // @[ReservationStation.scala 721:65]
    if (s1_out_fire_0) begin // @[Reg.scala 17:18]
      if (s1_issue_oldest_0) begin // @[ReservationStation.scala 518:30]
        data_uop_robIdx_flag <= payloadArray_io_read_1_data_robIdx_flag;
      end else if (select_io_grant_0_valid) begin // @[ReservationStation.scala 519:10]
        data_uop_robIdx_flag <= payloadArray_io_read_0_data_robIdx_flag;
      end else begin
        data_uop_robIdx_flag <= s1_dispatchUops_dup_0_0_bits_robIdx_flag;
      end
    end
    if (s1_out_fire_0) begin // @[Reg.scala 17:18]
      if (s1_issue_oldest_0) begin // @[ReservationStation.scala 518:30]
        data_uop_robIdx_value <= payloadArray_io_read_1_data_robIdx_value;
      end else if (select_io_grant_0_valid) begin // @[ReservationStation.scala 519:10]
        data_uop_robIdx_value <= payloadArray_io_read_0_data_robIdx_value;
      end else begin
        data_uop_robIdx_value <= s1_dispatchUops_dup_0_0_bits_robIdx_value;
      end
    end
    if (s1_out_fire_0) begin // @[Reg.scala 17:18]
      if (s1_issue_oldest_0) begin // @[ReservationStation.scala 518:30]
        data_uop_ctrl_fuType <= payloadArray_io_read_1_data_ctrl_fuType;
      end else if (select_io_grant_0_valid) begin // @[ReservationStation.scala 519:10]
        data_uop_ctrl_fuType <= payloadArray_io_read_0_data_ctrl_fuType;
      end else begin
        data_uop_ctrl_fuType <= s1_dispatchUops_dup_0_0_bits_ctrl_fuType;
      end
    end
    if (s1_out_fire_0) begin // @[Reg.scala 17:18]
      if (s1_issue_oldest_0) begin // @[ReservationStation.scala 518:30]
        data_uop_ctrl_fuOpType <= payloadArray_io_read_1_data_ctrl_fuOpType;
      end else if (select_io_grant_0_valid) begin // @[ReservationStation.scala 519:10]
        data_uop_ctrl_fuOpType <= payloadArray_io_read_0_data_ctrl_fuOpType;
      end else begin
        data_uop_ctrl_fuOpType <= s1_dispatchUops_dup_0_0_bits_ctrl_fuOpType;
      end
    end
    if (s1_out_fire_0) begin // @[Reg.scala 17:18]
      if (s1_issue_oldest_0) begin // @[ReservationStation.scala 518:30]
        data_uop_ctrl_rfWen <= payloadArray_io_read_1_data_ctrl_rfWen;
      end else if (select_io_grant_0_valid) begin // @[ReservationStation.scala 519:10]
        data_uop_ctrl_rfWen <= payloadArray_io_read_0_data_ctrl_rfWen;
      end else begin
        data_uop_ctrl_rfWen <= s1_dispatchUops_dup_0_0_bits_ctrl_rfWen;
      end
    end
    if (s1_out_fire_0) begin // @[Reg.scala 17:18]
      if (s1_issue_oldest_0) begin // @[ReservationStation.scala 518:30]
        data_uop_ctrl_fpWen <= payloadArray_io_read_1_data_ctrl_fpWen;
      end else if (select_io_grant_0_valid) begin // @[ReservationStation.scala 519:10]
        data_uop_ctrl_fpWen <= payloadArray_io_read_0_data_ctrl_fpWen;
      end else begin
        data_uop_ctrl_fpWen <= s1_dispatchUops_dup_0_0_bits_ctrl_fpWen;
      end
    end
    if (s1_out_fire_0) begin // @[Reg.scala 17:18]
      if (s1_issue_oldest_0) begin // @[ReservationStation.scala 518:30]
        data_uop_pdest <= payloadArray_io_read_1_data_pdest;
      end else if (select_io_grant_0_valid) begin // @[ReservationStation.scala 519:10]
        data_uop_pdest <= payloadArray_io_read_0_data_pdest;
      end else begin
        data_uop_pdest <= s1_dispatchUops_dup_0_0_bits_pdest;
      end
    end
    io_perf_0_value_REG <= &statusArray_io_isValid; // @[ReservationStation.scala 966:56]
    io_perf_0_value_REG_1 <= io_perf_0_value_REG; // @[PerfCounterUtils.scala 188:27]
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ReservationStation.scala 284:52]
      validAfterAllocate <= 8'h0;
    end else begin
      validAfterAllocate <= statusArray_io_isValidNext | validUpdateByAllocate;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PipelineConnect.scala 111:21]
      valid <= 1'h0; // @[PipelineConnect.scala 111:29]
    end else begin
      valid <= s1_out_fire_0 | _GEN_657;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  validAfterAllocate = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  emptyThisCycle = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  allocateThisCycle = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  allocateThisCycle_1 = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  enqVec_REG = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  enqVec_REG_1 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  s1_dispatchUops_dup_0_0_valid = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  s1_dispatchUops_dup_0_0_bits_ctrl_srcType_0 = _RAND_7[1:0];
  _RAND_8 = {1{`RANDOM}};
  s1_dispatchUops_dup_0_0_bits_ctrl_srcType_1 = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  s1_dispatchUops_dup_0_0_bits_ctrl_fuType = _RAND_9[3:0];
  _RAND_10 = {1{`RANDOM}};
  s1_dispatchUops_dup_0_0_bits_ctrl_fuOpType = _RAND_10[6:0];
  _RAND_11 = {1{`RANDOM}};
  s1_dispatchUops_dup_0_0_bits_ctrl_rfWen = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  s1_dispatchUops_dup_0_0_bits_ctrl_fpWen = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  s1_dispatchUops_dup_0_0_bits_srcState_0 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  s1_dispatchUops_dup_0_0_bits_srcState_1 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  s1_dispatchUops_dup_0_0_bits_psrc_0 = _RAND_15[5:0];
  _RAND_16 = {1{`RANDOM}};
  s1_dispatchUops_dup_0_0_bits_psrc_1 = _RAND_16[5:0];
  _RAND_17 = {1{`RANDOM}};
  s1_dispatchUops_dup_0_0_bits_pdest = _RAND_17[5:0];
  _RAND_18 = {1{`RANDOM}};
  s1_dispatchUops_dup_0_0_bits_robIdx_flag = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  s1_dispatchUops_dup_0_0_bits_robIdx_value = _RAND_19[4:0];
  _RAND_20 = {1{`RANDOM}};
  s1_dispatchUops_dup_0_1_valid = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  s1_dispatchUops_dup_0_1_bits_ctrl_srcType_0 = _RAND_21[1:0];
  _RAND_22 = {1{`RANDOM}};
  s1_dispatchUops_dup_0_1_bits_ctrl_srcType_1 = _RAND_22[1:0];
  _RAND_23 = {1{`RANDOM}};
  s1_dispatchUops_dup_0_1_bits_srcState_0 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  s1_dispatchUops_dup_0_1_bits_srcState_1 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  s1_dispatchUops_dup_0_1_bits_psrc_0 = _RAND_25[5:0];
  _RAND_26 = {1{`RANDOM}};
  s1_dispatchUops_dup_0_1_bits_psrc_1 = _RAND_26[5:0];
  _RAND_27 = {1{`RANDOM}};
  s1_dispatchUops_dup_0_1_bits_robIdx_flag = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  s1_dispatchUops_dup_0_1_bits_robIdx_value = _RAND_28[4:0];
  _RAND_29 = {1{`RANDOM}};
  s1_dispatchUops_dup_1_0_valid = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  s1_dispatchUops_dup_1_0_bits_ctrl_fuType = _RAND_30[3:0];
  _RAND_31 = {1{`RANDOM}};
  s1_dispatchUops_dup_1_0_bits_ctrl_fuOpType = _RAND_31[6:0];
  _RAND_32 = {1{`RANDOM}};
  s1_dispatchUops_dup_1_0_bits_ctrl_rfWen = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  s1_dispatchUops_dup_1_0_bits_ctrl_fpWen = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  s1_dispatchUops_dup_1_0_bits_pdest = _RAND_34[5:0];
  _RAND_35 = {1{`RANDOM}};
  s1_dispatchUops_dup_1_0_bits_robIdx_flag = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  s1_dispatchUops_dup_1_0_bits_robIdx_value = _RAND_36[4:0];
  _RAND_37 = {1{`RANDOM}};
  s1_dispatchUops_dup_1_1_valid = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  s1_dispatchUops_dup_1_1_bits_ctrl_fuType = _RAND_38[3:0];
  _RAND_39 = {1{`RANDOM}};
  s1_dispatchUops_dup_1_1_bits_ctrl_fuOpType = _RAND_39[6:0];
  _RAND_40 = {1{`RANDOM}};
  s1_dispatchUops_dup_1_1_bits_ctrl_rfWen = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  s1_dispatchUops_dup_1_1_bits_ctrl_fpWen = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  s1_dispatchUops_dup_1_1_bits_pdest = _RAND_42[5:0];
  _RAND_43 = {1{`RANDOM}};
  s1_dispatchUops_dup_1_1_bits_robIdx_flag = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  s1_dispatchUops_dup_1_1_bits_robIdx_value = _RAND_44[4:0];
  _RAND_45 = {1{`RANDOM}};
  s1_dispatchUops_dup_2_0_valid = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  s1_dispatchUops_dup_2_0_bits_ctrl_srcType_0 = _RAND_46[1:0];
  _RAND_47 = {1{`RANDOM}};
  s1_dispatchUops_dup_2_0_bits_ctrl_srcType_1 = _RAND_47[1:0];
  _RAND_48 = {1{`RANDOM}};
  s1_dispatchUops_dup_2_0_bits_ctrl_imm = _RAND_48[19:0];
  _RAND_49 = {1{`RANDOM}};
  s1_dispatchUops_dup_2_0_bits_srcState_0 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  s1_dispatchUops_dup_2_0_bits_srcState_1 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  s1_dispatchUops_dup_2_1_valid = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  s1_dispatchUops_dup_2_1_bits_ctrl_srcType_0 = _RAND_52[1:0];
  _RAND_53 = {1{`RANDOM}};
  s1_dispatchUops_dup_2_1_bits_ctrl_srcType_1 = _RAND_53[1:0];
  _RAND_54 = {1{`RANDOM}};
  s1_dispatchUops_dup_2_1_bits_ctrl_imm = _RAND_54[19:0];
  _RAND_55 = {1{`RANDOM}};
  s1_dispatchUops_dup_2_1_bits_srcState_0 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  s1_dispatchUops_dup_2_1_bits_srcState_1 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  s1_allocatePtrOH_dup_0_0 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  s1_allocatePtrOH_dup_0_1 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  s1_allocatePtrOH_dup_1_0 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  s1_allocatePtrOH_dup_1_1 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  s1_allocatePtrOH_dup_2_0 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  s1_allocatePtrOH_dup_2_1 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  s1_enqWakeup_0_0 = _RAND_63[4:0];
  _RAND_64 = {1{`RANDOM}};
  s1_enqWakeup_0_1 = _RAND_64[4:0];
  _RAND_65 = {1{`RANDOM}};
  s1_enqWakeup_1_0 = _RAND_65[4:0];
  _RAND_66 = {1{`RANDOM}};
  s1_enqWakeup_1_1 = _RAND_66[4:0];
  _RAND_67 = {1{`RANDOM}};
  s1_enqDataCapture_0_0 = _RAND_67[4:0];
  _RAND_68 = {1{`RANDOM}};
  s1_enqDataCapture_0_1 = _RAND_68[4:0];
  _RAND_69 = {1{`RANDOM}};
  s1_enqDataCapture_1_0 = _RAND_69[4:0];
  _RAND_70 = {1{`RANDOM}};
  s1_enqDataCapture_1_1 = _RAND_70[4:0];
  _RAND_71 = {1{`RANDOM}};
  s1_fastWakeup_0_0_0 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  s1_fastWakeup_0_1_0 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  s1_fastWakeup_1_0_0 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  s1_fastWakeup_1_1_0 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  valid = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  slowWakeupMatchVec_0_0 = _RAND_76[4:0];
  _RAND_77 = {1{`RANDOM}};
  slowWakeupMatchVec_0_1 = _RAND_77[4:0];
  _RAND_78 = {1{`RANDOM}};
  slowWakeupMatchVec_1_0 = _RAND_78[4:0];
  _RAND_79 = {1{`RANDOM}};
  slowWakeupMatchVec_1_1 = _RAND_79[4:0];
  _RAND_80 = {1{`RANDOM}};
  slowWakeupMatchVec_2_0 = _RAND_80[4:0];
  _RAND_81 = {1{`RANDOM}};
  slowWakeupMatchVec_2_1 = _RAND_81[4:0];
  _RAND_82 = {1{`RANDOM}};
  slowWakeupMatchVec_3_0 = _RAND_82[4:0];
  _RAND_83 = {1{`RANDOM}};
  slowWakeupMatchVec_3_1 = _RAND_83[4:0];
  _RAND_84 = {1{`RANDOM}};
  slowWakeupMatchVec_4_0 = _RAND_84[4:0];
  _RAND_85 = {1{`RANDOM}};
  slowWakeupMatchVec_4_1 = _RAND_85[4:0];
  _RAND_86 = {1{`RANDOM}};
  slowWakeupMatchVec_5_0 = _RAND_86[4:0];
  _RAND_87 = {1{`RANDOM}};
  slowWakeupMatchVec_5_1 = _RAND_87[4:0];
  _RAND_88 = {1{`RANDOM}};
  slowWakeupMatchVec_6_0 = _RAND_88[4:0];
  _RAND_89 = {1{`RANDOM}};
  slowWakeupMatchVec_6_1 = _RAND_89[4:0];
  _RAND_90 = {1{`RANDOM}};
  slowWakeupMatchVec_7_0 = _RAND_90[4:0];
  _RAND_91 = {1{`RANDOM}};
  slowWakeupMatchVec_7_1 = _RAND_91[4:0];
  _RAND_92 = {1{`RANDOM}};
  dataArray_io_multiWrite_0_enable_REG = _RAND_92[0:0];
  _RAND_93 = {2{`RANDOM}};
  dataArray_io_multiWrite_0_data_r = _RAND_93[63:0];
  _RAND_94 = {1{`RANDOM}};
  dataArray_io_multiWrite_1_enable_REG = _RAND_94[0:0];
  _RAND_95 = {2{`RANDOM}};
  dataArray_io_multiWrite_1_data_r = _RAND_95[63:0];
  _RAND_96 = {1{`RANDOM}};
  dataArray_io_multiWrite_2_enable_REG = _RAND_96[0:0];
  _RAND_97 = {2{`RANDOM}};
  dataArray_io_multiWrite_2_data_r = _RAND_97[63:0];
  _RAND_98 = {1{`RANDOM}};
  dataArray_io_multiWrite_3_enable_REG = _RAND_98[0:0];
  _RAND_99 = {2{`RANDOM}};
  dataArray_io_multiWrite_3_data_r = _RAND_99[63:0];
  _RAND_100 = {1{`RANDOM}};
  dataArray_io_multiWrite_4_enable_REG = _RAND_100[0:0];
  _RAND_101 = {2{`RANDOM}};
  dataArray_io_multiWrite_4_data_r = _RAND_101[63:0];
  _RAND_102 = {1{`RANDOM}};
  fastWakeupMatch_0_0_0 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  fastWakeupMatch_0_1_0 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  fastWakeupMatch_1_0_0 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  fastWakeupMatch_1_1_0 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  fastWakeupMatch_2_0_0 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  fastWakeupMatch_2_1_0 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  fastWakeupMatch_3_0_0 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  fastWakeupMatch_3_1_0 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  fastWakeupMatch_4_0_0 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  fastWakeupMatch_4_1_0 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  fastWakeupMatch_5_0_0 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  fastWakeupMatch_5_1_0 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  fastWakeupMatch_6_0_0 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  fastWakeupMatch_6_1_0 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  fastWakeupMatch_7_0_0 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  fastWakeupMatch_7_1_0 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  data_uop_robIdx_flag = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  data_uop_robIdx_value = _RAND_119[4:0];
  _RAND_120 = {1{`RANDOM}};
  data_uop_ctrl_fuType = _RAND_120[3:0];
  _RAND_121 = {1{`RANDOM}};
  data_uop_ctrl_fuOpType = _RAND_121[6:0];
  _RAND_122 = {1{`RANDOM}};
  data_uop_ctrl_rfWen = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  data_uop_ctrl_fpWen = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  data_uop_pdest = _RAND_124[5:0];
  _RAND_125 = {1{`RANDOM}};
  io_perf_0_value_REG = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  io_perf_0_value_REG_1 = _RAND_126[0:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    validAfterAllocate = 8'h0;
  end
  if (reset) begin
    valid = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule

