module CSA3_2_3358(
  input  [7:0] io_in_0,
  input  [7:0] io_in_1,
  input  [7:0] io_in_2,
  output [7:0] io_out_0,
  output [7:0] io_out_1
);
  wire  a = io_in_0[0]; // @[FDIV.scala 677:32]
  wire  b = io_in_1[0]; // @[FDIV.scala 677:45]
  wire  cin = io_in_2[0]; // @[FDIV.scala 677:58]
  wire  a_xor_b = a ^ b; // @[FDIV.scala 678:21]
  wire  a_and_b = a & b; // @[FDIV.scala 679:21]
  wire  sum = a_xor_b ^ cin; // @[FDIV.scala 680:23]
  wire  cout = a_and_b | a_xor_b & cin; // @[FDIV.scala 681:24]
  wire [1:0] temp_0 = {cout,sum}; // @[Cat.scala 31:58]
  wire  a_1 = io_in_0[1]; // @[FDIV.scala 677:32]
  wire  b_1 = io_in_1[1]; // @[FDIV.scala 677:45]
  wire  cin_1 = io_in_2[1]; // @[FDIV.scala 677:58]
  wire  a_xor_b1 = a_1 ^ b_1; // @[FDIV.scala 678:21]
  wire  a_and_b1 = a_1 & b_1; // @[FDIV.scala 679:21]
  wire  sum_1 = a_xor_b1 ^ cin_1; // @[FDIV.scala 680:23]
  wire  cout_1 = a_and_b1 | a_xor_b1 & cin_1; // @[FDIV.scala 681:24]
  wire [1:0] temp_1 = {cout_1,sum_1}; // @[Cat.scala 31:58]
  wire  a_2 = io_in_0[2]; // @[FDIV.scala 677:32]
  wire  b_2 = io_in_1[2]; // @[FDIV.scala 677:45]
  wire  cin_2 = io_in_2[2]; // @[FDIV.scala 677:58]
  wire  a_xor_b2 = a_2 ^ b_2; // @[FDIV.scala 678:21]
  wire  a_and_b2 = a_2 & b_2; // @[FDIV.scala 679:21]
  wire  sum_2 = a_xor_b2 ^ cin_2; // @[FDIV.scala 680:23]
  wire  cout_2 = a_and_b2 | a_xor_b2 & cin_2; // @[FDIV.scala 681:24]
  wire [1:0] temp_2 = {cout_2,sum_2}; // @[Cat.scala 31:58]
  wire  a_3 = io_in_0[3]; // @[FDIV.scala 677:32]
  wire  b_3 = io_in_1[3]; // @[FDIV.scala 677:45]
  wire  cin_3 = io_in_2[3]; // @[FDIV.scala 677:58]
  wire  a_xor_b3 = a_3 ^ b_3; // @[FDIV.scala 678:21]
  wire  a_and_b3 = a_3 & b_3; // @[FDIV.scala 679:21]
  wire  sum_3 = a_xor_b3 ^ cin_3; // @[FDIV.scala 680:23]
  wire  cout_3 = a_and_b3 | a_xor_b3 & cin_3; // @[FDIV.scala 681:24]
  wire [1:0] temp_3 = {cout_3,sum_3}; // @[Cat.scala 31:58]
  wire  a_4 = io_in_0[4]; // @[FDIV.scala 677:32]
  wire  b_4 = io_in_1[4]; // @[FDIV.scala 677:45]
  wire  cin_4 = io_in_2[4]; // @[FDIV.scala 677:58]
  wire  a_xor_b4 = a_4 ^ b_4; // @[FDIV.scala 678:21]
  wire  a_and_b4 = a_4 & b_4; // @[FDIV.scala 679:21]
  wire  sum_4 = a_xor_b4 ^ cin_4; // @[FDIV.scala 680:23]
  wire  cout_4 = a_and_b4 | a_xor_b4 & cin_4; // @[FDIV.scala 681:24]
  wire [1:0] temp_4 = {cout_4,sum_4}; // @[Cat.scala 31:58]
  wire  a_5 = io_in_0[5]; // @[FDIV.scala 677:32]
  wire  b_5 = io_in_1[5]; // @[FDIV.scala 677:45]
  wire  cin_5 = io_in_2[5]; // @[FDIV.scala 677:58]
  wire  a_xor_b5 = a_5 ^ b_5; // @[FDIV.scala 678:21]
  wire  a_and_b5 = a_5 & b_5; // @[FDIV.scala 679:21]
  wire  sum_5 = a_xor_b5 ^ cin_5; // @[FDIV.scala 680:23]
  wire  cout_5 = a_and_b5 | a_xor_b5 & cin_5; // @[FDIV.scala 681:24]
  wire [1:0] temp_5 = {cout_5,sum_5}; // @[Cat.scala 31:58]
  wire  a_6 = io_in_0[6]; // @[FDIV.scala 677:32]
  wire  b_6 = io_in_1[6]; // @[FDIV.scala 677:45]
  wire  cin_6 = io_in_2[6]; // @[FDIV.scala 677:58]
  wire  a_xor_b6 = a_6 ^ b_6; // @[FDIV.scala 678:21]
  wire  a_and_b6 = a_6 & b_6; // @[FDIV.scala 679:21]
  wire  sum_6 = a_xor_b6 ^ cin_6; // @[FDIV.scala 680:23]
  wire  cout_6 = a_and_b6 | a_xor_b6 & cin_6; // @[FDIV.scala 681:24]
  wire [1:0] temp_6 = {cout_6,sum_6}; // @[Cat.scala 31:58]
  wire  a_7 = io_in_0[7]; // @[FDIV.scala 677:32]
  wire  b_7 = io_in_1[7]; // @[FDIV.scala 677:45]
  wire  cin_7 = io_in_2[7]; // @[FDIV.scala 677:58]
  wire  a_xor_b7 = a_7 ^ b_7; // @[FDIV.scala 678:21]
  wire  a_and_b7 = a_7 & b_7; // @[FDIV.scala 679:21]
  wire  sum_7 = a_xor_b7 ^ cin_7; // @[FDIV.scala 680:23]
  wire  cout_7 = a_and_b7 | a_xor_b7 & cin_7; // @[FDIV.scala 681:24]
  wire [1:0] temp_7 = {cout_7,sum_7}; // @[Cat.scala 31:58]
  wire [3:0] io_out_0_lo = {temp_3[0],temp_2[0],temp_1[0],temp_0[0]}; // @[Cat.scala 31:58]
  wire [3:0] io_out_0_hi = {temp_7[0],temp_6[0],temp_5[0],temp_4[0]}; // @[Cat.scala 31:58]
  wire [3:0] io_out_1_lo = {temp_3[1],temp_2[1],temp_1[1],temp_0[1]}; // @[Cat.scala 31:58]
  wire [3:0] io_out_1_hi = {temp_7[1],temp_6[1],temp_5[1],temp_4[1]}; // @[Cat.scala 31:58]
  assign io_out_0 = {io_out_0_hi,io_out_0_lo}; // @[Cat.scala 31:58]
  assign io_out_1 = {io_out_1_hi,io_out_1_lo}; // @[Cat.scala 31:58]
endmodule

