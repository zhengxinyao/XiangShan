module PMP(
  input         clock,
  input         reset,
  input         io_distribute_csr_wvalid,
  input  [11:0] io_distribute_csr_waddr,
  input  [63:0] io_distribute_csr_wdata,
  output        io_pmp_0_cfg_l,
  output [1:0]  io_pmp_0_cfg_a,
  output        io_pmp_0_cfg_x,
  output        io_pmp_0_cfg_w,
  output        io_pmp_0_cfg_r,
  output [33:0] io_pmp_0_addr,
  output [35:0] io_pmp_0_mask,
  output        io_pmp_1_cfg_l,
  output [1:0]  io_pmp_1_cfg_a,
  output        io_pmp_1_cfg_x,
  output        io_pmp_1_cfg_w,
  output        io_pmp_1_cfg_r,
  output [33:0] io_pmp_1_addr,
  output [35:0] io_pmp_1_mask,
  output        io_pmp_2_cfg_l,
  output [1:0]  io_pmp_2_cfg_a,
  output        io_pmp_2_cfg_x,
  output        io_pmp_2_cfg_w,
  output        io_pmp_2_cfg_r,
  output [33:0] io_pmp_2_addr,
  output [35:0] io_pmp_2_mask,
  output        io_pmp_3_cfg_l,
  output [1:0]  io_pmp_3_cfg_a,
  output        io_pmp_3_cfg_x,
  output        io_pmp_3_cfg_w,
  output        io_pmp_3_cfg_r,
  output [33:0] io_pmp_3_addr,
  output [35:0] io_pmp_3_mask,
  output        io_pmp_4_cfg_l,
  output [1:0]  io_pmp_4_cfg_a,
  output        io_pmp_4_cfg_x,
  output        io_pmp_4_cfg_w,
  output        io_pmp_4_cfg_r,
  output [33:0] io_pmp_4_addr,
  output [35:0] io_pmp_4_mask,
  output        io_pmp_5_cfg_l,
  output [1:0]  io_pmp_5_cfg_a,
  output        io_pmp_5_cfg_x,
  output        io_pmp_5_cfg_w,
  output        io_pmp_5_cfg_r,
  output [33:0] io_pmp_5_addr,
  output [35:0] io_pmp_5_mask,
  output        io_pmp_6_cfg_l,
  output [1:0]  io_pmp_6_cfg_a,
  output        io_pmp_6_cfg_x,
  output        io_pmp_6_cfg_w,
  output        io_pmp_6_cfg_r,
  output [33:0] io_pmp_6_addr,
  output [35:0] io_pmp_6_mask,
  output        io_pmp_7_cfg_l,
  output [1:0]  io_pmp_7_cfg_a,
  output        io_pmp_7_cfg_x,
  output        io_pmp_7_cfg_w,
  output        io_pmp_7_cfg_r,
  output [33:0] io_pmp_7_addr,
  output [35:0] io_pmp_7_mask,
  output        io_pmp_8_cfg_l,
  output [1:0]  io_pmp_8_cfg_a,
  output        io_pmp_8_cfg_x,
  output        io_pmp_8_cfg_w,
  output        io_pmp_8_cfg_r,
  output [33:0] io_pmp_8_addr,
  output [35:0] io_pmp_8_mask,
  output        io_pmp_9_cfg_l,
  output [1:0]  io_pmp_9_cfg_a,
  output        io_pmp_9_cfg_x,
  output        io_pmp_9_cfg_w,
  output        io_pmp_9_cfg_r,
  output [33:0] io_pmp_9_addr,
  output [35:0] io_pmp_9_mask,
  output        io_pmp_10_cfg_l,
  output [1:0]  io_pmp_10_cfg_a,
  output        io_pmp_10_cfg_x,
  output        io_pmp_10_cfg_w,
  output        io_pmp_10_cfg_r,
  output [33:0] io_pmp_10_addr,
  output [35:0] io_pmp_10_mask,
  output        io_pmp_11_cfg_l,
  output [1:0]  io_pmp_11_cfg_a,
  output        io_pmp_11_cfg_x,
  output        io_pmp_11_cfg_w,
  output        io_pmp_11_cfg_r,
  output [33:0] io_pmp_11_addr,
  output [35:0] io_pmp_11_mask,
  output        io_pmp_12_cfg_l,
  output [1:0]  io_pmp_12_cfg_a,
  output        io_pmp_12_cfg_x,
  output        io_pmp_12_cfg_w,
  output        io_pmp_12_cfg_r,
  output [33:0] io_pmp_12_addr,
  output [35:0] io_pmp_12_mask,
  output        io_pmp_13_cfg_l,
  output [1:0]  io_pmp_13_cfg_a,
  output        io_pmp_13_cfg_x,
  output        io_pmp_13_cfg_w,
  output        io_pmp_13_cfg_r,
  output [33:0] io_pmp_13_addr,
  output [35:0] io_pmp_13_mask,
  output        io_pmp_14_cfg_l,
  output [1:0]  io_pmp_14_cfg_a,
  output        io_pmp_14_cfg_x,
  output        io_pmp_14_cfg_w,
  output        io_pmp_14_cfg_r,
  output [33:0] io_pmp_14_addr,
  output [35:0] io_pmp_14_mask,
  output        io_pmp_15_cfg_l,
  output [1:0]  io_pmp_15_cfg_a,
  output        io_pmp_15_cfg_x,
  output        io_pmp_15_cfg_w,
  output        io_pmp_15_cfg_r,
  output [33:0] io_pmp_15_addr,
  output [35:0] io_pmp_15_mask,
  output        io_pma_0_cfg_c,
  output        io_pma_0_cfg_atomic,
  output [1:0]  io_pma_0_cfg_a,
  output        io_pma_0_cfg_x,
  output        io_pma_0_cfg_w,
  output        io_pma_0_cfg_r,
  output [33:0] io_pma_0_addr,
  output [35:0] io_pma_0_mask,
  output        io_pma_1_cfg_c,
  output        io_pma_1_cfg_atomic,
  output [1:0]  io_pma_1_cfg_a,
  output        io_pma_1_cfg_x,
  output        io_pma_1_cfg_w,
  output        io_pma_1_cfg_r,
  output [33:0] io_pma_1_addr,
  output [35:0] io_pma_1_mask,
  output        io_pma_2_cfg_c,
  output        io_pma_2_cfg_atomic,
  output [1:0]  io_pma_2_cfg_a,
  output        io_pma_2_cfg_x,
  output        io_pma_2_cfg_w,
  output        io_pma_2_cfg_r,
  output [33:0] io_pma_2_addr,
  output [35:0] io_pma_2_mask,
  output        io_pma_3_cfg_c,
  output        io_pma_3_cfg_atomic,
  output [1:0]  io_pma_3_cfg_a,
  output        io_pma_3_cfg_x,
  output        io_pma_3_cfg_w,
  output        io_pma_3_cfg_r,
  output [33:0] io_pma_3_addr,
  output [35:0] io_pma_3_mask,
  output        io_pma_4_cfg_c,
  output        io_pma_4_cfg_atomic,
  output [1:0]  io_pma_4_cfg_a,
  output        io_pma_4_cfg_x,
  output        io_pma_4_cfg_w,
  output        io_pma_4_cfg_r,
  output [33:0] io_pma_4_addr,
  output [35:0] io_pma_4_mask,
  output        io_pma_5_cfg_c,
  output        io_pma_5_cfg_atomic,
  output [1:0]  io_pma_5_cfg_a,
  output        io_pma_5_cfg_x,
  output        io_pma_5_cfg_w,
  output        io_pma_5_cfg_r,
  output [33:0] io_pma_5_addr,
  output [35:0] io_pma_5_mask,
  output        io_pma_6_cfg_c,
  output        io_pma_6_cfg_atomic,
  output [1:0]  io_pma_6_cfg_a,
  output        io_pma_6_cfg_x,
  output        io_pma_6_cfg_w,
  output        io_pma_6_cfg_r,
  output [33:0] io_pma_6_addr,
  output [35:0] io_pma_6_mask,
  output        io_pma_7_cfg_c,
  output        io_pma_7_cfg_atomic,
  output [1:0]  io_pma_7_cfg_a,
  output        io_pma_7_cfg_x,
  output        io_pma_7_cfg_w,
  output        io_pma_7_cfg_r,
  output [33:0] io_pma_7_addr,
  output [35:0] io_pma_7_mask,
  output        io_pma_8_cfg_c,
  output        io_pma_8_cfg_atomic,
  output [1:0]  io_pma_8_cfg_a,
  output        io_pma_8_cfg_x,
  output        io_pma_8_cfg_w,
  output        io_pma_8_cfg_r,
  output [33:0] io_pma_8_addr,
  output [35:0] io_pma_8_mask,
  output        io_pma_9_cfg_c,
  output        io_pma_9_cfg_atomic,
  output [1:0]  io_pma_9_cfg_a,
  output        io_pma_9_cfg_x,
  output        io_pma_9_cfg_w,
  output        io_pma_9_cfg_r,
  output [33:0] io_pma_9_addr,
  output [35:0] io_pma_9_mask,
  output        io_pma_10_cfg_c,
  output        io_pma_10_cfg_atomic,
  output [1:0]  io_pma_10_cfg_a,
  output        io_pma_10_cfg_x,
  output        io_pma_10_cfg_w,
  output        io_pma_10_cfg_r,
  output [33:0] io_pma_10_addr,
  output [35:0] io_pma_10_mask,
  output        io_pma_11_cfg_c,
  output        io_pma_11_cfg_atomic,
  output [1:0]  io_pma_11_cfg_a,
  output        io_pma_11_cfg_x,
  output        io_pma_11_cfg_w,
  output        io_pma_11_cfg_r,
  output [33:0] io_pma_11_addr,
  output [35:0] io_pma_11_mask,
  output        io_pma_12_cfg_c,
  output        io_pma_12_cfg_atomic,
  output [1:0]  io_pma_12_cfg_a,
  output        io_pma_12_cfg_x,
  output        io_pma_12_cfg_w,
  output        io_pma_12_cfg_r,
  output [33:0] io_pma_12_addr,
  output [35:0] io_pma_12_mask,
  output        io_pma_13_cfg_c,
  output        io_pma_13_cfg_atomic,
  output [1:0]  io_pma_13_cfg_a,
  output        io_pma_13_cfg_x,
  output        io_pma_13_cfg_w,
  output        io_pma_13_cfg_r,
  output [33:0] io_pma_13_addr,
  output [35:0] io_pma_13_mask,
  output        io_pma_14_cfg_c,
  output        io_pma_14_cfg_atomic,
  output [1:0]  io_pma_14_cfg_a,
  output        io_pma_14_cfg_x,
  output        io_pma_14_cfg_w,
  output        io_pma_14_cfg_r,
  output [33:0] io_pma_14_addr,
  output [35:0] io_pma_14_mask,
  output        io_pma_15_cfg_c,
  output        io_pma_15_cfg_atomic,
  output [1:0]  io_pma_15_cfg_a,
  output        io_pma_15_cfg_x,
  output        io_pma_15_cfg_w,
  output        io_pma_15_cfg_r,
  output [33:0] io_pma_15_addr,
  output [35:0] io_pma_15_mask
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [63:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [63:0] _RAND_39;
  reg [63:0] _RAND_40;
  reg [63:0] _RAND_41;
  reg [63:0] _RAND_42;
  reg [63:0] _RAND_43;
  reg [63:0] _RAND_44;
  reg [63:0] _RAND_45;
  reg [63:0] _RAND_46;
  reg [63:0] _RAND_47;
  reg [63:0] _RAND_48;
  reg [63:0] _RAND_49;
  reg [63:0] _RAND_50;
  reg [63:0] _RAND_51;
  reg [63:0] _RAND_52;
  reg [63:0] _RAND_53;
  reg [63:0] _RAND_54;
  reg [63:0] _RAND_55;
  reg [63:0] _RAND_56;
  reg [63:0] _RAND_57;
  reg [63:0] _RAND_58;
  reg [63:0] _RAND_59;
  reg [63:0] _RAND_60;
  reg [63:0] _RAND_61;
  reg [63:0] _RAND_62;
  reg [63:0] _RAND_63;
  reg [63:0] _RAND_64;
  reg [63:0] _RAND_65;
  reg [63:0] _RAND_66;
  reg [63:0] _RAND_67;
  reg [63:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] cfgMerged__0; // @[PMP.scala 310:28]
  reg [63:0] cfgMerged__1; // @[PMP.scala 310:28]
  wire [127:0] _cfgs_T = {cfgMerged__1,cfgMerged__0}; // @[PMP.scala 311:44]
  wire [1:0] cfgs__0_a = _cfgs_T[4:3]; // @[PMP.scala 311:44]
  wire  cfgs__0_l = _cfgs_T[7]; // @[PMP.scala 311:44]
  wire [1:0] cfgs__1_a = _cfgs_T[12:11]; // @[PMP.scala 311:44]
  wire  cfgs__1_l = _cfgs_T[15]; // @[PMP.scala 311:44]
  wire [1:0] cfgs__2_a = _cfgs_T[20:19]; // @[PMP.scala 311:44]
  wire  cfgs__2_l = _cfgs_T[23]; // @[PMP.scala 311:44]
  wire [1:0] cfgs__3_a = _cfgs_T[28:27]; // @[PMP.scala 311:44]
  wire  cfgs__3_l = _cfgs_T[31]; // @[PMP.scala 311:44]
  wire [1:0] cfgs__4_a = _cfgs_T[36:35]; // @[PMP.scala 311:44]
  wire  cfgs__4_l = _cfgs_T[39]; // @[PMP.scala 311:44]
  wire [1:0] cfgs__5_a = _cfgs_T[44:43]; // @[PMP.scala 311:44]
  wire  cfgs__5_l = _cfgs_T[47]; // @[PMP.scala 311:44]
  wire [1:0] cfgs__6_a = _cfgs_T[52:51]; // @[PMP.scala 311:44]
  wire  cfgs__6_l = _cfgs_T[55]; // @[PMP.scala 311:44]
  wire [1:0] cfgs__7_a = _cfgs_T[60:59]; // @[PMP.scala 311:44]
  wire  cfgs__7_l = _cfgs_T[63]; // @[PMP.scala 311:44]
  wire [1:0] cfgs__8_a = _cfgs_T[68:67]; // @[PMP.scala 311:44]
  wire  cfgs__8_l = _cfgs_T[71]; // @[PMP.scala 311:44]
  wire [1:0] cfgs__9_a = _cfgs_T[76:75]; // @[PMP.scala 311:44]
  wire  cfgs__9_l = _cfgs_T[79]; // @[PMP.scala 311:44]
  wire [1:0] cfgs__10_a = _cfgs_T[84:83]; // @[PMP.scala 311:44]
  wire  cfgs__10_l = _cfgs_T[87]; // @[PMP.scala 311:44]
  wire [1:0] cfgs__11_a = _cfgs_T[92:91]; // @[PMP.scala 311:44]
  wire  cfgs__11_l = _cfgs_T[95]; // @[PMP.scala 311:44]
  wire [1:0] cfgs__12_a = _cfgs_T[100:99]; // @[PMP.scala 311:44]
  wire  cfgs__12_l = _cfgs_T[103]; // @[PMP.scala 311:44]
  wire [1:0] cfgs__13_a = _cfgs_T[108:107]; // @[PMP.scala 311:44]
  wire  cfgs__13_l = _cfgs_T[111]; // @[PMP.scala 311:44]
  wire [1:0] cfgs__14_a = _cfgs_T[116:115]; // @[PMP.scala 311:44]
  wire  cfgs__14_l = _cfgs_T[119]; // @[PMP.scala 311:44]
  wire [1:0] cfgs__15_a = _cfgs_T[124:123]; // @[PMP.scala 311:44]
  wire  cfgs__15_l = _cfgs_T[127]; // @[PMP.scala 311:44]
  reg [33:0] addr_1_0; // @[PMP.scala 312:23]
  reg [33:0] addr_1_1; // @[PMP.scala 312:23]
  reg [33:0] addr_1_2; // @[PMP.scala 312:23]
  reg [33:0] addr_1_3; // @[PMP.scala 312:23]
  reg [33:0] addr_1_4; // @[PMP.scala 312:23]
  reg [33:0] addr_1_5; // @[PMP.scala 312:23]
  reg [33:0] addr_1_6; // @[PMP.scala 312:23]
  reg [33:0] addr_1_7; // @[PMP.scala 312:23]
  reg [33:0] addr_1_8; // @[PMP.scala 312:23]
  reg [33:0] addr_1_9; // @[PMP.scala 312:23]
  reg [33:0] addr_1_10; // @[PMP.scala 312:23]
  reg [33:0] addr_1_11; // @[PMP.scala 312:23]
  reg [33:0] addr_1_12; // @[PMP.scala 312:23]
  reg [33:0] addr_1_13; // @[PMP.scala 312:23]
  reg [33:0] addr_1_14; // @[PMP.scala 312:23]
  reg [33:0] addr_1_15; // @[PMP.scala 312:23]
  reg [35:0] mask_1_0; // @[PMP.scala 313:23]
  reg [35:0] mask_1_1; // @[PMP.scala 313:23]
  reg [35:0] mask_1_2; // @[PMP.scala 313:23]
  reg [35:0] mask_1_3; // @[PMP.scala 313:23]
  reg [35:0] mask_1_4; // @[PMP.scala 313:23]
  reg [35:0] mask_1_5; // @[PMP.scala 313:23]
  reg [35:0] mask_1_6; // @[PMP.scala 313:23]
  reg [35:0] mask_1_7; // @[PMP.scala 313:23]
  reg [35:0] mask_1_8; // @[PMP.scala 313:23]
  reg [35:0] mask_1_9; // @[PMP.scala 313:23]
  reg [35:0] mask_1_10; // @[PMP.scala 313:23]
  reg [35:0] mask_1_11; // @[PMP.scala 313:23]
  reg [35:0] mask_1_12; // @[PMP.scala 313:23]
  reg [35:0] mask_1_13; // @[PMP.scala 313:23]
  reg [35:0] mask_1_14; // @[PMP.scala 313:23]
  reg [35:0] mask_1_15; // @[PMP.scala 313:23]
  reg [63:0] cfgMerged_1_0; // @[PMP.scala 310:28]
  reg [63:0] cfgMerged_1_1; // @[PMP.scala 310:28]
  wire [127:0] _cfgs_T_113 = {cfgMerged_1_1,cfgMerged_1_0}; // @[PMP.scala 311:44]
  wire [1:0] cfgs_1_0_a = _cfgs_T_113[4:3]; // @[PMP.scala 311:44]
  wire  cfgs_1_0_l = _cfgs_T_113[7]; // @[PMP.scala 311:44]
  wire [1:0] cfgs_1_1_a = _cfgs_T_113[12:11]; // @[PMP.scala 311:44]
  wire  cfgs_1_1_l = _cfgs_T_113[15]; // @[PMP.scala 311:44]
  wire [1:0] cfgs_1_2_a = _cfgs_T_113[20:19]; // @[PMP.scala 311:44]
  wire  cfgs_1_2_l = _cfgs_T_113[23]; // @[PMP.scala 311:44]
  wire [1:0] cfgs_1_3_a = _cfgs_T_113[28:27]; // @[PMP.scala 311:44]
  wire  cfgs_1_3_l = _cfgs_T_113[31]; // @[PMP.scala 311:44]
  wire [1:0] cfgs_1_4_a = _cfgs_T_113[36:35]; // @[PMP.scala 311:44]
  wire  cfgs_1_4_l = _cfgs_T_113[39]; // @[PMP.scala 311:44]
  wire [1:0] cfgs_1_5_a = _cfgs_T_113[44:43]; // @[PMP.scala 311:44]
  wire  cfgs_1_5_l = _cfgs_T_113[47]; // @[PMP.scala 311:44]
  wire [1:0] cfgs_1_6_a = _cfgs_T_113[52:51]; // @[PMP.scala 311:44]
  wire  cfgs_1_6_l = _cfgs_T_113[55]; // @[PMP.scala 311:44]
  wire [1:0] cfgs_1_7_a = _cfgs_T_113[60:59]; // @[PMP.scala 311:44]
  wire  cfgs_1_7_l = _cfgs_T_113[63]; // @[PMP.scala 311:44]
  wire [1:0] cfgs_1_8_a = _cfgs_T_113[68:67]; // @[PMP.scala 311:44]
  wire  cfgs_1_8_l = _cfgs_T_113[71]; // @[PMP.scala 311:44]
  wire [1:0] cfgs_1_9_a = _cfgs_T_113[76:75]; // @[PMP.scala 311:44]
  wire  cfgs_1_9_l = _cfgs_T_113[79]; // @[PMP.scala 311:44]
  wire [1:0] cfgs_1_10_a = _cfgs_T_113[84:83]; // @[PMP.scala 311:44]
  wire  cfgs_1_10_l = _cfgs_T_113[87]; // @[PMP.scala 311:44]
  wire [1:0] cfgs_1_11_a = _cfgs_T_113[92:91]; // @[PMP.scala 311:44]
  wire  cfgs_1_11_l = _cfgs_T_113[95]; // @[PMP.scala 311:44]
  wire [1:0] cfgs_1_12_a = _cfgs_T_113[100:99]; // @[PMP.scala 311:44]
  wire  cfgs_1_12_l = _cfgs_T_113[103]; // @[PMP.scala 311:44]
  wire [1:0] cfgs_1_13_a = _cfgs_T_113[108:107]; // @[PMP.scala 311:44]
  wire  cfgs_1_13_l = _cfgs_T_113[111]; // @[PMP.scala 311:44]
  wire [1:0] cfgs_1_14_a = _cfgs_T_113[116:115]; // @[PMP.scala 311:44]
  wire  cfgs_1_14_l = _cfgs_T_113[119]; // @[PMP.scala 311:44]
  wire [1:0] cfgs_1_15_a = _cfgs_T_113[124:123]; // @[PMP.scala 311:44]
  wire  cfgs_1_15_l = _cfgs_T_113[127]; // @[PMP.scala 311:44]
  reg [33:0] addr_2_0; // @[PMP.scala 312:23]
  reg [33:0] addr_2_1; // @[PMP.scala 312:23]
  reg [33:0] addr_2_2; // @[PMP.scala 312:23]
  reg [33:0] addr_2_3; // @[PMP.scala 312:23]
  reg [33:0] addr_2_4; // @[PMP.scala 312:23]
  reg [33:0] addr_2_5; // @[PMP.scala 312:23]
  reg [33:0] addr_2_6; // @[PMP.scala 312:23]
  reg [33:0] addr_2_7; // @[PMP.scala 312:23]
  reg [33:0] addr_2_8; // @[PMP.scala 312:23]
  reg [33:0] addr_2_9; // @[PMP.scala 312:23]
  reg [33:0] addr_2_10; // @[PMP.scala 312:23]
  reg [33:0] addr_2_11; // @[PMP.scala 312:23]
  reg [33:0] addr_2_12; // @[PMP.scala 312:23]
  reg [33:0] addr_2_13; // @[PMP.scala 312:23]
  reg [33:0] addr_2_14; // @[PMP.scala 312:23]
  reg [33:0] addr_2_15; // @[PMP.scala 312:23]
  reg [35:0] mask_2_0; // @[PMP.scala 313:23]
  reg [35:0] mask_2_1; // @[PMP.scala 313:23]
  reg [35:0] mask_2_2; // @[PMP.scala 313:23]
  reg [35:0] mask_2_3; // @[PMP.scala 313:23]
  reg [35:0] mask_2_4; // @[PMP.scala 313:23]
  reg [35:0] mask_2_5; // @[PMP.scala 313:23]
  reg [35:0] mask_2_6; // @[PMP.scala 313:23]
  reg [35:0] mask_2_7; // @[PMP.scala 313:23]
  reg [35:0] mask_2_8; // @[PMP.scala 313:23]
  reg [35:0] mask_2_9; // @[PMP.scala 313:23]
  reg [35:0] mask_2_10; // @[PMP.scala 313:23]
  reg [35:0] mask_2_11; // @[PMP.scala 313:23]
  reg [35:0] mask_2_12; // @[PMP.scala 313:23]
  reg [35:0] mask_2_13; // @[PMP.scala 313:23]
  reg [35:0] mask_2_14; // @[PMP.scala 313:23]
  reg [35:0] mask_2_15; // @[PMP.scala 313:23]
  reg [63:0] wdata_reg; // @[Reg.scala 16:16]
  reg  wen_reg; // @[RegMap.scala 55:30]
  wire  _addr_3_mask_3_T = cfgs_1_4_a == 2'h1; // @[PMP.scala 53:15]
  wire  _addr_3_mask_3_T_2 = cfgs_1_3_l | cfgs_1_4_l & _addr_3_mask_3_T; // @[PMP.scala 61:51]
  wire  _addr_3_mask_3_T_3 = ~_addr_3_mask_3_T_2; // @[PMP.scala 271:17]
  wire [64:0] _addr_3_mask_3_match_mask_c_addr_T_1 = {wdata_reg,cfgs_1_3_a[0]}; // @[Cat.scala 31:58]
  wire [64:0] addr_3_mask_3_match_mask_c_addr = _addr_3_mask_3_match_mask_c_addr_T_1 | 65'h3ff; // @[PMP.scala 86:50]
  wire [64:0] _addr_3_mask_3_T_5 = addr_3_mask_3_match_mask_c_addr + 65'h1; // @[PMP.scala 87:49]
  wire [64:0] _addr_3_mask_3_T_6 = ~_addr_3_mask_3_T_5; // @[PMP.scala 87:29]
  wire [64:0] _addr_3_mask_3_T_7 = addr_3_mask_3_match_mask_c_addr & _addr_3_mask_3_T_6; // @[PMP.scala 87:27]
  wire [66:0] _addr_3_mask_3_T_8 = {_addr_3_mask_3_T_7,2'h3}; // @[Cat.scala 31:58]
  wire [66:0] _addr_3_mask_3_T_9 = ~_addr_3_mask_3_T_2 ? _addr_3_mask_3_T_8 : {{31'd0}, mask_2_3}; // @[PMP.scala 271:16]
  wire [63:0] _addr_3_T_8 = _addr_3_mask_3_T_3 ? wdata_reg : {{30'd0}, addr_2_3}; // @[PMP.scala 272:8]
  wire [66:0] _GEN_1 = wen_reg ? _addr_3_mask_3_T_9 : {{31'd0}, mask_2_3}; // @[PMP.scala 271:10 313:23 RegMap.scala 56:24]
  wire [63:0] _GEN_2 = wen_reg ? _addr_3_T_8 : {{30'd0}, addr_2_3}; // @[PMP.scala 312:23 RegMap.scala 56:{24,28}]
  reg  wen_reg_1; // @[RegMap.scala 55:30]
  wire  _addr_7_mask_7_T = cfgs_1_8_a == 2'h1; // @[PMP.scala 53:15]
  wire  _addr_7_mask_7_T_2 = cfgs_1_7_l | cfgs_1_8_l & _addr_7_mask_7_T; // @[PMP.scala 61:51]
  wire  _addr_7_mask_7_T_3 = ~_addr_7_mask_7_T_2; // @[PMP.scala 271:17]
  wire [64:0] _addr_7_mask_7_match_mask_c_addr_T_1 = {wdata_reg,cfgs_1_7_a[0]}; // @[Cat.scala 31:58]
  wire [64:0] addr_7_mask_7_match_mask_c_addr = _addr_7_mask_7_match_mask_c_addr_T_1 | 65'h3ff; // @[PMP.scala 86:50]
  wire [64:0] _addr_7_mask_7_T_5 = addr_7_mask_7_match_mask_c_addr + 65'h1; // @[PMP.scala 87:49]
  wire [64:0] _addr_7_mask_7_T_6 = ~_addr_7_mask_7_T_5; // @[PMP.scala 87:29]
  wire [64:0] _addr_7_mask_7_T_7 = addr_7_mask_7_match_mask_c_addr & _addr_7_mask_7_T_6; // @[PMP.scala 87:27]
  wire [66:0] _addr_7_mask_7_T_8 = {_addr_7_mask_7_T_7,2'h3}; // @[Cat.scala 31:58]
  wire [66:0] _addr_7_mask_7_T_9 = ~_addr_7_mask_7_T_2 ? _addr_7_mask_7_T_8 : {{31'd0}, mask_2_7}; // @[PMP.scala 271:16]
  wire [63:0] _addr_7_T_8 = _addr_7_mask_7_T_3 ? wdata_reg : {{30'd0}, addr_2_7}; // @[PMP.scala 272:8]
  wire [66:0] _GEN_3 = wen_reg_1 ? _addr_7_mask_7_T_9 : {{31'd0}, mask_2_7}; // @[PMP.scala 271:10 313:23 RegMap.scala 56:24]
  wire [63:0] _GEN_4 = wen_reg_1 ? _addr_7_T_8 : {{30'd0}, addr_2_7}; // @[PMP.scala 312:23 RegMap.scala 56:{24,28}]
  reg  wen_reg_2; // @[RegMap.scala 55:30]
  wire  _addr_1_mask_1_T = cfgs__2_a == 2'h1; // @[PMP.scala 53:15]
  wire  _addr_1_mask_1_T_2 = cfgs__1_l | cfgs__2_l & _addr_1_mask_1_T; // @[PMP.scala 61:51]
  wire  _addr_1_mask_1_T_3 = ~_addr_1_mask_1_T_2; // @[PMP.scala 271:17]
  wire [64:0] _addr_1_mask_1_match_mask_c_addr_T_1 = {wdata_reg,cfgs__1_a[0]}; // @[Cat.scala 31:58]
  wire [64:0] addr_1_mask_1_match_mask_c_addr = _addr_1_mask_1_match_mask_c_addr_T_1 | 65'h3ff; // @[PMP.scala 86:50]
  wire [64:0] _addr_1_mask_1_T_5 = addr_1_mask_1_match_mask_c_addr + 65'h1; // @[PMP.scala 87:49]
  wire [64:0] _addr_1_mask_1_T_6 = ~_addr_1_mask_1_T_5; // @[PMP.scala 87:29]
  wire [64:0] _addr_1_mask_1_T_7 = addr_1_mask_1_match_mask_c_addr & _addr_1_mask_1_T_6; // @[PMP.scala 87:27]
  wire [66:0] _addr_1_mask_1_T_8 = {_addr_1_mask_1_T_7,2'h3}; // @[Cat.scala 31:58]
  wire [66:0] _addr_1_mask_1_T_9 = ~_addr_1_mask_1_T_2 ? _addr_1_mask_1_T_8 : {{31'd0}, mask_1_1}; // @[PMP.scala 271:16]
  wire [63:0] _addr_1_T_8 = _addr_1_mask_1_T_3 ? wdata_reg : {{30'd0}, addr_1_1}; // @[PMP.scala 272:8]
  wire [66:0] _GEN_5 = wen_reg_2 ? _addr_1_mask_1_T_9 : {{31'd0}, mask_1_1}; // @[PMP.scala 271:10 313:23 RegMap.scala 56:24]
  wire [63:0] _GEN_6 = wen_reg_2 ? _addr_1_T_8 : {{30'd0}, addr_1_1}; // @[PMP.scala 312:23 RegMap.scala 56:{24,28}]
  reg  wen_reg_3; // @[RegMap.scala 55:30]
  wire  cfgMerged_1_cfg_wm_tmp_r = wdata_reg[0]; // @[PMP.scala 93:61]
  wire  cfgMerged_1_cfg_wm_tmp_w = wdata_reg[1]; // @[PMP.scala 93:61]
  wire  cfgMerged_1_cfg_wm_tmp_x = wdata_reg[2]; // @[PMP.scala 93:61]
  wire [1:0] cfgMerged_1_cfg_wm_tmp_a = wdata_reg[4:3]; // @[PMP.scala 93:61]
  wire  cfgMerged_1_cfg_wm_tmp_atomic = wdata_reg[5]; // @[PMP.scala 93:61]
  wire  cfgMerged_1_cfg_wm_tmp_c = wdata_reg[6]; // @[PMP.scala 93:61]
  wire  cfgMerged_1_cfg_wm_tmp_l = wdata_reg[7]; // @[PMP.scala 93:61]
  wire  _cfgMerged_1_cfgVec_0_a_T_1 = |cfgMerged_1_cfg_wm_tmp_a; // @[PMP.scala 97:80]
  wire [1:0] _cfgMerged_1_cfgVec_0_a_T_2 = {cfgMerged_1_cfg_wm_tmp_a[1],_cfgMerged_1_cfgVec_0_a_T_1}; // @[Cat.scala 31:58]
  wire [1:0] cfgMerged_1_cfgVec__0_a = ~cfgMerged_1_cfg_wm_tmp_l ? _cfgMerged_1_cfgVec_0_a_T_2 :
    cfgMerged_1_cfg_wm_tmp_a; // @[PMP.scala 94:17 95:29 97:41]
  wire [34:0] _cfgMerged_1_mask_8_match_mask_c_addr_T_1 = {addr_1_8,cfgMerged_1_cfgVec__0_a[0]}; // @[Cat.scala 31:58]
  wire [34:0] cfgMerged_1_mask_8_match_mask_c_addr = _cfgMerged_1_mask_8_match_mask_c_addr_T_1 | 35'h3ff; // @[PMP.scala 86:50]
  wire [34:0] _cfgMerged_1_mask_8_T_1 = cfgMerged_1_mask_8_match_mask_c_addr + 35'h1; // @[PMP.scala 87:49]
  wire [34:0] _cfgMerged_1_mask_8_T_2 = ~_cfgMerged_1_mask_8_T_1; // @[PMP.scala 87:29]
  wire [34:0] _cfgMerged_1_mask_8_T_3 = cfgMerged_1_mask_8_match_mask_c_addr & _cfgMerged_1_mask_8_T_2; // @[PMP.scala 87:27]
  wire [36:0] _cfgMerged_1_mask_8_T_4 = {_cfgMerged_1_mask_8_T_3,2'h3}; // @[Cat.scala 31:58]
  wire [36:0] _GEN_7 = cfgMerged_1_cfgVec__0_a[1] ? _cfgMerged_1_mask_8_T_4 : {{1'd0}, mask_1_8}; // @[PMP.scala 313:23 98:36 99:27]
  wire  cfgMerged_1_cfgVec__0_w = ~cfgMerged_1_cfg_wm_tmp_l ? cfgMerged_1_cfg_wm_tmp_w & cfgMerged_1_cfg_wm_tmp_r :
    cfgMerged_1_cfg_wm_tmp_w; // @[PMP.scala 94:17 95:29 96:21]
  wire [36:0] _GEN_10 = ~cfgMerged_1_cfg_wm_tmp_l ? _GEN_7 : {{1'd0}, mask_1_8}; // @[PMP.scala 313:23 95:29]
  wire  cfgMerged_1_cfg_wm_tmp_1_r = wdata_reg[8]; // @[PMP.scala 93:61]
  wire  cfgMerged_1_cfg_wm_tmp_1_w = wdata_reg[9]; // @[PMP.scala 93:61]
  wire  cfgMerged_1_cfg_wm_tmp_1_x = wdata_reg[10]; // @[PMP.scala 93:61]
  wire [1:0] cfgMerged_1_cfg_wm_tmp_1_a = wdata_reg[12:11]; // @[PMP.scala 93:61]
  wire  cfgMerged_1_cfg_wm_tmp_1_atomic = wdata_reg[13]; // @[PMP.scala 93:61]
  wire  cfgMerged_1_cfg_wm_tmp_1_c = wdata_reg[14]; // @[PMP.scala 93:61]
  wire  cfgMerged_1_cfg_wm_tmp_1_l = wdata_reg[15]; // @[PMP.scala 93:61]
  wire  _cfgMerged_1_cfgVec_1_a_T_1 = |cfgMerged_1_cfg_wm_tmp_1_a; // @[PMP.scala 97:80]
  wire [1:0] _cfgMerged_1_cfgVec_1_a_T_2 = {cfgMerged_1_cfg_wm_tmp_1_a[1],_cfgMerged_1_cfgVec_1_a_T_1}; // @[Cat.scala 31:58]
  wire [1:0] cfgMerged_1_cfgVec__1_a = ~cfgMerged_1_cfg_wm_tmp_1_l ? _cfgMerged_1_cfgVec_1_a_T_2 :
    cfgMerged_1_cfg_wm_tmp_1_a; // @[PMP.scala 94:17 95:29 97:41]
  wire [34:0] _cfgMerged_1_mask_9_match_mask_c_addr_T_1 = {addr_1_9,cfgMerged_1_cfgVec__1_a[0]}; // @[Cat.scala 31:58]
  wire [34:0] cfgMerged_1_mask_9_match_mask_c_addr = _cfgMerged_1_mask_9_match_mask_c_addr_T_1 | 35'h3ff; // @[PMP.scala 86:50]
  wire [34:0] _cfgMerged_1_mask_9_T_1 = cfgMerged_1_mask_9_match_mask_c_addr + 35'h1; // @[PMP.scala 87:49]
  wire [34:0] _cfgMerged_1_mask_9_T_2 = ~_cfgMerged_1_mask_9_T_1; // @[PMP.scala 87:29]
  wire [34:0] _cfgMerged_1_mask_9_T_3 = cfgMerged_1_mask_9_match_mask_c_addr & _cfgMerged_1_mask_9_T_2; // @[PMP.scala 87:27]
  wire [36:0] _cfgMerged_1_mask_9_T_4 = {_cfgMerged_1_mask_9_T_3,2'h3}; // @[Cat.scala 31:58]
  wire [36:0] _GEN_11 = cfgMerged_1_cfgVec__1_a[1] ? _cfgMerged_1_mask_9_T_4 : {{1'd0}, mask_1_9}; // @[PMP.scala 313:23 98:36 99:27]
  wire  cfgMerged_1_cfgVec__1_w = ~cfgMerged_1_cfg_wm_tmp_1_l ? cfgMerged_1_cfg_wm_tmp_1_w &
    cfgMerged_1_cfg_wm_tmp_1_r : cfgMerged_1_cfg_wm_tmp_1_w; // @[PMP.scala 94:17 95:29 96:21]
  wire [36:0] _GEN_14 = ~cfgMerged_1_cfg_wm_tmp_1_l ? _GEN_11 : {{1'd0}, mask_1_9}; // @[PMP.scala 313:23 95:29]
  wire  cfgMerged_1_cfg_wm_tmp_2_r = wdata_reg[16]; // @[PMP.scala 93:61]
  wire  cfgMerged_1_cfg_wm_tmp_2_w = wdata_reg[17]; // @[PMP.scala 93:61]
  wire  cfgMerged_1_cfg_wm_tmp_2_x = wdata_reg[18]; // @[PMP.scala 93:61]
  wire [1:0] cfgMerged_1_cfg_wm_tmp_2_a = wdata_reg[20:19]; // @[PMP.scala 93:61]
  wire  cfgMerged_1_cfg_wm_tmp_2_atomic = wdata_reg[21]; // @[PMP.scala 93:61]
  wire  cfgMerged_1_cfg_wm_tmp_2_c = wdata_reg[22]; // @[PMP.scala 93:61]
  wire  cfgMerged_1_cfg_wm_tmp_2_l = wdata_reg[23]; // @[PMP.scala 93:61]
  wire  _cfgMerged_1_cfgVec_2_a_T_1 = |cfgMerged_1_cfg_wm_tmp_2_a; // @[PMP.scala 97:80]
  wire [1:0] _cfgMerged_1_cfgVec_2_a_T_2 = {cfgMerged_1_cfg_wm_tmp_2_a[1],_cfgMerged_1_cfgVec_2_a_T_1}; // @[Cat.scala 31:58]
  wire [1:0] cfgMerged_1_cfgVec__2_a = ~cfgMerged_1_cfg_wm_tmp_2_l ? _cfgMerged_1_cfgVec_2_a_T_2 :
    cfgMerged_1_cfg_wm_tmp_2_a; // @[PMP.scala 94:17 95:29 97:41]
  wire [34:0] _cfgMerged_1_mask_10_match_mask_c_addr_T_1 = {addr_1_10,cfgMerged_1_cfgVec__2_a[0]}; // @[Cat.scala 31:58]
  wire [34:0] cfgMerged_1_mask_10_match_mask_c_addr = _cfgMerged_1_mask_10_match_mask_c_addr_T_1 | 35'h3ff; // @[PMP.scala 86:50]
  wire [34:0] _cfgMerged_1_mask_10_T_1 = cfgMerged_1_mask_10_match_mask_c_addr + 35'h1; // @[PMP.scala 87:49]
  wire [34:0] _cfgMerged_1_mask_10_T_2 = ~_cfgMerged_1_mask_10_T_1; // @[PMP.scala 87:29]
  wire [34:0] _cfgMerged_1_mask_10_T_3 = cfgMerged_1_mask_10_match_mask_c_addr & _cfgMerged_1_mask_10_T_2; // @[PMP.scala 87:27]
  wire [36:0] _cfgMerged_1_mask_10_T_4 = {_cfgMerged_1_mask_10_T_3,2'h3}; // @[Cat.scala 31:58]
  wire [36:0] _GEN_15 = cfgMerged_1_cfgVec__2_a[1] ? _cfgMerged_1_mask_10_T_4 : {{1'd0}, mask_1_10}; // @[PMP.scala 313:23 98:36 99:27]
  wire  cfgMerged_1_cfgVec__2_w = ~cfgMerged_1_cfg_wm_tmp_2_l ? cfgMerged_1_cfg_wm_tmp_2_w &
    cfgMerged_1_cfg_wm_tmp_2_r : cfgMerged_1_cfg_wm_tmp_2_w; // @[PMP.scala 94:17 95:29 96:21]
  wire [36:0] _GEN_18 = ~cfgMerged_1_cfg_wm_tmp_2_l ? _GEN_15 : {{1'd0}, mask_1_10}; // @[PMP.scala 313:23 95:29]
  wire  cfgMerged_1_cfg_wm_tmp_3_r = wdata_reg[24]; // @[PMP.scala 93:61]
  wire  cfgMerged_1_cfg_wm_tmp_3_w = wdata_reg[25]; // @[PMP.scala 93:61]
  wire  cfgMerged_1_cfg_wm_tmp_3_x = wdata_reg[26]; // @[PMP.scala 93:61]
  wire [1:0] cfgMerged_1_cfg_wm_tmp_3_a = wdata_reg[28:27]; // @[PMP.scala 93:61]
  wire  cfgMerged_1_cfg_wm_tmp_3_atomic = wdata_reg[29]; // @[PMP.scala 93:61]
  wire  cfgMerged_1_cfg_wm_tmp_3_c = wdata_reg[30]; // @[PMP.scala 93:61]
  wire  cfgMerged_1_cfg_wm_tmp_3_l = wdata_reg[31]; // @[PMP.scala 93:61]
  wire  _cfgMerged_1_cfgVec_3_a_T_1 = |cfgMerged_1_cfg_wm_tmp_3_a; // @[PMP.scala 97:80]
  wire [1:0] _cfgMerged_1_cfgVec_3_a_T_2 = {cfgMerged_1_cfg_wm_tmp_3_a[1],_cfgMerged_1_cfgVec_3_a_T_1}; // @[Cat.scala 31:58]
  wire [1:0] cfgMerged_1_cfgVec__3_a = ~cfgMerged_1_cfg_wm_tmp_3_l ? _cfgMerged_1_cfgVec_3_a_T_2 :
    cfgMerged_1_cfg_wm_tmp_3_a; // @[PMP.scala 94:17 95:29 97:41]
  wire [34:0] _cfgMerged_1_mask_11_match_mask_c_addr_T_1 = {addr_1_11,cfgMerged_1_cfgVec__3_a[0]}; // @[Cat.scala 31:58]
  wire [34:0] cfgMerged_1_mask_11_match_mask_c_addr = _cfgMerged_1_mask_11_match_mask_c_addr_T_1 | 35'h3ff; // @[PMP.scala 86:50]
  wire [34:0] _cfgMerged_1_mask_11_T_1 = cfgMerged_1_mask_11_match_mask_c_addr + 35'h1; // @[PMP.scala 87:49]
  wire [34:0] _cfgMerged_1_mask_11_T_2 = ~_cfgMerged_1_mask_11_T_1; // @[PMP.scala 87:29]
  wire [34:0] _cfgMerged_1_mask_11_T_3 = cfgMerged_1_mask_11_match_mask_c_addr & _cfgMerged_1_mask_11_T_2; // @[PMP.scala 87:27]
  wire [36:0] _cfgMerged_1_mask_11_T_4 = {_cfgMerged_1_mask_11_T_3,2'h3}; // @[Cat.scala 31:58]
  wire [36:0] _GEN_19 = cfgMerged_1_cfgVec__3_a[1] ? _cfgMerged_1_mask_11_T_4 : {{1'd0}, mask_1_11}; // @[PMP.scala 313:23 98:36 99:27]
  wire  cfgMerged_1_cfgVec__3_w = ~cfgMerged_1_cfg_wm_tmp_3_l ? cfgMerged_1_cfg_wm_tmp_3_w &
    cfgMerged_1_cfg_wm_tmp_3_r : cfgMerged_1_cfg_wm_tmp_3_w; // @[PMP.scala 94:17 95:29 96:21]
  wire [36:0] _GEN_22 = ~cfgMerged_1_cfg_wm_tmp_3_l ? _GEN_19 : {{1'd0}, mask_1_11}; // @[PMP.scala 313:23 95:29]
  wire  cfgMerged_1_cfg_wm_tmp_4_r = wdata_reg[32]; // @[PMP.scala 93:61]
  wire  cfgMerged_1_cfg_wm_tmp_4_w = wdata_reg[33]; // @[PMP.scala 93:61]
  wire  cfgMerged_1_cfg_wm_tmp_4_x = wdata_reg[34]; // @[PMP.scala 93:61]
  wire [1:0] cfgMerged_1_cfg_wm_tmp_4_a = wdata_reg[36:35]; // @[PMP.scala 93:61]
  wire  cfgMerged_1_cfg_wm_tmp_4_atomic = wdata_reg[37]; // @[PMP.scala 93:61]
  wire  cfgMerged_1_cfg_wm_tmp_4_c = wdata_reg[38]; // @[PMP.scala 93:61]
  wire  cfgMerged_1_cfg_wm_tmp_4_l = wdata_reg[39]; // @[PMP.scala 93:61]
  wire  _cfgMerged_1_cfgVec_4_a_T_1 = |cfgMerged_1_cfg_wm_tmp_4_a; // @[PMP.scala 97:80]
  wire [1:0] _cfgMerged_1_cfgVec_4_a_T_2 = {cfgMerged_1_cfg_wm_tmp_4_a[1],_cfgMerged_1_cfgVec_4_a_T_1}; // @[Cat.scala 31:58]
  wire [1:0] cfgMerged_1_cfgVec__4_a = ~cfgMerged_1_cfg_wm_tmp_4_l ? _cfgMerged_1_cfgVec_4_a_T_2 :
    cfgMerged_1_cfg_wm_tmp_4_a; // @[PMP.scala 94:17 95:29 97:41]
  wire [34:0] _cfgMerged_1_mask_12_match_mask_c_addr_T_1 = {addr_1_12,cfgMerged_1_cfgVec__4_a[0]}; // @[Cat.scala 31:58]
  wire [34:0] cfgMerged_1_mask_12_match_mask_c_addr = _cfgMerged_1_mask_12_match_mask_c_addr_T_1 | 35'h3ff; // @[PMP.scala 86:50]
  wire [34:0] _cfgMerged_1_mask_12_T_1 = cfgMerged_1_mask_12_match_mask_c_addr + 35'h1; // @[PMP.scala 87:49]
  wire [34:0] _cfgMerged_1_mask_12_T_2 = ~_cfgMerged_1_mask_12_T_1; // @[PMP.scala 87:29]
  wire [34:0] _cfgMerged_1_mask_12_T_3 = cfgMerged_1_mask_12_match_mask_c_addr & _cfgMerged_1_mask_12_T_2; // @[PMP.scala 87:27]
  wire [36:0] _cfgMerged_1_mask_12_T_4 = {_cfgMerged_1_mask_12_T_3,2'h3}; // @[Cat.scala 31:58]
  wire [36:0] _GEN_23 = cfgMerged_1_cfgVec__4_a[1] ? _cfgMerged_1_mask_12_T_4 : {{1'd0}, mask_1_12}; // @[PMP.scala 313:23 98:36 99:27]
  wire  cfgMerged_1_cfgVec__4_w = ~cfgMerged_1_cfg_wm_tmp_4_l ? cfgMerged_1_cfg_wm_tmp_4_w &
    cfgMerged_1_cfg_wm_tmp_4_r : cfgMerged_1_cfg_wm_tmp_4_w; // @[PMP.scala 94:17 95:29 96:21]
  wire [36:0] _GEN_26 = ~cfgMerged_1_cfg_wm_tmp_4_l ? _GEN_23 : {{1'd0}, mask_1_12}; // @[PMP.scala 313:23 95:29]
  wire  cfgMerged_1_cfg_wm_tmp_5_r = wdata_reg[40]; // @[PMP.scala 93:61]
  wire  cfgMerged_1_cfg_wm_tmp_5_w = wdata_reg[41]; // @[PMP.scala 93:61]
  wire  cfgMerged_1_cfg_wm_tmp_5_x = wdata_reg[42]; // @[PMP.scala 93:61]
  wire [1:0] cfgMerged_1_cfg_wm_tmp_5_a = wdata_reg[44:43]; // @[PMP.scala 93:61]
  wire  cfgMerged_1_cfg_wm_tmp_5_atomic = wdata_reg[45]; // @[PMP.scala 93:61]
  wire  cfgMerged_1_cfg_wm_tmp_5_c = wdata_reg[46]; // @[PMP.scala 93:61]
  wire  cfgMerged_1_cfg_wm_tmp_5_l = wdata_reg[47]; // @[PMP.scala 93:61]
  wire  _cfgMerged_1_cfgVec_5_a_T_1 = |cfgMerged_1_cfg_wm_tmp_5_a; // @[PMP.scala 97:80]
  wire [1:0] _cfgMerged_1_cfgVec_5_a_T_2 = {cfgMerged_1_cfg_wm_tmp_5_a[1],_cfgMerged_1_cfgVec_5_a_T_1}; // @[Cat.scala 31:58]
  wire [1:0] cfgMerged_1_cfgVec__5_a = ~cfgMerged_1_cfg_wm_tmp_5_l ? _cfgMerged_1_cfgVec_5_a_T_2 :
    cfgMerged_1_cfg_wm_tmp_5_a; // @[PMP.scala 94:17 95:29 97:41]
  wire [34:0] _cfgMerged_1_mask_13_match_mask_c_addr_T_1 = {addr_1_13,cfgMerged_1_cfgVec__5_a[0]}; // @[Cat.scala 31:58]
  wire [34:0] cfgMerged_1_mask_13_match_mask_c_addr = _cfgMerged_1_mask_13_match_mask_c_addr_T_1 | 35'h3ff; // @[PMP.scala 86:50]
  wire [34:0] _cfgMerged_1_mask_13_T_1 = cfgMerged_1_mask_13_match_mask_c_addr + 35'h1; // @[PMP.scala 87:49]
  wire [34:0] _cfgMerged_1_mask_13_T_2 = ~_cfgMerged_1_mask_13_T_1; // @[PMP.scala 87:29]
  wire [34:0] _cfgMerged_1_mask_13_T_3 = cfgMerged_1_mask_13_match_mask_c_addr & _cfgMerged_1_mask_13_T_2; // @[PMP.scala 87:27]
  wire [36:0] _cfgMerged_1_mask_13_T_4 = {_cfgMerged_1_mask_13_T_3,2'h3}; // @[Cat.scala 31:58]
  wire [36:0] _GEN_27 = cfgMerged_1_cfgVec__5_a[1] ? _cfgMerged_1_mask_13_T_4 : {{1'd0}, mask_1_13}; // @[PMP.scala 313:23 98:36 99:27]
  wire  cfgMerged_1_cfgVec__5_w = ~cfgMerged_1_cfg_wm_tmp_5_l ? cfgMerged_1_cfg_wm_tmp_5_w &
    cfgMerged_1_cfg_wm_tmp_5_r : cfgMerged_1_cfg_wm_tmp_5_w; // @[PMP.scala 94:17 95:29 96:21]
  wire [36:0] _GEN_30 = ~cfgMerged_1_cfg_wm_tmp_5_l ? _GEN_27 : {{1'd0}, mask_1_13}; // @[PMP.scala 313:23 95:29]
  wire  cfgMerged_1_cfg_wm_tmp_6_r = wdata_reg[48]; // @[PMP.scala 93:61]
  wire  cfgMerged_1_cfg_wm_tmp_6_w = wdata_reg[49]; // @[PMP.scala 93:61]
  wire  cfgMerged_1_cfg_wm_tmp_6_x = wdata_reg[50]; // @[PMP.scala 93:61]
  wire [1:0] cfgMerged_1_cfg_wm_tmp_6_a = wdata_reg[52:51]; // @[PMP.scala 93:61]
  wire  cfgMerged_1_cfg_wm_tmp_6_atomic = wdata_reg[53]; // @[PMP.scala 93:61]
  wire  cfgMerged_1_cfg_wm_tmp_6_c = wdata_reg[54]; // @[PMP.scala 93:61]
  wire  cfgMerged_1_cfg_wm_tmp_6_l = wdata_reg[55]; // @[PMP.scala 93:61]
  wire  _cfgMerged_1_cfgVec_6_a_T_1 = |cfgMerged_1_cfg_wm_tmp_6_a; // @[PMP.scala 97:80]
  wire [1:0] _cfgMerged_1_cfgVec_6_a_T_2 = {cfgMerged_1_cfg_wm_tmp_6_a[1],_cfgMerged_1_cfgVec_6_a_T_1}; // @[Cat.scala 31:58]
  wire [1:0] cfgMerged_1_cfgVec__6_a = ~cfgMerged_1_cfg_wm_tmp_6_l ? _cfgMerged_1_cfgVec_6_a_T_2 :
    cfgMerged_1_cfg_wm_tmp_6_a; // @[PMP.scala 94:17 95:29 97:41]
  wire [34:0] _cfgMerged_1_mask_14_match_mask_c_addr_T_1 = {addr_1_14,cfgMerged_1_cfgVec__6_a[0]}; // @[Cat.scala 31:58]
  wire [34:0] cfgMerged_1_mask_14_match_mask_c_addr = _cfgMerged_1_mask_14_match_mask_c_addr_T_1 | 35'h3ff; // @[PMP.scala 86:50]
  wire [34:0] _cfgMerged_1_mask_14_T_1 = cfgMerged_1_mask_14_match_mask_c_addr + 35'h1; // @[PMP.scala 87:49]
  wire [34:0] _cfgMerged_1_mask_14_T_2 = ~_cfgMerged_1_mask_14_T_1; // @[PMP.scala 87:29]
  wire [34:0] _cfgMerged_1_mask_14_T_3 = cfgMerged_1_mask_14_match_mask_c_addr & _cfgMerged_1_mask_14_T_2; // @[PMP.scala 87:27]
  wire [36:0] _cfgMerged_1_mask_14_T_4 = {_cfgMerged_1_mask_14_T_3,2'h3}; // @[Cat.scala 31:58]
  wire [36:0] _GEN_31 = cfgMerged_1_cfgVec__6_a[1] ? _cfgMerged_1_mask_14_T_4 : {{1'd0}, mask_1_14}; // @[PMP.scala 313:23 98:36 99:27]
  wire  cfgMerged_1_cfgVec__6_w = ~cfgMerged_1_cfg_wm_tmp_6_l ? cfgMerged_1_cfg_wm_tmp_6_w &
    cfgMerged_1_cfg_wm_tmp_6_r : cfgMerged_1_cfg_wm_tmp_6_w; // @[PMP.scala 94:17 95:29 96:21]
  wire [36:0] _GEN_34 = ~cfgMerged_1_cfg_wm_tmp_6_l ? _GEN_31 : {{1'd0}, mask_1_14}; // @[PMP.scala 313:23 95:29]
  wire  cfgMerged_1_cfg_wm_tmp_7_r = wdata_reg[56]; // @[PMP.scala 93:61]
  wire  cfgMerged_1_cfg_wm_tmp_7_w = wdata_reg[57]; // @[PMP.scala 93:61]
  wire  cfgMerged_1_cfg_wm_tmp_7_x = wdata_reg[58]; // @[PMP.scala 93:61]
  wire [1:0] cfgMerged_1_cfg_wm_tmp_7_a = wdata_reg[60:59]; // @[PMP.scala 93:61]
  wire  cfgMerged_1_cfg_wm_tmp_7_atomic = wdata_reg[61]; // @[PMP.scala 93:61]
  wire  cfgMerged_1_cfg_wm_tmp_7_c = wdata_reg[62]; // @[PMP.scala 93:61]
  wire  cfgMerged_1_cfg_wm_tmp_7_l = wdata_reg[63]; // @[PMP.scala 93:61]
  wire  _cfgMerged_1_cfgVec_7_a_T_1 = |cfgMerged_1_cfg_wm_tmp_7_a; // @[PMP.scala 97:80]
  wire [1:0] _cfgMerged_1_cfgVec_7_a_T_2 = {cfgMerged_1_cfg_wm_tmp_7_a[1],_cfgMerged_1_cfgVec_7_a_T_1}; // @[Cat.scala 31:58]
  wire [1:0] cfgMerged_1_cfgVec__7_a = ~cfgMerged_1_cfg_wm_tmp_7_l ? _cfgMerged_1_cfgVec_7_a_T_2 :
    cfgMerged_1_cfg_wm_tmp_7_a; // @[PMP.scala 94:17 95:29 97:41]
  wire [34:0] _cfgMerged_1_mask_15_match_mask_c_addr_T_1 = {addr_1_15,cfgMerged_1_cfgVec__7_a[0]}; // @[Cat.scala 31:58]
  wire [34:0] cfgMerged_1_mask_15_match_mask_c_addr = _cfgMerged_1_mask_15_match_mask_c_addr_T_1 | 35'h3ff; // @[PMP.scala 86:50]
  wire [34:0] _cfgMerged_1_mask_15_T_1 = cfgMerged_1_mask_15_match_mask_c_addr + 35'h1; // @[PMP.scala 87:49]
  wire [34:0] _cfgMerged_1_mask_15_T_2 = ~_cfgMerged_1_mask_15_T_1; // @[PMP.scala 87:29]
  wire [34:0] _cfgMerged_1_mask_15_T_3 = cfgMerged_1_mask_15_match_mask_c_addr & _cfgMerged_1_mask_15_T_2; // @[PMP.scala 87:27]
  wire [36:0] _cfgMerged_1_mask_15_T_4 = {_cfgMerged_1_mask_15_T_3,2'h3}; // @[Cat.scala 31:58]
  wire [36:0] _GEN_35 = cfgMerged_1_cfgVec__7_a[1] ? _cfgMerged_1_mask_15_T_4 : {{1'd0}, mask_1_15}; // @[PMP.scala 313:23 98:36 99:27]
  wire  cfgMerged_1_cfgVec__7_w = ~cfgMerged_1_cfg_wm_tmp_7_l ? cfgMerged_1_cfg_wm_tmp_7_w &
    cfgMerged_1_cfg_wm_tmp_7_r : cfgMerged_1_cfg_wm_tmp_7_w; // @[PMP.scala 94:17 95:29 96:21]
  wire [36:0] _GEN_38 = ~cfgMerged_1_cfg_wm_tmp_7_l ? _GEN_35 : {{1'd0}, mask_1_15}; // @[PMP.scala 313:23 95:29]
  wire [7:0] cfgMerged_1_lo_lo_lo = {cfgMerged_1_cfg_wm_tmp_l,cfgMerged_1_cfg_wm_tmp_c,cfgMerged_1_cfg_wm_tmp_atomic,
    cfgMerged_1_cfgVec__0_a,cfgMerged_1_cfg_wm_tmp_x,cfgMerged_1_cfgVec__0_w,cfgMerged_1_cfg_wm_tmp_r}; // @[PMP.scala 103:12]
  wire [15:0] cfgMerged_1_lo_lo = {cfgMerged_1_cfg_wm_tmp_1_l,cfgMerged_1_cfg_wm_tmp_1_c,
    cfgMerged_1_cfg_wm_tmp_1_atomic,cfgMerged_1_cfgVec__1_a,cfgMerged_1_cfg_wm_tmp_1_x,cfgMerged_1_cfgVec__1_w,
    cfgMerged_1_cfg_wm_tmp_1_r,cfgMerged_1_lo_lo_lo}; // @[PMP.scala 103:12]
  wire [7:0] cfgMerged_1_lo_hi_lo = {cfgMerged_1_cfg_wm_tmp_2_l,cfgMerged_1_cfg_wm_tmp_2_c,
    cfgMerged_1_cfg_wm_tmp_2_atomic,cfgMerged_1_cfgVec__2_a,cfgMerged_1_cfg_wm_tmp_2_x,cfgMerged_1_cfgVec__2_w,
    cfgMerged_1_cfg_wm_tmp_2_r}; // @[PMP.scala 103:12]
  wire [31:0] cfgMerged_1_lo = {cfgMerged_1_cfg_wm_tmp_3_l,cfgMerged_1_cfg_wm_tmp_3_c,cfgMerged_1_cfg_wm_tmp_3_atomic
    ,cfgMerged_1_cfgVec__3_a,cfgMerged_1_cfg_wm_tmp_3_x,cfgMerged_1_cfgVec__3_w,cfgMerged_1_cfg_wm_tmp_3_r,
    cfgMerged_1_lo_hi_lo,cfgMerged_1_lo_lo}; // @[PMP.scala 103:12]
  wire [7:0] cfgMerged_1_hi_lo_lo = {cfgMerged_1_cfg_wm_tmp_4_l,cfgMerged_1_cfg_wm_tmp_4_c,
    cfgMerged_1_cfg_wm_tmp_4_atomic,cfgMerged_1_cfgVec__4_a,cfgMerged_1_cfg_wm_tmp_4_x,cfgMerged_1_cfgVec__4_w,
    cfgMerged_1_cfg_wm_tmp_4_r}; // @[PMP.scala 103:12]
  wire [15:0] cfgMerged_1_hi_lo = {cfgMerged_1_cfg_wm_tmp_5_l,cfgMerged_1_cfg_wm_tmp_5_c,
    cfgMerged_1_cfg_wm_tmp_5_atomic,cfgMerged_1_cfgVec__5_a,cfgMerged_1_cfg_wm_tmp_5_x,cfgMerged_1_cfgVec__5_w,
    cfgMerged_1_cfg_wm_tmp_5_r,cfgMerged_1_hi_lo_lo}; // @[PMP.scala 103:12]
  wire [7:0] cfgMerged_1_hi_hi_lo = {cfgMerged_1_cfg_wm_tmp_6_l,cfgMerged_1_cfg_wm_tmp_6_c,
    cfgMerged_1_cfg_wm_tmp_6_atomic,cfgMerged_1_cfgVec__6_a,cfgMerged_1_cfg_wm_tmp_6_x,cfgMerged_1_cfgVec__6_w,
    cfgMerged_1_cfg_wm_tmp_6_r}; // @[PMP.scala 103:12]
  wire [63:0] _cfgMerged_1_T_20 = {cfgMerged_1_cfg_wm_tmp_7_l,cfgMerged_1_cfg_wm_tmp_7_c,
    cfgMerged_1_cfg_wm_tmp_7_atomic,cfgMerged_1_cfgVec__7_a,cfgMerged_1_cfg_wm_tmp_7_x,cfgMerged_1_cfgVec__7_w,
    cfgMerged_1_cfg_wm_tmp_7_r,cfgMerged_1_hi_hi_lo,cfgMerged_1_hi_lo,cfgMerged_1_lo}; // @[PMP.scala 103:12]
  wire [36:0] _GEN_39 = wen_reg_3 ? _GEN_10 : {{1'd0}, mask_1_8}; // @[PMP.scala 313:23 RegMap.scala 56:24]
  wire [36:0] _GEN_40 = wen_reg_3 ? _GEN_14 : {{1'd0}, mask_1_9}; // @[PMP.scala 313:23 RegMap.scala 56:24]
  wire [36:0] _GEN_41 = wen_reg_3 ? _GEN_18 : {{1'd0}, mask_1_10}; // @[PMP.scala 313:23 RegMap.scala 56:24]
  wire [36:0] _GEN_42 = wen_reg_3 ? _GEN_22 : {{1'd0}, mask_1_11}; // @[PMP.scala 313:23 RegMap.scala 56:24]
  wire [36:0] _GEN_43 = wen_reg_3 ? _GEN_26 : {{1'd0}, mask_1_12}; // @[PMP.scala 313:23 RegMap.scala 56:24]
  wire [36:0] _GEN_44 = wen_reg_3 ? _GEN_30 : {{1'd0}, mask_1_13}; // @[PMP.scala 313:23 RegMap.scala 56:24]
  wire [36:0] _GEN_45 = wen_reg_3 ? _GEN_34 : {{1'd0}, mask_1_14}; // @[PMP.scala 313:23 RegMap.scala 56:24]
  wire [36:0] _GEN_46 = wen_reg_3 ? _GEN_38 : {{1'd0}, mask_1_15}; // @[PMP.scala 313:23 RegMap.scala 56:24]
  reg  wen_reg_4; // @[RegMap.scala 55:30]
  wire  _addr_0_mask_0_T = cfgs_1_1_a == 2'h1; // @[PMP.scala 53:15]
  wire  _addr_0_mask_0_T_2 = cfgs_1_0_l | cfgs_1_1_l & _addr_0_mask_0_T; // @[PMP.scala 61:51]
  wire  _addr_0_mask_0_T_3 = ~_addr_0_mask_0_T_2; // @[PMP.scala 271:17]
  wire [64:0] _addr_0_mask_0_match_mask_c_addr_T_1 = {wdata_reg,cfgs_1_0_a[0]}; // @[Cat.scala 31:58]
  wire [64:0] addr_0_mask_0_match_mask_c_addr = _addr_0_mask_0_match_mask_c_addr_T_1 | 65'h3ff; // @[PMP.scala 86:50]
  wire [64:0] _addr_0_mask_0_T_5 = addr_0_mask_0_match_mask_c_addr + 65'h1; // @[PMP.scala 87:49]
  wire [64:0] _addr_0_mask_0_T_6 = ~_addr_0_mask_0_T_5; // @[PMP.scala 87:29]
  wire [64:0] _addr_0_mask_0_T_7 = addr_0_mask_0_match_mask_c_addr & _addr_0_mask_0_T_6; // @[PMP.scala 87:27]
  wire [66:0] _addr_0_mask_0_T_8 = {_addr_0_mask_0_T_7,2'h3}; // @[Cat.scala 31:58]
  wire [66:0] _addr_0_mask_0_T_9 = ~_addr_0_mask_0_T_2 ? _addr_0_mask_0_T_8 : {{31'd0}, mask_2_0}; // @[PMP.scala 271:16]
  wire [63:0] _addr_0_T_8 = _addr_0_mask_0_T_3 ? wdata_reg : {{30'd0}, addr_2_0}; // @[PMP.scala 272:8]
  wire [66:0] _GEN_48 = wen_reg_4 ? _addr_0_mask_0_T_9 : {{31'd0}, mask_2_0}; // @[PMP.scala 271:10 313:23 RegMap.scala 56:24]
  wire [63:0] _GEN_49 = wen_reg_4 ? _addr_0_T_8 : {{30'd0}, addr_2_0}; // @[PMP.scala 312:23 RegMap.scala 56:{24,28}]
  reg  wen_reg_5; // @[RegMap.scala 55:30]
  wire  _addr_5_mask_5_T = cfgs__6_a == 2'h1; // @[PMP.scala 53:15]
  wire  _addr_5_mask_5_T_2 = cfgs__5_l | cfgs__6_l & _addr_5_mask_5_T; // @[PMP.scala 61:51]
  wire  _addr_5_mask_5_T_3 = ~_addr_5_mask_5_T_2; // @[PMP.scala 271:17]
  wire [64:0] _addr_5_mask_5_match_mask_c_addr_T_1 = {wdata_reg,cfgs__5_a[0]}; // @[Cat.scala 31:58]
  wire [64:0] addr_5_mask_5_match_mask_c_addr = _addr_5_mask_5_match_mask_c_addr_T_1 | 65'h3ff; // @[PMP.scala 86:50]
  wire [64:0] _addr_5_mask_5_T_5 = addr_5_mask_5_match_mask_c_addr + 65'h1; // @[PMP.scala 87:49]
  wire [64:0] _addr_5_mask_5_T_6 = ~_addr_5_mask_5_T_5; // @[PMP.scala 87:29]
  wire [64:0] _addr_5_mask_5_T_7 = addr_5_mask_5_match_mask_c_addr & _addr_5_mask_5_T_6; // @[PMP.scala 87:27]
  wire [66:0] _addr_5_mask_5_T_8 = {_addr_5_mask_5_T_7,2'h3}; // @[Cat.scala 31:58]
  wire [66:0] _addr_5_mask_5_T_9 = ~_addr_5_mask_5_T_2 ? _addr_5_mask_5_T_8 : {{31'd0}, mask_1_5}; // @[PMP.scala 271:16]
  wire [63:0] _addr_5_T_8 = _addr_5_mask_5_T_3 ? wdata_reg : {{30'd0}, addr_1_5}; // @[PMP.scala 272:8]
  wire [66:0] _GEN_50 = wen_reg_5 ? _addr_5_mask_5_T_9 : {{31'd0}, mask_1_5}; // @[PMP.scala 271:10 313:23 RegMap.scala 56:24]
  wire [63:0] _GEN_51 = wen_reg_5 ? _addr_5_T_8 : {{30'd0}, addr_1_5}; // @[PMP.scala 312:23 RegMap.scala 56:{24,28}]
  reg  wen_reg_6; // @[RegMap.scala 55:30]
  wire  _addr_15_mask_15_T = ~cfgs_1_15_l; // @[PMP.scala 276:17]
  wire [64:0] _addr_15_mask_15_match_mask_c_addr_T_1 = {wdata_reg,cfgs_1_15_a[0]}; // @[Cat.scala 31:58]
  wire [64:0] addr_15_mask_15_match_mask_c_addr = _addr_15_mask_15_match_mask_c_addr_T_1 | 65'h3ff; // @[PMP.scala 86:50]
  wire [64:0] _addr_15_mask_15_T_2 = addr_15_mask_15_match_mask_c_addr + 65'h1; // @[PMP.scala 87:49]
  wire [64:0] _addr_15_mask_15_T_3 = ~_addr_15_mask_15_T_2; // @[PMP.scala 87:29]
  wire [64:0] _addr_15_mask_15_T_4 = addr_15_mask_15_match_mask_c_addr & _addr_15_mask_15_T_3; // @[PMP.scala 87:27]
  wire [66:0] _addr_15_mask_15_T_5 = {_addr_15_mask_15_T_4,2'h3}; // @[Cat.scala 31:58]
  wire [66:0] _addr_15_mask_15_T_6 = ~cfgs_1_15_l ? _addr_15_mask_15_T_5 : {{31'd0}, mask_2_15}; // @[PMP.scala 276:16]
  wire [63:0] _addr_15_T_5 = _addr_15_mask_15_T ? wdata_reg : {{30'd0}, addr_2_15}; // @[PMP.scala 277:8]
  wire [66:0] _GEN_52 = wen_reg_6 ? _addr_15_mask_15_T_6 : {{31'd0}, mask_2_15}; // @[PMP.scala 276:10 313:23 RegMap.scala 56:24]
  wire [63:0] _GEN_53 = wen_reg_6 ? _addr_15_T_5 : {{30'd0}, addr_2_15}; // @[PMP.scala 312:23 RegMap.scala 56:{24,28}]
  reg  wen_reg_7; // @[RegMap.scala 55:30]
  wire  _addr_12_mask_12_T = cfgs__13_a == 2'h1; // @[PMP.scala 53:15]
  wire  _addr_12_mask_12_T_2 = cfgs__12_l | cfgs__13_l & _addr_12_mask_12_T; // @[PMP.scala 61:51]
  wire  _addr_12_mask_12_T_3 = ~_addr_12_mask_12_T_2; // @[PMP.scala 271:17]
  wire [64:0] _addr_12_mask_12_match_mask_c_addr_T_1 = {wdata_reg,cfgs__12_a[0]}; // @[Cat.scala 31:58]
  wire [64:0] addr_12_mask_12_match_mask_c_addr = _addr_12_mask_12_match_mask_c_addr_T_1 | 65'h3ff; // @[PMP.scala 86:50]
  wire [64:0] _addr_12_mask_12_T_5 = addr_12_mask_12_match_mask_c_addr + 65'h1; // @[PMP.scala 87:49]
  wire [64:0] _addr_12_mask_12_T_6 = ~_addr_12_mask_12_T_5; // @[PMP.scala 87:29]
  wire [64:0] _addr_12_mask_12_T_7 = addr_12_mask_12_match_mask_c_addr & _addr_12_mask_12_T_6; // @[PMP.scala 87:27]
  wire [66:0] _addr_12_mask_12_T_8 = {_addr_12_mask_12_T_7,2'h3}; // @[Cat.scala 31:58]
  wire [66:0] _addr_12_mask_12_T_9 = ~_addr_12_mask_12_T_2 ? _addr_12_mask_12_T_8 : {{31'd0}, mask_1_12}; // @[PMP.scala 271:16]
  wire [63:0] _addr_12_T_8 = _addr_12_mask_12_T_3 ? wdata_reg : {{30'd0}, addr_1_12}; // @[PMP.scala 272:8]
  wire [66:0] _GEN_54 = wen_reg_7 ? _addr_12_mask_12_T_9 : {{30'd0}, _GEN_43}; // @[PMP.scala 271:10 RegMap.scala 56:24]
  wire [63:0] _GEN_55 = wen_reg_7 ? _addr_12_T_8 : {{30'd0}, addr_1_12}; // @[PMP.scala 312:23 RegMap.scala 56:{24,28}]
  reg  wen_reg_8; // @[RegMap.scala 55:30]
  wire  _addr_10_mask_10_T = cfgs_1_11_a == 2'h1; // @[PMP.scala 53:15]
  wire  _addr_10_mask_10_T_2 = cfgs_1_10_l | cfgs_1_11_l & _addr_10_mask_10_T; // @[PMP.scala 61:51]
  wire  _addr_10_mask_10_T_3 = ~_addr_10_mask_10_T_2; // @[PMP.scala 271:17]
  wire [64:0] _addr_10_mask_10_match_mask_c_addr_T_1 = {wdata_reg,cfgs_1_10_a[0]}; // @[Cat.scala 31:58]
  wire [64:0] addr_10_mask_10_match_mask_c_addr = _addr_10_mask_10_match_mask_c_addr_T_1 | 65'h3ff; // @[PMP.scala 86:50]
  wire [64:0] _addr_10_mask_10_T_5 = addr_10_mask_10_match_mask_c_addr + 65'h1; // @[PMP.scala 87:49]
  wire [64:0] _addr_10_mask_10_T_6 = ~_addr_10_mask_10_T_5; // @[PMP.scala 87:29]
  wire [64:0] _addr_10_mask_10_T_7 = addr_10_mask_10_match_mask_c_addr & _addr_10_mask_10_T_6; // @[PMP.scala 87:27]
  wire [66:0] _addr_10_mask_10_T_8 = {_addr_10_mask_10_T_7,2'h3}; // @[Cat.scala 31:58]
  wire [66:0] _addr_10_mask_10_T_9 = ~_addr_10_mask_10_T_2 ? _addr_10_mask_10_T_8 : {{31'd0}, mask_2_10}; // @[PMP.scala 271:16]
  wire [63:0] _addr_10_T_8 = _addr_10_mask_10_T_3 ? wdata_reg : {{30'd0}, addr_2_10}; // @[PMP.scala 272:8]
  wire [66:0] _GEN_56 = wen_reg_8 ? _addr_10_mask_10_T_9 : {{31'd0}, mask_2_10}; // @[PMP.scala 271:10 313:23 RegMap.scala 56:24]
  wire [63:0] _GEN_57 = wen_reg_8 ? _addr_10_T_8 : {{30'd0}, addr_2_10}; // @[PMP.scala 312:23 RegMap.scala 56:{24,28}]
  reg  wen_reg_9; // @[RegMap.scala 55:30]
  wire  _addr_8_mask_8_T = cfgs_1_9_a == 2'h1; // @[PMP.scala 53:15]
  wire  _addr_8_mask_8_T_2 = cfgs_1_8_l | cfgs_1_9_l & _addr_8_mask_8_T; // @[PMP.scala 61:51]
  wire  _addr_8_mask_8_T_3 = ~_addr_8_mask_8_T_2; // @[PMP.scala 271:17]
  wire [64:0] _addr_8_mask_8_match_mask_c_addr_T_1 = {wdata_reg,cfgs_1_8_a[0]}; // @[Cat.scala 31:58]
  wire [64:0] addr_8_mask_8_match_mask_c_addr = _addr_8_mask_8_match_mask_c_addr_T_1 | 65'h3ff; // @[PMP.scala 86:50]
  wire [64:0] _addr_8_mask_8_T_5 = addr_8_mask_8_match_mask_c_addr + 65'h1; // @[PMP.scala 87:49]
  wire [64:0] _addr_8_mask_8_T_6 = ~_addr_8_mask_8_T_5; // @[PMP.scala 87:29]
  wire [64:0] _addr_8_mask_8_T_7 = addr_8_mask_8_match_mask_c_addr & _addr_8_mask_8_T_6; // @[PMP.scala 87:27]
  wire [66:0] _addr_8_mask_8_T_8 = {_addr_8_mask_8_T_7,2'h3}; // @[Cat.scala 31:58]
  wire [66:0] _addr_8_mask_8_T_9 = ~_addr_8_mask_8_T_2 ? _addr_8_mask_8_T_8 : {{31'd0}, mask_2_8}; // @[PMP.scala 271:16]
  wire [63:0] _addr_8_T_8 = _addr_8_mask_8_T_3 ? wdata_reg : {{30'd0}, addr_2_8}; // @[PMP.scala 272:8]
  wire [66:0] _GEN_58 = wen_reg_9 ? _addr_8_mask_8_T_9 : {{31'd0}, mask_2_8}; // @[PMP.scala 271:10 313:23 RegMap.scala 56:24]
  wire [63:0] _GEN_59 = wen_reg_9 ? _addr_8_T_8 : {{30'd0}, addr_2_8}; // @[PMP.scala 312:23 RegMap.scala 56:{24,28}]
  reg  wen_reg_10; // @[RegMap.scala 55:30]
  wire  _addr_13_mask_13_T = cfgs__14_a == 2'h1; // @[PMP.scala 53:15]
  wire  _addr_13_mask_13_T_2 = cfgs__13_l | cfgs__14_l & _addr_13_mask_13_T; // @[PMP.scala 61:51]
  wire  _addr_13_mask_13_T_3 = ~_addr_13_mask_13_T_2; // @[PMP.scala 271:17]
  wire [64:0] _addr_13_mask_13_match_mask_c_addr_T_1 = {wdata_reg,cfgs__13_a[0]}; // @[Cat.scala 31:58]
  wire [64:0] addr_13_mask_13_match_mask_c_addr = _addr_13_mask_13_match_mask_c_addr_T_1 | 65'h3ff; // @[PMP.scala 86:50]
  wire [64:0] _addr_13_mask_13_T_5 = addr_13_mask_13_match_mask_c_addr + 65'h1; // @[PMP.scala 87:49]
  wire [64:0] _addr_13_mask_13_T_6 = ~_addr_13_mask_13_T_5; // @[PMP.scala 87:29]
  wire [64:0] _addr_13_mask_13_T_7 = addr_13_mask_13_match_mask_c_addr & _addr_13_mask_13_T_6; // @[PMP.scala 87:27]
  wire [66:0] _addr_13_mask_13_T_8 = {_addr_13_mask_13_T_7,2'h3}; // @[Cat.scala 31:58]
  wire [66:0] _addr_13_mask_13_T_9 = ~_addr_13_mask_13_T_2 ? _addr_13_mask_13_T_8 : {{31'd0}, mask_1_13}; // @[PMP.scala 271:16]
  wire [63:0] _addr_13_T_8 = _addr_13_mask_13_T_3 ? wdata_reg : {{30'd0}, addr_1_13}; // @[PMP.scala 272:8]
  wire [66:0] _GEN_60 = wen_reg_10 ? _addr_13_mask_13_T_9 : {{30'd0}, _GEN_44}; // @[PMP.scala 271:10 RegMap.scala 56:24]
  wire [63:0] _GEN_61 = wen_reg_10 ? _addr_13_T_8 : {{30'd0}, addr_1_13}; // @[PMP.scala 312:23 RegMap.scala 56:{24,28}]
  reg  wen_reg_11; // @[RegMap.scala 55:30]
  wire  _addr_8_mask_8_T_10 = cfgs__9_a == 2'h1; // @[PMP.scala 53:15]
  wire  _addr_8_mask_8_T_12 = cfgs__8_l | cfgs__9_l & _addr_8_mask_8_T_10; // @[PMP.scala 61:51]
  wire  _addr_8_mask_8_T_13 = ~_addr_8_mask_8_T_12; // @[PMP.scala 271:17]
  wire [64:0] _addr_8_mask_8_match_mask_c_addr_T_3 = {wdata_reg,cfgs__8_a[0]}; // @[Cat.scala 31:58]
  wire [64:0] addr_8_mask_8_match_mask_c_addr_1 = _addr_8_mask_8_match_mask_c_addr_T_3 | 65'h3ff; // @[PMP.scala 86:50]
  wire [64:0] _addr_8_mask_8_T_15 = addr_8_mask_8_match_mask_c_addr_1 + 65'h1; // @[PMP.scala 87:49]
  wire [64:0] _addr_8_mask_8_T_16 = ~_addr_8_mask_8_T_15; // @[PMP.scala 87:29]
  wire [64:0] _addr_8_mask_8_T_17 = addr_8_mask_8_match_mask_c_addr_1 & _addr_8_mask_8_T_16; // @[PMP.scala 87:27]
  wire [66:0] _addr_8_mask_8_T_18 = {_addr_8_mask_8_T_17,2'h3}; // @[Cat.scala 31:58]
  wire [66:0] _addr_8_mask_8_T_19 = ~_addr_8_mask_8_T_12 ? _addr_8_mask_8_T_18 : {{31'd0}, mask_1_8}; // @[PMP.scala 271:16]
  wire [63:0] _addr_8_T_17 = _addr_8_mask_8_T_13 ? wdata_reg : {{30'd0}, addr_1_8}; // @[PMP.scala 272:8]
  wire [66:0] _GEN_62 = wen_reg_11 ? _addr_8_mask_8_T_19 : {{30'd0}, _GEN_39}; // @[PMP.scala 271:10 RegMap.scala 56:24]
  wire [63:0] _GEN_63 = wen_reg_11 ? _addr_8_T_17 : {{30'd0}, addr_1_8}; // @[PMP.scala 312:23 RegMap.scala 56:{24,28}]
  reg  wen_reg_12; // @[RegMap.scala 55:30]
  wire  _addr_4_mask_4_T = cfgs__5_a == 2'h1; // @[PMP.scala 53:15]
  wire  _addr_4_mask_4_T_2 = cfgs__4_l | cfgs__5_l & _addr_4_mask_4_T; // @[PMP.scala 61:51]
  wire  _addr_4_mask_4_T_3 = ~_addr_4_mask_4_T_2; // @[PMP.scala 271:17]
  wire [64:0] _addr_4_mask_4_match_mask_c_addr_T_1 = {wdata_reg,cfgs__4_a[0]}; // @[Cat.scala 31:58]
  wire [64:0] addr_4_mask_4_match_mask_c_addr = _addr_4_mask_4_match_mask_c_addr_T_1 | 65'h3ff; // @[PMP.scala 86:50]
  wire [64:0] _addr_4_mask_4_T_5 = addr_4_mask_4_match_mask_c_addr + 65'h1; // @[PMP.scala 87:49]
  wire [64:0] _addr_4_mask_4_T_6 = ~_addr_4_mask_4_T_5; // @[PMP.scala 87:29]
  wire [64:0] _addr_4_mask_4_T_7 = addr_4_mask_4_match_mask_c_addr & _addr_4_mask_4_T_6; // @[PMP.scala 87:27]
  wire [66:0] _addr_4_mask_4_T_8 = {_addr_4_mask_4_T_7,2'h3}; // @[Cat.scala 31:58]
  wire [66:0] _addr_4_mask_4_T_9 = ~_addr_4_mask_4_T_2 ? _addr_4_mask_4_T_8 : {{31'd0}, mask_1_4}; // @[PMP.scala 271:16]
  wire [63:0] _addr_4_T_8 = _addr_4_mask_4_T_3 ? wdata_reg : {{30'd0}, addr_1_4}; // @[PMP.scala 272:8]
  wire [66:0] _GEN_64 = wen_reg_12 ? _addr_4_mask_4_T_9 : {{31'd0}, mask_1_4}; // @[PMP.scala 271:10 313:23 RegMap.scala 56:24]
  wire [63:0] _GEN_65 = wen_reg_12 ? _addr_4_T_8 : {{30'd0}, addr_1_4}; // @[PMP.scala 312:23 RegMap.scala 56:{24,28}]
  reg  wen_reg_13; // @[RegMap.scala 55:30]
  wire  _addr_14_mask_14_T = cfgs_1_15_a == 2'h1; // @[PMP.scala 53:15]
  wire  _addr_14_mask_14_T_2 = cfgs_1_14_l | cfgs_1_15_l & _addr_14_mask_14_T; // @[PMP.scala 61:51]
  wire  _addr_14_mask_14_T_3 = ~_addr_14_mask_14_T_2; // @[PMP.scala 271:17]
  wire [64:0] _addr_14_mask_14_match_mask_c_addr_T_1 = {wdata_reg,cfgs_1_14_a[0]}; // @[Cat.scala 31:58]
  wire [64:0] addr_14_mask_14_match_mask_c_addr = _addr_14_mask_14_match_mask_c_addr_T_1 | 65'h3ff; // @[PMP.scala 86:50]
  wire [64:0] _addr_14_mask_14_T_5 = addr_14_mask_14_match_mask_c_addr + 65'h1; // @[PMP.scala 87:49]
  wire [64:0] _addr_14_mask_14_T_6 = ~_addr_14_mask_14_T_5; // @[PMP.scala 87:29]
  wire [64:0] _addr_14_mask_14_T_7 = addr_14_mask_14_match_mask_c_addr & _addr_14_mask_14_T_6; // @[PMP.scala 87:27]
  wire [66:0] _addr_14_mask_14_T_8 = {_addr_14_mask_14_T_7,2'h3}; // @[Cat.scala 31:58]
  wire [66:0] _addr_14_mask_14_T_9 = ~_addr_14_mask_14_T_2 ? _addr_14_mask_14_T_8 : {{31'd0}, mask_2_14}; // @[PMP.scala 271:16]
  wire [63:0] _addr_14_T_8 = _addr_14_mask_14_T_3 ? wdata_reg : {{30'd0}, addr_2_14}; // @[PMP.scala 272:8]
  wire [66:0] _GEN_66 = wen_reg_13 ? _addr_14_mask_14_T_9 : {{31'd0}, mask_2_14}; // @[PMP.scala 271:10 313:23 RegMap.scala 56:24]
  wire [63:0] _GEN_67 = wen_reg_13 ? _addr_14_T_8 : {{30'd0}, addr_2_14}; // @[PMP.scala 312:23 RegMap.scala 56:{24,28}]
  reg  wen_reg_14; // @[RegMap.scala 55:30]
  wire [34:0] _cfgMerged_0_mask_0_match_mask_c_addr_T_1 = {addr_2_0,cfgMerged_1_cfgVec__0_a[0]}; // @[Cat.scala 31:58]
  wire [34:0] cfgMerged_0_mask_0_match_mask_c_addr = _cfgMerged_0_mask_0_match_mask_c_addr_T_1 | 35'h3ff; // @[PMP.scala 86:50]
  wire [34:0] _cfgMerged_0_mask_0_T_1 = cfgMerged_0_mask_0_match_mask_c_addr + 35'h1; // @[PMP.scala 87:49]
  wire [34:0] _cfgMerged_0_mask_0_T_2 = ~_cfgMerged_0_mask_0_T_1; // @[PMP.scala 87:29]
  wire [34:0] _cfgMerged_0_mask_0_T_3 = cfgMerged_0_mask_0_match_mask_c_addr & _cfgMerged_0_mask_0_T_2; // @[PMP.scala 87:27]
  wire [36:0] _cfgMerged_0_mask_0_T_4 = {_cfgMerged_0_mask_0_T_3,2'h3}; // @[Cat.scala 31:58]
  wire [66:0] _GEN_68 = cfgMerged_1_cfgVec__0_a[1] ? {{30'd0}, _cfgMerged_0_mask_0_T_4} : _GEN_48; // @[PMP.scala 98:36 99:27]
  wire [66:0] _GEN_71 = ~cfgMerged_1_cfg_wm_tmp_l ? _GEN_68 : _GEN_48; // @[PMP.scala 95:29]
  wire [34:0] _cfgMerged_0_mask_1_match_mask_c_addr_T_1 = {addr_2_1,cfgMerged_1_cfgVec__1_a[0]}; // @[Cat.scala 31:58]
  wire [34:0] cfgMerged_0_mask_1_match_mask_c_addr = _cfgMerged_0_mask_1_match_mask_c_addr_T_1 | 35'h3ff; // @[PMP.scala 86:50]
  wire [34:0] _cfgMerged_0_mask_1_T_1 = cfgMerged_0_mask_1_match_mask_c_addr + 35'h1; // @[PMP.scala 87:49]
  wire [34:0] _cfgMerged_0_mask_1_T_2 = ~_cfgMerged_0_mask_1_T_1; // @[PMP.scala 87:29]
  wire [34:0] _cfgMerged_0_mask_1_T_3 = cfgMerged_0_mask_1_match_mask_c_addr & _cfgMerged_0_mask_1_T_2; // @[PMP.scala 87:27]
  wire [36:0] _cfgMerged_0_mask_1_T_4 = {_cfgMerged_0_mask_1_T_3,2'h3}; // @[Cat.scala 31:58]
  wire [36:0] _GEN_72 = cfgMerged_1_cfgVec__1_a[1] ? _cfgMerged_0_mask_1_T_4 : {{1'd0}, mask_2_1}; // @[PMP.scala 313:23 98:36 99:27]
  wire [36:0] _GEN_75 = ~cfgMerged_1_cfg_wm_tmp_1_l ? _GEN_72 : {{1'd0}, mask_2_1}; // @[PMP.scala 313:23 95:29]
  wire [34:0] _cfgMerged_0_mask_2_match_mask_c_addr_T_1 = {addr_2_2,cfgMerged_1_cfgVec__2_a[0]}; // @[Cat.scala 31:58]
  wire [34:0] cfgMerged_0_mask_2_match_mask_c_addr = _cfgMerged_0_mask_2_match_mask_c_addr_T_1 | 35'h3ff; // @[PMP.scala 86:50]
  wire [34:0] _cfgMerged_0_mask_2_T_1 = cfgMerged_0_mask_2_match_mask_c_addr + 35'h1; // @[PMP.scala 87:49]
  wire [34:0] _cfgMerged_0_mask_2_T_2 = ~_cfgMerged_0_mask_2_T_1; // @[PMP.scala 87:29]
  wire [34:0] _cfgMerged_0_mask_2_T_3 = cfgMerged_0_mask_2_match_mask_c_addr & _cfgMerged_0_mask_2_T_2; // @[PMP.scala 87:27]
  wire [36:0] _cfgMerged_0_mask_2_T_4 = {_cfgMerged_0_mask_2_T_3,2'h3}; // @[Cat.scala 31:58]
  wire [36:0] _GEN_76 = cfgMerged_1_cfgVec__2_a[1] ? _cfgMerged_0_mask_2_T_4 : {{1'd0}, mask_2_2}; // @[PMP.scala 313:23 98:36 99:27]
  wire [36:0] _GEN_79 = ~cfgMerged_1_cfg_wm_tmp_2_l ? _GEN_76 : {{1'd0}, mask_2_2}; // @[PMP.scala 313:23 95:29]
  wire [34:0] _cfgMerged_0_mask_3_match_mask_c_addr_T_1 = {addr_2_3,cfgMerged_1_cfgVec__3_a[0]}; // @[Cat.scala 31:58]
  wire [34:0] cfgMerged_0_mask_3_match_mask_c_addr = _cfgMerged_0_mask_3_match_mask_c_addr_T_1 | 35'h3ff; // @[PMP.scala 86:50]
  wire [34:0] _cfgMerged_0_mask_3_T_1 = cfgMerged_0_mask_3_match_mask_c_addr + 35'h1; // @[PMP.scala 87:49]
  wire [34:0] _cfgMerged_0_mask_3_T_2 = ~_cfgMerged_0_mask_3_T_1; // @[PMP.scala 87:29]
  wire [34:0] _cfgMerged_0_mask_3_T_3 = cfgMerged_0_mask_3_match_mask_c_addr & _cfgMerged_0_mask_3_T_2; // @[PMP.scala 87:27]
  wire [36:0] _cfgMerged_0_mask_3_T_4 = {_cfgMerged_0_mask_3_T_3,2'h3}; // @[Cat.scala 31:58]
  wire [66:0] _GEN_80 = cfgMerged_1_cfgVec__3_a[1] ? {{30'd0}, _cfgMerged_0_mask_3_T_4} : _GEN_1; // @[PMP.scala 98:36 99:27]
  wire [66:0] _GEN_83 = ~cfgMerged_1_cfg_wm_tmp_3_l ? _GEN_80 : _GEN_1; // @[PMP.scala 95:29]
  wire [34:0] _cfgMerged_0_mask_4_match_mask_c_addr_T_1 = {addr_2_4,cfgMerged_1_cfgVec__4_a[0]}; // @[Cat.scala 31:58]
  wire [34:0] cfgMerged_0_mask_4_match_mask_c_addr = _cfgMerged_0_mask_4_match_mask_c_addr_T_1 | 35'h3ff; // @[PMP.scala 86:50]
  wire [34:0] _cfgMerged_0_mask_4_T_1 = cfgMerged_0_mask_4_match_mask_c_addr + 35'h1; // @[PMP.scala 87:49]
  wire [34:0] _cfgMerged_0_mask_4_T_2 = ~_cfgMerged_0_mask_4_T_1; // @[PMP.scala 87:29]
  wire [34:0] _cfgMerged_0_mask_4_T_3 = cfgMerged_0_mask_4_match_mask_c_addr & _cfgMerged_0_mask_4_T_2; // @[PMP.scala 87:27]
  wire [36:0] _cfgMerged_0_mask_4_T_4 = {_cfgMerged_0_mask_4_T_3,2'h3}; // @[Cat.scala 31:58]
  wire [36:0] _GEN_84 = cfgMerged_1_cfgVec__4_a[1] ? _cfgMerged_0_mask_4_T_4 : {{1'd0}, mask_2_4}; // @[PMP.scala 313:23 98:36 99:27]
  wire [36:0] _GEN_87 = ~cfgMerged_1_cfg_wm_tmp_4_l ? _GEN_84 : {{1'd0}, mask_2_4}; // @[PMP.scala 313:23 95:29]
  wire [34:0] _cfgMerged_0_mask_5_match_mask_c_addr_T_1 = {addr_2_5,cfgMerged_1_cfgVec__5_a[0]}; // @[Cat.scala 31:58]
  wire [34:0] cfgMerged_0_mask_5_match_mask_c_addr = _cfgMerged_0_mask_5_match_mask_c_addr_T_1 | 35'h3ff; // @[PMP.scala 86:50]
  wire [34:0] _cfgMerged_0_mask_5_T_1 = cfgMerged_0_mask_5_match_mask_c_addr + 35'h1; // @[PMP.scala 87:49]
  wire [34:0] _cfgMerged_0_mask_5_T_2 = ~_cfgMerged_0_mask_5_T_1; // @[PMP.scala 87:29]
  wire [34:0] _cfgMerged_0_mask_5_T_3 = cfgMerged_0_mask_5_match_mask_c_addr & _cfgMerged_0_mask_5_T_2; // @[PMP.scala 87:27]
  wire [36:0] _cfgMerged_0_mask_5_T_4 = {_cfgMerged_0_mask_5_T_3,2'h3}; // @[Cat.scala 31:58]
  wire [36:0] _GEN_88 = cfgMerged_1_cfgVec__5_a[1] ? _cfgMerged_0_mask_5_T_4 : {{1'd0}, mask_2_5}; // @[PMP.scala 313:23 98:36 99:27]
  wire [36:0] _GEN_91 = ~cfgMerged_1_cfg_wm_tmp_5_l ? _GEN_88 : {{1'd0}, mask_2_5}; // @[PMP.scala 313:23 95:29]
  wire [34:0] _cfgMerged_0_mask_6_match_mask_c_addr_T_1 = {addr_2_6,cfgMerged_1_cfgVec__6_a[0]}; // @[Cat.scala 31:58]
  wire [34:0] cfgMerged_0_mask_6_match_mask_c_addr = _cfgMerged_0_mask_6_match_mask_c_addr_T_1 | 35'h3ff; // @[PMP.scala 86:50]
  wire [34:0] _cfgMerged_0_mask_6_T_1 = cfgMerged_0_mask_6_match_mask_c_addr + 35'h1; // @[PMP.scala 87:49]
  wire [34:0] _cfgMerged_0_mask_6_T_2 = ~_cfgMerged_0_mask_6_T_1; // @[PMP.scala 87:29]
  wire [34:0] _cfgMerged_0_mask_6_T_3 = cfgMerged_0_mask_6_match_mask_c_addr & _cfgMerged_0_mask_6_T_2; // @[PMP.scala 87:27]
  wire [36:0] _cfgMerged_0_mask_6_T_4 = {_cfgMerged_0_mask_6_T_3,2'h3}; // @[Cat.scala 31:58]
  wire [36:0] _GEN_92 = cfgMerged_1_cfgVec__6_a[1] ? _cfgMerged_0_mask_6_T_4 : {{1'd0}, mask_2_6}; // @[PMP.scala 313:23 98:36 99:27]
  wire [36:0] _GEN_95 = ~cfgMerged_1_cfg_wm_tmp_6_l ? _GEN_92 : {{1'd0}, mask_2_6}; // @[PMP.scala 313:23 95:29]
  wire [34:0] _cfgMerged_0_mask_7_match_mask_c_addr_T_1 = {addr_2_7,cfgMerged_1_cfgVec__7_a[0]}; // @[Cat.scala 31:58]
  wire [34:0] cfgMerged_0_mask_7_match_mask_c_addr = _cfgMerged_0_mask_7_match_mask_c_addr_T_1 | 35'h3ff; // @[PMP.scala 86:50]
  wire [34:0] _cfgMerged_0_mask_7_T_1 = cfgMerged_0_mask_7_match_mask_c_addr + 35'h1; // @[PMP.scala 87:49]
  wire [34:0] _cfgMerged_0_mask_7_T_2 = ~_cfgMerged_0_mask_7_T_1; // @[PMP.scala 87:29]
  wire [34:0] _cfgMerged_0_mask_7_T_3 = cfgMerged_0_mask_7_match_mask_c_addr & _cfgMerged_0_mask_7_T_2; // @[PMP.scala 87:27]
  wire [36:0] _cfgMerged_0_mask_7_T_4 = {_cfgMerged_0_mask_7_T_3,2'h3}; // @[Cat.scala 31:58]
  wire [66:0] _GEN_96 = cfgMerged_1_cfgVec__7_a[1] ? {{30'd0}, _cfgMerged_0_mask_7_T_4} : _GEN_3; // @[PMP.scala 98:36 99:27]
  wire [66:0] _GEN_99 = ~cfgMerged_1_cfg_wm_tmp_7_l ? _GEN_96 : _GEN_3; // @[PMP.scala 95:29]
  wire [66:0] _GEN_100 = wen_reg_14 ? _GEN_71 : _GEN_48; // @[RegMap.scala 56:24]
  wire [36:0] _GEN_101 = wen_reg_14 ? _GEN_75 : {{1'd0}, mask_2_1}; // @[PMP.scala 313:23 RegMap.scala 56:24]
  wire [36:0] _GEN_102 = wen_reg_14 ? _GEN_79 : {{1'd0}, mask_2_2}; // @[PMP.scala 313:23 RegMap.scala 56:24]
  wire [66:0] _GEN_103 = wen_reg_14 ? _GEN_83 : _GEN_1; // @[RegMap.scala 56:24]
  wire [36:0] _GEN_104 = wen_reg_14 ? _GEN_87 : {{1'd0}, mask_2_4}; // @[PMP.scala 313:23 RegMap.scala 56:24]
  wire [36:0] _GEN_105 = wen_reg_14 ? _GEN_91 : {{1'd0}, mask_2_5}; // @[PMP.scala 313:23 RegMap.scala 56:24]
  wire [36:0] _GEN_106 = wen_reg_14 ? _GEN_95 : {{1'd0}, mask_2_6}; // @[PMP.scala 313:23 RegMap.scala 56:24]
  wire [66:0] _GEN_107 = wen_reg_14 ? _GEN_99 : _GEN_3; // @[RegMap.scala 56:24]
  reg  wen_reg_15; // @[RegMap.scala 55:30]
  wire  _addr_9_mask_9_T = cfgs__10_a == 2'h1; // @[PMP.scala 53:15]
  wire  _addr_9_mask_9_T_2 = cfgs__9_l | cfgs__10_l & _addr_9_mask_9_T; // @[PMP.scala 61:51]
  wire  _addr_9_mask_9_T_3 = ~_addr_9_mask_9_T_2; // @[PMP.scala 271:17]
  wire [64:0] _addr_9_mask_9_match_mask_c_addr_T_1 = {wdata_reg,cfgs__9_a[0]}; // @[Cat.scala 31:58]
  wire [64:0] addr_9_mask_9_match_mask_c_addr = _addr_9_mask_9_match_mask_c_addr_T_1 | 65'h3ff; // @[PMP.scala 86:50]
  wire [64:0] _addr_9_mask_9_T_5 = addr_9_mask_9_match_mask_c_addr + 65'h1; // @[PMP.scala 87:49]
  wire [64:0] _addr_9_mask_9_T_6 = ~_addr_9_mask_9_T_5; // @[PMP.scala 87:29]
  wire [64:0] _addr_9_mask_9_T_7 = addr_9_mask_9_match_mask_c_addr & _addr_9_mask_9_T_6; // @[PMP.scala 87:27]
  wire [66:0] _addr_9_mask_9_T_8 = {_addr_9_mask_9_T_7,2'h3}; // @[Cat.scala 31:58]
  wire [66:0] _addr_9_mask_9_T_9 = ~_addr_9_mask_9_T_2 ? _addr_9_mask_9_T_8 : {{31'd0}, mask_1_9}; // @[PMP.scala 271:16]
  wire [63:0] _addr_9_T_8 = _addr_9_mask_9_T_3 ? wdata_reg : {{30'd0}, addr_1_9}; // @[PMP.scala 272:8]
  wire [66:0] _GEN_109 = wen_reg_15 ? _addr_9_mask_9_T_9 : {{30'd0}, _GEN_40}; // @[PMP.scala 271:10 RegMap.scala 56:24]
  wire [63:0] _GEN_110 = wen_reg_15 ? _addr_9_T_8 : {{30'd0}, addr_1_9}; // @[PMP.scala 312:23 RegMap.scala 56:{24,28}]
  reg  wen_reg_16; // @[RegMap.scala 55:30]
  wire  _addr_4_mask_4_T_10 = cfgs_1_5_a == 2'h1; // @[PMP.scala 53:15]
  wire  _addr_4_mask_4_T_12 = cfgs_1_4_l | cfgs_1_5_l & _addr_4_mask_4_T_10; // @[PMP.scala 61:51]
  wire  _addr_4_mask_4_T_13 = ~_addr_4_mask_4_T_12; // @[PMP.scala 271:17]
  wire [64:0] _addr_4_mask_4_match_mask_c_addr_T_3 = {wdata_reg,cfgs_1_4_a[0]}; // @[Cat.scala 31:58]
  wire [64:0] addr_4_mask_4_match_mask_c_addr_1 = _addr_4_mask_4_match_mask_c_addr_T_3 | 65'h3ff; // @[PMP.scala 86:50]
  wire [64:0] _addr_4_mask_4_T_15 = addr_4_mask_4_match_mask_c_addr_1 + 65'h1; // @[PMP.scala 87:49]
  wire [64:0] _addr_4_mask_4_T_16 = ~_addr_4_mask_4_T_15; // @[PMP.scala 87:29]
  wire [64:0] _addr_4_mask_4_T_17 = addr_4_mask_4_match_mask_c_addr_1 & _addr_4_mask_4_T_16; // @[PMP.scala 87:27]
  wire [66:0] _addr_4_mask_4_T_18 = {_addr_4_mask_4_T_17,2'h3}; // @[Cat.scala 31:58]
  wire [66:0] _addr_4_mask_4_T_19 = ~_addr_4_mask_4_T_12 ? _addr_4_mask_4_T_18 : {{31'd0}, mask_2_4}; // @[PMP.scala 271:16]
  wire [63:0] _addr_4_T_17 = _addr_4_mask_4_T_13 ? wdata_reg : {{30'd0}, addr_2_4}; // @[PMP.scala 272:8]
  wire [66:0] _GEN_111 = wen_reg_16 ? _addr_4_mask_4_T_19 : {{30'd0}, _GEN_104}; // @[PMP.scala 271:10 RegMap.scala 56:24]
  wire [63:0] _GEN_112 = wen_reg_16 ? _addr_4_T_17 : {{30'd0}, addr_2_4}; // @[PMP.scala 312:23 RegMap.scala 56:{24,28}]
  reg  wen_reg_17; // @[RegMap.scala 55:30]
  wire  _addr_9_mask_9_T_10 = cfgs_1_10_a == 2'h1; // @[PMP.scala 53:15]
  wire  _addr_9_mask_9_T_12 = cfgs_1_9_l | cfgs_1_10_l & _addr_9_mask_9_T_10; // @[PMP.scala 61:51]
  wire  _addr_9_mask_9_T_13 = ~_addr_9_mask_9_T_12; // @[PMP.scala 271:17]
  wire [64:0] _addr_9_mask_9_match_mask_c_addr_T_3 = {wdata_reg,cfgs_1_9_a[0]}; // @[Cat.scala 31:58]
  wire [64:0] addr_9_mask_9_match_mask_c_addr_1 = _addr_9_mask_9_match_mask_c_addr_T_3 | 65'h3ff; // @[PMP.scala 86:50]
  wire [64:0] _addr_9_mask_9_T_15 = addr_9_mask_9_match_mask_c_addr_1 + 65'h1; // @[PMP.scala 87:49]
  wire [64:0] _addr_9_mask_9_T_16 = ~_addr_9_mask_9_T_15; // @[PMP.scala 87:29]
  wire [64:0] _addr_9_mask_9_T_17 = addr_9_mask_9_match_mask_c_addr_1 & _addr_9_mask_9_T_16; // @[PMP.scala 87:27]
  wire [66:0] _addr_9_mask_9_T_18 = {_addr_9_mask_9_T_17,2'h3}; // @[Cat.scala 31:58]
  wire [66:0] _addr_9_mask_9_T_19 = ~_addr_9_mask_9_T_12 ? _addr_9_mask_9_T_18 : {{31'd0}, mask_2_9}; // @[PMP.scala 271:16]
  wire [63:0] _addr_9_T_17 = _addr_9_mask_9_T_13 ? wdata_reg : {{30'd0}, addr_2_9}; // @[PMP.scala 272:8]
  wire [66:0] _GEN_113 = wen_reg_17 ? _addr_9_mask_9_T_19 : {{31'd0}, mask_2_9}; // @[PMP.scala 271:10 313:23 RegMap.scala 56:24]
  wire [63:0] _GEN_114 = wen_reg_17 ? _addr_9_T_17 : {{30'd0}, addr_2_9}; // @[PMP.scala 312:23 RegMap.scala 56:{24,28}]
  reg  wen_reg_18; // @[RegMap.scala 55:30]
  wire  _addr_14_mask_14_T_10 = cfgs__15_a == 2'h1; // @[PMP.scala 53:15]
  wire  _addr_14_mask_14_T_12 = cfgs__14_l | cfgs__15_l & _addr_14_mask_14_T_10; // @[PMP.scala 61:51]
  wire  _addr_14_mask_14_T_13 = ~_addr_14_mask_14_T_12; // @[PMP.scala 271:17]
  wire [64:0] _addr_14_mask_14_match_mask_c_addr_T_3 = {wdata_reg,cfgs__14_a[0]}; // @[Cat.scala 31:58]
  wire [64:0] addr_14_mask_14_match_mask_c_addr_1 = _addr_14_mask_14_match_mask_c_addr_T_3 | 65'h3ff; // @[PMP.scala 86:50]
  wire [64:0] _addr_14_mask_14_T_15 = addr_14_mask_14_match_mask_c_addr_1 + 65'h1; // @[PMP.scala 87:49]
  wire [64:0] _addr_14_mask_14_T_16 = ~_addr_14_mask_14_T_15; // @[PMP.scala 87:29]
  wire [64:0] _addr_14_mask_14_T_17 = addr_14_mask_14_match_mask_c_addr_1 & _addr_14_mask_14_T_16; // @[PMP.scala 87:27]
  wire [66:0] _addr_14_mask_14_T_18 = {_addr_14_mask_14_T_17,2'h3}; // @[Cat.scala 31:58]
  wire [66:0] _addr_14_mask_14_T_19 = ~_addr_14_mask_14_T_12 ? _addr_14_mask_14_T_18 : {{31'd0}, mask_1_14}; // @[PMP.scala 271:16]
  wire [63:0] _addr_14_T_17 = _addr_14_mask_14_T_13 ? wdata_reg : {{30'd0}, addr_1_14}; // @[PMP.scala 272:8]
  wire [66:0] _GEN_115 = wen_reg_18 ? _addr_14_mask_14_T_19 : {{30'd0}, _GEN_45}; // @[PMP.scala 271:10 RegMap.scala 56:24]
  wire [63:0] _GEN_116 = wen_reg_18 ? _addr_14_T_17 : {{30'd0}, addr_1_14}; // @[PMP.scala 312:23 RegMap.scala 56:{24,28}]
  reg  wen_reg_19; // @[RegMap.scala 55:30]
  wire  _addr_5_mask_5_T_10 = cfgs_1_6_a == 2'h1; // @[PMP.scala 53:15]
  wire  _addr_5_mask_5_T_12 = cfgs_1_5_l | cfgs_1_6_l & _addr_5_mask_5_T_10; // @[PMP.scala 61:51]
  wire  _addr_5_mask_5_T_13 = ~_addr_5_mask_5_T_12; // @[PMP.scala 271:17]
  wire [64:0] _addr_5_mask_5_match_mask_c_addr_T_3 = {wdata_reg,cfgs_1_5_a[0]}; // @[Cat.scala 31:58]
  wire [64:0] addr_5_mask_5_match_mask_c_addr_1 = _addr_5_mask_5_match_mask_c_addr_T_3 | 65'h3ff; // @[PMP.scala 86:50]
  wire [64:0] _addr_5_mask_5_T_15 = addr_5_mask_5_match_mask_c_addr_1 + 65'h1; // @[PMP.scala 87:49]
  wire [64:0] _addr_5_mask_5_T_16 = ~_addr_5_mask_5_T_15; // @[PMP.scala 87:29]
  wire [64:0] _addr_5_mask_5_T_17 = addr_5_mask_5_match_mask_c_addr_1 & _addr_5_mask_5_T_16; // @[PMP.scala 87:27]
  wire [66:0] _addr_5_mask_5_T_18 = {_addr_5_mask_5_T_17,2'h3}; // @[Cat.scala 31:58]
  wire [66:0] _addr_5_mask_5_T_19 = ~_addr_5_mask_5_T_12 ? _addr_5_mask_5_T_18 : {{31'd0}, mask_2_5}; // @[PMP.scala 271:16]
  wire [63:0] _addr_5_T_17 = _addr_5_mask_5_T_13 ? wdata_reg : {{30'd0}, addr_2_5}; // @[PMP.scala 272:8]
  wire [66:0] _GEN_117 = wen_reg_19 ? _addr_5_mask_5_T_19 : {{30'd0}, _GEN_105}; // @[PMP.scala 271:10 RegMap.scala 56:24]
  wire [63:0] _GEN_118 = wen_reg_19 ? _addr_5_T_17 : {{30'd0}, addr_2_5}; // @[PMP.scala 312:23 RegMap.scala 56:{24,28}]
  reg  wen_reg_20; // @[RegMap.scala 55:30]
  wire  _addr_3_mask_3_T_10 = cfgs__4_a == 2'h1; // @[PMP.scala 53:15]
  wire  _addr_3_mask_3_T_12 = cfgs__3_l | cfgs__4_l & _addr_3_mask_3_T_10; // @[PMP.scala 61:51]
  wire  _addr_3_mask_3_T_13 = ~_addr_3_mask_3_T_12; // @[PMP.scala 271:17]
  wire [64:0] _addr_3_mask_3_match_mask_c_addr_T_3 = {wdata_reg,cfgs__3_a[0]}; // @[Cat.scala 31:58]
  wire [64:0] addr_3_mask_3_match_mask_c_addr_1 = _addr_3_mask_3_match_mask_c_addr_T_3 | 65'h3ff; // @[PMP.scala 86:50]
  wire [64:0] _addr_3_mask_3_T_15 = addr_3_mask_3_match_mask_c_addr_1 + 65'h1; // @[PMP.scala 87:49]
  wire [64:0] _addr_3_mask_3_T_16 = ~_addr_3_mask_3_T_15; // @[PMP.scala 87:29]
  wire [64:0] _addr_3_mask_3_T_17 = addr_3_mask_3_match_mask_c_addr_1 & _addr_3_mask_3_T_16; // @[PMP.scala 87:27]
  wire [66:0] _addr_3_mask_3_T_18 = {_addr_3_mask_3_T_17,2'h3}; // @[Cat.scala 31:58]
  wire [66:0] _addr_3_mask_3_T_19 = ~_addr_3_mask_3_T_12 ? _addr_3_mask_3_T_18 : {{31'd0}, mask_1_3}; // @[PMP.scala 271:16]
  wire [63:0] _addr_3_T_17 = _addr_3_mask_3_T_13 ? wdata_reg : {{30'd0}, addr_1_3}; // @[PMP.scala 272:8]
  wire [66:0] _GEN_119 = wen_reg_20 ? _addr_3_mask_3_T_19 : {{31'd0}, mask_1_3}; // @[PMP.scala 271:10 313:23 RegMap.scala 56:24]
  wire [63:0] _GEN_120 = wen_reg_20 ? _addr_3_T_17 : {{30'd0}, addr_1_3}; // @[PMP.scala 312:23 RegMap.scala 56:{24,28}]
  reg  wen_reg_21; // @[RegMap.scala 55:30]
  wire  _addr_1_mask_1_T_10 = cfgs_1_2_a == 2'h1; // @[PMP.scala 53:15]
  wire  _addr_1_mask_1_T_12 = cfgs_1_1_l | cfgs_1_2_l & _addr_1_mask_1_T_10; // @[PMP.scala 61:51]
  wire  _addr_1_mask_1_T_13 = ~_addr_1_mask_1_T_12; // @[PMP.scala 271:17]
  wire [64:0] _addr_1_mask_1_match_mask_c_addr_T_3 = {wdata_reg,cfgs_1_1_a[0]}; // @[Cat.scala 31:58]
  wire [64:0] addr_1_mask_1_match_mask_c_addr_1 = _addr_1_mask_1_match_mask_c_addr_T_3 | 65'h3ff; // @[PMP.scala 86:50]
  wire [64:0] _addr_1_mask_1_T_15 = addr_1_mask_1_match_mask_c_addr_1 + 65'h1; // @[PMP.scala 87:49]
  wire [64:0] _addr_1_mask_1_T_16 = ~_addr_1_mask_1_T_15; // @[PMP.scala 87:29]
  wire [64:0] _addr_1_mask_1_T_17 = addr_1_mask_1_match_mask_c_addr_1 & _addr_1_mask_1_T_16; // @[PMP.scala 87:27]
  wire [66:0] _addr_1_mask_1_T_18 = {_addr_1_mask_1_T_17,2'h3}; // @[Cat.scala 31:58]
  wire [66:0] _addr_1_mask_1_T_19 = ~_addr_1_mask_1_T_12 ? _addr_1_mask_1_T_18 : {{31'd0}, mask_2_1}; // @[PMP.scala 271:16]
  wire [63:0] _addr_1_T_17 = _addr_1_mask_1_T_13 ? wdata_reg : {{30'd0}, addr_2_1}; // @[PMP.scala 272:8]
  wire [66:0] _GEN_121 = wen_reg_21 ? _addr_1_mask_1_T_19 : {{30'd0}, _GEN_101}; // @[PMP.scala 271:10 RegMap.scala 56:24]
  wire [63:0] _GEN_122 = wen_reg_21 ? _addr_1_T_17 : {{30'd0}, addr_2_1}; // @[PMP.scala 312:23 RegMap.scala 56:{24,28}]
  reg  wen_reg_22; // @[RegMap.scala 55:30]
  wire  _addr_15_mask_15_T_7 = ~cfgs__15_l; // @[PMP.scala 276:17]
  wire [64:0] _addr_15_mask_15_match_mask_c_addr_T_3 = {wdata_reg,cfgs__15_a[0]}; // @[Cat.scala 31:58]
  wire [64:0] addr_15_mask_15_match_mask_c_addr_1 = _addr_15_mask_15_match_mask_c_addr_T_3 | 65'h3ff; // @[PMP.scala 86:50]
  wire [64:0] _addr_15_mask_15_T_9 = addr_15_mask_15_match_mask_c_addr_1 + 65'h1; // @[PMP.scala 87:49]
  wire [64:0] _addr_15_mask_15_T_10 = ~_addr_15_mask_15_T_9; // @[PMP.scala 87:29]
  wire [64:0] _addr_15_mask_15_T_11 = addr_15_mask_15_match_mask_c_addr_1 & _addr_15_mask_15_T_10; // @[PMP.scala 87:27]
  wire [66:0] _addr_15_mask_15_T_12 = {_addr_15_mask_15_T_11,2'h3}; // @[Cat.scala 31:58]
  wire [66:0] _addr_15_mask_15_T_13 = ~cfgs__15_l ? _addr_15_mask_15_T_12 : {{31'd0}, mask_1_15}; // @[PMP.scala 276:16]
  wire [63:0] _addr_15_T_11 = _addr_15_mask_15_T_7 ? wdata_reg : {{30'd0}, addr_1_15}; // @[PMP.scala 277:8]
  wire [66:0] _GEN_123 = wen_reg_22 ? _addr_15_mask_15_T_13 : {{30'd0}, _GEN_46}; // @[PMP.scala 276:10 RegMap.scala 56:24]
  wire [63:0] _GEN_124 = wen_reg_22 ? _addr_15_T_11 : {{30'd0}, addr_1_15}; // @[PMP.scala 312:23 RegMap.scala 56:{24,28}]
  reg  wen_reg_23; // @[RegMap.scala 55:30]
  wire  _addr_13_mask_13_T_10 = cfgs_1_14_a == 2'h1; // @[PMP.scala 53:15]
  wire  _addr_13_mask_13_T_12 = cfgs_1_13_l | cfgs_1_14_l & _addr_13_mask_13_T_10; // @[PMP.scala 61:51]
  wire  _addr_13_mask_13_T_13 = ~_addr_13_mask_13_T_12; // @[PMP.scala 271:17]
  wire [64:0] _addr_13_mask_13_match_mask_c_addr_T_3 = {wdata_reg,cfgs_1_13_a[0]}; // @[Cat.scala 31:58]
  wire [64:0] addr_13_mask_13_match_mask_c_addr_1 = _addr_13_mask_13_match_mask_c_addr_T_3 | 65'h3ff; // @[PMP.scala 86:50]
  wire [64:0] _addr_13_mask_13_T_15 = addr_13_mask_13_match_mask_c_addr_1 + 65'h1; // @[PMP.scala 87:49]
  wire [64:0] _addr_13_mask_13_T_16 = ~_addr_13_mask_13_T_15; // @[PMP.scala 87:29]
  wire [64:0] _addr_13_mask_13_T_17 = addr_13_mask_13_match_mask_c_addr_1 & _addr_13_mask_13_T_16; // @[PMP.scala 87:27]
  wire [66:0] _addr_13_mask_13_T_18 = {_addr_13_mask_13_T_17,2'h3}; // @[Cat.scala 31:58]
  wire [66:0] _addr_13_mask_13_T_19 = ~_addr_13_mask_13_T_12 ? _addr_13_mask_13_T_18 : {{31'd0}, mask_2_13}; // @[PMP.scala 271:16]
  wire [63:0] _addr_13_T_17 = _addr_13_mask_13_T_13 ? wdata_reg : {{30'd0}, addr_2_13}; // @[PMP.scala 272:8]
  wire [66:0] _GEN_125 = wen_reg_23 ? _addr_13_mask_13_T_19 : {{31'd0}, mask_2_13}; // @[PMP.scala 271:10 313:23 RegMap.scala 56:24]
  wire [63:0] _GEN_126 = wen_reg_23 ? _addr_13_T_17 : {{30'd0}, addr_2_13}; // @[PMP.scala 312:23 RegMap.scala 56:{24,28}]
  reg  wen_reg_24; // @[RegMap.scala 55:30]
  wire  _addr_0_mask_0_T_10 = cfgs__1_a == 2'h1; // @[PMP.scala 53:15]
  wire  _addr_0_mask_0_T_12 = cfgs__0_l | cfgs__1_l & _addr_0_mask_0_T_10; // @[PMP.scala 61:51]
  wire  _addr_0_mask_0_T_13 = ~_addr_0_mask_0_T_12; // @[PMP.scala 271:17]
  wire [64:0] _addr_0_mask_0_match_mask_c_addr_T_3 = {wdata_reg,cfgs__0_a[0]}; // @[Cat.scala 31:58]
  wire [64:0] addr_0_mask_0_match_mask_c_addr_1 = _addr_0_mask_0_match_mask_c_addr_T_3 | 65'h3ff; // @[PMP.scala 86:50]
  wire [64:0] _addr_0_mask_0_T_15 = addr_0_mask_0_match_mask_c_addr_1 + 65'h1; // @[PMP.scala 87:49]
  wire [64:0] _addr_0_mask_0_T_16 = ~_addr_0_mask_0_T_15; // @[PMP.scala 87:29]
  wire [64:0] _addr_0_mask_0_T_17 = addr_0_mask_0_match_mask_c_addr_1 & _addr_0_mask_0_T_16; // @[PMP.scala 87:27]
  wire [66:0] _addr_0_mask_0_T_18 = {_addr_0_mask_0_T_17,2'h3}; // @[Cat.scala 31:58]
  wire [66:0] _addr_0_mask_0_T_19 = ~_addr_0_mask_0_T_12 ? _addr_0_mask_0_T_18 : {{31'd0}, mask_1_0}; // @[PMP.scala 271:16]
  wire [63:0] _addr_0_T_17 = _addr_0_mask_0_T_13 ? wdata_reg : {{30'd0}, addr_1_0}; // @[PMP.scala 272:8]
  wire [66:0] _GEN_127 = wen_reg_24 ? _addr_0_mask_0_T_19 : {{31'd0}, mask_1_0}; // @[PMP.scala 271:10 313:23 RegMap.scala 56:24]
  wire [63:0] _GEN_128 = wen_reg_24 ? _addr_0_T_17 : {{30'd0}, addr_1_0}; // @[PMP.scala 312:23 RegMap.scala 56:{24,28}]
  reg  wen_reg_25; // @[RegMap.scala 55:30]
  wire  _addr_10_mask_10_T_10 = cfgs__11_a == 2'h1; // @[PMP.scala 53:15]
  wire  _addr_10_mask_10_T_12 = cfgs__10_l | cfgs__11_l & _addr_10_mask_10_T_10; // @[PMP.scala 61:51]
  wire  _addr_10_mask_10_T_13 = ~_addr_10_mask_10_T_12; // @[PMP.scala 271:17]
  wire [64:0] _addr_10_mask_10_match_mask_c_addr_T_3 = {wdata_reg,cfgs__10_a[0]}; // @[Cat.scala 31:58]
  wire [64:0] addr_10_mask_10_match_mask_c_addr_1 = _addr_10_mask_10_match_mask_c_addr_T_3 | 65'h3ff; // @[PMP.scala 86:50]
  wire [64:0] _addr_10_mask_10_T_15 = addr_10_mask_10_match_mask_c_addr_1 + 65'h1; // @[PMP.scala 87:49]
  wire [64:0] _addr_10_mask_10_T_16 = ~_addr_10_mask_10_T_15; // @[PMP.scala 87:29]
  wire [64:0] _addr_10_mask_10_T_17 = addr_10_mask_10_match_mask_c_addr_1 & _addr_10_mask_10_T_16; // @[PMP.scala 87:27]
  wire [66:0] _addr_10_mask_10_T_18 = {_addr_10_mask_10_T_17,2'h3}; // @[Cat.scala 31:58]
  wire [66:0] _addr_10_mask_10_T_19 = ~_addr_10_mask_10_T_12 ? _addr_10_mask_10_T_18 : {{31'd0}, mask_1_10}; // @[PMP.scala 271:16]
  wire [63:0] _addr_10_T_17 = _addr_10_mask_10_T_13 ? wdata_reg : {{30'd0}, addr_1_10}; // @[PMP.scala 272:8]
  wire [66:0] _GEN_129 = wen_reg_25 ? _addr_10_mask_10_T_19 : {{30'd0}, _GEN_41}; // @[PMP.scala 271:10 RegMap.scala 56:24]
  wire [63:0] _GEN_130 = wen_reg_25 ? _addr_10_T_17 : {{30'd0}, addr_1_10}; // @[PMP.scala 312:23 RegMap.scala 56:{24,28}]
  reg  wen_reg_26; // @[RegMap.scala 55:30]
  wire  _addr_7_mask_7_T_10 = cfgs__8_a == 2'h1; // @[PMP.scala 53:15]
  wire  _addr_7_mask_7_T_12 = cfgs__7_l | cfgs__8_l & _addr_7_mask_7_T_10; // @[PMP.scala 61:51]
  wire  _addr_7_mask_7_T_13 = ~_addr_7_mask_7_T_12; // @[PMP.scala 271:17]
  wire [64:0] _addr_7_mask_7_match_mask_c_addr_T_3 = {wdata_reg,cfgs__7_a[0]}; // @[Cat.scala 31:58]
  wire [64:0] addr_7_mask_7_match_mask_c_addr_1 = _addr_7_mask_7_match_mask_c_addr_T_3 | 65'h3ff; // @[PMP.scala 86:50]
  wire [64:0] _addr_7_mask_7_T_15 = addr_7_mask_7_match_mask_c_addr_1 + 65'h1; // @[PMP.scala 87:49]
  wire [64:0] _addr_7_mask_7_T_16 = ~_addr_7_mask_7_T_15; // @[PMP.scala 87:29]
  wire [64:0] _addr_7_mask_7_T_17 = addr_7_mask_7_match_mask_c_addr_1 & _addr_7_mask_7_T_16; // @[PMP.scala 87:27]
  wire [66:0] _addr_7_mask_7_T_18 = {_addr_7_mask_7_T_17,2'h3}; // @[Cat.scala 31:58]
  wire [66:0] _addr_7_mask_7_T_19 = ~_addr_7_mask_7_T_12 ? _addr_7_mask_7_T_18 : {{31'd0}, mask_1_7}; // @[PMP.scala 271:16]
  wire [63:0] _addr_7_T_17 = _addr_7_mask_7_T_13 ? wdata_reg : {{30'd0}, addr_1_7}; // @[PMP.scala 272:8]
  wire [66:0] _GEN_131 = wen_reg_26 ? _addr_7_mask_7_T_19 : {{31'd0}, mask_1_7}; // @[PMP.scala 271:10 313:23 RegMap.scala 56:24]
  wire [63:0] _GEN_132 = wen_reg_26 ? _addr_7_T_17 : {{30'd0}, addr_1_7}; // @[PMP.scala 312:23 RegMap.scala 56:{24,28}]
  reg  wen_reg_27; // @[RegMap.scala 55:30]
  wire  _addr_6_mask_6_T = cfgs_1_7_a == 2'h1; // @[PMP.scala 53:15]
  wire  _addr_6_mask_6_T_2 = cfgs_1_6_l | cfgs_1_7_l & _addr_6_mask_6_T; // @[PMP.scala 61:51]
  wire  _addr_6_mask_6_T_3 = ~_addr_6_mask_6_T_2; // @[PMP.scala 271:17]
  wire [64:0] _addr_6_mask_6_match_mask_c_addr_T_1 = {wdata_reg,cfgs_1_6_a[0]}; // @[Cat.scala 31:58]
  wire [64:0] addr_6_mask_6_match_mask_c_addr = _addr_6_mask_6_match_mask_c_addr_T_1 | 65'h3ff; // @[PMP.scala 86:50]
  wire [64:0] _addr_6_mask_6_T_5 = addr_6_mask_6_match_mask_c_addr + 65'h1; // @[PMP.scala 87:49]
  wire [64:0] _addr_6_mask_6_T_6 = ~_addr_6_mask_6_T_5; // @[PMP.scala 87:29]
  wire [64:0] _addr_6_mask_6_T_7 = addr_6_mask_6_match_mask_c_addr & _addr_6_mask_6_T_6; // @[PMP.scala 87:27]
  wire [66:0] _addr_6_mask_6_T_8 = {_addr_6_mask_6_T_7,2'h3}; // @[Cat.scala 31:58]
  wire [66:0] _addr_6_mask_6_T_9 = ~_addr_6_mask_6_T_2 ? _addr_6_mask_6_T_8 : {{31'd0}, mask_2_6}; // @[PMP.scala 271:16]
  wire [63:0] _addr_6_T_8 = _addr_6_mask_6_T_3 ? wdata_reg : {{30'd0}, addr_2_6}; // @[PMP.scala 272:8]
  wire [66:0] _GEN_133 = wen_reg_27 ? _addr_6_mask_6_T_9 : {{30'd0}, _GEN_106}; // @[PMP.scala 271:10 RegMap.scala 56:24]
  wire [63:0] _GEN_134 = wen_reg_27 ? _addr_6_T_8 : {{30'd0}, addr_2_6}; // @[PMP.scala 312:23 RegMap.scala 56:{24,28}]
  reg  wen_reg_28; // @[RegMap.scala 55:30]
  wire  _addr_2_mask_2_T = cfgs__3_a == 2'h1; // @[PMP.scala 53:15]
  wire  _addr_2_mask_2_T_2 = cfgs__2_l | cfgs__3_l & _addr_2_mask_2_T; // @[PMP.scala 61:51]
  wire  _addr_2_mask_2_T_3 = ~_addr_2_mask_2_T_2; // @[PMP.scala 271:17]
  wire [64:0] _addr_2_mask_2_match_mask_c_addr_T_1 = {wdata_reg,cfgs__2_a[0]}; // @[Cat.scala 31:58]
  wire [64:0] addr_2_mask_2_match_mask_c_addr = _addr_2_mask_2_match_mask_c_addr_T_1 | 65'h3ff; // @[PMP.scala 86:50]
  wire [64:0] _addr_2_mask_2_T_5 = addr_2_mask_2_match_mask_c_addr + 65'h1; // @[PMP.scala 87:49]
  wire [64:0] _addr_2_mask_2_T_6 = ~_addr_2_mask_2_T_5; // @[PMP.scala 87:29]
  wire [64:0] _addr_2_mask_2_T_7 = addr_2_mask_2_match_mask_c_addr & _addr_2_mask_2_T_6; // @[PMP.scala 87:27]
  wire [66:0] _addr_2_mask_2_T_8 = {_addr_2_mask_2_T_7,2'h3}; // @[Cat.scala 31:58]
  wire [66:0] _addr_2_mask_2_T_9 = ~_addr_2_mask_2_T_2 ? _addr_2_mask_2_T_8 : {{31'd0}, mask_1_2}; // @[PMP.scala 271:16]
  wire [63:0] _addr_2_T_8 = _addr_2_mask_2_T_3 ? wdata_reg : {{30'd0}, addr_1_2}; // @[PMP.scala 272:8]
  wire [66:0] _GEN_135 = wen_reg_28 ? _addr_2_mask_2_T_9 : {{31'd0}, mask_1_2}; // @[PMP.scala 271:10 313:23 RegMap.scala 56:24]
  wire [63:0] _GEN_136 = wen_reg_28 ? _addr_2_T_8 : {{30'd0}, addr_1_2}; // @[PMP.scala 312:23 RegMap.scala 56:{24,28}]
  reg  wen_reg_29; // @[RegMap.scala 55:30]
  wire  _addr_12_mask_12_T_10 = cfgs_1_13_a == 2'h1; // @[PMP.scala 53:15]
  wire  _addr_12_mask_12_T_12 = cfgs_1_12_l | cfgs_1_13_l & _addr_12_mask_12_T_10; // @[PMP.scala 61:51]
  wire  _addr_12_mask_12_T_13 = ~_addr_12_mask_12_T_12; // @[PMP.scala 271:17]
  wire [64:0] _addr_12_mask_12_match_mask_c_addr_T_3 = {wdata_reg,cfgs_1_12_a[0]}; // @[Cat.scala 31:58]
  wire [64:0] addr_12_mask_12_match_mask_c_addr_1 = _addr_12_mask_12_match_mask_c_addr_T_3 | 65'h3ff; // @[PMP.scala 86:50]
  wire [64:0] _addr_12_mask_12_T_15 = addr_12_mask_12_match_mask_c_addr_1 + 65'h1; // @[PMP.scala 87:49]
  wire [64:0] _addr_12_mask_12_T_16 = ~_addr_12_mask_12_T_15; // @[PMP.scala 87:29]
  wire [64:0] _addr_12_mask_12_T_17 = addr_12_mask_12_match_mask_c_addr_1 & _addr_12_mask_12_T_16; // @[PMP.scala 87:27]
  wire [66:0] _addr_12_mask_12_T_18 = {_addr_12_mask_12_T_17,2'h3}; // @[Cat.scala 31:58]
  wire [66:0] _addr_12_mask_12_T_19 = ~_addr_12_mask_12_T_12 ? _addr_12_mask_12_T_18 : {{31'd0}, mask_2_12}; // @[PMP.scala 271:16]
  wire [63:0] _addr_12_T_17 = _addr_12_mask_12_T_13 ? wdata_reg : {{30'd0}, addr_2_12}; // @[PMP.scala 272:8]
  wire [66:0] _GEN_137 = wen_reg_29 ? _addr_12_mask_12_T_19 : {{31'd0}, mask_2_12}; // @[PMP.scala 271:10 313:23 RegMap.scala 56:24]
  wire [63:0] _GEN_138 = wen_reg_29 ? _addr_12_T_17 : {{30'd0}, addr_2_12}; // @[PMP.scala 312:23 RegMap.scala 56:{24,28}]
  reg  wen_reg_30; // @[RegMap.scala 55:30]
  wire  _addr_2_mask_2_T_10 = cfgs_1_3_a == 2'h1; // @[PMP.scala 53:15]
  wire  _addr_2_mask_2_T_12 = cfgs_1_2_l | cfgs_1_3_l & _addr_2_mask_2_T_10; // @[PMP.scala 61:51]
  wire  _addr_2_mask_2_T_13 = ~_addr_2_mask_2_T_12; // @[PMP.scala 271:17]
  wire [64:0] _addr_2_mask_2_match_mask_c_addr_T_3 = {wdata_reg,cfgs_1_2_a[0]}; // @[Cat.scala 31:58]
  wire [64:0] addr_2_mask_2_match_mask_c_addr_1 = _addr_2_mask_2_match_mask_c_addr_T_3 | 65'h3ff; // @[PMP.scala 86:50]
  wire [64:0] _addr_2_mask_2_T_15 = addr_2_mask_2_match_mask_c_addr_1 + 65'h1; // @[PMP.scala 87:49]
  wire [64:0] _addr_2_mask_2_T_16 = ~_addr_2_mask_2_T_15; // @[PMP.scala 87:29]
  wire [64:0] _addr_2_mask_2_T_17 = addr_2_mask_2_match_mask_c_addr_1 & _addr_2_mask_2_T_16; // @[PMP.scala 87:27]
  wire [66:0] _addr_2_mask_2_T_18 = {_addr_2_mask_2_T_17,2'h3}; // @[Cat.scala 31:58]
  wire [66:0] _addr_2_mask_2_T_19 = ~_addr_2_mask_2_T_12 ? _addr_2_mask_2_T_18 : {{31'd0}, mask_2_2}; // @[PMP.scala 271:16]
  wire [63:0] _addr_2_T_17 = _addr_2_mask_2_T_13 ? wdata_reg : {{30'd0}, addr_2_2}; // @[PMP.scala 272:8]
  wire [66:0] _GEN_139 = wen_reg_30 ? _addr_2_mask_2_T_19 : {{30'd0}, _GEN_102}; // @[PMP.scala 271:10 RegMap.scala 56:24]
  wire [63:0] _GEN_140 = wen_reg_30 ? _addr_2_T_17 : {{30'd0}, addr_2_2}; // @[PMP.scala 312:23 RegMap.scala 56:{24,28}]
  reg  wen_reg_31; // @[RegMap.scala 55:30]
  wire  _addr_11_mask_11_T = cfgs_1_12_a == 2'h1; // @[PMP.scala 53:15]
  wire  _addr_11_mask_11_T_2 = cfgs_1_11_l | cfgs_1_12_l & _addr_11_mask_11_T; // @[PMP.scala 61:51]
  wire  _addr_11_mask_11_T_3 = ~_addr_11_mask_11_T_2; // @[PMP.scala 271:17]
  wire [64:0] _addr_11_mask_11_match_mask_c_addr_T_1 = {wdata_reg,cfgs_1_11_a[0]}; // @[Cat.scala 31:58]
  wire [64:0] addr_11_mask_11_match_mask_c_addr = _addr_11_mask_11_match_mask_c_addr_T_1 | 65'h3ff; // @[PMP.scala 86:50]
  wire [64:0] _addr_11_mask_11_T_5 = addr_11_mask_11_match_mask_c_addr + 65'h1; // @[PMP.scala 87:49]
  wire [64:0] _addr_11_mask_11_T_6 = ~_addr_11_mask_11_T_5; // @[PMP.scala 87:29]
  wire [64:0] _addr_11_mask_11_T_7 = addr_11_mask_11_match_mask_c_addr & _addr_11_mask_11_T_6; // @[PMP.scala 87:27]
  wire [66:0] _addr_11_mask_11_T_8 = {_addr_11_mask_11_T_7,2'h3}; // @[Cat.scala 31:58]
  wire [66:0] _addr_11_mask_11_T_9 = ~_addr_11_mask_11_T_2 ? _addr_11_mask_11_T_8 : {{31'd0}, mask_2_11}; // @[PMP.scala 271:16]
  wire [63:0] _addr_11_T_8 = _addr_11_mask_11_T_3 ? wdata_reg : {{30'd0}, addr_2_11}; // @[PMP.scala 272:8]
  wire [66:0] _GEN_141 = wen_reg_31 ? _addr_11_mask_11_T_9 : {{31'd0}, mask_2_11}; // @[PMP.scala 271:10 313:23 RegMap.scala 56:24]
  wire [63:0] _GEN_142 = wen_reg_31 ? _addr_11_T_8 : {{30'd0}, addr_2_11}; // @[PMP.scala 312:23 RegMap.scala 56:{24,28}]
  reg  wen_reg_32; // @[RegMap.scala 55:30]
  wire  _addr_6_mask_6_T_10 = cfgs__7_a == 2'h1; // @[PMP.scala 53:15]
  wire  _addr_6_mask_6_T_12 = cfgs__6_l | cfgs__7_l & _addr_6_mask_6_T_10; // @[PMP.scala 61:51]
  wire  _addr_6_mask_6_T_13 = ~_addr_6_mask_6_T_12; // @[PMP.scala 271:17]
  wire [64:0] _addr_6_mask_6_match_mask_c_addr_T_3 = {wdata_reg,cfgs__6_a[0]}; // @[Cat.scala 31:58]
  wire [64:0] addr_6_mask_6_match_mask_c_addr_1 = _addr_6_mask_6_match_mask_c_addr_T_3 | 65'h3ff; // @[PMP.scala 86:50]
  wire [64:0] _addr_6_mask_6_T_15 = addr_6_mask_6_match_mask_c_addr_1 + 65'h1; // @[PMP.scala 87:49]
  wire [64:0] _addr_6_mask_6_T_16 = ~_addr_6_mask_6_T_15; // @[PMP.scala 87:29]
  wire [64:0] _addr_6_mask_6_T_17 = addr_6_mask_6_match_mask_c_addr_1 & _addr_6_mask_6_T_16; // @[PMP.scala 87:27]
  wire [66:0] _addr_6_mask_6_T_18 = {_addr_6_mask_6_T_17,2'h3}; // @[Cat.scala 31:58]
  wire [66:0] _addr_6_mask_6_T_19 = ~_addr_6_mask_6_T_12 ? _addr_6_mask_6_T_18 : {{31'd0}, mask_1_6}; // @[PMP.scala 271:16]
  wire [63:0] _addr_6_T_17 = _addr_6_mask_6_T_13 ? wdata_reg : {{30'd0}, addr_1_6}; // @[PMP.scala 272:8]
  wire [66:0] _GEN_143 = wen_reg_32 ? _addr_6_mask_6_T_19 : {{31'd0}, mask_1_6}; // @[PMP.scala 271:10 313:23 RegMap.scala 56:24]
  wire [63:0] _GEN_144 = wen_reg_32 ? _addr_6_T_17 : {{30'd0}, addr_1_6}; // @[PMP.scala 312:23 RegMap.scala 56:{24,28}]
  reg  wen_reg_33; // @[RegMap.scala 55:30]
  wire [34:0] _cfgMerged_1_mask_8_match_mask_c_addr_T_3 = {addr_2_8,cfgMerged_1_cfgVec__0_a[0]}; // @[Cat.scala 31:58]
  wire [34:0] cfgMerged_1_mask_8_match_mask_c_addr_1 = _cfgMerged_1_mask_8_match_mask_c_addr_T_3 | 35'h3ff; // @[PMP.scala 86:50]
  wire [34:0] _cfgMerged_1_mask_8_T_6 = cfgMerged_1_mask_8_match_mask_c_addr_1 + 35'h1; // @[PMP.scala 87:49]
  wire [34:0] _cfgMerged_1_mask_8_T_7 = ~_cfgMerged_1_mask_8_T_6; // @[PMP.scala 87:29]
  wire [34:0] _cfgMerged_1_mask_8_T_8 = cfgMerged_1_mask_8_match_mask_c_addr_1 & _cfgMerged_1_mask_8_T_7; // @[PMP.scala 87:27]
  wire [36:0] _cfgMerged_1_mask_8_T_9 = {_cfgMerged_1_mask_8_T_8,2'h3}; // @[Cat.scala 31:58]
  wire [66:0] _GEN_145 = cfgMerged_1_cfgVec__0_a[1] ? {{30'd0}, _cfgMerged_1_mask_8_T_9} : _GEN_58; // @[PMP.scala 98:36 99:27]
  wire [66:0] _GEN_148 = ~cfgMerged_1_cfg_wm_tmp_l ? _GEN_145 : _GEN_58; // @[PMP.scala 95:29]
  wire [34:0] _cfgMerged_1_mask_9_match_mask_c_addr_T_3 = {addr_2_9,cfgMerged_1_cfgVec__1_a[0]}; // @[Cat.scala 31:58]
  wire [34:0] cfgMerged_1_mask_9_match_mask_c_addr_1 = _cfgMerged_1_mask_9_match_mask_c_addr_T_3 | 35'h3ff; // @[PMP.scala 86:50]
  wire [34:0] _cfgMerged_1_mask_9_T_6 = cfgMerged_1_mask_9_match_mask_c_addr_1 + 35'h1; // @[PMP.scala 87:49]
  wire [34:0] _cfgMerged_1_mask_9_T_7 = ~_cfgMerged_1_mask_9_T_6; // @[PMP.scala 87:29]
  wire [34:0] _cfgMerged_1_mask_9_T_8 = cfgMerged_1_mask_9_match_mask_c_addr_1 & _cfgMerged_1_mask_9_T_7; // @[PMP.scala 87:27]
  wire [36:0] _cfgMerged_1_mask_9_T_9 = {_cfgMerged_1_mask_9_T_8,2'h3}; // @[Cat.scala 31:58]
  wire [66:0] _GEN_149 = cfgMerged_1_cfgVec__1_a[1] ? {{30'd0}, _cfgMerged_1_mask_9_T_9} : _GEN_113; // @[PMP.scala 98:36 99:27]
  wire [66:0] _GEN_152 = ~cfgMerged_1_cfg_wm_tmp_1_l ? _GEN_149 : _GEN_113; // @[PMP.scala 95:29]
  wire [34:0] _cfgMerged_1_mask_10_match_mask_c_addr_T_3 = {addr_2_10,cfgMerged_1_cfgVec__2_a[0]}; // @[Cat.scala 31:58]
  wire [34:0] cfgMerged_1_mask_10_match_mask_c_addr_1 = _cfgMerged_1_mask_10_match_mask_c_addr_T_3 | 35'h3ff; // @[PMP.scala 86:50]
  wire [34:0] _cfgMerged_1_mask_10_T_6 = cfgMerged_1_mask_10_match_mask_c_addr_1 + 35'h1; // @[PMP.scala 87:49]
  wire [34:0] _cfgMerged_1_mask_10_T_7 = ~_cfgMerged_1_mask_10_T_6; // @[PMP.scala 87:29]
  wire [34:0] _cfgMerged_1_mask_10_T_8 = cfgMerged_1_mask_10_match_mask_c_addr_1 & _cfgMerged_1_mask_10_T_7; // @[PMP.scala 87:27]
  wire [36:0] _cfgMerged_1_mask_10_T_9 = {_cfgMerged_1_mask_10_T_8,2'h3}; // @[Cat.scala 31:58]
  wire [66:0] _GEN_153 = cfgMerged_1_cfgVec__2_a[1] ? {{30'd0}, _cfgMerged_1_mask_10_T_9} : _GEN_56; // @[PMP.scala 98:36 99:27]
  wire [66:0] _GEN_156 = ~cfgMerged_1_cfg_wm_tmp_2_l ? _GEN_153 : _GEN_56; // @[PMP.scala 95:29]
  wire [34:0] _cfgMerged_1_mask_11_match_mask_c_addr_T_3 = {addr_2_11,cfgMerged_1_cfgVec__3_a[0]}; // @[Cat.scala 31:58]
  wire [34:0] cfgMerged_1_mask_11_match_mask_c_addr_1 = _cfgMerged_1_mask_11_match_mask_c_addr_T_3 | 35'h3ff; // @[PMP.scala 86:50]
  wire [34:0] _cfgMerged_1_mask_11_T_6 = cfgMerged_1_mask_11_match_mask_c_addr_1 + 35'h1; // @[PMP.scala 87:49]
  wire [34:0] _cfgMerged_1_mask_11_T_7 = ~_cfgMerged_1_mask_11_T_6; // @[PMP.scala 87:29]
  wire [34:0] _cfgMerged_1_mask_11_T_8 = cfgMerged_1_mask_11_match_mask_c_addr_1 & _cfgMerged_1_mask_11_T_7; // @[PMP.scala 87:27]
  wire [36:0] _cfgMerged_1_mask_11_T_9 = {_cfgMerged_1_mask_11_T_8,2'h3}; // @[Cat.scala 31:58]
  wire [66:0] _GEN_157 = cfgMerged_1_cfgVec__3_a[1] ? {{30'd0}, _cfgMerged_1_mask_11_T_9} : _GEN_141; // @[PMP.scala 98:36 99:27]
  wire [66:0] _GEN_160 = ~cfgMerged_1_cfg_wm_tmp_3_l ? _GEN_157 : _GEN_141; // @[PMP.scala 95:29]
  wire [34:0] _cfgMerged_1_mask_12_match_mask_c_addr_T_3 = {addr_2_12,cfgMerged_1_cfgVec__4_a[0]}; // @[Cat.scala 31:58]
  wire [34:0] cfgMerged_1_mask_12_match_mask_c_addr_1 = _cfgMerged_1_mask_12_match_mask_c_addr_T_3 | 35'h3ff; // @[PMP.scala 86:50]
  wire [34:0] _cfgMerged_1_mask_12_T_6 = cfgMerged_1_mask_12_match_mask_c_addr_1 + 35'h1; // @[PMP.scala 87:49]
  wire [34:0] _cfgMerged_1_mask_12_T_7 = ~_cfgMerged_1_mask_12_T_6; // @[PMP.scala 87:29]
  wire [34:0] _cfgMerged_1_mask_12_T_8 = cfgMerged_1_mask_12_match_mask_c_addr_1 & _cfgMerged_1_mask_12_T_7; // @[PMP.scala 87:27]
  wire [36:0] _cfgMerged_1_mask_12_T_9 = {_cfgMerged_1_mask_12_T_8,2'h3}; // @[Cat.scala 31:58]
  wire [66:0] _GEN_161 = cfgMerged_1_cfgVec__4_a[1] ? {{30'd0}, _cfgMerged_1_mask_12_T_9} : _GEN_137; // @[PMP.scala 98:36 99:27]
  wire [66:0] _GEN_164 = ~cfgMerged_1_cfg_wm_tmp_4_l ? _GEN_161 : _GEN_137; // @[PMP.scala 95:29]
  wire [34:0] _cfgMerged_1_mask_13_match_mask_c_addr_T_3 = {addr_2_13,cfgMerged_1_cfgVec__5_a[0]}; // @[Cat.scala 31:58]
  wire [34:0] cfgMerged_1_mask_13_match_mask_c_addr_1 = _cfgMerged_1_mask_13_match_mask_c_addr_T_3 | 35'h3ff; // @[PMP.scala 86:50]
  wire [34:0] _cfgMerged_1_mask_13_T_6 = cfgMerged_1_mask_13_match_mask_c_addr_1 + 35'h1; // @[PMP.scala 87:49]
  wire [34:0] _cfgMerged_1_mask_13_T_7 = ~_cfgMerged_1_mask_13_T_6; // @[PMP.scala 87:29]
  wire [34:0] _cfgMerged_1_mask_13_T_8 = cfgMerged_1_mask_13_match_mask_c_addr_1 & _cfgMerged_1_mask_13_T_7; // @[PMP.scala 87:27]
  wire [36:0] _cfgMerged_1_mask_13_T_9 = {_cfgMerged_1_mask_13_T_8,2'h3}; // @[Cat.scala 31:58]
  wire [66:0] _GEN_165 = cfgMerged_1_cfgVec__5_a[1] ? {{30'd0}, _cfgMerged_1_mask_13_T_9} : _GEN_125; // @[PMP.scala 98:36 99:27]
  wire [66:0] _GEN_168 = ~cfgMerged_1_cfg_wm_tmp_5_l ? _GEN_165 : _GEN_125; // @[PMP.scala 95:29]
  wire [34:0] _cfgMerged_1_mask_14_match_mask_c_addr_T_3 = {addr_2_14,cfgMerged_1_cfgVec__6_a[0]}; // @[Cat.scala 31:58]
  wire [34:0] cfgMerged_1_mask_14_match_mask_c_addr_1 = _cfgMerged_1_mask_14_match_mask_c_addr_T_3 | 35'h3ff; // @[PMP.scala 86:50]
  wire [34:0] _cfgMerged_1_mask_14_T_6 = cfgMerged_1_mask_14_match_mask_c_addr_1 + 35'h1; // @[PMP.scala 87:49]
  wire [34:0] _cfgMerged_1_mask_14_T_7 = ~_cfgMerged_1_mask_14_T_6; // @[PMP.scala 87:29]
  wire [34:0] _cfgMerged_1_mask_14_T_8 = cfgMerged_1_mask_14_match_mask_c_addr_1 & _cfgMerged_1_mask_14_T_7; // @[PMP.scala 87:27]
  wire [36:0] _cfgMerged_1_mask_14_T_9 = {_cfgMerged_1_mask_14_T_8,2'h3}; // @[Cat.scala 31:58]
  wire [66:0] _GEN_169 = cfgMerged_1_cfgVec__6_a[1] ? {{30'd0}, _cfgMerged_1_mask_14_T_9} : _GEN_66; // @[PMP.scala 98:36 99:27]
  wire [66:0] _GEN_172 = ~cfgMerged_1_cfg_wm_tmp_6_l ? _GEN_169 : _GEN_66; // @[PMP.scala 95:29]
  wire [34:0] _cfgMerged_1_mask_15_match_mask_c_addr_T_3 = {addr_2_15,cfgMerged_1_cfgVec__7_a[0]}; // @[Cat.scala 31:58]
  wire [34:0] cfgMerged_1_mask_15_match_mask_c_addr_1 = _cfgMerged_1_mask_15_match_mask_c_addr_T_3 | 35'h3ff; // @[PMP.scala 86:50]
  wire [34:0] _cfgMerged_1_mask_15_T_6 = cfgMerged_1_mask_15_match_mask_c_addr_1 + 35'h1; // @[PMP.scala 87:49]
  wire [34:0] _cfgMerged_1_mask_15_T_7 = ~_cfgMerged_1_mask_15_T_6; // @[PMP.scala 87:29]
  wire [34:0] _cfgMerged_1_mask_15_T_8 = cfgMerged_1_mask_15_match_mask_c_addr_1 & _cfgMerged_1_mask_15_T_7; // @[PMP.scala 87:27]
  wire [36:0] _cfgMerged_1_mask_15_T_9 = {_cfgMerged_1_mask_15_T_8,2'h3}; // @[Cat.scala 31:58]
  wire [66:0] _GEN_173 = cfgMerged_1_cfgVec__7_a[1] ? {{30'd0}, _cfgMerged_1_mask_15_T_9} : _GEN_52; // @[PMP.scala 98:36 99:27]
  wire [66:0] _GEN_176 = ~cfgMerged_1_cfg_wm_tmp_7_l ? _GEN_173 : _GEN_52; // @[PMP.scala 95:29]
  wire [66:0] _GEN_177 = wen_reg_33 ? _GEN_148 : _GEN_58; // @[RegMap.scala 56:24]
  wire [66:0] _GEN_178 = wen_reg_33 ? _GEN_152 : _GEN_113; // @[RegMap.scala 56:24]
  wire [66:0] _GEN_179 = wen_reg_33 ? _GEN_156 : _GEN_56; // @[RegMap.scala 56:24]
  wire [66:0] _GEN_180 = wen_reg_33 ? _GEN_160 : _GEN_141; // @[RegMap.scala 56:24]
  wire [66:0] _GEN_181 = wen_reg_33 ? _GEN_164 : _GEN_137; // @[RegMap.scala 56:24]
  wire [66:0] _GEN_182 = wen_reg_33 ? _GEN_168 : _GEN_125; // @[RegMap.scala 56:24]
  wire [66:0] _GEN_183 = wen_reg_33 ? _GEN_172 : _GEN_66; // @[RegMap.scala 56:24]
  wire [66:0] _GEN_184 = wen_reg_33 ? _GEN_176 : _GEN_52; // @[RegMap.scala 56:24]
  reg  wen_reg_34; // @[RegMap.scala 55:30]
  wire  _addr_11_mask_11_T_10 = cfgs__12_a == 2'h1; // @[PMP.scala 53:15]
  wire  _addr_11_mask_11_T_12 = cfgs__11_l | cfgs__12_l & _addr_11_mask_11_T_10; // @[PMP.scala 61:51]
  wire  _addr_11_mask_11_T_13 = ~_addr_11_mask_11_T_12; // @[PMP.scala 271:17]
  wire [64:0] _addr_11_mask_11_match_mask_c_addr_T_3 = {wdata_reg,cfgs__11_a[0]}; // @[Cat.scala 31:58]
  wire [64:0] addr_11_mask_11_match_mask_c_addr_1 = _addr_11_mask_11_match_mask_c_addr_T_3 | 65'h3ff; // @[PMP.scala 86:50]
  wire [64:0] _addr_11_mask_11_T_15 = addr_11_mask_11_match_mask_c_addr_1 + 65'h1; // @[PMP.scala 87:49]
  wire [64:0] _addr_11_mask_11_T_16 = ~_addr_11_mask_11_T_15; // @[PMP.scala 87:29]
  wire [64:0] _addr_11_mask_11_T_17 = addr_11_mask_11_match_mask_c_addr_1 & _addr_11_mask_11_T_16; // @[PMP.scala 87:27]
  wire [66:0] _addr_11_mask_11_T_18 = {_addr_11_mask_11_T_17,2'h3}; // @[Cat.scala 31:58]
  wire [66:0] _addr_11_mask_11_T_19 = ~_addr_11_mask_11_T_12 ? _addr_11_mask_11_T_18 : {{31'd0}, mask_1_11}; // @[PMP.scala 271:16]
  wire [63:0] _addr_11_T_17 = _addr_11_mask_11_T_13 ? wdata_reg : {{30'd0}, addr_1_11}; // @[PMP.scala 272:8]
  wire [66:0] _GEN_186 = wen_reg_34 ? _addr_11_mask_11_T_19 : {{30'd0}, _GEN_42}; // @[PMP.scala 271:10 RegMap.scala 56:24]
  wire [63:0] _GEN_187 = wen_reg_34 ? _addr_11_T_17 : {{30'd0}, addr_1_11}; // @[PMP.scala 312:23 RegMap.scala 56:{24,28}]
  reg  wen_reg_35; // @[RegMap.scala 55:30]
  wire [34:0] _cfgMerged_0_mask_0_match_mask_c_addr_T_3 = {addr_1_0,cfgMerged_1_cfgVec__0_a[0]}; // @[Cat.scala 31:58]
  wire [34:0] cfgMerged_0_mask_0_match_mask_c_addr_1 = _cfgMerged_0_mask_0_match_mask_c_addr_T_3 | 35'h3ff; // @[PMP.scala 86:50]
  wire [34:0] _cfgMerged_0_mask_0_T_6 = cfgMerged_0_mask_0_match_mask_c_addr_1 + 35'h1; // @[PMP.scala 87:49]
  wire [34:0] _cfgMerged_0_mask_0_T_7 = ~_cfgMerged_0_mask_0_T_6; // @[PMP.scala 87:29]
  wire [34:0] _cfgMerged_0_mask_0_T_8 = cfgMerged_0_mask_0_match_mask_c_addr_1 & _cfgMerged_0_mask_0_T_7; // @[PMP.scala 87:27]
  wire [36:0] _cfgMerged_0_mask_0_T_9 = {_cfgMerged_0_mask_0_T_8,2'h3}; // @[Cat.scala 31:58]
  wire [66:0] _GEN_188 = cfgMerged_1_cfgVec__0_a[1] ? {{30'd0}, _cfgMerged_0_mask_0_T_9} : _GEN_127; // @[PMP.scala 98:36 99:27]
  wire [66:0] _GEN_191 = ~cfgMerged_1_cfg_wm_tmp_l ? _GEN_188 : _GEN_127; // @[PMP.scala 95:29]
  wire [34:0] _cfgMerged_0_mask_1_match_mask_c_addr_T_3 = {addr_1_1,cfgMerged_1_cfgVec__1_a[0]}; // @[Cat.scala 31:58]
  wire [34:0] cfgMerged_0_mask_1_match_mask_c_addr_1 = _cfgMerged_0_mask_1_match_mask_c_addr_T_3 | 35'h3ff; // @[PMP.scala 86:50]
  wire [34:0] _cfgMerged_0_mask_1_T_6 = cfgMerged_0_mask_1_match_mask_c_addr_1 + 35'h1; // @[PMP.scala 87:49]
  wire [34:0] _cfgMerged_0_mask_1_T_7 = ~_cfgMerged_0_mask_1_T_6; // @[PMP.scala 87:29]
  wire [34:0] _cfgMerged_0_mask_1_T_8 = cfgMerged_0_mask_1_match_mask_c_addr_1 & _cfgMerged_0_mask_1_T_7; // @[PMP.scala 87:27]
  wire [36:0] _cfgMerged_0_mask_1_T_9 = {_cfgMerged_0_mask_1_T_8,2'h3}; // @[Cat.scala 31:58]
  wire [66:0] _GEN_192 = cfgMerged_1_cfgVec__1_a[1] ? {{30'd0}, _cfgMerged_0_mask_1_T_9} : _GEN_5; // @[PMP.scala 98:36 99:27]
  wire [66:0] _GEN_195 = ~cfgMerged_1_cfg_wm_tmp_1_l ? _GEN_192 : _GEN_5; // @[PMP.scala 95:29]
  wire [34:0] _cfgMerged_0_mask_2_match_mask_c_addr_T_3 = {addr_1_2,cfgMerged_1_cfgVec__2_a[0]}; // @[Cat.scala 31:58]
  wire [34:0] cfgMerged_0_mask_2_match_mask_c_addr_1 = _cfgMerged_0_mask_2_match_mask_c_addr_T_3 | 35'h3ff; // @[PMP.scala 86:50]
  wire [34:0] _cfgMerged_0_mask_2_T_6 = cfgMerged_0_mask_2_match_mask_c_addr_1 + 35'h1; // @[PMP.scala 87:49]
  wire [34:0] _cfgMerged_0_mask_2_T_7 = ~_cfgMerged_0_mask_2_T_6; // @[PMP.scala 87:29]
  wire [34:0] _cfgMerged_0_mask_2_T_8 = cfgMerged_0_mask_2_match_mask_c_addr_1 & _cfgMerged_0_mask_2_T_7; // @[PMP.scala 87:27]
  wire [36:0] _cfgMerged_0_mask_2_T_9 = {_cfgMerged_0_mask_2_T_8,2'h3}; // @[Cat.scala 31:58]
  wire [66:0] _GEN_196 = cfgMerged_1_cfgVec__2_a[1] ? {{30'd0}, _cfgMerged_0_mask_2_T_9} : _GEN_135; // @[PMP.scala 98:36 99:27]
  wire [66:0] _GEN_199 = ~cfgMerged_1_cfg_wm_tmp_2_l ? _GEN_196 : _GEN_135; // @[PMP.scala 95:29]
  wire [34:0] _cfgMerged_0_mask_3_match_mask_c_addr_T_3 = {addr_1_3,cfgMerged_1_cfgVec__3_a[0]}; // @[Cat.scala 31:58]
  wire [34:0] cfgMerged_0_mask_3_match_mask_c_addr_1 = _cfgMerged_0_mask_3_match_mask_c_addr_T_3 | 35'h3ff; // @[PMP.scala 86:50]
  wire [34:0] _cfgMerged_0_mask_3_T_6 = cfgMerged_0_mask_3_match_mask_c_addr_1 + 35'h1; // @[PMP.scala 87:49]
  wire [34:0] _cfgMerged_0_mask_3_T_7 = ~_cfgMerged_0_mask_3_T_6; // @[PMP.scala 87:29]
  wire [34:0] _cfgMerged_0_mask_3_T_8 = cfgMerged_0_mask_3_match_mask_c_addr_1 & _cfgMerged_0_mask_3_T_7; // @[PMP.scala 87:27]
  wire [36:0] _cfgMerged_0_mask_3_T_9 = {_cfgMerged_0_mask_3_T_8,2'h3}; // @[Cat.scala 31:58]
  wire [66:0] _GEN_200 = cfgMerged_1_cfgVec__3_a[1] ? {{30'd0}, _cfgMerged_0_mask_3_T_9} : _GEN_119; // @[PMP.scala 98:36 99:27]
  wire [66:0] _GEN_203 = ~cfgMerged_1_cfg_wm_tmp_3_l ? _GEN_200 : _GEN_119; // @[PMP.scala 95:29]
  wire [34:0] _cfgMerged_0_mask_4_match_mask_c_addr_T_3 = {addr_1_4,cfgMerged_1_cfgVec__4_a[0]}; // @[Cat.scala 31:58]
  wire [34:0] cfgMerged_0_mask_4_match_mask_c_addr_1 = _cfgMerged_0_mask_4_match_mask_c_addr_T_3 | 35'h3ff; // @[PMP.scala 86:50]
  wire [34:0] _cfgMerged_0_mask_4_T_6 = cfgMerged_0_mask_4_match_mask_c_addr_1 + 35'h1; // @[PMP.scala 87:49]
  wire [34:0] _cfgMerged_0_mask_4_T_7 = ~_cfgMerged_0_mask_4_T_6; // @[PMP.scala 87:29]
  wire [34:0] _cfgMerged_0_mask_4_T_8 = cfgMerged_0_mask_4_match_mask_c_addr_1 & _cfgMerged_0_mask_4_T_7; // @[PMP.scala 87:27]
  wire [36:0] _cfgMerged_0_mask_4_T_9 = {_cfgMerged_0_mask_4_T_8,2'h3}; // @[Cat.scala 31:58]
  wire [66:0] _GEN_204 = cfgMerged_1_cfgVec__4_a[1] ? {{30'd0}, _cfgMerged_0_mask_4_T_9} : _GEN_64; // @[PMP.scala 98:36 99:27]
  wire [66:0] _GEN_207 = ~cfgMerged_1_cfg_wm_tmp_4_l ? _GEN_204 : _GEN_64; // @[PMP.scala 95:29]
  wire [34:0] _cfgMerged_0_mask_5_match_mask_c_addr_T_3 = {addr_1_5,cfgMerged_1_cfgVec__5_a[0]}; // @[Cat.scala 31:58]
  wire [34:0] cfgMerged_0_mask_5_match_mask_c_addr_1 = _cfgMerged_0_mask_5_match_mask_c_addr_T_3 | 35'h3ff; // @[PMP.scala 86:50]
  wire [34:0] _cfgMerged_0_mask_5_T_6 = cfgMerged_0_mask_5_match_mask_c_addr_1 + 35'h1; // @[PMP.scala 87:49]
  wire [34:0] _cfgMerged_0_mask_5_T_7 = ~_cfgMerged_0_mask_5_T_6; // @[PMP.scala 87:29]
  wire [34:0] _cfgMerged_0_mask_5_T_8 = cfgMerged_0_mask_5_match_mask_c_addr_1 & _cfgMerged_0_mask_5_T_7; // @[PMP.scala 87:27]
  wire [36:0] _cfgMerged_0_mask_5_T_9 = {_cfgMerged_0_mask_5_T_8,2'h3}; // @[Cat.scala 31:58]
  wire [66:0] _GEN_208 = cfgMerged_1_cfgVec__5_a[1] ? {{30'd0}, _cfgMerged_0_mask_5_T_9} : _GEN_50; // @[PMP.scala 98:36 99:27]
  wire [66:0] _GEN_211 = ~cfgMerged_1_cfg_wm_tmp_5_l ? _GEN_208 : _GEN_50; // @[PMP.scala 95:29]
  wire [34:0] _cfgMerged_0_mask_6_match_mask_c_addr_T_3 = {addr_1_6,cfgMerged_1_cfgVec__6_a[0]}; // @[Cat.scala 31:58]
  wire [34:0] cfgMerged_0_mask_6_match_mask_c_addr_1 = _cfgMerged_0_mask_6_match_mask_c_addr_T_3 | 35'h3ff; // @[PMP.scala 86:50]
  wire [34:0] _cfgMerged_0_mask_6_T_6 = cfgMerged_0_mask_6_match_mask_c_addr_1 + 35'h1; // @[PMP.scala 87:49]
  wire [34:0] _cfgMerged_0_mask_6_T_7 = ~_cfgMerged_0_mask_6_T_6; // @[PMP.scala 87:29]
  wire [34:0] _cfgMerged_0_mask_6_T_8 = cfgMerged_0_mask_6_match_mask_c_addr_1 & _cfgMerged_0_mask_6_T_7; // @[PMP.scala 87:27]
  wire [36:0] _cfgMerged_0_mask_6_T_9 = {_cfgMerged_0_mask_6_T_8,2'h3}; // @[Cat.scala 31:58]
  wire [66:0] _GEN_212 = cfgMerged_1_cfgVec__6_a[1] ? {{30'd0}, _cfgMerged_0_mask_6_T_9} : _GEN_143; // @[PMP.scala 98:36 99:27]
  wire [66:0] _GEN_215 = ~cfgMerged_1_cfg_wm_tmp_6_l ? _GEN_212 : _GEN_143; // @[PMP.scala 95:29]
  wire [34:0] _cfgMerged_0_mask_7_match_mask_c_addr_T_3 = {addr_1_7,cfgMerged_1_cfgVec__7_a[0]}; // @[Cat.scala 31:58]
  wire [34:0] cfgMerged_0_mask_7_match_mask_c_addr_1 = _cfgMerged_0_mask_7_match_mask_c_addr_T_3 | 35'h3ff; // @[PMP.scala 86:50]
  wire [34:0] _cfgMerged_0_mask_7_T_6 = cfgMerged_0_mask_7_match_mask_c_addr_1 + 35'h1; // @[PMP.scala 87:49]
  wire [34:0] _cfgMerged_0_mask_7_T_7 = ~_cfgMerged_0_mask_7_T_6; // @[PMP.scala 87:29]
  wire [34:0] _cfgMerged_0_mask_7_T_8 = cfgMerged_0_mask_7_match_mask_c_addr_1 & _cfgMerged_0_mask_7_T_7; // @[PMP.scala 87:27]
  wire [36:0] _cfgMerged_0_mask_7_T_9 = {_cfgMerged_0_mask_7_T_8,2'h3}; // @[Cat.scala 31:58]
  wire [66:0] _GEN_216 = cfgMerged_1_cfgVec__7_a[1] ? {{30'd0}, _cfgMerged_0_mask_7_T_9} : _GEN_131; // @[PMP.scala 98:36 99:27]
  wire [66:0] _GEN_219 = ~cfgMerged_1_cfg_wm_tmp_7_l ? _GEN_216 : _GEN_131; // @[PMP.scala 95:29]
  wire [66:0] _GEN_220 = wen_reg_35 ? _GEN_191 : _GEN_127; // @[RegMap.scala 56:24]
  wire [66:0] _GEN_221 = wen_reg_35 ? _GEN_195 : _GEN_5; // @[RegMap.scala 56:24]
  wire [66:0] _GEN_222 = wen_reg_35 ? _GEN_199 : _GEN_135; // @[RegMap.scala 56:24]
  wire [66:0] _GEN_223 = wen_reg_35 ? _GEN_203 : _GEN_119; // @[RegMap.scala 56:24]
  wire [66:0] _GEN_224 = wen_reg_35 ? _GEN_207 : _GEN_64; // @[RegMap.scala 56:24]
  wire [66:0] _GEN_225 = wen_reg_35 ? _GEN_211 : _GEN_50; // @[RegMap.scala 56:24]
  wire [66:0] _GEN_226 = wen_reg_35 ? _GEN_215 : _GEN_143; // @[RegMap.scala 56:24]
  wire [66:0] _GEN_227 = wen_reg_35 ? _GEN_219 : _GEN_131; // @[RegMap.scala 56:24]
  assign io_pmp_0_cfg_l = _cfgs_T[7]; // @[PMP.scala 311:44]
  assign io_pmp_0_cfg_a = _cfgs_T[4:3]; // @[PMP.scala 311:44]
  assign io_pmp_0_cfg_x = _cfgs_T[2]; // @[PMP.scala 311:44]
  assign io_pmp_0_cfg_w = _cfgs_T[1]; // @[PMP.scala 311:44]
  assign io_pmp_0_cfg_r = _cfgs_T[0]; // @[PMP.scala 311:44]
  assign io_pmp_0_addr = addr_1_0; // @[PMP.scala 283:15 353:17]
  assign io_pmp_0_mask = mask_1_0; // @[PMP.scala 284:15 353:17]
  assign io_pmp_1_cfg_l = _cfgs_T[15]; // @[PMP.scala 311:44]
  assign io_pmp_1_cfg_a = _cfgs_T[12:11]; // @[PMP.scala 311:44]
  assign io_pmp_1_cfg_x = _cfgs_T[10]; // @[PMP.scala 311:44]
  assign io_pmp_1_cfg_w = _cfgs_T[9]; // @[PMP.scala 311:44]
  assign io_pmp_1_cfg_r = _cfgs_T[8]; // @[PMP.scala 311:44]
  assign io_pmp_1_addr = addr_1_1; // @[PMP.scala 283:15 353:17]
  assign io_pmp_1_mask = mask_1_1; // @[PMP.scala 284:15 353:17]
  assign io_pmp_2_cfg_l = _cfgs_T[23]; // @[PMP.scala 311:44]
  assign io_pmp_2_cfg_a = _cfgs_T[20:19]; // @[PMP.scala 311:44]
  assign io_pmp_2_cfg_x = _cfgs_T[18]; // @[PMP.scala 311:44]
  assign io_pmp_2_cfg_w = _cfgs_T[17]; // @[PMP.scala 311:44]
  assign io_pmp_2_cfg_r = _cfgs_T[16]; // @[PMP.scala 311:44]
  assign io_pmp_2_addr = addr_1_2; // @[PMP.scala 283:15 353:17]
  assign io_pmp_2_mask = mask_1_2; // @[PMP.scala 284:15 353:17]
  assign io_pmp_3_cfg_l = _cfgs_T[31]; // @[PMP.scala 311:44]
  assign io_pmp_3_cfg_a = _cfgs_T[28:27]; // @[PMP.scala 311:44]
  assign io_pmp_3_cfg_x = _cfgs_T[26]; // @[PMP.scala 311:44]
  assign io_pmp_3_cfg_w = _cfgs_T[25]; // @[PMP.scala 311:44]
  assign io_pmp_3_cfg_r = _cfgs_T[24]; // @[PMP.scala 311:44]
  assign io_pmp_3_addr = addr_1_3; // @[PMP.scala 283:15 353:17]
  assign io_pmp_3_mask = mask_1_3; // @[PMP.scala 284:15 353:17]
  assign io_pmp_4_cfg_l = _cfgs_T[39]; // @[PMP.scala 311:44]
  assign io_pmp_4_cfg_a = _cfgs_T[36:35]; // @[PMP.scala 311:44]
  assign io_pmp_4_cfg_x = _cfgs_T[34]; // @[PMP.scala 311:44]
  assign io_pmp_4_cfg_w = _cfgs_T[33]; // @[PMP.scala 311:44]
  assign io_pmp_4_cfg_r = _cfgs_T[32]; // @[PMP.scala 311:44]
  assign io_pmp_4_addr = addr_1_4; // @[PMP.scala 283:15 353:17]
  assign io_pmp_4_mask = mask_1_4; // @[PMP.scala 284:15 353:17]
  assign io_pmp_5_cfg_l = _cfgs_T[47]; // @[PMP.scala 311:44]
  assign io_pmp_5_cfg_a = _cfgs_T[44:43]; // @[PMP.scala 311:44]
  assign io_pmp_5_cfg_x = _cfgs_T[42]; // @[PMP.scala 311:44]
  assign io_pmp_5_cfg_w = _cfgs_T[41]; // @[PMP.scala 311:44]
  assign io_pmp_5_cfg_r = _cfgs_T[40]; // @[PMP.scala 311:44]
  assign io_pmp_5_addr = addr_1_5; // @[PMP.scala 283:15 353:17]
  assign io_pmp_5_mask = mask_1_5; // @[PMP.scala 284:15 353:17]
  assign io_pmp_6_cfg_l = _cfgs_T[55]; // @[PMP.scala 311:44]
  assign io_pmp_6_cfg_a = _cfgs_T[52:51]; // @[PMP.scala 311:44]
  assign io_pmp_6_cfg_x = _cfgs_T[50]; // @[PMP.scala 311:44]
  assign io_pmp_6_cfg_w = _cfgs_T[49]; // @[PMP.scala 311:44]
  assign io_pmp_6_cfg_r = _cfgs_T[48]; // @[PMP.scala 311:44]
  assign io_pmp_6_addr = addr_1_6; // @[PMP.scala 283:15 353:17]
  assign io_pmp_6_mask = mask_1_6; // @[PMP.scala 284:15 353:17]
  assign io_pmp_7_cfg_l = _cfgs_T[63]; // @[PMP.scala 311:44]
  assign io_pmp_7_cfg_a = _cfgs_T[60:59]; // @[PMP.scala 311:44]
  assign io_pmp_7_cfg_x = _cfgs_T[58]; // @[PMP.scala 311:44]
  assign io_pmp_7_cfg_w = _cfgs_T[57]; // @[PMP.scala 311:44]
  assign io_pmp_7_cfg_r = _cfgs_T[56]; // @[PMP.scala 311:44]
  assign io_pmp_7_addr = addr_1_7; // @[PMP.scala 283:15 353:17]
  assign io_pmp_7_mask = mask_1_7; // @[PMP.scala 284:15 353:17]
  assign io_pmp_8_cfg_l = _cfgs_T[71]; // @[PMP.scala 311:44]
  assign io_pmp_8_cfg_a = _cfgs_T[68:67]; // @[PMP.scala 311:44]
  assign io_pmp_8_cfg_x = _cfgs_T[66]; // @[PMP.scala 311:44]
  assign io_pmp_8_cfg_w = _cfgs_T[65]; // @[PMP.scala 311:44]
  assign io_pmp_8_cfg_r = _cfgs_T[64]; // @[PMP.scala 311:44]
  assign io_pmp_8_addr = addr_1_8; // @[PMP.scala 283:15 353:17]
  assign io_pmp_8_mask = mask_1_8; // @[PMP.scala 284:15 353:17]
  assign io_pmp_9_cfg_l = _cfgs_T[79]; // @[PMP.scala 311:44]
  assign io_pmp_9_cfg_a = _cfgs_T[76:75]; // @[PMP.scala 311:44]
  assign io_pmp_9_cfg_x = _cfgs_T[74]; // @[PMP.scala 311:44]
  assign io_pmp_9_cfg_w = _cfgs_T[73]; // @[PMP.scala 311:44]
  assign io_pmp_9_cfg_r = _cfgs_T[72]; // @[PMP.scala 311:44]
  assign io_pmp_9_addr = addr_1_9; // @[PMP.scala 283:15 353:17]
  assign io_pmp_9_mask = mask_1_9; // @[PMP.scala 284:15 353:17]
  assign io_pmp_10_cfg_l = _cfgs_T[87]; // @[PMP.scala 311:44]
  assign io_pmp_10_cfg_a = _cfgs_T[84:83]; // @[PMP.scala 311:44]
  assign io_pmp_10_cfg_x = _cfgs_T[82]; // @[PMP.scala 311:44]
  assign io_pmp_10_cfg_w = _cfgs_T[81]; // @[PMP.scala 311:44]
  assign io_pmp_10_cfg_r = _cfgs_T[80]; // @[PMP.scala 311:44]
  assign io_pmp_10_addr = addr_1_10; // @[PMP.scala 283:15 353:17]
  assign io_pmp_10_mask = mask_1_10; // @[PMP.scala 284:15 353:17]
  assign io_pmp_11_cfg_l = _cfgs_T[95]; // @[PMP.scala 311:44]
  assign io_pmp_11_cfg_a = _cfgs_T[92:91]; // @[PMP.scala 311:44]
  assign io_pmp_11_cfg_x = _cfgs_T[90]; // @[PMP.scala 311:44]
  assign io_pmp_11_cfg_w = _cfgs_T[89]; // @[PMP.scala 311:44]
  assign io_pmp_11_cfg_r = _cfgs_T[88]; // @[PMP.scala 311:44]
  assign io_pmp_11_addr = addr_1_11; // @[PMP.scala 283:15 353:17]
  assign io_pmp_11_mask = mask_1_11; // @[PMP.scala 284:15 353:17]
  assign io_pmp_12_cfg_l = _cfgs_T[103]; // @[PMP.scala 311:44]
  assign io_pmp_12_cfg_a = _cfgs_T[100:99]; // @[PMP.scala 311:44]
  assign io_pmp_12_cfg_x = _cfgs_T[98]; // @[PMP.scala 311:44]
  assign io_pmp_12_cfg_w = _cfgs_T[97]; // @[PMP.scala 311:44]
  assign io_pmp_12_cfg_r = _cfgs_T[96]; // @[PMP.scala 311:44]
  assign io_pmp_12_addr = addr_1_12; // @[PMP.scala 283:15 353:17]
  assign io_pmp_12_mask = mask_1_12; // @[PMP.scala 284:15 353:17]
  assign io_pmp_13_cfg_l = _cfgs_T[111]; // @[PMP.scala 311:44]
  assign io_pmp_13_cfg_a = _cfgs_T[108:107]; // @[PMP.scala 311:44]
  assign io_pmp_13_cfg_x = _cfgs_T[106]; // @[PMP.scala 311:44]
  assign io_pmp_13_cfg_w = _cfgs_T[105]; // @[PMP.scala 311:44]
  assign io_pmp_13_cfg_r = _cfgs_T[104]; // @[PMP.scala 311:44]
  assign io_pmp_13_addr = addr_1_13; // @[PMP.scala 283:15 353:17]
  assign io_pmp_13_mask = mask_1_13; // @[PMP.scala 284:15 353:17]
  assign io_pmp_14_cfg_l = _cfgs_T[119]; // @[PMP.scala 311:44]
  assign io_pmp_14_cfg_a = _cfgs_T[116:115]; // @[PMP.scala 311:44]
  assign io_pmp_14_cfg_x = _cfgs_T[114]; // @[PMP.scala 311:44]
  assign io_pmp_14_cfg_w = _cfgs_T[113]; // @[PMP.scala 311:44]
  assign io_pmp_14_cfg_r = _cfgs_T[112]; // @[PMP.scala 311:44]
  assign io_pmp_14_addr = addr_1_14; // @[PMP.scala 283:15 353:17]
  assign io_pmp_14_mask = mask_1_14; // @[PMP.scala 284:15 353:17]
  assign io_pmp_15_cfg_l = _cfgs_T[127]; // @[PMP.scala 311:44]
  assign io_pmp_15_cfg_a = _cfgs_T[124:123]; // @[PMP.scala 311:44]
  assign io_pmp_15_cfg_x = _cfgs_T[122]; // @[PMP.scala 311:44]
  assign io_pmp_15_cfg_w = _cfgs_T[121]; // @[PMP.scala 311:44]
  assign io_pmp_15_cfg_r = _cfgs_T[120]; // @[PMP.scala 311:44]
  assign io_pmp_15_addr = addr_1_15; // @[PMP.scala 283:15 353:17]
  assign io_pmp_15_mask = mask_1_15; // @[PMP.scala 284:15 353:17]
  assign io_pma_0_cfg_c = _cfgs_T_113[6]; // @[PMP.scala 311:44]
  assign io_pma_0_cfg_atomic = _cfgs_T_113[5]; // @[PMP.scala 311:44]
  assign io_pma_0_cfg_a = _cfgs_T_113[4:3]; // @[PMP.scala 311:44]
  assign io_pma_0_cfg_x = _cfgs_T_113[2]; // @[PMP.scala 311:44]
  assign io_pma_0_cfg_w = _cfgs_T_113[1]; // @[PMP.scala 311:44]
  assign io_pma_0_cfg_r = _cfgs_T_113[0]; // @[PMP.scala 311:44]
  assign io_pma_0_addr = addr_2_0; // @[PMP.scala 283:15 354:17]
  assign io_pma_0_mask = mask_2_0; // @[PMP.scala 284:15 354:17]
  assign io_pma_1_cfg_c = _cfgs_T_113[14]; // @[PMP.scala 311:44]
  assign io_pma_1_cfg_atomic = _cfgs_T_113[13]; // @[PMP.scala 311:44]
  assign io_pma_1_cfg_a = _cfgs_T_113[12:11]; // @[PMP.scala 311:44]
  assign io_pma_1_cfg_x = _cfgs_T_113[10]; // @[PMP.scala 311:44]
  assign io_pma_1_cfg_w = _cfgs_T_113[9]; // @[PMP.scala 311:44]
  assign io_pma_1_cfg_r = _cfgs_T_113[8]; // @[PMP.scala 311:44]
  assign io_pma_1_addr = addr_2_1; // @[PMP.scala 283:15 354:17]
  assign io_pma_1_mask = mask_2_1; // @[PMP.scala 284:15 354:17]
  assign io_pma_2_cfg_c = _cfgs_T_113[22]; // @[PMP.scala 311:44]
  assign io_pma_2_cfg_atomic = _cfgs_T_113[21]; // @[PMP.scala 311:44]
  assign io_pma_2_cfg_a = _cfgs_T_113[20:19]; // @[PMP.scala 311:44]
  assign io_pma_2_cfg_x = _cfgs_T_113[18]; // @[PMP.scala 311:44]
  assign io_pma_2_cfg_w = _cfgs_T_113[17]; // @[PMP.scala 311:44]
  assign io_pma_2_cfg_r = _cfgs_T_113[16]; // @[PMP.scala 311:44]
  assign io_pma_2_addr = addr_2_2; // @[PMP.scala 283:15 354:17]
  assign io_pma_2_mask = mask_2_2; // @[PMP.scala 284:15 354:17]
  assign io_pma_3_cfg_c = _cfgs_T_113[30]; // @[PMP.scala 311:44]
  assign io_pma_3_cfg_atomic = _cfgs_T_113[29]; // @[PMP.scala 311:44]
  assign io_pma_3_cfg_a = _cfgs_T_113[28:27]; // @[PMP.scala 311:44]
  assign io_pma_3_cfg_x = _cfgs_T_113[26]; // @[PMP.scala 311:44]
  assign io_pma_3_cfg_w = _cfgs_T_113[25]; // @[PMP.scala 311:44]
  assign io_pma_3_cfg_r = _cfgs_T_113[24]; // @[PMP.scala 311:44]
  assign io_pma_3_addr = addr_2_3; // @[PMP.scala 283:15 354:17]
  assign io_pma_3_mask = mask_2_3; // @[PMP.scala 284:15 354:17]
  assign io_pma_4_cfg_c = _cfgs_T_113[38]; // @[PMP.scala 311:44]
  assign io_pma_4_cfg_atomic = _cfgs_T_113[37]; // @[PMP.scala 311:44]
  assign io_pma_4_cfg_a = _cfgs_T_113[36:35]; // @[PMP.scala 311:44]
  assign io_pma_4_cfg_x = _cfgs_T_113[34]; // @[PMP.scala 311:44]
  assign io_pma_4_cfg_w = _cfgs_T_113[33]; // @[PMP.scala 311:44]
  assign io_pma_4_cfg_r = _cfgs_T_113[32]; // @[PMP.scala 311:44]
  assign io_pma_4_addr = addr_2_4; // @[PMP.scala 283:15 354:17]
  assign io_pma_4_mask = mask_2_4; // @[PMP.scala 284:15 354:17]
  assign io_pma_5_cfg_c = _cfgs_T_113[46]; // @[PMP.scala 311:44]
  assign io_pma_5_cfg_atomic = _cfgs_T_113[45]; // @[PMP.scala 311:44]
  assign io_pma_5_cfg_a = _cfgs_T_113[44:43]; // @[PMP.scala 311:44]
  assign io_pma_5_cfg_x = _cfgs_T_113[42]; // @[PMP.scala 311:44]
  assign io_pma_5_cfg_w = _cfgs_T_113[41]; // @[PMP.scala 311:44]
  assign io_pma_5_cfg_r = _cfgs_T_113[40]; // @[PMP.scala 311:44]
  assign io_pma_5_addr = addr_2_5; // @[PMP.scala 283:15 354:17]
  assign io_pma_5_mask = mask_2_5; // @[PMP.scala 284:15 354:17]
  assign io_pma_6_cfg_c = _cfgs_T_113[54]; // @[PMP.scala 311:44]
  assign io_pma_6_cfg_atomic = _cfgs_T_113[53]; // @[PMP.scala 311:44]
  assign io_pma_6_cfg_a = _cfgs_T_113[52:51]; // @[PMP.scala 311:44]
  assign io_pma_6_cfg_x = _cfgs_T_113[50]; // @[PMP.scala 311:44]
  assign io_pma_6_cfg_w = _cfgs_T_113[49]; // @[PMP.scala 311:44]
  assign io_pma_6_cfg_r = _cfgs_T_113[48]; // @[PMP.scala 311:44]
  assign io_pma_6_addr = addr_2_6; // @[PMP.scala 283:15 354:17]
  assign io_pma_6_mask = mask_2_6; // @[PMP.scala 284:15 354:17]
  assign io_pma_7_cfg_c = _cfgs_T_113[62]; // @[PMP.scala 311:44]
  assign io_pma_7_cfg_atomic = _cfgs_T_113[61]; // @[PMP.scala 311:44]
  assign io_pma_7_cfg_a = _cfgs_T_113[60:59]; // @[PMP.scala 311:44]
  assign io_pma_7_cfg_x = _cfgs_T_113[58]; // @[PMP.scala 311:44]
  assign io_pma_7_cfg_w = _cfgs_T_113[57]; // @[PMP.scala 311:44]
  assign io_pma_7_cfg_r = _cfgs_T_113[56]; // @[PMP.scala 311:44]
  assign io_pma_7_addr = addr_2_7; // @[PMP.scala 283:15 354:17]
  assign io_pma_7_mask = mask_2_7; // @[PMP.scala 284:15 354:17]
  assign io_pma_8_cfg_c = _cfgs_T_113[70]; // @[PMP.scala 311:44]
  assign io_pma_8_cfg_atomic = _cfgs_T_113[69]; // @[PMP.scala 311:44]
  assign io_pma_8_cfg_a = _cfgs_T_113[68:67]; // @[PMP.scala 311:44]
  assign io_pma_8_cfg_x = _cfgs_T_113[66]; // @[PMP.scala 311:44]
  assign io_pma_8_cfg_w = _cfgs_T_113[65]; // @[PMP.scala 311:44]
  assign io_pma_8_cfg_r = _cfgs_T_113[64]; // @[PMP.scala 311:44]
  assign io_pma_8_addr = addr_2_8; // @[PMP.scala 283:15 354:17]
  assign io_pma_8_mask = mask_2_8; // @[PMP.scala 284:15 354:17]
  assign io_pma_9_cfg_c = _cfgs_T_113[78]; // @[PMP.scala 311:44]
  assign io_pma_9_cfg_atomic = _cfgs_T_113[77]; // @[PMP.scala 311:44]
  assign io_pma_9_cfg_a = _cfgs_T_113[76:75]; // @[PMP.scala 311:44]
  assign io_pma_9_cfg_x = _cfgs_T_113[74]; // @[PMP.scala 311:44]
  assign io_pma_9_cfg_w = _cfgs_T_113[73]; // @[PMP.scala 311:44]
  assign io_pma_9_cfg_r = _cfgs_T_113[72]; // @[PMP.scala 311:44]
  assign io_pma_9_addr = addr_2_9; // @[PMP.scala 283:15 354:17]
  assign io_pma_9_mask = mask_2_9; // @[PMP.scala 284:15 354:17]
  assign io_pma_10_cfg_c = _cfgs_T_113[86]; // @[PMP.scala 311:44]
  assign io_pma_10_cfg_atomic = _cfgs_T_113[85]; // @[PMP.scala 311:44]
  assign io_pma_10_cfg_a = _cfgs_T_113[84:83]; // @[PMP.scala 311:44]
  assign io_pma_10_cfg_x = _cfgs_T_113[82]; // @[PMP.scala 311:44]
  assign io_pma_10_cfg_w = _cfgs_T_113[81]; // @[PMP.scala 311:44]
  assign io_pma_10_cfg_r = _cfgs_T_113[80]; // @[PMP.scala 311:44]
  assign io_pma_10_addr = addr_2_10; // @[PMP.scala 283:15 354:17]
  assign io_pma_10_mask = mask_2_10; // @[PMP.scala 284:15 354:17]
  assign io_pma_11_cfg_c = _cfgs_T_113[94]; // @[PMP.scala 311:44]
  assign io_pma_11_cfg_atomic = _cfgs_T_113[93]; // @[PMP.scala 311:44]
  assign io_pma_11_cfg_a = _cfgs_T_113[92:91]; // @[PMP.scala 311:44]
  assign io_pma_11_cfg_x = _cfgs_T_113[90]; // @[PMP.scala 311:44]
  assign io_pma_11_cfg_w = _cfgs_T_113[89]; // @[PMP.scala 311:44]
  assign io_pma_11_cfg_r = _cfgs_T_113[88]; // @[PMP.scala 311:44]
  assign io_pma_11_addr = addr_2_11; // @[PMP.scala 283:15 354:17]
  assign io_pma_11_mask = mask_2_11; // @[PMP.scala 284:15 354:17]
  assign io_pma_12_cfg_c = _cfgs_T_113[102]; // @[PMP.scala 311:44]
  assign io_pma_12_cfg_atomic = _cfgs_T_113[101]; // @[PMP.scala 311:44]
  assign io_pma_12_cfg_a = _cfgs_T_113[100:99]; // @[PMP.scala 311:44]
  assign io_pma_12_cfg_x = _cfgs_T_113[98]; // @[PMP.scala 311:44]
  assign io_pma_12_cfg_w = _cfgs_T_113[97]; // @[PMP.scala 311:44]
  assign io_pma_12_cfg_r = _cfgs_T_113[96]; // @[PMP.scala 311:44]
  assign io_pma_12_addr = addr_2_12; // @[PMP.scala 283:15 354:17]
  assign io_pma_12_mask = mask_2_12; // @[PMP.scala 284:15 354:17]
  assign io_pma_13_cfg_c = _cfgs_T_113[110]; // @[PMP.scala 311:44]
  assign io_pma_13_cfg_atomic = _cfgs_T_113[109]; // @[PMP.scala 311:44]
  assign io_pma_13_cfg_a = _cfgs_T_113[108:107]; // @[PMP.scala 311:44]
  assign io_pma_13_cfg_x = _cfgs_T_113[106]; // @[PMP.scala 311:44]
  assign io_pma_13_cfg_w = _cfgs_T_113[105]; // @[PMP.scala 311:44]
  assign io_pma_13_cfg_r = _cfgs_T_113[104]; // @[PMP.scala 311:44]
  assign io_pma_13_addr = addr_2_13; // @[PMP.scala 283:15 354:17]
  assign io_pma_13_mask = mask_2_13; // @[PMP.scala 284:15 354:17]
  assign io_pma_14_cfg_c = _cfgs_T_113[118]; // @[PMP.scala 311:44]
  assign io_pma_14_cfg_atomic = _cfgs_T_113[117]; // @[PMP.scala 311:44]
  assign io_pma_14_cfg_a = _cfgs_T_113[116:115]; // @[PMP.scala 311:44]
  assign io_pma_14_cfg_x = _cfgs_T_113[114]; // @[PMP.scala 311:44]
  assign io_pma_14_cfg_w = _cfgs_T_113[113]; // @[PMP.scala 311:44]
  assign io_pma_14_cfg_r = _cfgs_T_113[112]; // @[PMP.scala 311:44]
  assign io_pma_14_addr = addr_2_14; // @[PMP.scala 283:15 354:17]
  assign io_pma_14_mask = mask_2_14; // @[PMP.scala 284:15 354:17]
  assign io_pma_15_cfg_c = _cfgs_T_113[126]; // @[PMP.scala 311:44]
  assign io_pma_15_cfg_atomic = _cfgs_T_113[125]; // @[PMP.scala 311:44]
  assign io_pma_15_cfg_a = _cfgs_T_113[124:123]; // @[PMP.scala 311:44]
  assign io_pma_15_cfg_x = _cfgs_T_113[122]; // @[PMP.scala 311:44]
  assign io_pma_15_cfg_w = _cfgs_T_113[121]; // @[PMP.scala 311:44]
  assign io_pma_15_cfg_r = _cfgs_T_113[120]; // @[PMP.scala 311:44]
  assign io_pma_15_addr = addr_2_15; // @[PMP.scala 283:15 354:17]
  assign io_pma_15_mask = mask_2_15; // @[PMP.scala 284:15 354:17]
  always @(posedge clock) begin
    addr_1_0 <= _GEN_128[33:0];
    addr_1_1 <= _GEN_6[33:0];
    addr_1_2 <= _GEN_136[33:0];
    addr_1_3 <= _GEN_120[33:0];
    addr_1_4 <= _GEN_65[33:0];
    addr_1_5 <= _GEN_51[33:0];
    addr_1_6 <= _GEN_144[33:0];
    addr_1_7 <= _GEN_132[33:0];
    addr_1_8 <= _GEN_63[33:0];
    addr_1_9 <= _GEN_110[33:0];
    addr_1_10 <= _GEN_130[33:0];
    addr_1_11 <= _GEN_187[33:0];
    addr_1_12 <= _GEN_55[33:0];
    addr_1_13 <= _GEN_61[33:0];
    addr_1_14 <= _GEN_116[33:0];
    addr_1_15 <= _GEN_124[33:0];
    mask_1_0 <= _GEN_220[35:0];
    mask_1_1 <= _GEN_221[35:0];
    mask_1_2 <= _GEN_222[35:0];
    mask_1_3 <= _GEN_223[35:0];
    mask_1_4 <= _GEN_224[35:0];
    mask_1_5 <= _GEN_225[35:0];
    mask_1_6 <= _GEN_226[35:0];
    mask_1_7 <= _GEN_227[35:0];
    mask_1_8 <= _GEN_62[35:0];
    mask_1_9 <= _GEN_109[35:0];
    mask_1_10 <= _GEN_129[35:0];
    mask_1_11 <= _GEN_186[35:0];
    mask_1_12 <= _GEN_54[35:0];
    mask_1_13 <= _GEN_60[35:0];
    mask_1_14 <= _GEN_115[35:0];
    mask_1_15 <= _GEN_123[35:0];
    if (io_distribute_csr_wvalid) begin // @[Reg.scala 17:18]
      wdata_reg <= io_distribute_csr_wdata; // @[Reg.scala 17:22]
    end
    wen_reg <= io_distribute_csr_wvalid & io_distribute_csr_waddr == 12'h7cb; // @[RegMap.scala 55:35]
    wen_reg_1 <= io_distribute_csr_wvalid & io_distribute_csr_waddr == 12'h7cf; // @[RegMap.scala 55:35]
    wen_reg_2 <= io_distribute_csr_wvalid & io_distribute_csr_waddr == 12'h3b1; // @[RegMap.scala 55:35]
    wen_reg_3 <= io_distribute_csr_wvalid & io_distribute_csr_waddr == 12'h3a2; // @[RegMap.scala 55:35]
    wen_reg_4 <= io_distribute_csr_wvalid & io_distribute_csr_waddr == 12'h7c8; // @[RegMap.scala 55:35]
    wen_reg_5 <= io_distribute_csr_wvalid & io_distribute_csr_waddr == 12'h3b5; // @[RegMap.scala 55:35]
    wen_reg_6 <= io_distribute_csr_wvalid & io_distribute_csr_waddr == 12'h7d7; // @[RegMap.scala 55:35]
    wen_reg_7 <= io_distribute_csr_wvalid & io_distribute_csr_waddr == 12'h3bc; // @[RegMap.scala 55:35]
    wen_reg_8 <= io_distribute_csr_wvalid & io_distribute_csr_waddr == 12'h7d2; // @[RegMap.scala 55:35]
    wen_reg_9 <= io_distribute_csr_wvalid & io_distribute_csr_waddr == 12'h7d0; // @[RegMap.scala 55:35]
    wen_reg_10 <= io_distribute_csr_wvalid & io_distribute_csr_waddr == 12'h3bd; // @[RegMap.scala 55:35]
    wen_reg_11 <= io_distribute_csr_wvalid & io_distribute_csr_waddr == 12'h3b8; // @[RegMap.scala 55:35]
    wen_reg_12 <= io_distribute_csr_wvalid & io_distribute_csr_waddr == 12'h3b4; // @[RegMap.scala 55:35]
    wen_reg_13 <= io_distribute_csr_wvalid & io_distribute_csr_waddr == 12'h7d6; // @[RegMap.scala 55:35]
    wen_reg_14 <= io_distribute_csr_wvalid & io_distribute_csr_waddr == 12'h7c0; // @[RegMap.scala 55:35]
    wen_reg_15 <= io_distribute_csr_wvalid & io_distribute_csr_waddr == 12'h3b9; // @[RegMap.scala 55:35]
    wen_reg_16 <= io_distribute_csr_wvalid & io_distribute_csr_waddr == 12'h7cc; // @[RegMap.scala 55:35]
    wen_reg_17 <= io_distribute_csr_wvalid & io_distribute_csr_waddr == 12'h7d1; // @[RegMap.scala 55:35]
    wen_reg_18 <= io_distribute_csr_wvalid & io_distribute_csr_waddr == 12'h3be; // @[RegMap.scala 55:35]
    wen_reg_19 <= io_distribute_csr_wvalid & io_distribute_csr_waddr == 12'h7cd; // @[RegMap.scala 55:35]
    wen_reg_20 <= io_distribute_csr_wvalid & io_distribute_csr_waddr == 12'h3b3; // @[RegMap.scala 55:35]
    wen_reg_21 <= io_distribute_csr_wvalid & io_distribute_csr_waddr == 12'h7c9; // @[RegMap.scala 55:35]
    wen_reg_22 <= io_distribute_csr_wvalid & io_distribute_csr_waddr == 12'h3bf; // @[RegMap.scala 55:35]
    wen_reg_23 <= io_distribute_csr_wvalid & io_distribute_csr_waddr == 12'h7d5; // @[RegMap.scala 55:35]
    wen_reg_24 <= io_distribute_csr_wvalid & io_distribute_csr_waddr == 12'h3b0; // @[RegMap.scala 55:35]
    wen_reg_25 <= io_distribute_csr_wvalid & io_distribute_csr_waddr == 12'h3ba; // @[RegMap.scala 55:35]
    wen_reg_26 <= io_distribute_csr_wvalid & io_distribute_csr_waddr == 12'h3b7; // @[RegMap.scala 55:35]
    wen_reg_27 <= io_distribute_csr_wvalid & io_distribute_csr_waddr == 12'h7ce; // @[RegMap.scala 55:35]
    wen_reg_28 <= io_distribute_csr_wvalid & io_distribute_csr_waddr == 12'h3b2; // @[RegMap.scala 55:35]
    wen_reg_29 <= io_distribute_csr_wvalid & io_distribute_csr_waddr == 12'h7d4; // @[RegMap.scala 55:35]
    wen_reg_30 <= io_distribute_csr_wvalid & io_distribute_csr_waddr == 12'h7ca; // @[RegMap.scala 55:35]
    wen_reg_31 <= io_distribute_csr_wvalid & io_distribute_csr_waddr == 12'h7d3; // @[RegMap.scala 55:35]
    wen_reg_32 <= io_distribute_csr_wvalid & io_distribute_csr_waddr == 12'h3b6; // @[RegMap.scala 55:35]
    wen_reg_33 <= io_distribute_csr_wvalid & io_distribute_csr_waddr == 12'h7c2; // @[RegMap.scala 55:35]
    wen_reg_34 <= io_distribute_csr_wvalid & io_distribute_csr_waddr == 12'h3bb; // @[RegMap.scala 55:35]
    wen_reg_35 <= io_distribute_csr_wvalid & io_distribute_csr_waddr == 12'h3a0; // @[RegMap.scala 55:35]
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[RegMap.scala 56:24]
      cfgMerged__0 <= 64'h0; // @[RegMap.scala 56:28]
    end else if (wen_reg_35) begin // @[PMP.scala 310:28]
      cfgMerged__0 <= _cfgMerged_1_T_20;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[RegMap.scala 56:24]
      cfgMerged__1 <= 64'h0; // @[RegMap.scala 56:28]
    end else if (wen_reg_3) begin // @[PMP.scala 310:28]
      cfgMerged__1 <= _cfgMerged_1_T_20;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[RegMap.scala 56:24]
      cfgMerged_1_0 <= 64'hf0b0b0b0f0b0000; // @[RegMap.scala 56:28]
    end else if (wen_reg_14) begin // @[PMP.scala 310:28]
      cfgMerged_1_0 <= _cfgMerged_1_T_20;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[RegMap.scala 56:24]
      cfgMerged_1_1 <= 64'h7f1b080b080b080b; // @[RegMap.scala 56:28]
    end else if (wen_reg_33) begin // @[PMP.scala 310:28]
      cfgMerged_1_1 <= _cfgMerged_1_T_20;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PMP.scala 312:23]
      addr_2_0 <= 34'h0; // @[PMP.scala 312:23]
    end else begin
      addr_2_0 <= _GEN_49[33:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PMP.scala 312:23]
      addr_2_1 <= 34'h0; // @[PMP.scala 312:23]
    end else begin
      addr_2_1 <= _GEN_122[33:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PMP.scala 312:23]
      addr_2_2 <= 34'h4000000; // @[PMP.scala 312:23]
    end else begin
      addr_2_2 <= _GEN_140[33:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PMP.scala 312:23]
      addr_2_3 <= 34'h8000000; // @[PMP.scala 312:23]
    end else begin
      addr_2_3 <= _GEN_2[33:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PMP.scala 312:23]
      addr_2_4 <= 34'hc004000; // @[PMP.scala 312:23]
    end else begin
      addr_2_4 <= _GEN_112[33:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PMP.scala 312:23]
      addr_2_5 <= 34'hc014000; // @[PMP.scala 312:23]
    end else begin
      addr_2_5 <= _GEN_118[33:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PMP.scala 312:23]
      addr_2_6 <= 34'he008000; // @[PMP.scala 312:23]
    end else begin
      addr_2_6 <= _GEN_134[33:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PMP.scala 312:23]
      addr_2_7 <= 34'he008400; // @[PMP.scala 312:23]
    end else begin
      addr_2_7 <= _GEN_4[33:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PMP.scala 312:23]
      addr_2_8 <= 34'he008800; // @[PMP.scala 312:23]
    end else begin
      addr_2_8 <= _GEN_59[33:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PMP.scala 312:23]
      addr_2_9 <= 34'he400000; // @[PMP.scala 312:23]
    end else begin
      addr_2_9 <= _GEN_114[33:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PMP.scala 312:23]
      addr_2_10 <= 34'he400800; // @[PMP.scala 312:23]
    end else begin
      addr_2_10 <= _GEN_57[33:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PMP.scala 312:23]
      addr_2_11 <= 34'he800000; // @[PMP.scala 312:23]
    end else begin
      addr_2_11 <= _GEN_142[33:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PMP.scala 312:23]
      addr_2_12 <= 34'he800400; // @[PMP.scala 312:23]
    end else begin
      addr_2_12 <= _GEN_138[33:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PMP.scala 312:23]
      addr_2_13 <= 34'hf000000; // @[PMP.scala 312:23]
    end else begin
      addr_2_13 <= _GEN_126[33:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PMP.scala 312:23]
      addr_2_14 <= 34'hfffffff; // @[PMP.scala 312:23]
    end else begin
      addr_2_14 <= _GEN_67[33:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PMP.scala 312:23]
      addr_2_15 <= 34'h1ffffffff; // @[PMP.scala 312:23]
    end else begin
      addr_2_15 <= _GEN_53[33:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PMP.scala 313:23]
      mask_2_0 <= 36'hfff; // @[PMP.scala 313:23]
    end else begin
      mask_2_0 <= _GEN_100[35:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PMP.scala 313:23]
      mask_2_1 <= 36'hfff; // @[PMP.scala 313:23]
    end else begin
      mask_2_1 <= _GEN_121[35:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PMP.scala 313:23]
      mask_2_2 <= 36'hfff; // @[PMP.scala 313:23]
    end else begin
      mask_2_2 <= _GEN_139[35:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PMP.scala 313:23]
      mask_2_3 <= 36'hfff; // @[PMP.scala 313:23]
    end else begin
      mask_2_3 <= _GEN_103[35:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PMP.scala 313:23]
      mask_2_4 <= 36'hfff; // @[PMP.scala 313:23]
    end else begin
      mask_2_4 <= _GEN_111[35:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PMP.scala 313:23]
      mask_2_5 <= 36'hfff; // @[PMP.scala 313:23]
    end else begin
      mask_2_5 <= _GEN_117[35:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PMP.scala 313:23]
      mask_2_6 <= 36'hfff; // @[PMP.scala 313:23]
    end else begin
      mask_2_6 <= _GEN_133[35:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PMP.scala 313:23]
      mask_2_7 <= 36'hfff; // @[PMP.scala 313:23]
    end else begin
      mask_2_7 <= _GEN_107[35:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PMP.scala 313:23]
      mask_2_8 <= 36'hfff; // @[PMP.scala 313:23]
    end else begin
      mask_2_8 <= _GEN_177[35:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PMP.scala 313:23]
      mask_2_9 <= 36'hfff; // @[PMP.scala 313:23]
    end else begin
      mask_2_9 <= _GEN_178[35:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PMP.scala 313:23]
      mask_2_10 <= 36'hfff; // @[PMP.scala 313:23]
    end else begin
      mask_2_10 <= _GEN_179[35:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PMP.scala 313:23]
      mask_2_11 <= 36'hfff; // @[PMP.scala 313:23]
    end else begin
      mask_2_11 <= _GEN_180[35:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PMP.scala 313:23]
      mask_2_12 <= 36'hfff; // @[PMP.scala 313:23]
    end else begin
      mask_2_12 <= _GEN_181[35:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PMP.scala 313:23]
      mask_2_13 <= 36'hfff; // @[PMP.scala 313:23]
    end else begin
      mask_2_13 <= _GEN_182[35:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PMP.scala 313:23]
      mask_2_14 <= 36'h7fffffff; // @[PMP.scala 313:23]
    end else begin
      mask_2_14 <= _GEN_183[35:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PMP.scala 313:23]
      mask_2_15 <= 36'hfffffffff; // @[PMP.scala 313:23]
    end else begin
      mask_2_15 <= _GEN_184[35:0];
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  cfgMerged__0 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  cfgMerged__1 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  addr_1_0 = _RAND_2[33:0];
  _RAND_3 = {2{`RANDOM}};
  addr_1_1 = _RAND_3[33:0];
  _RAND_4 = {2{`RANDOM}};
  addr_1_2 = _RAND_4[33:0];
  _RAND_5 = {2{`RANDOM}};
  addr_1_3 = _RAND_5[33:0];
  _RAND_6 = {2{`RANDOM}};
  addr_1_4 = _RAND_6[33:0];
  _RAND_7 = {2{`RANDOM}};
  addr_1_5 = _RAND_7[33:0];
  _RAND_8 = {2{`RANDOM}};
  addr_1_6 = _RAND_8[33:0];
  _RAND_9 = {2{`RANDOM}};
  addr_1_7 = _RAND_9[33:0];
  _RAND_10 = {2{`RANDOM}};
  addr_1_8 = _RAND_10[33:0];
  _RAND_11 = {2{`RANDOM}};
  addr_1_9 = _RAND_11[33:0];
  _RAND_12 = {2{`RANDOM}};
  addr_1_10 = _RAND_12[33:0];
  _RAND_13 = {2{`RANDOM}};
  addr_1_11 = _RAND_13[33:0];
  _RAND_14 = {2{`RANDOM}};
  addr_1_12 = _RAND_14[33:0];
  _RAND_15 = {2{`RANDOM}};
  addr_1_13 = _RAND_15[33:0];
  _RAND_16 = {2{`RANDOM}};
  addr_1_14 = _RAND_16[33:0];
  _RAND_17 = {2{`RANDOM}};
  addr_1_15 = _RAND_17[33:0];
  _RAND_18 = {2{`RANDOM}};
  mask_1_0 = _RAND_18[35:0];
  _RAND_19 = {2{`RANDOM}};
  mask_1_1 = _RAND_19[35:0];
  _RAND_20 = {2{`RANDOM}};
  mask_1_2 = _RAND_20[35:0];
  _RAND_21 = {2{`RANDOM}};
  mask_1_3 = _RAND_21[35:0];
  _RAND_22 = {2{`RANDOM}};
  mask_1_4 = _RAND_22[35:0];
  _RAND_23 = {2{`RANDOM}};
  mask_1_5 = _RAND_23[35:0];
  _RAND_24 = {2{`RANDOM}};
  mask_1_6 = _RAND_24[35:0];
  _RAND_25 = {2{`RANDOM}};
  mask_1_7 = _RAND_25[35:0];
  _RAND_26 = {2{`RANDOM}};
  mask_1_8 = _RAND_26[35:0];
  _RAND_27 = {2{`RANDOM}};
  mask_1_9 = _RAND_27[35:0];
  _RAND_28 = {2{`RANDOM}};
  mask_1_10 = _RAND_28[35:0];
  _RAND_29 = {2{`RANDOM}};
  mask_1_11 = _RAND_29[35:0];
  _RAND_30 = {2{`RANDOM}};
  mask_1_12 = _RAND_30[35:0];
  _RAND_31 = {2{`RANDOM}};
  mask_1_13 = _RAND_31[35:0];
  _RAND_32 = {2{`RANDOM}};
  mask_1_14 = _RAND_32[35:0];
  _RAND_33 = {2{`RANDOM}};
  mask_1_15 = _RAND_33[35:0];
  _RAND_34 = {2{`RANDOM}};
  cfgMerged_1_0 = _RAND_34[63:0];
  _RAND_35 = {2{`RANDOM}};
  cfgMerged_1_1 = _RAND_35[63:0];
  _RAND_36 = {2{`RANDOM}};
  addr_2_0 = _RAND_36[33:0];
  _RAND_37 = {2{`RANDOM}};
  addr_2_1 = _RAND_37[33:0];
  _RAND_38 = {2{`RANDOM}};
  addr_2_2 = _RAND_38[33:0];
  _RAND_39 = {2{`RANDOM}};
  addr_2_3 = _RAND_39[33:0];
  _RAND_40 = {2{`RANDOM}};
  addr_2_4 = _RAND_40[33:0];
  _RAND_41 = {2{`RANDOM}};
  addr_2_5 = _RAND_41[33:0];
  _RAND_42 = {2{`RANDOM}};
  addr_2_6 = _RAND_42[33:0];
  _RAND_43 = {2{`RANDOM}};
  addr_2_7 = _RAND_43[33:0];
  _RAND_44 = {2{`RANDOM}};
  addr_2_8 = _RAND_44[33:0];
  _RAND_45 = {2{`RANDOM}};
  addr_2_9 = _RAND_45[33:0];
  _RAND_46 = {2{`RANDOM}};
  addr_2_10 = _RAND_46[33:0];
  _RAND_47 = {2{`RANDOM}};
  addr_2_11 = _RAND_47[33:0];
  _RAND_48 = {2{`RANDOM}};
  addr_2_12 = _RAND_48[33:0];
  _RAND_49 = {2{`RANDOM}};
  addr_2_13 = _RAND_49[33:0];
  _RAND_50 = {2{`RANDOM}};
  addr_2_14 = _RAND_50[33:0];
  _RAND_51 = {2{`RANDOM}};
  addr_2_15 = _RAND_51[33:0];
  _RAND_52 = {2{`RANDOM}};
  mask_2_0 = _RAND_52[35:0];
  _RAND_53 = {2{`RANDOM}};
  mask_2_1 = _RAND_53[35:0];
  _RAND_54 = {2{`RANDOM}};
  mask_2_2 = _RAND_54[35:0];
  _RAND_55 = {2{`RANDOM}};
  mask_2_3 = _RAND_55[35:0];
  _RAND_56 = {2{`RANDOM}};
  mask_2_4 = _RAND_56[35:0];
  _RAND_57 = {2{`RANDOM}};
  mask_2_5 = _RAND_57[35:0];
  _RAND_58 = {2{`RANDOM}};
  mask_2_6 = _RAND_58[35:0];
  _RAND_59 = {2{`RANDOM}};
  mask_2_7 = _RAND_59[35:0];
  _RAND_60 = {2{`RANDOM}};
  mask_2_8 = _RAND_60[35:0];
  _RAND_61 = {2{`RANDOM}};
  mask_2_9 = _RAND_61[35:0];
  _RAND_62 = {2{`RANDOM}};
  mask_2_10 = _RAND_62[35:0];
  _RAND_63 = {2{`RANDOM}};
  mask_2_11 = _RAND_63[35:0];
  _RAND_64 = {2{`RANDOM}};
  mask_2_12 = _RAND_64[35:0];
  _RAND_65 = {2{`RANDOM}};
  mask_2_13 = _RAND_65[35:0];
  _RAND_66 = {2{`RANDOM}};
  mask_2_14 = _RAND_66[35:0];
  _RAND_67 = {2{`RANDOM}};
  mask_2_15 = _RAND_67[35:0];
  _RAND_68 = {2{`RANDOM}};
  wdata_reg = _RAND_68[63:0];
  _RAND_69 = {1{`RANDOM}};
  wen_reg = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  wen_reg_1 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  wen_reg_2 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  wen_reg_3 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  wen_reg_4 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  wen_reg_5 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  wen_reg_6 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  wen_reg_7 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  wen_reg_8 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  wen_reg_9 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  wen_reg_10 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  wen_reg_11 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  wen_reg_12 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  wen_reg_13 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  wen_reg_14 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  wen_reg_15 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  wen_reg_16 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  wen_reg_17 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  wen_reg_18 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  wen_reg_19 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  wen_reg_20 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  wen_reg_21 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  wen_reg_22 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  wen_reg_23 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  wen_reg_24 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  wen_reg_25 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  wen_reg_26 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  wen_reg_27 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  wen_reg_28 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  wen_reg_29 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  wen_reg_30 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  wen_reg_31 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  wen_reg_32 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  wen_reg_33 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  wen_reg_34 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  wen_reg_35 = _RAND_104[0:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    cfgMerged__0 = 64'h0;
  end
  if (reset) begin
    cfgMerged__1 = 64'h0;
  end
  if (reset) begin
    cfgMerged_1_0 = 64'hf0b0b0b0f0b0000;
  end
  if (reset) begin
    cfgMerged_1_1 = 64'h7f1b080b080b080b;
  end
  if (reset) begin
    addr_2_0 = 34'h0;
  end
  if (reset) begin
    addr_2_1 = 34'h0;
  end
  if (reset) begin
    addr_2_2 = 34'h4000000;
  end
  if (reset) begin
    addr_2_3 = 34'h8000000;
  end
  if (reset) begin
    addr_2_4 = 34'hc004000;
  end
  if (reset) begin
    addr_2_5 = 34'hc014000;
  end
  if (reset) begin
    addr_2_6 = 34'he008000;
  end
  if (reset) begin
    addr_2_7 = 34'he008400;
  end
  if (reset) begin
    addr_2_8 = 34'he008800;
  end
  if (reset) begin
    addr_2_9 = 34'he400000;
  end
  if (reset) begin
    addr_2_10 = 34'he400800;
  end
  if (reset) begin
    addr_2_11 = 34'he800000;
  end
  if (reset) begin
    addr_2_12 = 34'he800400;
  end
  if (reset) begin
    addr_2_13 = 34'hf000000;
  end
  if (reset) begin
    addr_2_14 = 34'hfffffff;
  end
  if (reset) begin
    addr_2_15 = 34'h1ffffffff;
  end
  if (reset) begin
    mask_2_0 = 36'hfff;
  end
  if (reset) begin
    mask_2_1 = 36'hfff;
  end
  if (reset) begin
    mask_2_2 = 36'hfff;
  end
  if (reset) begin
    mask_2_3 = 36'hfff;
  end
  if (reset) begin
    mask_2_4 = 36'hfff;
  end
  if (reset) begin
    mask_2_5 = 36'hfff;
  end
  if (reset) begin
    mask_2_6 = 36'hfff;
  end
  if (reset) begin
    mask_2_7 = 36'hfff;
  end
  if (reset) begin
    mask_2_8 = 36'hfff;
  end
  if (reset) begin
    mask_2_9 = 36'hfff;
  end
  if (reset) begin
    mask_2_10 = 36'hfff;
  end
  if (reset) begin
    mask_2_11 = 36'hfff;
  end
  if (reset) begin
    mask_2_12 = 36'hfff;
  end
  if (reset) begin
    mask_2_13 = 36'hfff;
  end
  if (reset) begin
    mask_2_14 = 36'h7fffffff;
  end
  if (reset) begin
    mask_2_15 = 36'hfffffffff;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule

