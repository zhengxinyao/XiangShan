module CSA3_2_1978(
  input  [9:0] io_in_0,
  input  [9:0] io_in_1,
  input  [9:0] io_in_2,
  output [9:0] io_out_0,
  output [9:0] io_out_1
);
  wire  a = io_in_0[0]; // @[CSA.scala 43:32]
  wire  b = io_in_1[0]; // @[CSA.scala 43:45]
  wire  cin = io_in_2[0]; // @[CSA.scala 43:58]
  wire  a_xor_b = a ^ b; // @[CSA.scala 44:21]
  wire  a_and_b = a & b; // @[CSA.scala 45:21]
  wire  sum = a_xor_b ^ cin; // @[CSA.scala 46:23]
  wire  cout = a_and_b | a_xor_b & cin; // @[CSA.scala 47:24]
  wire [1:0] temp_0 = {cout,sum}; // @[Cat.scala 31:58]
  wire  a_1 = io_in_0[1]; // @[CSA.scala 43:32]
  wire  b_1 = io_in_1[1]; // @[CSA.scala 43:45]
  wire  cin_1 = io_in_2[1]; // @[CSA.scala 43:58]
  wire  a_xor_b1 = a_1 ^ b_1; // @[CSA.scala 44:21]
  wire  a_and_b1 = a_1 & b_1; // @[CSA.scala 45:21]
  wire  sum_1 = a_xor_b1 ^ cin_1; // @[CSA.scala 46:23]
  wire  cout_1 = a_and_b1 | a_xor_b1 & cin_1; // @[CSA.scala 47:24]
  wire [1:0] temp_1 = {cout_1,sum_1}; // @[Cat.scala 31:58]
  wire  a_2 = io_in_0[2]; // @[CSA.scala 43:32]
  wire  b_2 = io_in_1[2]; // @[CSA.scala 43:45]
  wire  cin_2 = io_in_2[2]; // @[CSA.scala 43:58]
  wire  a_xor_b2 = a_2 ^ b_2; // @[CSA.scala 44:21]
  wire  a_and_b2 = a_2 & b_2; // @[CSA.scala 45:21]
  wire  sum_2 = a_xor_b2 ^ cin_2; // @[CSA.scala 46:23]
  wire  cout_2 = a_and_b2 | a_xor_b2 & cin_2; // @[CSA.scala 47:24]
  wire [1:0] temp_2 = {cout_2,sum_2}; // @[Cat.scala 31:58]
  wire  a_3 = io_in_0[3]; // @[CSA.scala 43:32]
  wire  b_3 = io_in_1[3]; // @[CSA.scala 43:45]
  wire  cin_3 = io_in_2[3]; // @[CSA.scala 43:58]
  wire  a_xor_b3 = a_3 ^ b_3; // @[CSA.scala 44:21]
  wire  a_and_b3 = a_3 & b_3; // @[CSA.scala 45:21]
  wire  sum_3 = a_xor_b3 ^ cin_3; // @[CSA.scala 46:23]
  wire  cout_3 = a_and_b3 | a_xor_b3 & cin_3; // @[CSA.scala 47:24]
  wire [1:0] temp_3 = {cout_3,sum_3}; // @[Cat.scala 31:58]
  wire  a_4 = io_in_0[4]; // @[CSA.scala 43:32]
  wire  b_4 = io_in_1[4]; // @[CSA.scala 43:45]
  wire  cin_4 = io_in_2[4]; // @[CSA.scala 43:58]
  wire  a_xor_b4 = a_4 ^ b_4; // @[CSA.scala 44:21]
  wire  a_and_b4 = a_4 & b_4; // @[CSA.scala 45:21]
  wire  sum_4 = a_xor_b4 ^ cin_4; // @[CSA.scala 46:23]
  wire  cout_4 = a_and_b4 | a_xor_b4 & cin_4; // @[CSA.scala 47:24]
  wire [1:0] temp_4 = {cout_4,sum_4}; // @[Cat.scala 31:58]
  wire  a_5 = io_in_0[5]; // @[CSA.scala 43:32]
  wire  b_5 = io_in_1[5]; // @[CSA.scala 43:45]
  wire  cin_5 = io_in_2[5]; // @[CSA.scala 43:58]
  wire  a_xor_b5 = a_5 ^ b_5; // @[CSA.scala 44:21]
  wire  a_and_b5 = a_5 & b_5; // @[CSA.scala 45:21]
  wire  sum_5 = a_xor_b5 ^ cin_5; // @[CSA.scala 46:23]
  wire  cout_5 = a_and_b5 | a_xor_b5 & cin_5; // @[CSA.scala 47:24]
  wire [1:0] temp_5 = {cout_5,sum_5}; // @[Cat.scala 31:58]
  wire  a_6 = io_in_0[6]; // @[CSA.scala 43:32]
  wire  b_6 = io_in_1[6]; // @[CSA.scala 43:45]
  wire  cin_6 = io_in_2[6]; // @[CSA.scala 43:58]
  wire  a_xor_b6 = a_6 ^ b_6; // @[CSA.scala 44:21]
  wire  a_and_b6 = a_6 & b_6; // @[CSA.scala 45:21]
  wire  sum_6 = a_xor_b6 ^ cin_6; // @[CSA.scala 46:23]
  wire  cout_6 = a_and_b6 | a_xor_b6 & cin_6; // @[CSA.scala 47:24]
  wire [1:0] temp_6 = {cout_6,sum_6}; // @[Cat.scala 31:58]
  wire  a_7 = io_in_0[7]; // @[CSA.scala 43:32]
  wire  b_7 = io_in_1[7]; // @[CSA.scala 43:45]
  wire  cin_7 = io_in_2[7]; // @[CSA.scala 43:58]
  wire  a_xor_b7 = a_7 ^ b_7; // @[CSA.scala 44:21]
  wire  a_and_b7 = a_7 & b_7; // @[CSA.scala 45:21]
  wire  sum_7 = a_xor_b7 ^ cin_7; // @[CSA.scala 46:23]
  wire  cout_7 = a_and_b7 | a_xor_b7 & cin_7; // @[CSA.scala 47:24]
  wire [1:0] temp_7 = {cout_7,sum_7}; // @[Cat.scala 31:58]
  wire  a_8 = io_in_0[8]; // @[CSA.scala 43:32]
  wire  b_8 = io_in_1[8]; // @[CSA.scala 43:45]
  wire  cin_8 = io_in_2[8]; // @[CSA.scala 43:58]
  wire  a_xor_b8 = a_8 ^ b_8; // @[CSA.scala 44:21]
  wire  a_and_b8 = a_8 & b_8; // @[CSA.scala 45:21]
  wire  sum_8 = a_xor_b8 ^ cin_8; // @[CSA.scala 46:23]
  wire  cout_8 = a_and_b8 | a_xor_b8 & cin_8; // @[CSA.scala 47:24]
  wire [1:0] temp_8 = {cout_8,sum_8}; // @[Cat.scala 31:58]
  wire  a_9 = io_in_0[9]; // @[CSA.scala 43:32]
  wire  b_9 = io_in_1[9]; // @[CSA.scala 43:45]
  wire  cin_9 = io_in_2[9]; // @[CSA.scala 43:58]
  wire  a_xor_b9 = a_9 ^ b_9; // @[CSA.scala 44:21]
  wire  a_and_b9 = a_9 & b_9; // @[CSA.scala 45:21]
  wire  sum_9 = a_xor_b9 ^ cin_9; // @[CSA.scala 46:23]
  wire  cout_9 = a_and_b9 | a_xor_b9 & cin_9; // @[CSA.scala 47:24]
  wire [1:0] temp_9 = {cout_9,sum_9}; // @[Cat.scala 31:58]
  wire [4:0] io_out_0_lo = {temp_4[0],temp_3[0],temp_2[0],temp_1[0],temp_0[0]}; // @[Cat.scala 31:58]
  wire [4:0] io_out_0_hi = {temp_9[0],temp_8[0],temp_7[0],temp_6[0],temp_5[0]}; // @[Cat.scala 31:58]
  wire [4:0] io_out_1_lo = {temp_4[1],temp_3[1],temp_2[1],temp_1[1],temp_0[1]}; // @[Cat.scala 31:58]
  wire [4:0] io_out_1_hi = {temp_9[1],temp_8[1],temp_7[1],temp_6[1],temp_5[1]}; // @[Cat.scala 31:58]
  assign io_out_0 = {io_out_0_hi,io_out_0_lo}; // @[Cat.scala 31:58]
  assign io_out_1 = {io_out_1_hi,io_out_1_lo}; // @[Cat.scala 31:58]
endmodule

