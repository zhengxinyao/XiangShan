module DelayN_44(
  input   io_in,
  output  io_out
);
  assign io_out = io_in; // @[Hold.scala 92:10]
endmodule

