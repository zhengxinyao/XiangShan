module VlflowQueue(
  input         clock,
  input         reset,
  input         io_loadRegIn_0_valid,
  input  [4:0]  io_loadRegIn_0_bits_uop_robIdx_value,
  input  [38:0] io_loadRegIn_0_bits_baseaddr,
  input         io_loadRegIn_1_valid,
  input  [4:0]  io_loadRegIn_1_bits_uop_robIdx_value,
  input  [38:0] io_loadRegIn_1_bits_baseaddr,
  input         io_loadPipeOut_0_ready,
  output        io_loadPipeOut_0_valid,
  output [38:0] io_loadPipeOut_0_bits_vaddr,
  input         io_loadPipeOut_1_ready,
  output        io_loadPipeOut_1_valid,
  output [38:0] io_loadPipeOut_1_bits_vaddr
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [63:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [63:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [63:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [63:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [63:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [63:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [63:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [63:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [63:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [63:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [63:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [63:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [63:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [63:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [63:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [63:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [63:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [63:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [63:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [63:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [63:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [63:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [63:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [63:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [63:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [63:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [63:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [63:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [63:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [63:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [63:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [63:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [63:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [63:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [63:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [63:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [63:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [63:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [63:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [63:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [63:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [63:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [63:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [63:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [63:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [63:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
`endif // RANDOMIZE_REG_INIT
  reg [4:0] flow_entry_0_0_uop_robIdx_value; // @[Vlflowqueue.scala 134:29]
  reg [38:0] flow_entry_0_0_vaddr; // @[Vlflowqueue.scala 134:29]
  reg [4:0] flow_entry_0_1_uop_robIdx_value; // @[Vlflowqueue.scala 134:29]
  reg [38:0] flow_entry_0_1_vaddr; // @[Vlflowqueue.scala 134:29]
  reg [4:0] flow_entry_0_2_uop_robIdx_value; // @[Vlflowqueue.scala 134:29]
  reg [38:0] flow_entry_0_2_vaddr; // @[Vlflowqueue.scala 134:29]
  reg [4:0] flow_entry_0_3_uop_robIdx_value; // @[Vlflowqueue.scala 134:29]
  reg [38:0] flow_entry_0_3_vaddr; // @[Vlflowqueue.scala 134:29]
  reg [4:0] flow_entry_0_4_uop_robIdx_value; // @[Vlflowqueue.scala 134:29]
  reg [38:0] flow_entry_0_4_vaddr; // @[Vlflowqueue.scala 134:29]
  reg [4:0] flow_entry_0_5_uop_robIdx_value; // @[Vlflowqueue.scala 134:29]
  reg [38:0] flow_entry_0_5_vaddr; // @[Vlflowqueue.scala 134:29]
  reg [4:0] flow_entry_0_6_uop_robIdx_value; // @[Vlflowqueue.scala 134:29]
  reg [38:0] flow_entry_0_6_vaddr; // @[Vlflowqueue.scala 134:29]
  reg [4:0] flow_entry_0_7_uop_robIdx_value; // @[Vlflowqueue.scala 134:29]
  reg [38:0] flow_entry_0_7_vaddr; // @[Vlflowqueue.scala 134:29]
  reg [4:0] flow_entry_0_8_uop_robIdx_value; // @[Vlflowqueue.scala 134:29]
  reg [38:0] flow_entry_0_8_vaddr; // @[Vlflowqueue.scala 134:29]
  reg [4:0] flow_entry_0_9_uop_robIdx_value; // @[Vlflowqueue.scala 134:29]
  reg [38:0] flow_entry_0_9_vaddr; // @[Vlflowqueue.scala 134:29]
  reg [4:0] flow_entry_0_10_uop_robIdx_value; // @[Vlflowqueue.scala 134:29]
  reg [38:0] flow_entry_0_10_vaddr; // @[Vlflowqueue.scala 134:29]
  reg [4:0] flow_entry_0_11_uop_robIdx_value; // @[Vlflowqueue.scala 134:29]
  reg [38:0] flow_entry_0_11_vaddr; // @[Vlflowqueue.scala 134:29]
  reg [4:0] flow_entry_0_12_uop_robIdx_value; // @[Vlflowqueue.scala 134:29]
  reg [38:0] flow_entry_0_12_vaddr; // @[Vlflowqueue.scala 134:29]
  reg [4:0] flow_entry_0_13_uop_robIdx_value; // @[Vlflowqueue.scala 134:29]
  reg [38:0] flow_entry_0_13_vaddr; // @[Vlflowqueue.scala 134:29]
  reg [4:0] flow_entry_0_14_uop_robIdx_value; // @[Vlflowqueue.scala 134:29]
  reg [38:0] flow_entry_0_14_vaddr; // @[Vlflowqueue.scala 134:29]
  reg [4:0] flow_entry_0_15_uop_robIdx_value; // @[Vlflowqueue.scala 134:29]
  reg [38:0] flow_entry_0_15_vaddr; // @[Vlflowqueue.scala 134:29]
  reg [4:0] flow_entry_0_16_uop_robIdx_value; // @[Vlflowqueue.scala 134:29]
  reg [38:0] flow_entry_0_16_vaddr; // @[Vlflowqueue.scala 134:29]
  reg [4:0] flow_entry_0_17_uop_robIdx_value; // @[Vlflowqueue.scala 134:29]
  reg [38:0] flow_entry_0_17_vaddr; // @[Vlflowqueue.scala 134:29]
  reg [4:0] flow_entry_0_18_uop_robIdx_value; // @[Vlflowqueue.scala 134:29]
  reg [38:0] flow_entry_0_18_vaddr; // @[Vlflowqueue.scala 134:29]
  reg [4:0] flow_entry_0_19_uop_robIdx_value; // @[Vlflowqueue.scala 134:29]
  reg [38:0] flow_entry_0_19_vaddr; // @[Vlflowqueue.scala 134:29]
  reg [4:0] flow_entry_0_20_uop_robIdx_value; // @[Vlflowqueue.scala 134:29]
  reg [38:0] flow_entry_0_20_vaddr; // @[Vlflowqueue.scala 134:29]
  reg [4:0] flow_entry_0_21_uop_robIdx_value; // @[Vlflowqueue.scala 134:29]
  reg [38:0] flow_entry_0_21_vaddr; // @[Vlflowqueue.scala 134:29]
  reg [4:0] flow_entry_0_22_uop_robIdx_value; // @[Vlflowqueue.scala 134:29]
  reg [38:0] flow_entry_0_22_vaddr; // @[Vlflowqueue.scala 134:29]
  reg [4:0] flow_entry_0_23_uop_robIdx_value; // @[Vlflowqueue.scala 134:29]
  reg [38:0] flow_entry_0_23_vaddr; // @[Vlflowqueue.scala 134:29]
  reg [4:0] flow_entry_0_24_uop_robIdx_value; // @[Vlflowqueue.scala 134:29]
  reg [38:0] flow_entry_0_24_vaddr; // @[Vlflowqueue.scala 134:29]
  reg [4:0] flow_entry_0_25_uop_robIdx_value; // @[Vlflowqueue.scala 134:29]
  reg [38:0] flow_entry_0_25_vaddr; // @[Vlflowqueue.scala 134:29]
  reg [4:0] flow_entry_0_26_uop_robIdx_value; // @[Vlflowqueue.scala 134:29]
  reg [38:0] flow_entry_0_26_vaddr; // @[Vlflowqueue.scala 134:29]
  reg [4:0] flow_entry_0_27_uop_robIdx_value; // @[Vlflowqueue.scala 134:29]
  reg [38:0] flow_entry_0_27_vaddr; // @[Vlflowqueue.scala 134:29]
  reg [4:0] flow_entry_0_28_uop_robIdx_value; // @[Vlflowqueue.scala 134:29]
  reg [38:0] flow_entry_0_28_vaddr; // @[Vlflowqueue.scala 134:29]
  reg [4:0] flow_entry_0_29_uop_robIdx_value; // @[Vlflowqueue.scala 134:29]
  reg [38:0] flow_entry_0_29_vaddr; // @[Vlflowqueue.scala 134:29]
  reg [4:0] flow_entry_0_30_uop_robIdx_value; // @[Vlflowqueue.scala 134:29]
  reg [38:0] flow_entry_0_30_vaddr; // @[Vlflowqueue.scala 134:29]
  reg [4:0] flow_entry_0_31_uop_robIdx_value; // @[Vlflowqueue.scala 134:29]
  reg [38:0] flow_entry_0_31_vaddr; // @[Vlflowqueue.scala 134:29]
  reg [4:0] flow_entry_1_0_uop_robIdx_value; // @[Vlflowqueue.scala 134:29]
  reg [38:0] flow_entry_1_0_vaddr; // @[Vlflowqueue.scala 134:29]
  reg [4:0] flow_entry_1_1_uop_robIdx_value; // @[Vlflowqueue.scala 134:29]
  reg [38:0] flow_entry_1_1_vaddr; // @[Vlflowqueue.scala 134:29]
  reg [4:0] flow_entry_1_2_uop_robIdx_value; // @[Vlflowqueue.scala 134:29]
  reg [38:0] flow_entry_1_2_vaddr; // @[Vlflowqueue.scala 134:29]
  reg [4:0] flow_entry_1_3_uop_robIdx_value; // @[Vlflowqueue.scala 134:29]
  reg [38:0] flow_entry_1_3_vaddr; // @[Vlflowqueue.scala 134:29]
  reg [4:0] flow_entry_1_4_uop_robIdx_value; // @[Vlflowqueue.scala 134:29]
  reg [38:0] flow_entry_1_4_vaddr; // @[Vlflowqueue.scala 134:29]
  reg [4:0] flow_entry_1_5_uop_robIdx_value; // @[Vlflowqueue.scala 134:29]
  reg [38:0] flow_entry_1_5_vaddr; // @[Vlflowqueue.scala 134:29]
  reg [4:0] flow_entry_1_6_uop_robIdx_value; // @[Vlflowqueue.scala 134:29]
  reg [38:0] flow_entry_1_6_vaddr; // @[Vlflowqueue.scala 134:29]
  reg [4:0] flow_entry_1_7_uop_robIdx_value; // @[Vlflowqueue.scala 134:29]
  reg [38:0] flow_entry_1_7_vaddr; // @[Vlflowqueue.scala 134:29]
  reg [4:0] flow_entry_1_8_uop_robIdx_value; // @[Vlflowqueue.scala 134:29]
  reg [38:0] flow_entry_1_8_vaddr; // @[Vlflowqueue.scala 134:29]
  reg [4:0] flow_entry_1_9_uop_robIdx_value; // @[Vlflowqueue.scala 134:29]
  reg [38:0] flow_entry_1_9_vaddr; // @[Vlflowqueue.scala 134:29]
  reg [4:0] flow_entry_1_10_uop_robIdx_value; // @[Vlflowqueue.scala 134:29]
  reg [38:0] flow_entry_1_10_vaddr; // @[Vlflowqueue.scala 134:29]
  reg [4:0] flow_entry_1_11_uop_robIdx_value; // @[Vlflowqueue.scala 134:29]
  reg [38:0] flow_entry_1_11_vaddr; // @[Vlflowqueue.scala 134:29]
  reg [4:0] flow_entry_1_12_uop_robIdx_value; // @[Vlflowqueue.scala 134:29]
  reg [38:0] flow_entry_1_12_vaddr; // @[Vlflowqueue.scala 134:29]
  reg [4:0] flow_entry_1_13_uop_robIdx_value; // @[Vlflowqueue.scala 134:29]
  reg [38:0] flow_entry_1_13_vaddr; // @[Vlflowqueue.scala 134:29]
  reg [4:0] flow_entry_1_14_uop_robIdx_value; // @[Vlflowqueue.scala 134:29]
  reg [38:0] flow_entry_1_14_vaddr; // @[Vlflowqueue.scala 134:29]
  reg [4:0] flow_entry_1_15_uop_robIdx_value; // @[Vlflowqueue.scala 134:29]
  reg [38:0] flow_entry_1_15_vaddr; // @[Vlflowqueue.scala 134:29]
  reg [4:0] flow_entry_1_16_uop_robIdx_value; // @[Vlflowqueue.scala 134:29]
  reg [38:0] flow_entry_1_16_vaddr; // @[Vlflowqueue.scala 134:29]
  reg [4:0] flow_entry_1_17_uop_robIdx_value; // @[Vlflowqueue.scala 134:29]
  reg [38:0] flow_entry_1_17_vaddr; // @[Vlflowqueue.scala 134:29]
  reg [4:0] flow_entry_1_18_uop_robIdx_value; // @[Vlflowqueue.scala 134:29]
  reg [38:0] flow_entry_1_18_vaddr; // @[Vlflowqueue.scala 134:29]
  reg [4:0] flow_entry_1_19_uop_robIdx_value; // @[Vlflowqueue.scala 134:29]
  reg [38:0] flow_entry_1_19_vaddr; // @[Vlflowqueue.scala 134:29]
  reg [4:0] flow_entry_1_20_uop_robIdx_value; // @[Vlflowqueue.scala 134:29]
  reg [38:0] flow_entry_1_20_vaddr; // @[Vlflowqueue.scala 134:29]
  reg [4:0] flow_entry_1_21_uop_robIdx_value; // @[Vlflowqueue.scala 134:29]
  reg [38:0] flow_entry_1_21_vaddr; // @[Vlflowqueue.scala 134:29]
  reg [4:0] flow_entry_1_22_uop_robIdx_value; // @[Vlflowqueue.scala 134:29]
  reg [38:0] flow_entry_1_22_vaddr; // @[Vlflowqueue.scala 134:29]
  reg [4:0] flow_entry_1_23_uop_robIdx_value; // @[Vlflowqueue.scala 134:29]
  reg [38:0] flow_entry_1_23_vaddr; // @[Vlflowqueue.scala 134:29]
  reg [4:0] flow_entry_1_24_uop_robIdx_value; // @[Vlflowqueue.scala 134:29]
  reg [38:0] flow_entry_1_24_vaddr; // @[Vlflowqueue.scala 134:29]
  reg [4:0] flow_entry_1_25_uop_robIdx_value; // @[Vlflowqueue.scala 134:29]
  reg [38:0] flow_entry_1_25_vaddr; // @[Vlflowqueue.scala 134:29]
  reg [4:0] flow_entry_1_26_uop_robIdx_value; // @[Vlflowqueue.scala 134:29]
  reg [38:0] flow_entry_1_26_vaddr; // @[Vlflowqueue.scala 134:29]
  reg [4:0] flow_entry_1_27_uop_robIdx_value; // @[Vlflowqueue.scala 134:29]
  reg [38:0] flow_entry_1_27_vaddr; // @[Vlflowqueue.scala 134:29]
  reg [4:0] flow_entry_1_28_uop_robIdx_value; // @[Vlflowqueue.scala 134:29]
  reg [38:0] flow_entry_1_28_vaddr; // @[Vlflowqueue.scala 134:29]
  reg [4:0] flow_entry_1_29_uop_robIdx_value; // @[Vlflowqueue.scala 134:29]
  reg [38:0] flow_entry_1_29_vaddr; // @[Vlflowqueue.scala 134:29]
  reg [4:0] flow_entry_1_30_uop_robIdx_value; // @[Vlflowqueue.scala 134:29]
  reg [38:0] flow_entry_1_30_vaddr; // @[Vlflowqueue.scala 134:29]
  reg [4:0] flow_entry_1_31_uop_robIdx_value; // @[Vlflowqueue.scala 134:29]
  reg [38:0] flow_entry_1_31_vaddr; // @[Vlflowqueue.scala 134:29]
  reg  flow_entry_valid_0_0; // @[Vlflowqueue.scala 135:33]
  reg  flow_entry_valid_0_1; // @[Vlflowqueue.scala 135:33]
  reg  flow_entry_valid_0_2; // @[Vlflowqueue.scala 135:33]
  reg  flow_entry_valid_0_3; // @[Vlflowqueue.scala 135:33]
  reg  flow_entry_valid_0_4; // @[Vlflowqueue.scala 135:33]
  reg  flow_entry_valid_0_5; // @[Vlflowqueue.scala 135:33]
  reg  flow_entry_valid_0_6; // @[Vlflowqueue.scala 135:33]
  reg  flow_entry_valid_0_7; // @[Vlflowqueue.scala 135:33]
  reg  flow_entry_valid_0_8; // @[Vlflowqueue.scala 135:33]
  reg  flow_entry_valid_0_9; // @[Vlflowqueue.scala 135:33]
  reg  flow_entry_valid_0_10; // @[Vlflowqueue.scala 135:33]
  reg  flow_entry_valid_0_11; // @[Vlflowqueue.scala 135:33]
  reg  flow_entry_valid_0_12; // @[Vlflowqueue.scala 135:33]
  reg  flow_entry_valid_0_13; // @[Vlflowqueue.scala 135:33]
  reg  flow_entry_valid_0_14; // @[Vlflowqueue.scala 135:33]
  reg  flow_entry_valid_0_15; // @[Vlflowqueue.scala 135:33]
  reg  flow_entry_valid_0_16; // @[Vlflowqueue.scala 135:33]
  reg  flow_entry_valid_0_17; // @[Vlflowqueue.scala 135:33]
  reg  flow_entry_valid_0_18; // @[Vlflowqueue.scala 135:33]
  reg  flow_entry_valid_0_19; // @[Vlflowqueue.scala 135:33]
  reg  flow_entry_valid_0_20; // @[Vlflowqueue.scala 135:33]
  reg  flow_entry_valid_0_21; // @[Vlflowqueue.scala 135:33]
  reg  flow_entry_valid_0_22; // @[Vlflowqueue.scala 135:33]
  reg  flow_entry_valid_0_23; // @[Vlflowqueue.scala 135:33]
  reg  flow_entry_valid_0_24; // @[Vlflowqueue.scala 135:33]
  reg  flow_entry_valid_0_25; // @[Vlflowqueue.scala 135:33]
  reg  flow_entry_valid_0_26; // @[Vlflowqueue.scala 135:33]
  reg  flow_entry_valid_0_27; // @[Vlflowqueue.scala 135:33]
  reg  flow_entry_valid_0_28; // @[Vlflowqueue.scala 135:33]
  reg  flow_entry_valid_0_29; // @[Vlflowqueue.scala 135:33]
  reg  flow_entry_valid_0_30; // @[Vlflowqueue.scala 135:33]
  reg  flow_entry_valid_0_31; // @[Vlflowqueue.scala 135:33]
  reg  flow_entry_valid_1_0; // @[Vlflowqueue.scala 135:33]
  reg  flow_entry_valid_1_1; // @[Vlflowqueue.scala 135:33]
  reg  flow_entry_valid_1_2; // @[Vlflowqueue.scala 135:33]
  reg  flow_entry_valid_1_3; // @[Vlflowqueue.scala 135:33]
  reg  flow_entry_valid_1_4; // @[Vlflowqueue.scala 135:33]
  reg  flow_entry_valid_1_5; // @[Vlflowqueue.scala 135:33]
  reg  flow_entry_valid_1_6; // @[Vlflowqueue.scala 135:33]
  reg  flow_entry_valid_1_7; // @[Vlflowqueue.scala 135:33]
  reg  flow_entry_valid_1_8; // @[Vlflowqueue.scala 135:33]
  reg  flow_entry_valid_1_9; // @[Vlflowqueue.scala 135:33]
  reg  flow_entry_valid_1_10; // @[Vlflowqueue.scala 135:33]
  reg  flow_entry_valid_1_11; // @[Vlflowqueue.scala 135:33]
  reg  flow_entry_valid_1_12; // @[Vlflowqueue.scala 135:33]
  reg  flow_entry_valid_1_13; // @[Vlflowqueue.scala 135:33]
  reg  flow_entry_valid_1_14; // @[Vlflowqueue.scala 135:33]
  reg  flow_entry_valid_1_15; // @[Vlflowqueue.scala 135:33]
  reg  flow_entry_valid_1_16; // @[Vlflowqueue.scala 135:33]
  reg  flow_entry_valid_1_17; // @[Vlflowqueue.scala 135:33]
  reg  flow_entry_valid_1_18; // @[Vlflowqueue.scala 135:33]
  reg  flow_entry_valid_1_19; // @[Vlflowqueue.scala 135:33]
  reg  flow_entry_valid_1_20; // @[Vlflowqueue.scala 135:33]
  reg  flow_entry_valid_1_21; // @[Vlflowqueue.scala 135:33]
  reg  flow_entry_valid_1_22; // @[Vlflowqueue.scala 135:33]
  reg  flow_entry_valid_1_23; // @[Vlflowqueue.scala 135:33]
  reg  flow_entry_valid_1_24; // @[Vlflowqueue.scala 135:33]
  reg  flow_entry_valid_1_25; // @[Vlflowqueue.scala 135:33]
  reg  flow_entry_valid_1_26; // @[Vlflowqueue.scala 135:33]
  reg  flow_entry_valid_1_27; // @[Vlflowqueue.scala 135:33]
  reg  flow_entry_valid_1_28; // @[Vlflowqueue.scala 135:33]
  reg  flow_entry_valid_1_29; // @[Vlflowqueue.scala 135:33]
  reg  flow_entry_valid_1_30; // @[Vlflowqueue.scala 135:33]
  reg  flow_entry_valid_1_31; // @[Vlflowqueue.scala 135:33]
  wire  _needAlloc_0_T_15 = flow_entry_0_15_uop_robIdx_value == io_loadRegIn_0_bits_uop_robIdx_value; // @[Vlflowqueue.scala 161:65]
  wire  _needAlloc_0_T_46 = flow_entry_0_0_uop_robIdx_value == io_loadRegIn_0_bits_uop_robIdx_value |
    flow_entry_0_1_uop_robIdx_value == io_loadRegIn_0_bits_uop_robIdx_value | flow_entry_0_2_uop_robIdx_value ==
    io_loadRegIn_0_bits_uop_robIdx_value | flow_entry_0_3_uop_robIdx_value == io_loadRegIn_0_bits_uop_robIdx_value |
    flow_entry_0_4_uop_robIdx_value == io_loadRegIn_0_bits_uop_robIdx_value | flow_entry_0_5_uop_robIdx_value ==
    io_loadRegIn_0_bits_uop_robIdx_value | flow_entry_0_6_uop_robIdx_value == io_loadRegIn_0_bits_uop_robIdx_value |
    flow_entry_0_7_uop_robIdx_value == io_loadRegIn_0_bits_uop_robIdx_value | flow_entry_0_8_uop_robIdx_value ==
    io_loadRegIn_0_bits_uop_robIdx_value | flow_entry_0_9_uop_robIdx_value == io_loadRegIn_0_bits_uop_robIdx_value |
    flow_entry_0_10_uop_robIdx_value == io_loadRegIn_0_bits_uop_robIdx_value | flow_entry_0_11_uop_robIdx_value ==
    io_loadRegIn_0_bits_uop_robIdx_value | flow_entry_0_12_uop_robIdx_value == io_loadRegIn_0_bits_uop_robIdx_value |
    flow_entry_0_13_uop_robIdx_value == io_loadRegIn_0_bits_uop_robIdx_value | flow_entry_0_14_uop_robIdx_value ==
    io_loadRegIn_0_bits_uop_robIdx_value | _needAlloc_0_T_15; // @[Vlflowqueue.scala 161:117]
  wire  _needAlloc_0_T_61 = _needAlloc_0_T_46 | flow_entry_0_16_uop_robIdx_value == io_loadRegIn_0_bits_uop_robIdx_value
     | flow_entry_0_17_uop_robIdx_value == io_loadRegIn_0_bits_uop_robIdx_value | flow_entry_0_18_uop_robIdx_value ==
    io_loadRegIn_0_bits_uop_robIdx_value | flow_entry_0_19_uop_robIdx_value == io_loadRegIn_0_bits_uop_robIdx_value |
    flow_entry_0_20_uop_robIdx_value == io_loadRegIn_0_bits_uop_robIdx_value | flow_entry_0_21_uop_robIdx_value ==
    io_loadRegIn_0_bits_uop_robIdx_value | flow_entry_0_22_uop_robIdx_value == io_loadRegIn_0_bits_uop_robIdx_value |
    flow_entry_0_23_uop_robIdx_value == io_loadRegIn_0_bits_uop_robIdx_value | flow_entry_0_24_uop_robIdx_value ==
    io_loadRegIn_0_bits_uop_robIdx_value | flow_entry_0_25_uop_robIdx_value == io_loadRegIn_0_bits_uop_robIdx_value |
    flow_entry_0_26_uop_robIdx_value == io_loadRegIn_0_bits_uop_robIdx_value | flow_entry_0_27_uop_robIdx_value ==
    io_loadRegIn_0_bits_uop_robIdx_value | flow_entry_0_28_uop_robIdx_value == io_loadRegIn_0_bits_uop_robIdx_value |
    flow_entry_0_29_uop_robIdx_value == io_loadRegIn_0_bits_uop_robIdx_value | flow_entry_0_30_uop_robIdx_value ==
    io_loadRegIn_0_bits_uop_robIdx_value; // @[Vlflowqueue.scala 161:117]
  wire  _needAlloc_0_T_78 = flow_entry_1_15_uop_robIdx_value == io_loadRegIn_0_bits_uop_robIdx_value; // @[Vlflowqueue.scala 161:65]
  wire  _needAlloc_0_T_109 = flow_entry_1_0_uop_robIdx_value == io_loadRegIn_0_bits_uop_robIdx_value |
    flow_entry_1_1_uop_robIdx_value == io_loadRegIn_0_bits_uop_robIdx_value | flow_entry_1_2_uop_robIdx_value ==
    io_loadRegIn_0_bits_uop_robIdx_value | flow_entry_1_3_uop_robIdx_value == io_loadRegIn_0_bits_uop_robIdx_value |
    flow_entry_1_4_uop_robIdx_value == io_loadRegIn_0_bits_uop_robIdx_value | flow_entry_1_5_uop_robIdx_value ==
    io_loadRegIn_0_bits_uop_robIdx_value | flow_entry_1_6_uop_robIdx_value == io_loadRegIn_0_bits_uop_robIdx_value |
    flow_entry_1_7_uop_robIdx_value == io_loadRegIn_0_bits_uop_robIdx_value | flow_entry_1_8_uop_robIdx_value ==
    io_loadRegIn_0_bits_uop_robIdx_value | flow_entry_1_9_uop_robIdx_value == io_loadRegIn_0_bits_uop_robIdx_value |
    flow_entry_1_10_uop_robIdx_value == io_loadRegIn_0_bits_uop_robIdx_value | flow_entry_1_11_uop_robIdx_value ==
    io_loadRegIn_0_bits_uop_robIdx_value | flow_entry_1_12_uop_robIdx_value == io_loadRegIn_0_bits_uop_robIdx_value |
    flow_entry_1_13_uop_robIdx_value == io_loadRegIn_0_bits_uop_robIdx_value | flow_entry_1_14_uop_robIdx_value ==
    io_loadRegIn_0_bits_uop_robIdx_value | _needAlloc_0_T_78; // @[Vlflowqueue.scala 161:117]
  wire  _needAlloc_0_T_124 = _needAlloc_0_T_109 | flow_entry_1_16_uop_robIdx_value ==
    io_loadRegIn_0_bits_uop_robIdx_value | flow_entry_1_17_uop_robIdx_value == io_loadRegIn_0_bits_uop_robIdx_value |
    flow_entry_1_18_uop_robIdx_value == io_loadRegIn_0_bits_uop_robIdx_value | flow_entry_1_19_uop_robIdx_value ==
    io_loadRegIn_0_bits_uop_robIdx_value | flow_entry_1_20_uop_robIdx_value == io_loadRegIn_0_bits_uop_robIdx_value |
    flow_entry_1_21_uop_robIdx_value == io_loadRegIn_0_bits_uop_robIdx_value | flow_entry_1_22_uop_robIdx_value ==
    io_loadRegIn_0_bits_uop_robIdx_value | flow_entry_1_23_uop_robIdx_value == io_loadRegIn_0_bits_uop_robIdx_value |
    flow_entry_1_24_uop_robIdx_value == io_loadRegIn_0_bits_uop_robIdx_value | flow_entry_1_25_uop_robIdx_value ==
    io_loadRegIn_0_bits_uop_robIdx_value | flow_entry_1_26_uop_robIdx_value == io_loadRegIn_0_bits_uop_robIdx_value |
    flow_entry_1_27_uop_robIdx_value == io_loadRegIn_0_bits_uop_robIdx_value | flow_entry_1_28_uop_robIdx_value ==
    io_loadRegIn_0_bits_uop_robIdx_value | flow_entry_1_29_uop_robIdx_value == io_loadRegIn_0_bits_uop_robIdx_value |
    flow_entry_1_30_uop_robIdx_value == io_loadRegIn_0_bits_uop_robIdx_value; // @[Vlflowqueue.scala 161:117]
  wire  needAlloc_0 = ~(_needAlloc_0_T_61 | flow_entry_0_31_uop_robIdx_value == io_loadRegIn_0_bits_uop_robIdx_value | (
    _needAlloc_0_T_124 | flow_entry_1_31_uop_robIdx_value == io_loadRegIn_0_bits_uop_robIdx_value)) &
    io_loadRegIn_0_valid; // @[Vlflowqueue.scala 161:139]
  wire [4:0] _vend_0_0_T_2 = {{1'd0}, io_loadRegIn_0_bits_baseaddr[3:0]}; // @[Vlflowqueue.scala 164:41]
  wire [5:0] _vend_1_0_T_2 = {{1'd0}, io_loadRegIn_0_bits_baseaddr[4:0]}; // @[Vlflowqueue.scala 165:41]
  wire [6:0] _vend_2_0_T_2 = {{1'd0}, io_loadRegIn_0_bits_baseaddr[5:0]}; // @[Vlflowqueue.scala 166:41]
  wire [7:0] _vend_3_0_T_2 = {{1'd0}, io_loadRegIn_0_bits_baseaddr[6:0]}; // @[Vlflowqueue.scala 167:41]
  wire [7:0] vend_3_0 = {{1'd0}, _vend_3_0_T_2[6:0]}; // @[Vlflowqueue.scala 144:29 167:21]
  wire [6:0] vend_2_0 = {{1'd0}, _vend_2_0_T_2[5:0]}; // @[Vlflowqueue.scala 143:29 166:21]
  wire [5:0] vend_1_0 = {{1'd0}, _vend_1_0_T_2[4:0]}; // @[Vlflowqueue.scala 142:29 165:21]
  wire [4:0] vend_0_0 = {{1'd0}, _vend_0_0_T_2[3:0]}; // @[Vlflowqueue.scala 141:29 164:21]
  wire [1:0] _flowWriteNumber_0_T_10 = vend_1_0[5] ? vend_1_0[5:4] : {{1'd0}, vend_0_0[4]}; // @[Vlflowqueue.scala 168:114]
  wire [2:0] _flowWriteNumber_0_T_11 = vend_2_0[6] ? vend_2_0[6:4] : {{1'd0}, _flowWriteNumber_0_T_10}; // @[Vlflowqueue.scala 168:72]
  wire [3:0] _flowWriteNumber_0_T_12 = vend_3_0[7] ? vend_3_0[7:4] : {{1'd0}, _flowWriteNumber_0_T_11}; // @[Vlflowqueue.scala 168:30]
  wire  _needAlloc_1_T_15 = flow_entry_0_15_uop_robIdx_value == io_loadRegIn_1_bits_uop_robIdx_value; // @[Vlflowqueue.scala 161:65]
  wire  _needAlloc_1_T_46 = flow_entry_0_0_uop_robIdx_value == io_loadRegIn_1_bits_uop_robIdx_value |
    flow_entry_0_1_uop_robIdx_value == io_loadRegIn_1_bits_uop_robIdx_value | flow_entry_0_2_uop_robIdx_value ==
    io_loadRegIn_1_bits_uop_robIdx_value | flow_entry_0_3_uop_robIdx_value == io_loadRegIn_1_bits_uop_robIdx_value |
    flow_entry_0_4_uop_robIdx_value == io_loadRegIn_1_bits_uop_robIdx_value | flow_entry_0_5_uop_robIdx_value ==
    io_loadRegIn_1_bits_uop_robIdx_value | flow_entry_0_6_uop_robIdx_value == io_loadRegIn_1_bits_uop_robIdx_value |
    flow_entry_0_7_uop_robIdx_value == io_loadRegIn_1_bits_uop_robIdx_value | flow_entry_0_8_uop_robIdx_value ==
    io_loadRegIn_1_bits_uop_robIdx_value | flow_entry_0_9_uop_robIdx_value == io_loadRegIn_1_bits_uop_robIdx_value |
    flow_entry_0_10_uop_robIdx_value == io_loadRegIn_1_bits_uop_robIdx_value | flow_entry_0_11_uop_robIdx_value ==
    io_loadRegIn_1_bits_uop_robIdx_value | flow_entry_0_12_uop_robIdx_value == io_loadRegIn_1_bits_uop_robIdx_value |
    flow_entry_0_13_uop_robIdx_value == io_loadRegIn_1_bits_uop_robIdx_value | flow_entry_0_14_uop_robIdx_value ==
    io_loadRegIn_1_bits_uop_robIdx_value | _needAlloc_1_T_15; // @[Vlflowqueue.scala 161:117]
  wire  _needAlloc_1_T_61 = _needAlloc_1_T_46 | flow_entry_0_16_uop_robIdx_value == io_loadRegIn_1_bits_uop_robIdx_value
     | flow_entry_0_17_uop_robIdx_value == io_loadRegIn_1_bits_uop_robIdx_value | flow_entry_0_18_uop_robIdx_value ==
    io_loadRegIn_1_bits_uop_robIdx_value | flow_entry_0_19_uop_robIdx_value == io_loadRegIn_1_bits_uop_robIdx_value |
    flow_entry_0_20_uop_robIdx_value == io_loadRegIn_1_bits_uop_robIdx_value | flow_entry_0_21_uop_robIdx_value ==
    io_loadRegIn_1_bits_uop_robIdx_value | flow_entry_0_22_uop_robIdx_value == io_loadRegIn_1_bits_uop_robIdx_value |
    flow_entry_0_23_uop_robIdx_value == io_loadRegIn_1_bits_uop_robIdx_value | flow_entry_0_24_uop_robIdx_value ==
    io_loadRegIn_1_bits_uop_robIdx_value | flow_entry_0_25_uop_robIdx_value == io_loadRegIn_1_bits_uop_robIdx_value |
    flow_entry_0_26_uop_robIdx_value == io_loadRegIn_1_bits_uop_robIdx_value | flow_entry_0_27_uop_robIdx_value ==
    io_loadRegIn_1_bits_uop_robIdx_value | flow_entry_0_28_uop_robIdx_value == io_loadRegIn_1_bits_uop_robIdx_value |
    flow_entry_0_29_uop_robIdx_value == io_loadRegIn_1_bits_uop_robIdx_value | flow_entry_0_30_uop_robIdx_value ==
    io_loadRegIn_1_bits_uop_robIdx_value; // @[Vlflowqueue.scala 161:117]
  wire  _needAlloc_1_T_78 = flow_entry_1_15_uop_robIdx_value == io_loadRegIn_1_bits_uop_robIdx_value; // @[Vlflowqueue.scala 161:65]
  wire  _needAlloc_1_T_109 = flow_entry_1_0_uop_robIdx_value == io_loadRegIn_1_bits_uop_robIdx_value |
    flow_entry_1_1_uop_robIdx_value == io_loadRegIn_1_bits_uop_robIdx_value | flow_entry_1_2_uop_robIdx_value ==
    io_loadRegIn_1_bits_uop_robIdx_value | flow_entry_1_3_uop_robIdx_value == io_loadRegIn_1_bits_uop_robIdx_value |
    flow_entry_1_4_uop_robIdx_value == io_loadRegIn_1_bits_uop_robIdx_value | flow_entry_1_5_uop_robIdx_value ==
    io_loadRegIn_1_bits_uop_robIdx_value | flow_entry_1_6_uop_robIdx_value == io_loadRegIn_1_bits_uop_robIdx_value |
    flow_entry_1_7_uop_robIdx_value == io_loadRegIn_1_bits_uop_robIdx_value | flow_entry_1_8_uop_robIdx_value ==
    io_loadRegIn_1_bits_uop_robIdx_value | flow_entry_1_9_uop_robIdx_value == io_loadRegIn_1_bits_uop_robIdx_value |
    flow_entry_1_10_uop_robIdx_value == io_loadRegIn_1_bits_uop_robIdx_value | flow_entry_1_11_uop_robIdx_value ==
    io_loadRegIn_1_bits_uop_robIdx_value | flow_entry_1_12_uop_robIdx_value == io_loadRegIn_1_bits_uop_robIdx_value |
    flow_entry_1_13_uop_robIdx_value == io_loadRegIn_1_bits_uop_robIdx_value | flow_entry_1_14_uop_robIdx_value ==
    io_loadRegIn_1_bits_uop_robIdx_value | _needAlloc_1_T_78; // @[Vlflowqueue.scala 161:117]
  wire  _needAlloc_1_T_124 = _needAlloc_1_T_109 | flow_entry_1_16_uop_robIdx_value ==
    io_loadRegIn_1_bits_uop_robIdx_value | flow_entry_1_17_uop_robIdx_value == io_loadRegIn_1_bits_uop_robIdx_value |
    flow_entry_1_18_uop_robIdx_value == io_loadRegIn_1_bits_uop_robIdx_value | flow_entry_1_19_uop_robIdx_value ==
    io_loadRegIn_1_bits_uop_robIdx_value | flow_entry_1_20_uop_robIdx_value == io_loadRegIn_1_bits_uop_robIdx_value |
    flow_entry_1_21_uop_robIdx_value == io_loadRegIn_1_bits_uop_robIdx_value | flow_entry_1_22_uop_robIdx_value ==
    io_loadRegIn_1_bits_uop_robIdx_value | flow_entry_1_23_uop_robIdx_value == io_loadRegIn_1_bits_uop_robIdx_value |
    flow_entry_1_24_uop_robIdx_value == io_loadRegIn_1_bits_uop_robIdx_value | flow_entry_1_25_uop_robIdx_value ==
    io_loadRegIn_1_bits_uop_robIdx_value | flow_entry_1_26_uop_robIdx_value == io_loadRegIn_1_bits_uop_robIdx_value |
    flow_entry_1_27_uop_robIdx_value == io_loadRegIn_1_bits_uop_robIdx_value | flow_entry_1_28_uop_robIdx_value ==
    io_loadRegIn_1_bits_uop_robIdx_value | flow_entry_1_29_uop_robIdx_value == io_loadRegIn_1_bits_uop_robIdx_value |
    flow_entry_1_30_uop_robIdx_value == io_loadRegIn_1_bits_uop_robIdx_value; // @[Vlflowqueue.scala 161:117]
  wire  needAlloc_1 = ~(_needAlloc_1_T_61 | flow_entry_0_31_uop_robIdx_value == io_loadRegIn_1_bits_uop_robIdx_value | (
    _needAlloc_1_T_124 | flow_entry_1_31_uop_robIdx_value == io_loadRegIn_1_bits_uop_robIdx_value)) &
    io_loadRegIn_1_valid; // @[Vlflowqueue.scala 161:139]
  wire [4:0] _vend_0_1_T_2 = {{1'd0}, io_loadRegIn_1_bits_baseaddr[3:0]}; // @[Vlflowqueue.scala 164:41]
  wire [5:0] _vend_1_1_T_2 = {{1'd0}, io_loadRegIn_1_bits_baseaddr[4:0]}; // @[Vlflowqueue.scala 165:41]
  wire [6:0] _vend_2_1_T_2 = {{1'd0}, io_loadRegIn_1_bits_baseaddr[5:0]}; // @[Vlflowqueue.scala 166:41]
  wire [7:0] _vend_3_1_T_2 = {{1'd0}, io_loadRegIn_1_bits_baseaddr[6:0]}; // @[Vlflowqueue.scala 167:41]
  wire [7:0] vend_3_1 = {{1'd0}, _vend_3_1_T_2[6:0]}; // @[Vlflowqueue.scala 144:29 167:21]
  wire [6:0] vend_2_1 = {{1'd0}, _vend_2_1_T_2[5:0]}; // @[Vlflowqueue.scala 143:29 166:21]
  wire [5:0] vend_1_1 = {{1'd0}, _vend_1_1_T_2[4:0]}; // @[Vlflowqueue.scala 142:29 165:21]
  wire [4:0] vend_0_1 = {{1'd0}, _vend_0_1_T_2[3:0]}; // @[Vlflowqueue.scala 141:29 164:21]
  wire [1:0] _flowWriteNumber_1_T_10 = vend_1_1[5] ? vend_1_1[5:4] : {{1'd0}, vend_0_1[4]}; // @[Vlflowqueue.scala 168:114]
  wire [2:0] _flowWriteNumber_1_T_11 = vend_2_1[6] ? vend_2_1[6:4] : {{1'd0}, _flowWriteNumber_1_T_10}; // @[Vlflowqueue.scala 168:72]
  wire [3:0] _flowWriteNumber_1_T_12 = vend_3_1[7] ? vend_3_1[7:4] : {{1'd0}, _flowWriteNumber_1_T_11}; // @[Vlflowqueue.scala 168:30]
  reg [4:0] enqPtr_0_value; // @[Vlflowqueue.scala 171:23]
  reg [4:0] enqPtr_1_value; // @[Vlflowqueue.scala 171:23]
  reg  deqPtr_0_flag; // @[Vlflowqueue.scala 172:23]
  reg [4:0] deqPtr_0_value; // @[Vlflowqueue.scala 172:23]
  reg  deqPtr_1_flag; // @[Vlflowqueue.scala 172:23]
  reg [4:0] deqPtr_1_value; // @[Vlflowqueue.scala 172:23]
  wire  cross128_0 = io_loadRegIn_0_bits_baseaddr[3:0] != 4'h0; // @[Vlflowqueue.scala 176:42]
  wire [2:0] flowWriteNumber_0 = _flowWriteNumber_0_T_12[2:0]; // @[Vlflowqueue.scala 145:29 168:24]
  wire [2:0] _GEN_161414 = {{2'd0}, cross128_0}; // @[Vlflowqueue.scala 177:50]
  wire [2:0] _realFlowNum_0_T_1 = flowWriteNumber_0 + _GEN_161414; // @[Vlflowqueue.scala 177:50]
  wire [3:0] realFlowNum_0 = {{1'd0}, _realFlowNum_0_T_1}; // @[Vlflowqueue.scala 146:29 177:21]
  wire [4:0] _GEN_161415 = {{1'd0}, realFlowNum_0}; // @[Vlflowqueue.scala 178:40]
  wire  cross128_1 = io_loadRegIn_1_bits_baseaddr[3:0] != 4'h0; // @[Vlflowqueue.scala 176:42]
  wire [2:0] flowWriteNumber_1 = _flowWriteNumber_1_T_12[2:0]; // @[Vlflowqueue.scala 145:29 168:24]
  wire [2:0] _GEN_161416 = {{2'd0}, cross128_1}; // @[Vlflowqueue.scala 177:50]
  wire [2:0] _realFlowNum_1_T_1 = flowWriteNumber_1 + _GEN_161416; // @[Vlflowqueue.scala 177:50]
  wire [3:0] realFlowNum_1 = {{1'd0}, _realFlowNum_1_T_1}; // @[Vlflowqueue.scala 146:29 177:21]
  wire [4:0] _GEN_161417 = {{1'd0}, realFlowNum_1}; // @[Vlflowqueue.scala 178:40]
  wire [5:0] _GEN_161418 = {{1'd0}, enqPtr_0_value}; // @[CircularQueuePtr.scala 82:25]
  wire [5:0] _GEN_161420 = {{1'd0}, enqPtr_1_value}; // @[CircularQueuePtr.scala 82:25]
  wire [4:0] _index_0_T_17 = enqPtr_0_value + 5'h8; // @[Vlflowqueue.scala 195:39]
  wire [4:0] _index_0_T_15 = enqPtr_0_value + 5'h7; // @[Vlflowqueue.scala 195:39]
  wire [4:0] _index_0_T_13 = enqPtr_0_value + 5'h6; // @[Vlflowqueue.scala 195:39]
  wire [4:0] _index_0_T_11 = enqPtr_0_value + 5'h5; // @[Vlflowqueue.scala 195:39]
  wire [4:0] _index_0_T_9 = enqPtr_0_value + 5'h4; // @[Vlflowqueue.scala 195:39]
  wire [4:0] _index_0_T_7 = enqPtr_0_value + 5'h3; // @[Vlflowqueue.scala 195:39]
  wire [4:0] _index_0_T_5 = enqPtr_0_value + 5'h2; // @[Vlflowqueue.scala 195:39]
  wire [4:0] _index_0_T_3 = enqPtr_0_value + 5'h1; // @[Vlflowqueue.scala 195:39]
  wire [4:0] _GEN_16098 = 4'h1 < realFlowNum_0 ? _index_0_T_3 : _GEN_161418[4:0]; // @[Vlflowqueue.scala 194:37 195:20]
  wire [4:0] _GEN_24164 = 4'h2 < realFlowNum_0 ? _index_0_T_5 : _GEN_16098; // @[Vlflowqueue.scala 194:37 195:20]
  wire [4:0] _GEN_32230 = 4'h3 < realFlowNum_0 ? _index_0_T_7 : _GEN_24164; // @[Vlflowqueue.scala 194:37 195:20]
  wire [4:0] _GEN_40296 = 4'h4 < realFlowNum_0 ? _index_0_T_9 : _GEN_32230; // @[Vlflowqueue.scala 194:37 195:20]
  wire [4:0] _GEN_48362 = 4'h5 < realFlowNum_0 ? _index_0_T_11 : _GEN_40296; // @[Vlflowqueue.scala 194:37 195:20]
  wire [4:0] _GEN_56428 = 4'h6 < realFlowNum_0 ? _index_0_T_13 : _GEN_48362; // @[Vlflowqueue.scala 194:37 195:20]
  wire [4:0] _GEN_64494 = 4'h7 < realFlowNum_0 ? _index_0_T_15 : _GEN_56428; // @[Vlflowqueue.scala 194:37 195:20]
  wire [4:0] index_0 = 4'h8 < realFlowNum_0 ? _index_0_T_17 : _GEN_64494; // @[Vlflowqueue.scala 194:37 195:20]
  wire  _GEN_161423 = 5'h0 == index_0; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_3808 = 5'h0 == index_0 | flow_entry_valid_0_0; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_161424 = 5'h1 == index_0; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_3809 = 5'h1 == index_0 | flow_entry_valid_0_1; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_161425 = 5'h2 == index_0; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_3810 = 5'h2 == index_0 | flow_entry_valid_0_2; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_161426 = 5'h3 == index_0; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_3811 = 5'h3 == index_0 | flow_entry_valid_0_3; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_161427 = 5'h4 == index_0; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_3812 = 5'h4 == index_0 | flow_entry_valid_0_4; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_161428 = 5'h5 == index_0; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_3813 = 5'h5 == index_0 | flow_entry_valid_0_5; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_161429 = 5'h6 == index_0; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_3814 = 5'h6 == index_0 | flow_entry_valid_0_6; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_161430 = 5'h7 == index_0; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_3815 = 5'h7 == index_0 | flow_entry_valid_0_7; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_161431 = 5'h8 == index_0; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_3816 = 5'h8 == index_0 | flow_entry_valid_0_8; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_161432 = 5'h9 == index_0; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_3817 = 5'h9 == index_0 | flow_entry_valid_0_9; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_161433 = 5'ha == index_0; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_3818 = 5'ha == index_0 | flow_entry_valid_0_10; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_161434 = 5'hb == index_0; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_3819 = 5'hb == index_0 | flow_entry_valid_0_11; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_161435 = 5'hc == index_0; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_3820 = 5'hc == index_0 | flow_entry_valid_0_12; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_161436 = 5'hd == index_0; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_3821 = 5'hd == index_0 | flow_entry_valid_0_13; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_161437 = 5'he == index_0; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_3822 = 5'he == index_0 | flow_entry_valid_0_14; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_161438 = 5'hf == index_0; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_3823 = 5'hf == index_0 | flow_entry_valid_0_15; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_161439 = 5'h10 == index_0; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_3824 = 5'h10 == index_0 | flow_entry_valid_0_16; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_161440 = 5'h11 == index_0; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_3825 = 5'h11 == index_0 | flow_entry_valid_0_17; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_161441 = 5'h12 == index_0; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_3826 = 5'h12 == index_0 | flow_entry_valid_0_18; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_161442 = 5'h13 == index_0; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_3827 = 5'h13 == index_0 | flow_entry_valid_0_19; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_161443 = 5'h14 == index_0; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_3828 = 5'h14 == index_0 | flow_entry_valid_0_20; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_161444 = 5'h15 == index_0; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_3829 = 5'h15 == index_0 | flow_entry_valid_0_21; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_161445 = 5'h16 == index_0; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_3830 = 5'h16 == index_0 | flow_entry_valid_0_22; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_161446 = 5'h17 == index_0; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_3831 = 5'h17 == index_0 | flow_entry_valid_0_23; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_161447 = 5'h18 == index_0; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_3832 = 5'h18 == index_0 | flow_entry_valid_0_24; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_161448 = 5'h19 == index_0; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_3833 = 5'h19 == index_0 | flow_entry_valid_0_25; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_161449 = 5'h1a == index_0; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_3834 = 5'h1a == index_0 | flow_entry_valid_0_26; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_161450 = 5'h1b == index_0; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_3835 = 5'h1b == index_0 | flow_entry_valid_0_27; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_161451 = 5'h1c == index_0; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_3836 = 5'h1c == index_0 | flow_entry_valid_0_28; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_161452 = 5'h1d == index_0; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_3837 = 5'h1d == index_0 | flow_entry_valid_0_29; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_161453 = 5'h1e == index_0; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_3838 = 5'h1e == index_0 | flow_entry_valid_0_30; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_161454 = 5'h1f == index_0; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_3839 = 5'h1f == index_0 | flow_entry_valid_0_31; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire [4:0] _GEN_6784 = 5'h0 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : flow_entry_0_0_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 198:{51,51}]
  wire [4:0] _GEN_6785 = 5'h1 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : flow_entry_0_1_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 198:{51,51}]
  wire [4:0] _GEN_6786 = 5'h2 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : flow_entry_0_2_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 198:{51,51}]
  wire [4:0] _GEN_6787 = 5'h3 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : flow_entry_0_3_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 198:{51,51}]
  wire [4:0] _GEN_6788 = 5'h4 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : flow_entry_0_4_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 198:{51,51}]
  wire [4:0] _GEN_6789 = 5'h5 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : flow_entry_0_5_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 198:{51,51}]
  wire [4:0] _GEN_6790 = 5'h6 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : flow_entry_0_6_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 198:{51,51}]
  wire [4:0] _GEN_6791 = 5'h7 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : flow_entry_0_7_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 198:{51,51}]
  wire [4:0] _GEN_6792 = 5'h8 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : flow_entry_0_8_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 198:{51,51}]
  wire [4:0] _GEN_6793 = 5'h9 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : flow_entry_0_9_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 198:{51,51}]
  wire [4:0] _GEN_6794 = 5'ha == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : flow_entry_0_10_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 198:{51,51}]
  wire [4:0] _GEN_6795 = 5'hb == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : flow_entry_0_11_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 198:{51,51}]
  wire [4:0] _GEN_6796 = 5'hc == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : flow_entry_0_12_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 198:{51,51}]
  wire [4:0] _GEN_6797 = 5'hd == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : flow_entry_0_13_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 198:{51,51}]
  wire [4:0] _GEN_6798 = 5'he == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : flow_entry_0_14_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 198:{51,51}]
  wire [4:0] _GEN_6799 = 5'hf == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : flow_entry_0_15_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 198:{51,51}]
  wire [4:0] _GEN_6800 = 5'h10 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : flow_entry_0_16_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 198:{51,51}]
  wire [4:0] _GEN_6801 = 5'h11 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : flow_entry_0_17_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 198:{51,51}]
  wire [4:0] _GEN_6802 = 5'h12 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : flow_entry_0_18_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 198:{51,51}]
  wire [4:0] _GEN_6803 = 5'h13 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : flow_entry_0_19_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 198:{51,51}]
  wire [4:0] _GEN_6804 = 5'h14 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : flow_entry_0_20_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 198:{51,51}]
  wire [4:0] _GEN_6805 = 5'h15 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : flow_entry_0_21_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 198:{51,51}]
  wire [4:0] _GEN_6806 = 5'h16 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : flow_entry_0_22_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 198:{51,51}]
  wire [4:0] _GEN_6807 = 5'h17 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : flow_entry_0_23_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 198:{51,51}]
  wire [4:0] _GEN_6808 = 5'h18 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : flow_entry_0_24_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 198:{51,51}]
  wire [4:0] _GEN_6809 = 5'h19 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : flow_entry_0_25_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 198:{51,51}]
  wire [4:0] _GEN_6810 = 5'h1a == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : flow_entry_0_26_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 198:{51,51}]
  wire [4:0] _GEN_6811 = 5'h1b == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : flow_entry_0_27_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 198:{51,51}]
  wire [4:0] _GEN_6812 = 5'h1c == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : flow_entry_0_28_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 198:{51,51}]
  wire [4:0] _GEN_6813 = 5'h1d == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : flow_entry_0_29_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 198:{51,51}]
  wire [4:0] _GEN_6814 = 5'h1e == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : flow_entry_0_30_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 198:{51,51}]
  wire [4:0] _GEN_6815 = 5'h1f == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : flow_entry_0_31_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 198:{51,51}]
  wire [39:0] _vaddr_0_T_1 = {{1'd0}, io_loadRegIn_0_bits_baseaddr}; // @[Vlflowqueue.scala 91:32]
  wire [38:0] _vaddr_0_T_162 = io_loadRegIn_0_bits_baseaddr + 39'h80; // @[Vlflowqueue.scala 91:32]
  wire [38:0] _vaddr_0_T_142 = io_loadRegIn_0_bits_baseaddr + 39'h70; // @[Vlflowqueue.scala 91:32]
  wire [38:0] _vaddr_0_T_122 = io_loadRegIn_0_bits_baseaddr + 39'h60; // @[Vlflowqueue.scala 91:32]
  wire [38:0] _vaddr_0_T_102 = io_loadRegIn_0_bits_baseaddr + 39'h50; // @[Vlflowqueue.scala 91:32]
  wire [38:0] _vaddr_0_T_82 = io_loadRegIn_0_bits_baseaddr + 39'h40; // @[Vlflowqueue.scala 91:32]
  wire [38:0] _vaddr_0_T_62 = io_loadRegIn_0_bits_baseaddr + 39'h30; // @[Vlflowqueue.scala 91:32]
  wire [38:0] _vaddr_0_T_42 = io_loadRegIn_0_bits_baseaddr + 39'h20; // @[Vlflowqueue.scala 91:32]
  wire [38:0] _vaddr_0_T_22 = io_loadRegIn_0_bits_baseaddr + 39'h10; // @[Vlflowqueue.scala 91:32]
  wire [38:0] _GEN_19619 = 4'h1 < realFlowNum_0 ? _vaddr_0_T_22 : _vaddr_0_T_1[38:0]; // @[Vlflowqueue.scala 194:37 201:51]
  wire [38:0] _GEN_27685 = 4'h2 < realFlowNum_0 ? _vaddr_0_T_42 : _GEN_19619; // @[Vlflowqueue.scala 194:37 201:51]
  wire [38:0] _GEN_35751 = 4'h3 < realFlowNum_0 ? _vaddr_0_T_62 : _GEN_27685; // @[Vlflowqueue.scala 194:37 201:51]
  wire [38:0] _GEN_43817 = 4'h4 < realFlowNum_0 ? _vaddr_0_T_82 : _GEN_35751; // @[Vlflowqueue.scala 194:37 201:51]
  wire [38:0] _GEN_51883 = 4'h5 < realFlowNum_0 ? _vaddr_0_T_102 : _GEN_43817; // @[Vlflowqueue.scala 194:37 201:51]
  wire [38:0] _GEN_59949 = 4'h6 < realFlowNum_0 ? _vaddr_0_T_122 : _GEN_51883; // @[Vlflowqueue.scala 194:37 201:51]
  wire [38:0] _GEN_68015 = 4'h7 < realFlowNum_0 ? _vaddr_0_T_142 : _GEN_59949; // @[Vlflowqueue.scala 194:37 201:51]
  wire [38:0] vaddr_0 = 4'h8 < realFlowNum_0 ? _vaddr_0_T_162 : _GEN_68015; // @[Vlflowqueue.scala 194:37 201:51]
  wire [38:0] _GEN_7360 = 5'h0 == index_0 ? vaddr_0 : flow_entry_0_0_vaddr; // @[Vlflowqueue.scala 134:29 203:{51,51}]
  wire [38:0] _GEN_7361 = 5'h1 == index_0 ? vaddr_0 : flow_entry_0_1_vaddr; // @[Vlflowqueue.scala 134:29 203:{51,51}]
  wire [38:0] _GEN_7362 = 5'h2 == index_0 ? vaddr_0 : flow_entry_0_2_vaddr; // @[Vlflowqueue.scala 134:29 203:{51,51}]
  wire [38:0] _GEN_7363 = 5'h3 == index_0 ? vaddr_0 : flow_entry_0_3_vaddr; // @[Vlflowqueue.scala 134:29 203:{51,51}]
  wire [38:0] _GEN_7364 = 5'h4 == index_0 ? vaddr_0 : flow_entry_0_4_vaddr; // @[Vlflowqueue.scala 134:29 203:{51,51}]
  wire [38:0] _GEN_7365 = 5'h5 == index_0 ? vaddr_0 : flow_entry_0_5_vaddr; // @[Vlflowqueue.scala 134:29 203:{51,51}]
  wire [38:0] _GEN_7366 = 5'h6 == index_0 ? vaddr_0 : flow_entry_0_6_vaddr; // @[Vlflowqueue.scala 134:29 203:{51,51}]
  wire [38:0] _GEN_7367 = 5'h7 == index_0 ? vaddr_0 : flow_entry_0_7_vaddr; // @[Vlflowqueue.scala 134:29 203:{51,51}]
  wire [38:0] _GEN_7368 = 5'h8 == index_0 ? vaddr_0 : flow_entry_0_8_vaddr; // @[Vlflowqueue.scala 134:29 203:{51,51}]
  wire [38:0] _GEN_7369 = 5'h9 == index_0 ? vaddr_0 : flow_entry_0_9_vaddr; // @[Vlflowqueue.scala 134:29 203:{51,51}]
  wire [38:0] _GEN_7370 = 5'ha == index_0 ? vaddr_0 : flow_entry_0_10_vaddr; // @[Vlflowqueue.scala 134:29 203:{51,51}]
  wire [38:0] _GEN_7371 = 5'hb == index_0 ? vaddr_0 : flow_entry_0_11_vaddr; // @[Vlflowqueue.scala 134:29 203:{51,51}]
  wire [38:0] _GEN_7372 = 5'hc == index_0 ? vaddr_0 : flow_entry_0_12_vaddr; // @[Vlflowqueue.scala 134:29 203:{51,51}]
  wire [38:0] _GEN_7373 = 5'hd == index_0 ? vaddr_0 : flow_entry_0_13_vaddr; // @[Vlflowqueue.scala 134:29 203:{51,51}]
  wire [38:0] _GEN_7374 = 5'he == index_0 ? vaddr_0 : flow_entry_0_14_vaddr; // @[Vlflowqueue.scala 134:29 203:{51,51}]
  wire [38:0] _GEN_7375 = 5'hf == index_0 ? vaddr_0 : flow_entry_0_15_vaddr; // @[Vlflowqueue.scala 134:29 203:{51,51}]
  wire [38:0] _GEN_7376 = 5'h10 == index_0 ? vaddr_0 : flow_entry_0_16_vaddr; // @[Vlflowqueue.scala 134:29 203:{51,51}]
  wire [38:0] _GEN_7377 = 5'h11 == index_0 ? vaddr_0 : flow_entry_0_17_vaddr; // @[Vlflowqueue.scala 134:29 203:{51,51}]
  wire [38:0] _GEN_7378 = 5'h12 == index_0 ? vaddr_0 : flow_entry_0_18_vaddr; // @[Vlflowqueue.scala 134:29 203:{51,51}]
  wire [38:0] _GEN_7379 = 5'h13 == index_0 ? vaddr_0 : flow_entry_0_19_vaddr; // @[Vlflowqueue.scala 134:29 203:{51,51}]
  wire [38:0] _GEN_7380 = 5'h14 == index_0 ? vaddr_0 : flow_entry_0_20_vaddr; // @[Vlflowqueue.scala 134:29 203:{51,51}]
  wire [38:0] _GEN_7381 = 5'h15 == index_0 ? vaddr_0 : flow_entry_0_21_vaddr; // @[Vlflowqueue.scala 134:29 203:{51,51}]
  wire [38:0] _GEN_7382 = 5'h16 == index_0 ? vaddr_0 : flow_entry_0_22_vaddr; // @[Vlflowqueue.scala 134:29 203:{51,51}]
  wire [38:0] _GEN_7383 = 5'h17 == index_0 ? vaddr_0 : flow_entry_0_23_vaddr; // @[Vlflowqueue.scala 134:29 203:{51,51}]
  wire [38:0] _GEN_7384 = 5'h18 == index_0 ? vaddr_0 : flow_entry_0_24_vaddr; // @[Vlflowqueue.scala 134:29 203:{51,51}]
  wire [38:0] _GEN_7385 = 5'h19 == index_0 ? vaddr_0 : flow_entry_0_25_vaddr; // @[Vlflowqueue.scala 134:29 203:{51,51}]
  wire [38:0] _GEN_7386 = 5'h1a == index_0 ? vaddr_0 : flow_entry_0_26_vaddr; // @[Vlflowqueue.scala 134:29 203:{51,51}]
  wire [38:0] _GEN_7387 = 5'h1b == index_0 ? vaddr_0 : flow_entry_0_27_vaddr; // @[Vlflowqueue.scala 134:29 203:{51,51}]
  wire [38:0] _GEN_7388 = 5'h1c == index_0 ? vaddr_0 : flow_entry_0_28_vaddr; // @[Vlflowqueue.scala 134:29 203:{51,51}]
  wire [38:0] _GEN_7389 = 5'h1d == index_0 ? vaddr_0 : flow_entry_0_29_vaddr; // @[Vlflowqueue.scala 134:29 203:{51,51}]
  wire [38:0] _GEN_7390 = 5'h1e == index_0 ? vaddr_0 : flow_entry_0_30_vaddr; // @[Vlflowqueue.scala 134:29 203:{51,51}]
  wire [38:0] _GEN_7391 = 5'h1f == index_0 ? vaddr_0 : flow_entry_0_31_vaddr; // @[Vlflowqueue.scala 134:29 203:{51,51}]
  wire  _GEN_8033 = 4'h0 < realFlowNum_0 ? _GEN_3808 : flow_entry_valid_0_0; // @[Vlflowqueue.scala 135:33 194:37]
  wire  _GEN_8034 = 4'h0 < realFlowNum_0 ? _GEN_3809 : flow_entry_valid_0_1; // @[Vlflowqueue.scala 135:33 194:37]
  wire  _GEN_8035 = 4'h0 < realFlowNum_0 ? _GEN_3810 : flow_entry_valid_0_2; // @[Vlflowqueue.scala 135:33 194:37]
  wire  _GEN_8036 = 4'h0 < realFlowNum_0 ? _GEN_3811 : flow_entry_valid_0_3; // @[Vlflowqueue.scala 135:33 194:37]
  wire  _GEN_8037 = 4'h0 < realFlowNum_0 ? _GEN_3812 : flow_entry_valid_0_4; // @[Vlflowqueue.scala 135:33 194:37]
  wire  _GEN_8038 = 4'h0 < realFlowNum_0 ? _GEN_3813 : flow_entry_valid_0_5; // @[Vlflowqueue.scala 135:33 194:37]
  wire  _GEN_8039 = 4'h0 < realFlowNum_0 ? _GEN_3814 : flow_entry_valid_0_6; // @[Vlflowqueue.scala 135:33 194:37]
  wire  _GEN_8040 = 4'h0 < realFlowNum_0 ? _GEN_3815 : flow_entry_valid_0_7; // @[Vlflowqueue.scala 135:33 194:37]
  wire  _GEN_8041 = 4'h0 < realFlowNum_0 ? _GEN_3816 : flow_entry_valid_0_8; // @[Vlflowqueue.scala 135:33 194:37]
  wire  _GEN_8042 = 4'h0 < realFlowNum_0 ? _GEN_3817 : flow_entry_valid_0_9; // @[Vlflowqueue.scala 135:33 194:37]
  wire  _GEN_8043 = 4'h0 < realFlowNum_0 ? _GEN_3818 : flow_entry_valid_0_10; // @[Vlflowqueue.scala 135:33 194:37]
  wire  _GEN_8044 = 4'h0 < realFlowNum_0 ? _GEN_3819 : flow_entry_valid_0_11; // @[Vlflowqueue.scala 135:33 194:37]
  wire  _GEN_8045 = 4'h0 < realFlowNum_0 ? _GEN_3820 : flow_entry_valid_0_12; // @[Vlflowqueue.scala 135:33 194:37]
  wire  _GEN_8046 = 4'h0 < realFlowNum_0 ? _GEN_3821 : flow_entry_valid_0_13; // @[Vlflowqueue.scala 135:33 194:37]
  wire  _GEN_8047 = 4'h0 < realFlowNum_0 ? _GEN_3822 : flow_entry_valid_0_14; // @[Vlflowqueue.scala 135:33 194:37]
  wire  _GEN_8048 = 4'h0 < realFlowNum_0 ? _GEN_3823 : flow_entry_valid_0_15; // @[Vlflowqueue.scala 135:33 194:37]
  wire  _GEN_8049 = 4'h0 < realFlowNum_0 ? _GEN_3824 : flow_entry_valid_0_16; // @[Vlflowqueue.scala 135:33 194:37]
  wire  _GEN_8050 = 4'h0 < realFlowNum_0 ? _GEN_3825 : flow_entry_valid_0_17; // @[Vlflowqueue.scala 135:33 194:37]
  wire  _GEN_8051 = 4'h0 < realFlowNum_0 ? _GEN_3826 : flow_entry_valid_0_18; // @[Vlflowqueue.scala 135:33 194:37]
  wire  _GEN_8052 = 4'h0 < realFlowNum_0 ? _GEN_3827 : flow_entry_valid_0_19; // @[Vlflowqueue.scala 135:33 194:37]
  wire  _GEN_8053 = 4'h0 < realFlowNum_0 ? _GEN_3828 : flow_entry_valid_0_20; // @[Vlflowqueue.scala 135:33 194:37]
  wire  _GEN_8054 = 4'h0 < realFlowNum_0 ? _GEN_3829 : flow_entry_valid_0_21; // @[Vlflowqueue.scala 135:33 194:37]
  wire  _GEN_8055 = 4'h0 < realFlowNum_0 ? _GEN_3830 : flow_entry_valid_0_22; // @[Vlflowqueue.scala 135:33 194:37]
  wire  _GEN_8056 = 4'h0 < realFlowNum_0 ? _GEN_3831 : flow_entry_valid_0_23; // @[Vlflowqueue.scala 135:33 194:37]
  wire  _GEN_8057 = 4'h0 < realFlowNum_0 ? _GEN_3832 : flow_entry_valid_0_24; // @[Vlflowqueue.scala 135:33 194:37]
  wire  _GEN_8058 = 4'h0 < realFlowNum_0 ? _GEN_3833 : flow_entry_valid_0_25; // @[Vlflowqueue.scala 135:33 194:37]
  wire  _GEN_8059 = 4'h0 < realFlowNum_0 ? _GEN_3834 : flow_entry_valid_0_26; // @[Vlflowqueue.scala 135:33 194:37]
  wire  _GEN_8060 = 4'h0 < realFlowNum_0 ? _GEN_3835 : flow_entry_valid_0_27; // @[Vlflowqueue.scala 135:33 194:37]
  wire  _GEN_8061 = 4'h0 < realFlowNum_0 ? _GEN_3836 : flow_entry_valid_0_28; // @[Vlflowqueue.scala 135:33 194:37]
  wire  _GEN_8062 = 4'h0 < realFlowNum_0 ? _GEN_3837 : flow_entry_valid_0_29; // @[Vlflowqueue.scala 135:33 194:37]
  wire  _GEN_8063 = 4'h0 < realFlowNum_0 ? _GEN_3838 : flow_entry_valid_0_30; // @[Vlflowqueue.scala 135:33 194:37]
  wire  _GEN_8064 = 4'h0 < realFlowNum_0 ? _GEN_3839 : flow_entry_valid_0_31; // @[Vlflowqueue.scala 135:33 194:37]
  wire [4:0] _GEN_11009 = 4'h0 < realFlowNum_0 ? _GEN_6784 : flow_entry_0_0_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 194:37]
  wire [4:0] _GEN_11010 = 4'h0 < realFlowNum_0 ? _GEN_6785 : flow_entry_0_1_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 194:37]
  wire [4:0] _GEN_11011 = 4'h0 < realFlowNum_0 ? _GEN_6786 : flow_entry_0_2_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 194:37]
  wire [4:0] _GEN_11012 = 4'h0 < realFlowNum_0 ? _GEN_6787 : flow_entry_0_3_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 194:37]
  wire [4:0] _GEN_11013 = 4'h0 < realFlowNum_0 ? _GEN_6788 : flow_entry_0_4_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 194:37]
  wire [4:0] _GEN_11014 = 4'h0 < realFlowNum_0 ? _GEN_6789 : flow_entry_0_5_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 194:37]
  wire [4:0] _GEN_11015 = 4'h0 < realFlowNum_0 ? _GEN_6790 : flow_entry_0_6_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 194:37]
  wire [4:0] _GEN_11016 = 4'h0 < realFlowNum_0 ? _GEN_6791 : flow_entry_0_7_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 194:37]
  wire [4:0] _GEN_11017 = 4'h0 < realFlowNum_0 ? _GEN_6792 : flow_entry_0_8_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 194:37]
  wire [4:0] _GEN_11018 = 4'h0 < realFlowNum_0 ? _GEN_6793 : flow_entry_0_9_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 194:37]
  wire [4:0] _GEN_11019 = 4'h0 < realFlowNum_0 ? _GEN_6794 : flow_entry_0_10_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 194:37]
  wire [4:0] _GEN_11020 = 4'h0 < realFlowNum_0 ? _GEN_6795 : flow_entry_0_11_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 194:37]
  wire [4:0] _GEN_11021 = 4'h0 < realFlowNum_0 ? _GEN_6796 : flow_entry_0_12_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 194:37]
  wire [4:0] _GEN_11022 = 4'h0 < realFlowNum_0 ? _GEN_6797 : flow_entry_0_13_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 194:37]
  wire [4:0] _GEN_11023 = 4'h0 < realFlowNum_0 ? _GEN_6798 : flow_entry_0_14_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 194:37]
  wire [4:0] _GEN_11024 = 4'h0 < realFlowNum_0 ? _GEN_6799 : flow_entry_0_15_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 194:37]
  wire [4:0] _GEN_11025 = 4'h0 < realFlowNum_0 ? _GEN_6800 : flow_entry_0_16_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 194:37]
  wire [4:0] _GEN_11026 = 4'h0 < realFlowNum_0 ? _GEN_6801 : flow_entry_0_17_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 194:37]
  wire [4:0] _GEN_11027 = 4'h0 < realFlowNum_0 ? _GEN_6802 : flow_entry_0_18_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 194:37]
  wire [4:0] _GEN_11028 = 4'h0 < realFlowNum_0 ? _GEN_6803 : flow_entry_0_19_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 194:37]
  wire [4:0] _GEN_11029 = 4'h0 < realFlowNum_0 ? _GEN_6804 : flow_entry_0_20_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 194:37]
  wire [4:0] _GEN_11030 = 4'h0 < realFlowNum_0 ? _GEN_6805 : flow_entry_0_21_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 194:37]
  wire [4:0] _GEN_11031 = 4'h0 < realFlowNum_0 ? _GEN_6806 : flow_entry_0_22_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 194:37]
  wire [4:0] _GEN_11032 = 4'h0 < realFlowNum_0 ? _GEN_6807 : flow_entry_0_23_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 194:37]
  wire [4:0] _GEN_11033 = 4'h0 < realFlowNum_0 ? _GEN_6808 : flow_entry_0_24_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 194:37]
  wire [4:0] _GEN_11034 = 4'h0 < realFlowNum_0 ? _GEN_6809 : flow_entry_0_25_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 194:37]
  wire [4:0] _GEN_11035 = 4'h0 < realFlowNum_0 ? _GEN_6810 : flow_entry_0_26_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 194:37]
  wire [4:0] _GEN_11036 = 4'h0 < realFlowNum_0 ? _GEN_6811 : flow_entry_0_27_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 194:37]
  wire [4:0] _GEN_11037 = 4'h0 < realFlowNum_0 ? _GEN_6812 : flow_entry_0_28_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 194:37]
  wire [4:0] _GEN_11038 = 4'h0 < realFlowNum_0 ? _GEN_6813 : flow_entry_0_29_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 194:37]
  wire [4:0] _GEN_11039 = 4'h0 < realFlowNum_0 ? _GEN_6814 : flow_entry_0_30_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 194:37]
  wire [4:0] _GEN_11040 = 4'h0 < realFlowNum_0 ? _GEN_6815 : flow_entry_0_31_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 194:37]
  wire [38:0] _GEN_11586 = 4'h0 < realFlowNum_0 ? _GEN_7360 : flow_entry_0_0_vaddr; // @[Vlflowqueue.scala 134:29 194:37]
  wire [38:0] _GEN_11587 = 4'h0 < realFlowNum_0 ? _GEN_7361 : flow_entry_0_1_vaddr; // @[Vlflowqueue.scala 134:29 194:37]
  wire [38:0] _GEN_11588 = 4'h0 < realFlowNum_0 ? _GEN_7362 : flow_entry_0_2_vaddr; // @[Vlflowqueue.scala 134:29 194:37]
  wire [38:0] _GEN_11589 = 4'h0 < realFlowNum_0 ? _GEN_7363 : flow_entry_0_3_vaddr; // @[Vlflowqueue.scala 134:29 194:37]
  wire [38:0] _GEN_11590 = 4'h0 < realFlowNum_0 ? _GEN_7364 : flow_entry_0_4_vaddr; // @[Vlflowqueue.scala 134:29 194:37]
  wire [38:0] _GEN_11591 = 4'h0 < realFlowNum_0 ? _GEN_7365 : flow_entry_0_5_vaddr; // @[Vlflowqueue.scala 134:29 194:37]
  wire [38:0] _GEN_11592 = 4'h0 < realFlowNum_0 ? _GEN_7366 : flow_entry_0_6_vaddr; // @[Vlflowqueue.scala 134:29 194:37]
  wire [38:0] _GEN_11593 = 4'h0 < realFlowNum_0 ? _GEN_7367 : flow_entry_0_7_vaddr; // @[Vlflowqueue.scala 134:29 194:37]
  wire [38:0] _GEN_11594 = 4'h0 < realFlowNum_0 ? _GEN_7368 : flow_entry_0_8_vaddr; // @[Vlflowqueue.scala 134:29 194:37]
  wire [38:0] _GEN_11595 = 4'h0 < realFlowNum_0 ? _GEN_7369 : flow_entry_0_9_vaddr; // @[Vlflowqueue.scala 134:29 194:37]
  wire [38:0] _GEN_11596 = 4'h0 < realFlowNum_0 ? _GEN_7370 : flow_entry_0_10_vaddr; // @[Vlflowqueue.scala 134:29 194:37]
  wire [38:0] _GEN_11597 = 4'h0 < realFlowNum_0 ? _GEN_7371 : flow_entry_0_11_vaddr; // @[Vlflowqueue.scala 134:29 194:37]
  wire [38:0] _GEN_11598 = 4'h0 < realFlowNum_0 ? _GEN_7372 : flow_entry_0_12_vaddr; // @[Vlflowqueue.scala 134:29 194:37]
  wire [38:0] _GEN_11599 = 4'h0 < realFlowNum_0 ? _GEN_7373 : flow_entry_0_13_vaddr; // @[Vlflowqueue.scala 134:29 194:37]
  wire [38:0] _GEN_11600 = 4'h0 < realFlowNum_0 ? _GEN_7374 : flow_entry_0_14_vaddr; // @[Vlflowqueue.scala 134:29 194:37]
  wire [38:0] _GEN_11601 = 4'h0 < realFlowNum_0 ? _GEN_7375 : flow_entry_0_15_vaddr; // @[Vlflowqueue.scala 134:29 194:37]
  wire [38:0] _GEN_11602 = 4'h0 < realFlowNum_0 ? _GEN_7376 : flow_entry_0_16_vaddr; // @[Vlflowqueue.scala 134:29 194:37]
  wire [38:0] _GEN_11603 = 4'h0 < realFlowNum_0 ? _GEN_7377 : flow_entry_0_17_vaddr; // @[Vlflowqueue.scala 134:29 194:37]
  wire [38:0] _GEN_11604 = 4'h0 < realFlowNum_0 ? _GEN_7378 : flow_entry_0_18_vaddr; // @[Vlflowqueue.scala 134:29 194:37]
  wire [38:0] _GEN_11605 = 4'h0 < realFlowNum_0 ? _GEN_7379 : flow_entry_0_19_vaddr; // @[Vlflowqueue.scala 134:29 194:37]
  wire [38:0] _GEN_11606 = 4'h0 < realFlowNum_0 ? _GEN_7380 : flow_entry_0_20_vaddr; // @[Vlflowqueue.scala 134:29 194:37]
  wire [38:0] _GEN_11607 = 4'h0 < realFlowNum_0 ? _GEN_7381 : flow_entry_0_21_vaddr; // @[Vlflowqueue.scala 134:29 194:37]
  wire [38:0] _GEN_11608 = 4'h0 < realFlowNum_0 ? _GEN_7382 : flow_entry_0_22_vaddr; // @[Vlflowqueue.scala 134:29 194:37]
  wire [38:0] _GEN_11609 = 4'h0 < realFlowNum_0 ? _GEN_7383 : flow_entry_0_23_vaddr; // @[Vlflowqueue.scala 134:29 194:37]
  wire [38:0] _GEN_11610 = 4'h0 < realFlowNum_0 ? _GEN_7384 : flow_entry_0_24_vaddr; // @[Vlflowqueue.scala 134:29 194:37]
  wire [38:0] _GEN_11611 = 4'h0 < realFlowNum_0 ? _GEN_7385 : flow_entry_0_25_vaddr; // @[Vlflowqueue.scala 134:29 194:37]
  wire [38:0] _GEN_11612 = 4'h0 < realFlowNum_0 ? _GEN_7386 : flow_entry_0_26_vaddr; // @[Vlflowqueue.scala 134:29 194:37]
  wire [38:0] _GEN_11613 = 4'h0 < realFlowNum_0 ? _GEN_7387 : flow_entry_0_27_vaddr; // @[Vlflowqueue.scala 134:29 194:37]
  wire [38:0] _GEN_11614 = 4'h0 < realFlowNum_0 ? _GEN_7388 : flow_entry_0_28_vaddr; // @[Vlflowqueue.scala 134:29 194:37]
  wire [38:0] _GEN_11615 = 4'h0 < realFlowNum_0 ? _GEN_7389 : flow_entry_0_29_vaddr; // @[Vlflowqueue.scala 134:29 194:37]
  wire [38:0] _GEN_11616 = 4'h0 < realFlowNum_0 ? _GEN_7390 : flow_entry_0_30_vaddr; // @[Vlflowqueue.scala 134:29 194:37]
  wire [38:0] _GEN_11617 = 4'h0 < realFlowNum_0 ? _GEN_7391 : flow_entry_0_31_vaddr; // @[Vlflowqueue.scala 134:29 194:37]
  wire  _GEN_11874 = _GEN_161423 | _GEN_8033; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_11875 = _GEN_161424 | _GEN_8034; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_11876 = _GEN_161425 | _GEN_8035; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_11877 = _GEN_161426 | _GEN_8036; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_11878 = _GEN_161427 | _GEN_8037; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_11879 = _GEN_161428 | _GEN_8038; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_11880 = _GEN_161429 | _GEN_8039; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_11881 = _GEN_161430 | _GEN_8040; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_11882 = _GEN_161431 | _GEN_8041; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_11883 = _GEN_161432 | _GEN_8042; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_11884 = _GEN_161433 | _GEN_8043; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_11885 = _GEN_161434 | _GEN_8044; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_11886 = _GEN_161435 | _GEN_8045; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_11887 = _GEN_161436 | _GEN_8046; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_11888 = _GEN_161437 | _GEN_8047; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_11889 = _GEN_161438 | _GEN_8048; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_11890 = _GEN_161439 | _GEN_8049; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_11891 = _GEN_161440 | _GEN_8050; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_11892 = _GEN_161441 | _GEN_8051; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_11893 = _GEN_161442 | _GEN_8052; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_11894 = _GEN_161443 | _GEN_8053; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_11895 = _GEN_161444 | _GEN_8054; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_11896 = _GEN_161445 | _GEN_8055; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_11897 = _GEN_161446 | _GEN_8056; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_11898 = _GEN_161447 | _GEN_8057; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_11899 = _GEN_161448 | _GEN_8058; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_11900 = _GEN_161449 | _GEN_8059; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_11901 = _GEN_161450 | _GEN_8060; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_11902 = _GEN_161451 | _GEN_8061; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_11903 = _GEN_161452 | _GEN_8062; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_11904 = _GEN_161453 | _GEN_8063; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_11905 = _GEN_161454 | _GEN_8064; // @[Vlflowqueue.scala 197:{51,51}]
  wire [4:0] _GEN_14850 = 5'h0 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_11009; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_14851 = 5'h1 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_11010; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_14852 = 5'h2 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_11011; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_14853 = 5'h3 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_11012; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_14854 = 5'h4 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_11013; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_14855 = 5'h5 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_11014; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_14856 = 5'h6 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_11015; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_14857 = 5'h7 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_11016; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_14858 = 5'h8 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_11017; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_14859 = 5'h9 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_11018; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_14860 = 5'ha == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_11019; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_14861 = 5'hb == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_11020; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_14862 = 5'hc == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_11021; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_14863 = 5'hd == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_11022; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_14864 = 5'he == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_11023; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_14865 = 5'hf == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_11024; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_14866 = 5'h10 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_11025; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_14867 = 5'h11 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_11026; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_14868 = 5'h12 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_11027; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_14869 = 5'h13 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_11028; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_14870 = 5'h14 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_11029; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_14871 = 5'h15 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_11030; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_14872 = 5'h16 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_11031; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_14873 = 5'h17 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_11032; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_14874 = 5'h18 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_11033; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_14875 = 5'h19 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_11034; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_14876 = 5'h1a == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_11035; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_14877 = 5'h1b == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_11036; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_14878 = 5'h1c == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_11037; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_14879 = 5'h1d == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_11038; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_14880 = 5'h1e == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_11039; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_14881 = 5'h1f == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_11040; // @[Vlflowqueue.scala 198:{51,51}]
  wire [38:0] _GEN_15426 = 5'h0 == index_0 ? vaddr_0 : _GEN_11586; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_15427 = 5'h1 == index_0 ? vaddr_0 : _GEN_11587; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_15428 = 5'h2 == index_0 ? vaddr_0 : _GEN_11588; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_15429 = 5'h3 == index_0 ? vaddr_0 : _GEN_11589; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_15430 = 5'h4 == index_0 ? vaddr_0 : _GEN_11590; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_15431 = 5'h5 == index_0 ? vaddr_0 : _GEN_11591; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_15432 = 5'h6 == index_0 ? vaddr_0 : _GEN_11592; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_15433 = 5'h7 == index_0 ? vaddr_0 : _GEN_11593; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_15434 = 5'h8 == index_0 ? vaddr_0 : _GEN_11594; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_15435 = 5'h9 == index_0 ? vaddr_0 : _GEN_11595; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_15436 = 5'ha == index_0 ? vaddr_0 : _GEN_11596; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_15437 = 5'hb == index_0 ? vaddr_0 : _GEN_11597; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_15438 = 5'hc == index_0 ? vaddr_0 : _GEN_11598; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_15439 = 5'hd == index_0 ? vaddr_0 : _GEN_11599; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_15440 = 5'he == index_0 ? vaddr_0 : _GEN_11600; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_15441 = 5'hf == index_0 ? vaddr_0 : _GEN_11601; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_15442 = 5'h10 == index_0 ? vaddr_0 : _GEN_11602; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_15443 = 5'h11 == index_0 ? vaddr_0 : _GEN_11603; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_15444 = 5'h12 == index_0 ? vaddr_0 : _GEN_11604; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_15445 = 5'h13 == index_0 ? vaddr_0 : _GEN_11605; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_15446 = 5'h14 == index_0 ? vaddr_0 : _GEN_11606; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_15447 = 5'h15 == index_0 ? vaddr_0 : _GEN_11607; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_15448 = 5'h16 == index_0 ? vaddr_0 : _GEN_11608; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_15449 = 5'h17 == index_0 ? vaddr_0 : _GEN_11609; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_15450 = 5'h18 == index_0 ? vaddr_0 : _GEN_11610; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_15451 = 5'h19 == index_0 ? vaddr_0 : _GEN_11611; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_15452 = 5'h1a == index_0 ? vaddr_0 : _GEN_11612; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_15453 = 5'h1b == index_0 ? vaddr_0 : _GEN_11613; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_15454 = 5'h1c == index_0 ? vaddr_0 : _GEN_11614; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_15455 = 5'h1d == index_0 ? vaddr_0 : _GEN_11615; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_15456 = 5'h1e == index_0 ? vaddr_0 : _GEN_11616; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_15457 = 5'h1f == index_0 ? vaddr_0 : _GEN_11617; // @[Vlflowqueue.scala 203:{51,51}]
  wire  _GEN_16099 = 4'h1 < realFlowNum_0 ? _GEN_11874 : _GEN_8033; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_16100 = 4'h1 < realFlowNum_0 ? _GEN_11875 : _GEN_8034; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_16101 = 4'h1 < realFlowNum_0 ? _GEN_11876 : _GEN_8035; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_16102 = 4'h1 < realFlowNum_0 ? _GEN_11877 : _GEN_8036; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_16103 = 4'h1 < realFlowNum_0 ? _GEN_11878 : _GEN_8037; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_16104 = 4'h1 < realFlowNum_0 ? _GEN_11879 : _GEN_8038; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_16105 = 4'h1 < realFlowNum_0 ? _GEN_11880 : _GEN_8039; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_16106 = 4'h1 < realFlowNum_0 ? _GEN_11881 : _GEN_8040; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_16107 = 4'h1 < realFlowNum_0 ? _GEN_11882 : _GEN_8041; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_16108 = 4'h1 < realFlowNum_0 ? _GEN_11883 : _GEN_8042; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_16109 = 4'h1 < realFlowNum_0 ? _GEN_11884 : _GEN_8043; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_16110 = 4'h1 < realFlowNum_0 ? _GEN_11885 : _GEN_8044; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_16111 = 4'h1 < realFlowNum_0 ? _GEN_11886 : _GEN_8045; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_16112 = 4'h1 < realFlowNum_0 ? _GEN_11887 : _GEN_8046; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_16113 = 4'h1 < realFlowNum_0 ? _GEN_11888 : _GEN_8047; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_16114 = 4'h1 < realFlowNum_0 ? _GEN_11889 : _GEN_8048; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_16115 = 4'h1 < realFlowNum_0 ? _GEN_11890 : _GEN_8049; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_16116 = 4'h1 < realFlowNum_0 ? _GEN_11891 : _GEN_8050; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_16117 = 4'h1 < realFlowNum_0 ? _GEN_11892 : _GEN_8051; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_16118 = 4'h1 < realFlowNum_0 ? _GEN_11893 : _GEN_8052; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_16119 = 4'h1 < realFlowNum_0 ? _GEN_11894 : _GEN_8053; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_16120 = 4'h1 < realFlowNum_0 ? _GEN_11895 : _GEN_8054; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_16121 = 4'h1 < realFlowNum_0 ? _GEN_11896 : _GEN_8055; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_16122 = 4'h1 < realFlowNum_0 ? _GEN_11897 : _GEN_8056; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_16123 = 4'h1 < realFlowNum_0 ? _GEN_11898 : _GEN_8057; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_16124 = 4'h1 < realFlowNum_0 ? _GEN_11899 : _GEN_8058; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_16125 = 4'h1 < realFlowNum_0 ? _GEN_11900 : _GEN_8059; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_16126 = 4'h1 < realFlowNum_0 ? _GEN_11901 : _GEN_8060; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_16127 = 4'h1 < realFlowNum_0 ? _GEN_11902 : _GEN_8061; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_16128 = 4'h1 < realFlowNum_0 ? _GEN_11903 : _GEN_8062; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_16129 = 4'h1 < realFlowNum_0 ? _GEN_11904 : _GEN_8063; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_16130 = 4'h1 < realFlowNum_0 ? _GEN_11905 : _GEN_8064; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_19075 = 4'h1 < realFlowNum_0 ? _GEN_14850 : _GEN_11009; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_19076 = 4'h1 < realFlowNum_0 ? _GEN_14851 : _GEN_11010; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_19077 = 4'h1 < realFlowNum_0 ? _GEN_14852 : _GEN_11011; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_19078 = 4'h1 < realFlowNum_0 ? _GEN_14853 : _GEN_11012; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_19079 = 4'h1 < realFlowNum_0 ? _GEN_14854 : _GEN_11013; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_19080 = 4'h1 < realFlowNum_0 ? _GEN_14855 : _GEN_11014; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_19081 = 4'h1 < realFlowNum_0 ? _GEN_14856 : _GEN_11015; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_19082 = 4'h1 < realFlowNum_0 ? _GEN_14857 : _GEN_11016; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_19083 = 4'h1 < realFlowNum_0 ? _GEN_14858 : _GEN_11017; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_19084 = 4'h1 < realFlowNum_0 ? _GEN_14859 : _GEN_11018; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_19085 = 4'h1 < realFlowNum_0 ? _GEN_14860 : _GEN_11019; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_19086 = 4'h1 < realFlowNum_0 ? _GEN_14861 : _GEN_11020; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_19087 = 4'h1 < realFlowNum_0 ? _GEN_14862 : _GEN_11021; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_19088 = 4'h1 < realFlowNum_0 ? _GEN_14863 : _GEN_11022; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_19089 = 4'h1 < realFlowNum_0 ? _GEN_14864 : _GEN_11023; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_19090 = 4'h1 < realFlowNum_0 ? _GEN_14865 : _GEN_11024; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_19091 = 4'h1 < realFlowNum_0 ? _GEN_14866 : _GEN_11025; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_19092 = 4'h1 < realFlowNum_0 ? _GEN_14867 : _GEN_11026; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_19093 = 4'h1 < realFlowNum_0 ? _GEN_14868 : _GEN_11027; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_19094 = 4'h1 < realFlowNum_0 ? _GEN_14869 : _GEN_11028; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_19095 = 4'h1 < realFlowNum_0 ? _GEN_14870 : _GEN_11029; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_19096 = 4'h1 < realFlowNum_0 ? _GEN_14871 : _GEN_11030; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_19097 = 4'h1 < realFlowNum_0 ? _GEN_14872 : _GEN_11031; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_19098 = 4'h1 < realFlowNum_0 ? _GEN_14873 : _GEN_11032; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_19099 = 4'h1 < realFlowNum_0 ? _GEN_14874 : _GEN_11033; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_19100 = 4'h1 < realFlowNum_0 ? _GEN_14875 : _GEN_11034; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_19101 = 4'h1 < realFlowNum_0 ? _GEN_14876 : _GEN_11035; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_19102 = 4'h1 < realFlowNum_0 ? _GEN_14877 : _GEN_11036; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_19103 = 4'h1 < realFlowNum_0 ? _GEN_14878 : _GEN_11037; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_19104 = 4'h1 < realFlowNum_0 ? _GEN_14879 : _GEN_11038; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_19105 = 4'h1 < realFlowNum_0 ? _GEN_14880 : _GEN_11039; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_19106 = 4'h1 < realFlowNum_0 ? _GEN_14881 : _GEN_11040; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_19652 = 4'h1 < realFlowNum_0 ? _GEN_15426 : _GEN_11586; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_19653 = 4'h1 < realFlowNum_0 ? _GEN_15427 : _GEN_11587; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_19654 = 4'h1 < realFlowNum_0 ? _GEN_15428 : _GEN_11588; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_19655 = 4'h1 < realFlowNum_0 ? _GEN_15429 : _GEN_11589; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_19656 = 4'h1 < realFlowNum_0 ? _GEN_15430 : _GEN_11590; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_19657 = 4'h1 < realFlowNum_0 ? _GEN_15431 : _GEN_11591; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_19658 = 4'h1 < realFlowNum_0 ? _GEN_15432 : _GEN_11592; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_19659 = 4'h1 < realFlowNum_0 ? _GEN_15433 : _GEN_11593; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_19660 = 4'h1 < realFlowNum_0 ? _GEN_15434 : _GEN_11594; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_19661 = 4'h1 < realFlowNum_0 ? _GEN_15435 : _GEN_11595; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_19662 = 4'h1 < realFlowNum_0 ? _GEN_15436 : _GEN_11596; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_19663 = 4'h1 < realFlowNum_0 ? _GEN_15437 : _GEN_11597; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_19664 = 4'h1 < realFlowNum_0 ? _GEN_15438 : _GEN_11598; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_19665 = 4'h1 < realFlowNum_0 ? _GEN_15439 : _GEN_11599; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_19666 = 4'h1 < realFlowNum_0 ? _GEN_15440 : _GEN_11600; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_19667 = 4'h1 < realFlowNum_0 ? _GEN_15441 : _GEN_11601; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_19668 = 4'h1 < realFlowNum_0 ? _GEN_15442 : _GEN_11602; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_19669 = 4'h1 < realFlowNum_0 ? _GEN_15443 : _GEN_11603; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_19670 = 4'h1 < realFlowNum_0 ? _GEN_15444 : _GEN_11604; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_19671 = 4'h1 < realFlowNum_0 ? _GEN_15445 : _GEN_11605; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_19672 = 4'h1 < realFlowNum_0 ? _GEN_15446 : _GEN_11606; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_19673 = 4'h1 < realFlowNum_0 ? _GEN_15447 : _GEN_11607; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_19674 = 4'h1 < realFlowNum_0 ? _GEN_15448 : _GEN_11608; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_19675 = 4'h1 < realFlowNum_0 ? _GEN_15449 : _GEN_11609; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_19676 = 4'h1 < realFlowNum_0 ? _GEN_15450 : _GEN_11610; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_19677 = 4'h1 < realFlowNum_0 ? _GEN_15451 : _GEN_11611; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_19678 = 4'h1 < realFlowNum_0 ? _GEN_15452 : _GEN_11612; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_19679 = 4'h1 < realFlowNum_0 ? _GEN_15453 : _GEN_11613; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_19680 = 4'h1 < realFlowNum_0 ? _GEN_15454 : _GEN_11614; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_19681 = 4'h1 < realFlowNum_0 ? _GEN_15455 : _GEN_11615; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_19682 = 4'h1 < realFlowNum_0 ? _GEN_15456 : _GEN_11616; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_19683 = 4'h1 < realFlowNum_0 ? _GEN_15457 : _GEN_11617; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_19940 = _GEN_161423 | _GEN_16099; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_19941 = _GEN_161424 | _GEN_16100; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_19942 = _GEN_161425 | _GEN_16101; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_19943 = _GEN_161426 | _GEN_16102; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_19944 = _GEN_161427 | _GEN_16103; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_19945 = _GEN_161428 | _GEN_16104; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_19946 = _GEN_161429 | _GEN_16105; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_19947 = _GEN_161430 | _GEN_16106; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_19948 = _GEN_161431 | _GEN_16107; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_19949 = _GEN_161432 | _GEN_16108; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_19950 = _GEN_161433 | _GEN_16109; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_19951 = _GEN_161434 | _GEN_16110; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_19952 = _GEN_161435 | _GEN_16111; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_19953 = _GEN_161436 | _GEN_16112; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_19954 = _GEN_161437 | _GEN_16113; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_19955 = _GEN_161438 | _GEN_16114; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_19956 = _GEN_161439 | _GEN_16115; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_19957 = _GEN_161440 | _GEN_16116; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_19958 = _GEN_161441 | _GEN_16117; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_19959 = _GEN_161442 | _GEN_16118; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_19960 = _GEN_161443 | _GEN_16119; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_19961 = _GEN_161444 | _GEN_16120; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_19962 = _GEN_161445 | _GEN_16121; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_19963 = _GEN_161446 | _GEN_16122; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_19964 = _GEN_161447 | _GEN_16123; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_19965 = _GEN_161448 | _GEN_16124; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_19966 = _GEN_161449 | _GEN_16125; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_19967 = _GEN_161450 | _GEN_16126; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_19968 = _GEN_161451 | _GEN_16127; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_19969 = _GEN_161452 | _GEN_16128; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_19970 = _GEN_161453 | _GEN_16129; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_19971 = _GEN_161454 | _GEN_16130; // @[Vlflowqueue.scala 197:{51,51}]
  wire [4:0] _GEN_22916 = 5'h0 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_19075; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_22917 = 5'h1 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_19076; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_22918 = 5'h2 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_19077; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_22919 = 5'h3 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_19078; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_22920 = 5'h4 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_19079; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_22921 = 5'h5 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_19080; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_22922 = 5'h6 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_19081; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_22923 = 5'h7 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_19082; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_22924 = 5'h8 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_19083; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_22925 = 5'h9 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_19084; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_22926 = 5'ha == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_19085; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_22927 = 5'hb == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_19086; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_22928 = 5'hc == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_19087; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_22929 = 5'hd == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_19088; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_22930 = 5'he == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_19089; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_22931 = 5'hf == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_19090; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_22932 = 5'h10 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_19091; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_22933 = 5'h11 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_19092; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_22934 = 5'h12 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_19093; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_22935 = 5'h13 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_19094; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_22936 = 5'h14 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_19095; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_22937 = 5'h15 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_19096; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_22938 = 5'h16 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_19097; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_22939 = 5'h17 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_19098; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_22940 = 5'h18 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_19099; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_22941 = 5'h19 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_19100; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_22942 = 5'h1a == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_19101; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_22943 = 5'h1b == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_19102; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_22944 = 5'h1c == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_19103; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_22945 = 5'h1d == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_19104; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_22946 = 5'h1e == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_19105; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_22947 = 5'h1f == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_19106; // @[Vlflowqueue.scala 198:{51,51}]
  wire [38:0] _GEN_23492 = 5'h0 == index_0 ? vaddr_0 : _GEN_19652; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_23493 = 5'h1 == index_0 ? vaddr_0 : _GEN_19653; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_23494 = 5'h2 == index_0 ? vaddr_0 : _GEN_19654; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_23495 = 5'h3 == index_0 ? vaddr_0 : _GEN_19655; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_23496 = 5'h4 == index_0 ? vaddr_0 : _GEN_19656; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_23497 = 5'h5 == index_0 ? vaddr_0 : _GEN_19657; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_23498 = 5'h6 == index_0 ? vaddr_0 : _GEN_19658; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_23499 = 5'h7 == index_0 ? vaddr_0 : _GEN_19659; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_23500 = 5'h8 == index_0 ? vaddr_0 : _GEN_19660; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_23501 = 5'h9 == index_0 ? vaddr_0 : _GEN_19661; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_23502 = 5'ha == index_0 ? vaddr_0 : _GEN_19662; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_23503 = 5'hb == index_0 ? vaddr_0 : _GEN_19663; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_23504 = 5'hc == index_0 ? vaddr_0 : _GEN_19664; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_23505 = 5'hd == index_0 ? vaddr_0 : _GEN_19665; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_23506 = 5'he == index_0 ? vaddr_0 : _GEN_19666; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_23507 = 5'hf == index_0 ? vaddr_0 : _GEN_19667; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_23508 = 5'h10 == index_0 ? vaddr_0 : _GEN_19668; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_23509 = 5'h11 == index_0 ? vaddr_0 : _GEN_19669; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_23510 = 5'h12 == index_0 ? vaddr_0 : _GEN_19670; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_23511 = 5'h13 == index_0 ? vaddr_0 : _GEN_19671; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_23512 = 5'h14 == index_0 ? vaddr_0 : _GEN_19672; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_23513 = 5'h15 == index_0 ? vaddr_0 : _GEN_19673; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_23514 = 5'h16 == index_0 ? vaddr_0 : _GEN_19674; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_23515 = 5'h17 == index_0 ? vaddr_0 : _GEN_19675; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_23516 = 5'h18 == index_0 ? vaddr_0 : _GEN_19676; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_23517 = 5'h19 == index_0 ? vaddr_0 : _GEN_19677; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_23518 = 5'h1a == index_0 ? vaddr_0 : _GEN_19678; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_23519 = 5'h1b == index_0 ? vaddr_0 : _GEN_19679; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_23520 = 5'h1c == index_0 ? vaddr_0 : _GEN_19680; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_23521 = 5'h1d == index_0 ? vaddr_0 : _GEN_19681; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_23522 = 5'h1e == index_0 ? vaddr_0 : _GEN_19682; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_23523 = 5'h1f == index_0 ? vaddr_0 : _GEN_19683; // @[Vlflowqueue.scala 203:{51,51}]
  wire  _GEN_24165 = 4'h2 < realFlowNum_0 ? _GEN_19940 : _GEN_16099; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_24166 = 4'h2 < realFlowNum_0 ? _GEN_19941 : _GEN_16100; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_24167 = 4'h2 < realFlowNum_0 ? _GEN_19942 : _GEN_16101; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_24168 = 4'h2 < realFlowNum_0 ? _GEN_19943 : _GEN_16102; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_24169 = 4'h2 < realFlowNum_0 ? _GEN_19944 : _GEN_16103; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_24170 = 4'h2 < realFlowNum_0 ? _GEN_19945 : _GEN_16104; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_24171 = 4'h2 < realFlowNum_0 ? _GEN_19946 : _GEN_16105; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_24172 = 4'h2 < realFlowNum_0 ? _GEN_19947 : _GEN_16106; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_24173 = 4'h2 < realFlowNum_0 ? _GEN_19948 : _GEN_16107; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_24174 = 4'h2 < realFlowNum_0 ? _GEN_19949 : _GEN_16108; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_24175 = 4'h2 < realFlowNum_0 ? _GEN_19950 : _GEN_16109; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_24176 = 4'h2 < realFlowNum_0 ? _GEN_19951 : _GEN_16110; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_24177 = 4'h2 < realFlowNum_0 ? _GEN_19952 : _GEN_16111; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_24178 = 4'h2 < realFlowNum_0 ? _GEN_19953 : _GEN_16112; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_24179 = 4'h2 < realFlowNum_0 ? _GEN_19954 : _GEN_16113; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_24180 = 4'h2 < realFlowNum_0 ? _GEN_19955 : _GEN_16114; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_24181 = 4'h2 < realFlowNum_0 ? _GEN_19956 : _GEN_16115; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_24182 = 4'h2 < realFlowNum_0 ? _GEN_19957 : _GEN_16116; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_24183 = 4'h2 < realFlowNum_0 ? _GEN_19958 : _GEN_16117; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_24184 = 4'h2 < realFlowNum_0 ? _GEN_19959 : _GEN_16118; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_24185 = 4'h2 < realFlowNum_0 ? _GEN_19960 : _GEN_16119; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_24186 = 4'h2 < realFlowNum_0 ? _GEN_19961 : _GEN_16120; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_24187 = 4'h2 < realFlowNum_0 ? _GEN_19962 : _GEN_16121; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_24188 = 4'h2 < realFlowNum_0 ? _GEN_19963 : _GEN_16122; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_24189 = 4'h2 < realFlowNum_0 ? _GEN_19964 : _GEN_16123; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_24190 = 4'h2 < realFlowNum_0 ? _GEN_19965 : _GEN_16124; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_24191 = 4'h2 < realFlowNum_0 ? _GEN_19966 : _GEN_16125; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_24192 = 4'h2 < realFlowNum_0 ? _GEN_19967 : _GEN_16126; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_24193 = 4'h2 < realFlowNum_0 ? _GEN_19968 : _GEN_16127; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_24194 = 4'h2 < realFlowNum_0 ? _GEN_19969 : _GEN_16128; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_24195 = 4'h2 < realFlowNum_0 ? _GEN_19970 : _GEN_16129; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_24196 = 4'h2 < realFlowNum_0 ? _GEN_19971 : _GEN_16130; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_27141 = 4'h2 < realFlowNum_0 ? _GEN_22916 : _GEN_19075; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_27142 = 4'h2 < realFlowNum_0 ? _GEN_22917 : _GEN_19076; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_27143 = 4'h2 < realFlowNum_0 ? _GEN_22918 : _GEN_19077; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_27144 = 4'h2 < realFlowNum_0 ? _GEN_22919 : _GEN_19078; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_27145 = 4'h2 < realFlowNum_0 ? _GEN_22920 : _GEN_19079; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_27146 = 4'h2 < realFlowNum_0 ? _GEN_22921 : _GEN_19080; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_27147 = 4'h2 < realFlowNum_0 ? _GEN_22922 : _GEN_19081; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_27148 = 4'h2 < realFlowNum_0 ? _GEN_22923 : _GEN_19082; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_27149 = 4'h2 < realFlowNum_0 ? _GEN_22924 : _GEN_19083; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_27150 = 4'h2 < realFlowNum_0 ? _GEN_22925 : _GEN_19084; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_27151 = 4'h2 < realFlowNum_0 ? _GEN_22926 : _GEN_19085; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_27152 = 4'h2 < realFlowNum_0 ? _GEN_22927 : _GEN_19086; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_27153 = 4'h2 < realFlowNum_0 ? _GEN_22928 : _GEN_19087; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_27154 = 4'h2 < realFlowNum_0 ? _GEN_22929 : _GEN_19088; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_27155 = 4'h2 < realFlowNum_0 ? _GEN_22930 : _GEN_19089; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_27156 = 4'h2 < realFlowNum_0 ? _GEN_22931 : _GEN_19090; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_27157 = 4'h2 < realFlowNum_0 ? _GEN_22932 : _GEN_19091; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_27158 = 4'h2 < realFlowNum_0 ? _GEN_22933 : _GEN_19092; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_27159 = 4'h2 < realFlowNum_0 ? _GEN_22934 : _GEN_19093; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_27160 = 4'h2 < realFlowNum_0 ? _GEN_22935 : _GEN_19094; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_27161 = 4'h2 < realFlowNum_0 ? _GEN_22936 : _GEN_19095; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_27162 = 4'h2 < realFlowNum_0 ? _GEN_22937 : _GEN_19096; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_27163 = 4'h2 < realFlowNum_0 ? _GEN_22938 : _GEN_19097; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_27164 = 4'h2 < realFlowNum_0 ? _GEN_22939 : _GEN_19098; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_27165 = 4'h2 < realFlowNum_0 ? _GEN_22940 : _GEN_19099; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_27166 = 4'h2 < realFlowNum_0 ? _GEN_22941 : _GEN_19100; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_27167 = 4'h2 < realFlowNum_0 ? _GEN_22942 : _GEN_19101; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_27168 = 4'h2 < realFlowNum_0 ? _GEN_22943 : _GEN_19102; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_27169 = 4'h2 < realFlowNum_0 ? _GEN_22944 : _GEN_19103; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_27170 = 4'h2 < realFlowNum_0 ? _GEN_22945 : _GEN_19104; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_27171 = 4'h2 < realFlowNum_0 ? _GEN_22946 : _GEN_19105; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_27172 = 4'h2 < realFlowNum_0 ? _GEN_22947 : _GEN_19106; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_27718 = 4'h2 < realFlowNum_0 ? _GEN_23492 : _GEN_19652; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_27719 = 4'h2 < realFlowNum_0 ? _GEN_23493 : _GEN_19653; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_27720 = 4'h2 < realFlowNum_0 ? _GEN_23494 : _GEN_19654; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_27721 = 4'h2 < realFlowNum_0 ? _GEN_23495 : _GEN_19655; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_27722 = 4'h2 < realFlowNum_0 ? _GEN_23496 : _GEN_19656; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_27723 = 4'h2 < realFlowNum_0 ? _GEN_23497 : _GEN_19657; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_27724 = 4'h2 < realFlowNum_0 ? _GEN_23498 : _GEN_19658; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_27725 = 4'h2 < realFlowNum_0 ? _GEN_23499 : _GEN_19659; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_27726 = 4'h2 < realFlowNum_0 ? _GEN_23500 : _GEN_19660; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_27727 = 4'h2 < realFlowNum_0 ? _GEN_23501 : _GEN_19661; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_27728 = 4'h2 < realFlowNum_0 ? _GEN_23502 : _GEN_19662; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_27729 = 4'h2 < realFlowNum_0 ? _GEN_23503 : _GEN_19663; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_27730 = 4'h2 < realFlowNum_0 ? _GEN_23504 : _GEN_19664; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_27731 = 4'h2 < realFlowNum_0 ? _GEN_23505 : _GEN_19665; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_27732 = 4'h2 < realFlowNum_0 ? _GEN_23506 : _GEN_19666; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_27733 = 4'h2 < realFlowNum_0 ? _GEN_23507 : _GEN_19667; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_27734 = 4'h2 < realFlowNum_0 ? _GEN_23508 : _GEN_19668; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_27735 = 4'h2 < realFlowNum_0 ? _GEN_23509 : _GEN_19669; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_27736 = 4'h2 < realFlowNum_0 ? _GEN_23510 : _GEN_19670; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_27737 = 4'h2 < realFlowNum_0 ? _GEN_23511 : _GEN_19671; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_27738 = 4'h2 < realFlowNum_0 ? _GEN_23512 : _GEN_19672; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_27739 = 4'h2 < realFlowNum_0 ? _GEN_23513 : _GEN_19673; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_27740 = 4'h2 < realFlowNum_0 ? _GEN_23514 : _GEN_19674; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_27741 = 4'h2 < realFlowNum_0 ? _GEN_23515 : _GEN_19675; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_27742 = 4'h2 < realFlowNum_0 ? _GEN_23516 : _GEN_19676; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_27743 = 4'h2 < realFlowNum_0 ? _GEN_23517 : _GEN_19677; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_27744 = 4'h2 < realFlowNum_0 ? _GEN_23518 : _GEN_19678; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_27745 = 4'h2 < realFlowNum_0 ? _GEN_23519 : _GEN_19679; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_27746 = 4'h2 < realFlowNum_0 ? _GEN_23520 : _GEN_19680; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_27747 = 4'h2 < realFlowNum_0 ? _GEN_23521 : _GEN_19681; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_27748 = 4'h2 < realFlowNum_0 ? _GEN_23522 : _GEN_19682; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_27749 = 4'h2 < realFlowNum_0 ? _GEN_23523 : _GEN_19683; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_28006 = _GEN_161423 | _GEN_24165; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_28007 = _GEN_161424 | _GEN_24166; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_28008 = _GEN_161425 | _GEN_24167; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_28009 = _GEN_161426 | _GEN_24168; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_28010 = _GEN_161427 | _GEN_24169; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_28011 = _GEN_161428 | _GEN_24170; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_28012 = _GEN_161429 | _GEN_24171; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_28013 = _GEN_161430 | _GEN_24172; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_28014 = _GEN_161431 | _GEN_24173; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_28015 = _GEN_161432 | _GEN_24174; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_28016 = _GEN_161433 | _GEN_24175; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_28017 = _GEN_161434 | _GEN_24176; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_28018 = _GEN_161435 | _GEN_24177; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_28019 = _GEN_161436 | _GEN_24178; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_28020 = _GEN_161437 | _GEN_24179; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_28021 = _GEN_161438 | _GEN_24180; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_28022 = _GEN_161439 | _GEN_24181; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_28023 = _GEN_161440 | _GEN_24182; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_28024 = _GEN_161441 | _GEN_24183; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_28025 = _GEN_161442 | _GEN_24184; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_28026 = _GEN_161443 | _GEN_24185; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_28027 = _GEN_161444 | _GEN_24186; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_28028 = _GEN_161445 | _GEN_24187; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_28029 = _GEN_161446 | _GEN_24188; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_28030 = _GEN_161447 | _GEN_24189; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_28031 = _GEN_161448 | _GEN_24190; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_28032 = _GEN_161449 | _GEN_24191; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_28033 = _GEN_161450 | _GEN_24192; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_28034 = _GEN_161451 | _GEN_24193; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_28035 = _GEN_161452 | _GEN_24194; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_28036 = _GEN_161453 | _GEN_24195; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_28037 = _GEN_161454 | _GEN_24196; // @[Vlflowqueue.scala 197:{51,51}]
  wire [4:0] _GEN_30982 = 5'h0 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_27141; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_30983 = 5'h1 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_27142; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_30984 = 5'h2 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_27143; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_30985 = 5'h3 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_27144; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_30986 = 5'h4 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_27145; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_30987 = 5'h5 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_27146; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_30988 = 5'h6 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_27147; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_30989 = 5'h7 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_27148; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_30990 = 5'h8 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_27149; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_30991 = 5'h9 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_27150; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_30992 = 5'ha == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_27151; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_30993 = 5'hb == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_27152; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_30994 = 5'hc == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_27153; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_30995 = 5'hd == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_27154; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_30996 = 5'he == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_27155; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_30997 = 5'hf == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_27156; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_30998 = 5'h10 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_27157; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_30999 = 5'h11 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_27158; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_31000 = 5'h12 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_27159; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_31001 = 5'h13 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_27160; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_31002 = 5'h14 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_27161; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_31003 = 5'h15 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_27162; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_31004 = 5'h16 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_27163; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_31005 = 5'h17 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_27164; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_31006 = 5'h18 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_27165; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_31007 = 5'h19 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_27166; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_31008 = 5'h1a == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_27167; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_31009 = 5'h1b == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_27168; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_31010 = 5'h1c == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_27169; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_31011 = 5'h1d == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_27170; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_31012 = 5'h1e == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_27171; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_31013 = 5'h1f == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_27172; // @[Vlflowqueue.scala 198:{51,51}]
  wire [38:0] _GEN_31558 = 5'h0 == index_0 ? vaddr_0 : _GEN_27718; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_31559 = 5'h1 == index_0 ? vaddr_0 : _GEN_27719; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_31560 = 5'h2 == index_0 ? vaddr_0 : _GEN_27720; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_31561 = 5'h3 == index_0 ? vaddr_0 : _GEN_27721; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_31562 = 5'h4 == index_0 ? vaddr_0 : _GEN_27722; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_31563 = 5'h5 == index_0 ? vaddr_0 : _GEN_27723; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_31564 = 5'h6 == index_0 ? vaddr_0 : _GEN_27724; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_31565 = 5'h7 == index_0 ? vaddr_0 : _GEN_27725; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_31566 = 5'h8 == index_0 ? vaddr_0 : _GEN_27726; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_31567 = 5'h9 == index_0 ? vaddr_0 : _GEN_27727; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_31568 = 5'ha == index_0 ? vaddr_0 : _GEN_27728; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_31569 = 5'hb == index_0 ? vaddr_0 : _GEN_27729; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_31570 = 5'hc == index_0 ? vaddr_0 : _GEN_27730; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_31571 = 5'hd == index_0 ? vaddr_0 : _GEN_27731; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_31572 = 5'he == index_0 ? vaddr_0 : _GEN_27732; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_31573 = 5'hf == index_0 ? vaddr_0 : _GEN_27733; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_31574 = 5'h10 == index_0 ? vaddr_0 : _GEN_27734; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_31575 = 5'h11 == index_0 ? vaddr_0 : _GEN_27735; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_31576 = 5'h12 == index_0 ? vaddr_0 : _GEN_27736; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_31577 = 5'h13 == index_0 ? vaddr_0 : _GEN_27737; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_31578 = 5'h14 == index_0 ? vaddr_0 : _GEN_27738; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_31579 = 5'h15 == index_0 ? vaddr_0 : _GEN_27739; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_31580 = 5'h16 == index_0 ? vaddr_0 : _GEN_27740; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_31581 = 5'h17 == index_0 ? vaddr_0 : _GEN_27741; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_31582 = 5'h18 == index_0 ? vaddr_0 : _GEN_27742; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_31583 = 5'h19 == index_0 ? vaddr_0 : _GEN_27743; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_31584 = 5'h1a == index_0 ? vaddr_0 : _GEN_27744; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_31585 = 5'h1b == index_0 ? vaddr_0 : _GEN_27745; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_31586 = 5'h1c == index_0 ? vaddr_0 : _GEN_27746; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_31587 = 5'h1d == index_0 ? vaddr_0 : _GEN_27747; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_31588 = 5'h1e == index_0 ? vaddr_0 : _GEN_27748; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_31589 = 5'h1f == index_0 ? vaddr_0 : _GEN_27749; // @[Vlflowqueue.scala 203:{51,51}]
  wire  _GEN_32231 = 4'h3 < realFlowNum_0 ? _GEN_28006 : _GEN_24165; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_32232 = 4'h3 < realFlowNum_0 ? _GEN_28007 : _GEN_24166; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_32233 = 4'h3 < realFlowNum_0 ? _GEN_28008 : _GEN_24167; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_32234 = 4'h3 < realFlowNum_0 ? _GEN_28009 : _GEN_24168; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_32235 = 4'h3 < realFlowNum_0 ? _GEN_28010 : _GEN_24169; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_32236 = 4'h3 < realFlowNum_0 ? _GEN_28011 : _GEN_24170; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_32237 = 4'h3 < realFlowNum_0 ? _GEN_28012 : _GEN_24171; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_32238 = 4'h3 < realFlowNum_0 ? _GEN_28013 : _GEN_24172; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_32239 = 4'h3 < realFlowNum_0 ? _GEN_28014 : _GEN_24173; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_32240 = 4'h3 < realFlowNum_0 ? _GEN_28015 : _GEN_24174; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_32241 = 4'h3 < realFlowNum_0 ? _GEN_28016 : _GEN_24175; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_32242 = 4'h3 < realFlowNum_0 ? _GEN_28017 : _GEN_24176; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_32243 = 4'h3 < realFlowNum_0 ? _GEN_28018 : _GEN_24177; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_32244 = 4'h3 < realFlowNum_0 ? _GEN_28019 : _GEN_24178; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_32245 = 4'h3 < realFlowNum_0 ? _GEN_28020 : _GEN_24179; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_32246 = 4'h3 < realFlowNum_0 ? _GEN_28021 : _GEN_24180; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_32247 = 4'h3 < realFlowNum_0 ? _GEN_28022 : _GEN_24181; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_32248 = 4'h3 < realFlowNum_0 ? _GEN_28023 : _GEN_24182; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_32249 = 4'h3 < realFlowNum_0 ? _GEN_28024 : _GEN_24183; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_32250 = 4'h3 < realFlowNum_0 ? _GEN_28025 : _GEN_24184; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_32251 = 4'h3 < realFlowNum_0 ? _GEN_28026 : _GEN_24185; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_32252 = 4'h3 < realFlowNum_0 ? _GEN_28027 : _GEN_24186; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_32253 = 4'h3 < realFlowNum_0 ? _GEN_28028 : _GEN_24187; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_32254 = 4'h3 < realFlowNum_0 ? _GEN_28029 : _GEN_24188; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_32255 = 4'h3 < realFlowNum_0 ? _GEN_28030 : _GEN_24189; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_32256 = 4'h3 < realFlowNum_0 ? _GEN_28031 : _GEN_24190; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_32257 = 4'h3 < realFlowNum_0 ? _GEN_28032 : _GEN_24191; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_32258 = 4'h3 < realFlowNum_0 ? _GEN_28033 : _GEN_24192; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_32259 = 4'h3 < realFlowNum_0 ? _GEN_28034 : _GEN_24193; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_32260 = 4'h3 < realFlowNum_0 ? _GEN_28035 : _GEN_24194; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_32261 = 4'h3 < realFlowNum_0 ? _GEN_28036 : _GEN_24195; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_32262 = 4'h3 < realFlowNum_0 ? _GEN_28037 : _GEN_24196; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_35207 = 4'h3 < realFlowNum_0 ? _GEN_30982 : _GEN_27141; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_35208 = 4'h3 < realFlowNum_0 ? _GEN_30983 : _GEN_27142; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_35209 = 4'h3 < realFlowNum_0 ? _GEN_30984 : _GEN_27143; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_35210 = 4'h3 < realFlowNum_0 ? _GEN_30985 : _GEN_27144; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_35211 = 4'h3 < realFlowNum_0 ? _GEN_30986 : _GEN_27145; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_35212 = 4'h3 < realFlowNum_0 ? _GEN_30987 : _GEN_27146; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_35213 = 4'h3 < realFlowNum_0 ? _GEN_30988 : _GEN_27147; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_35214 = 4'h3 < realFlowNum_0 ? _GEN_30989 : _GEN_27148; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_35215 = 4'h3 < realFlowNum_0 ? _GEN_30990 : _GEN_27149; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_35216 = 4'h3 < realFlowNum_0 ? _GEN_30991 : _GEN_27150; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_35217 = 4'h3 < realFlowNum_0 ? _GEN_30992 : _GEN_27151; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_35218 = 4'h3 < realFlowNum_0 ? _GEN_30993 : _GEN_27152; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_35219 = 4'h3 < realFlowNum_0 ? _GEN_30994 : _GEN_27153; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_35220 = 4'h3 < realFlowNum_0 ? _GEN_30995 : _GEN_27154; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_35221 = 4'h3 < realFlowNum_0 ? _GEN_30996 : _GEN_27155; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_35222 = 4'h3 < realFlowNum_0 ? _GEN_30997 : _GEN_27156; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_35223 = 4'h3 < realFlowNum_0 ? _GEN_30998 : _GEN_27157; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_35224 = 4'h3 < realFlowNum_0 ? _GEN_30999 : _GEN_27158; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_35225 = 4'h3 < realFlowNum_0 ? _GEN_31000 : _GEN_27159; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_35226 = 4'h3 < realFlowNum_0 ? _GEN_31001 : _GEN_27160; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_35227 = 4'h3 < realFlowNum_0 ? _GEN_31002 : _GEN_27161; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_35228 = 4'h3 < realFlowNum_0 ? _GEN_31003 : _GEN_27162; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_35229 = 4'h3 < realFlowNum_0 ? _GEN_31004 : _GEN_27163; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_35230 = 4'h3 < realFlowNum_0 ? _GEN_31005 : _GEN_27164; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_35231 = 4'h3 < realFlowNum_0 ? _GEN_31006 : _GEN_27165; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_35232 = 4'h3 < realFlowNum_0 ? _GEN_31007 : _GEN_27166; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_35233 = 4'h3 < realFlowNum_0 ? _GEN_31008 : _GEN_27167; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_35234 = 4'h3 < realFlowNum_0 ? _GEN_31009 : _GEN_27168; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_35235 = 4'h3 < realFlowNum_0 ? _GEN_31010 : _GEN_27169; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_35236 = 4'h3 < realFlowNum_0 ? _GEN_31011 : _GEN_27170; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_35237 = 4'h3 < realFlowNum_0 ? _GEN_31012 : _GEN_27171; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_35238 = 4'h3 < realFlowNum_0 ? _GEN_31013 : _GEN_27172; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_35784 = 4'h3 < realFlowNum_0 ? _GEN_31558 : _GEN_27718; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_35785 = 4'h3 < realFlowNum_0 ? _GEN_31559 : _GEN_27719; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_35786 = 4'h3 < realFlowNum_0 ? _GEN_31560 : _GEN_27720; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_35787 = 4'h3 < realFlowNum_0 ? _GEN_31561 : _GEN_27721; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_35788 = 4'h3 < realFlowNum_0 ? _GEN_31562 : _GEN_27722; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_35789 = 4'h3 < realFlowNum_0 ? _GEN_31563 : _GEN_27723; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_35790 = 4'h3 < realFlowNum_0 ? _GEN_31564 : _GEN_27724; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_35791 = 4'h3 < realFlowNum_0 ? _GEN_31565 : _GEN_27725; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_35792 = 4'h3 < realFlowNum_0 ? _GEN_31566 : _GEN_27726; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_35793 = 4'h3 < realFlowNum_0 ? _GEN_31567 : _GEN_27727; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_35794 = 4'h3 < realFlowNum_0 ? _GEN_31568 : _GEN_27728; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_35795 = 4'h3 < realFlowNum_0 ? _GEN_31569 : _GEN_27729; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_35796 = 4'h3 < realFlowNum_0 ? _GEN_31570 : _GEN_27730; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_35797 = 4'h3 < realFlowNum_0 ? _GEN_31571 : _GEN_27731; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_35798 = 4'h3 < realFlowNum_0 ? _GEN_31572 : _GEN_27732; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_35799 = 4'h3 < realFlowNum_0 ? _GEN_31573 : _GEN_27733; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_35800 = 4'h3 < realFlowNum_0 ? _GEN_31574 : _GEN_27734; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_35801 = 4'h3 < realFlowNum_0 ? _GEN_31575 : _GEN_27735; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_35802 = 4'h3 < realFlowNum_0 ? _GEN_31576 : _GEN_27736; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_35803 = 4'h3 < realFlowNum_0 ? _GEN_31577 : _GEN_27737; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_35804 = 4'h3 < realFlowNum_0 ? _GEN_31578 : _GEN_27738; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_35805 = 4'h3 < realFlowNum_0 ? _GEN_31579 : _GEN_27739; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_35806 = 4'h3 < realFlowNum_0 ? _GEN_31580 : _GEN_27740; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_35807 = 4'h3 < realFlowNum_0 ? _GEN_31581 : _GEN_27741; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_35808 = 4'h3 < realFlowNum_0 ? _GEN_31582 : _GEN_27742; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_35809 = 4'h3 < realFlowNum_0 ? _GEN_31583 : _GEN_27743; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_35810 = 4'h3 < realFlowNum_0 ? _GEN_31584 : _GEN_27744; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_35811 = 4'h3 < realFlowNum_0 ? _GEN_31585 : _GEN_27745; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_35812 = 4'h3 < realFlowNum_0 ? _GEN_31586 : _GEN_27746; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_35813 = 4'h3 < realFlowNum_0 ? _GEN_31587 : _GEN_27747; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_35814 = 4'h3 < realFlowNum_0 ? _GEN_31588 : _GEN_27748; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_35815 = 4'h3 < realFlowNum_0 ? _GEN_31589 : _GEN_27749; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_36072 = _GEN_161423 | _GEN_32231; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_36073 = _GEN_161424 | _GEN_32232; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_36074 = _GEN_161425 | _GEN_32233; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_36075 = _GEN_161426 | _GEN_32234; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_36076 = _GEN_161427 | _GEN_32235; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_36077 = _GEN_161428 | _GEN_32236; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_36078 = _GEN_161429 | _GEN_32237; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_36079 = _GEN_161430 | _GEN_32238; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_36080 = _GEN_161431 | _GEN_32239; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_36081 = _GEN_161432 | _GEN_32240; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_36082 = _GEN_161433 | _GEN_32241; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_36083 = _GEN_161434 | _GEN_32242; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_36084 = _GEN_161435 | _GEN_32243; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_36085 = _GEN_161436 | _GEN_32244; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_36086 = _GEN_161437 | _GEN_32245; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_36087 = _GEN_161438 | _GEN_32246; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_36088 = _GEN_161439 | _GEN_32247; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_36089 = _GEN_161440 | _GEN_32248; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_36090 = _GEN_161441 | _GEN_32249; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_36091 = _GEN_161442 | _GEN_32250; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_36092 = _GEN_161443 | _GEN_32251; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_36093 = _GEN_161444 | _GEN_32252; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_36094 = _GEN_161445 | _GEN_32253; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_36095 = _GEN_161446 | _GEN_32254; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_36096 = _GEN_161447 | _GEN_32255; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_36097 = _GEN_161448 | _GEN_32256; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_36098 = _GEN_161449 | _GEN_32257; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_36099 = _GEN_161450 | _GEN_32258; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_36100 = _GEN_161451 | _GEN_32259; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_36101 = _GEN_161452 | _GEN_32260; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_36102 = _GEN_161453 | _GEN_32261; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_36103 = _GEN_161454 | _GEN_32262; // @[Vlflowqueue.scala 197:{51,51}]
  wire [4:0] _GEN_39048 = 5'h0 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_35207; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_39049 = 5'h1 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_35208; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_39050 = 5'h2 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_35209; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_39051 = 5'h3 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_35210; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_39052 = 5'h4 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_35211; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_39053 = 5'h5 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_35212; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_39054 = 5'h6 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_35213; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_39055 = 5'h7 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_35214; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_39056 = 5'h8 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_35215; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_39057 = 5'h9 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_35216; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_39058 = 5'ha == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_35217; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_39059 = 5'hb == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_35218; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_39060 = 5'hc == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_35219; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_39061 = 5'hd == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_35220; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_39062 = 5'he == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_35221; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_39063 = 5'hf == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_35222; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_39064 = 5'h10 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_35223; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_39065 = 5'h11 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_35224; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_39066 = 5'h12 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_35225; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_39067 = 5'h13 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_35226; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_39068 = 5'h14 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_35227; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_39069 = 5'h15 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_35228; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_39070 = 5'h16 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_35229; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_39071 = 5'h17 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_35230; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_39072 = 5'h18 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_35231; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_39073 = 5'h19 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_35232; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_39074 = 5'h1a == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_35233; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_39075 = 5'h1b == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_35234; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_39076 = 5'h1c == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_35235; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_39077 = 5'h1d == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_35236; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_39078 = 5'h1e == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_35237; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_39079 = 5'h1f == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_35238; // @[Vlflowqueue.scala 198:{51,51}]
  wire [38:0] _GEN_39624 = 5'h0 == index_0 ? vaddr_0 : _GEN_35784; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_39625 = 5'h1 == index_0 ? vaddr_0 : _GEN_35785; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_39626 = 5'h2 == index_0 ? vaddr_0 : _GEN_35786; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_39627 = 5'h3 == index_0 ? vaddr_0 : _GEN_35787; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_39628 = 5'h4 == index_0 ? vaddr_0 : _GEN_35788; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_39629 = 5'h5 == index_0 ? vaddr_0 : _GEN_35789; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_39630 = 5'h6 == index_0 ? vaddr_0 : _GEN_35790; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_39631 = 5'h7 == index_0 ? vaddr_0 : _GEN_35791; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_39632 = 5'h8 == index_0 ? vaddr_0 : _GEN_35792; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_39633 = 5'h9 == index_0 ? vaddr_0 : _GEN_35793; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_39634 = 5'ha == index_0 ? vaddr_0 : _GEN_35794; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_39635 = 5'hb == index_0 ? vaddr_0 : _GEN_35795; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_39636 = 5'hc == index_0 ? vaddr_0 : _GEN_35796; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_39637 = 5'hd == index_0 ? vaddr_0 : _GEN_35797; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_39638 = 5'he == index_0 ? vaddr_0 : _GEN_35798; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_39639 = 5'hf == index_0 ? vaddr_0 : _GEN_35799; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_39640 = 5'h10 == index_0 ? vaddr_0 : _GEN_35800; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_39641 = 5'h11 == index_0 ? vaddr_0 : _GEN_35801; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_39642 = 5'h12 == index_0 ? vaddr_0 : _GEN_35802; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_39643 = 5'h13 == index_0 ? vaddr_0 : _GEN_35803; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_39644 = 5'h14 == index_0 ? vaddr_0 : _GEN_35804; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_39645 = 5'h15 == index_0 ? vaddr_0 : _GEN_35805; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_39646 = 5'h16 == index_0 ? vaddr_0 : _GEN_35806; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_39647 = 5'h17 == index_0 ? vaddr_0 : _GEN_35807; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_39648 = 5'h18 == index_0 ? vaddr_0 : _GEN_35808; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_39649 = 5'h19 == index_0 ? vaddr_0 : _GEN_35809; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_39650 = 5'h1a == index_0 ? vaddr_0 : _GEN_35810; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_39651 = 5'h1b == index_0 ? vaddr_0 : _GEN_35811; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_39652 = 5'h1c == index_0 ? vaddr_0 : _GEN_35812; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_39653 = 5'h1d == index_0 ? vaddr_0 : _GEN_35813; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_39654 = 5'h1e == index_0 ? vaddr_0 : _GEN_35814; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_39655 = 5'h1f == index_0 ? vaddr_0 : _GEN_35815; // @[Vlflowqueue.scala 203:{51,51}]
  wire  _GEN_40297 = 4'h4 < realFlowNum_0 ? _GEN_36072 : _GEN_32231; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_40298 = 4'h4 < realFlowNum_0 ? _GEN_36073 : _GEN_32232; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_40299 = 4'h4 < realFlowNum_0 ? _GEN_36074 : _GEN_32233; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_40300 = 4'h4 < realFlowNum_0 ? _GEN_36075 : _GEN_32234; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_40301 = 4'h4 < realFlowNum_0 ? _GEN_36076 : _GEN_32235; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_40302 = 4'h4 < realFlowNum_0 ? _GEN_36077 : _GEN_32236; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_40303 = 4'h4 < realFlowNum_0 ? _GEN_36078 : _GEN_32237; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_40304 = 4'h4 < realFlowNum_0 ? _GEN_36079 : _GEN_32238; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_40305 = 4'h4 < realFlowNum_0 ? _GEN_36080 : _GEN_32239; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_40306 = 4'h4 < realFlowNum_0 ? _GEN_36081 : _GEN_32240; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_40307 = 4'h4 < realFlowNum_0 ? _GEN_36082 : _GEN_32241; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_40308 = 4'h4 < realFlowNum_0 ? _GEN_36083 : _GEN_32242; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_40309 = 4'h4 < realFlowNum_0 ? _GEN_36084 : _GEN_32243; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_40310 = 4'h4 < realFlowNum_0 ? _GEN_36085 : _GEN_32244; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_40311 = 4'h4 < realFlowNum_0 ? _GEN_36086 : _GEN_32245; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_40312 = 4'h4 < realFlowNum_0 ? _GEN_36087 : _GEN_32246; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_40313 = 4'h4 < realFlowNum_0 ? _GEN_36088 : _GEN_32247; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_40314 = 4'h4 < realFlowNum_0 ? _GEN_36089 : _GEN_32248; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_40315 = 4'h4 < realFlowNum_0 ? _GEN_36090 : _GEN_32249; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_40316 = 4'h4 < realFlowNum_0 ? _GEN_36091 : _GEN_32250; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_40317 = 4'h4 < realFlowNum_0 ? _GEN_36092 : _GEN_32251; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_40318 = 4'h4 < realFlowNum_0 ? _GEN_36093 : _GEN_32252; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_40319 = 4'h4 < realFlowNum_0 ? _GEN_36094 : _GEN_32253; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_40320 = 4'h4 < realFlowNum_0 ? _GEN_36095 : _GEN_32254; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_40321 = 4'h4 < realFlowNum_0 ? _GEN_36096 : _GEN_32255; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_40322 = 4'h4 < realFlowNum_0 ? _GEN_36097 : _GEN_32256; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_40323 = 4'h4 < realFlowNum_0 ? _GEN_36098 : _GEN_32257; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_40324 = 4'h4 < realFlowNum_0 ? _GEN_36099 : _GEN_32258; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_40325 = 4'h4 < realFlowNum_0 ? _GEN_36100 : _GEN_32259; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_40326 = 4'h4 < realFlowNum_0 ? _GEN_36101 : _GEN_32260; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_40327 = 4'h4 < realFlowNum_0 ? _GEN_36102 : _GEN_32261; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_40328 = 4'h4 < realFlowNum_0 ? _GEN_36103 : _GEN_32262; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_43273 = 4'h4 < realFlowNum_0 ? _GEN_39048 : _GEN_35207; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_43274 = 4'h4 < realFlowNum_0 ? _GEN_39049 : _GEN_35208; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_43275 = 4'h4 < realFlowNum_0 ? _GEN_39050 : _GEN_35209; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_43276 = 4'h4 < realFlowNum_0 ? _GEN_39051 : _GEN_35210; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_43277 = 4'h4 < realFlowNum_0 ? _GEN_39052 : _GEN_35211; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_43278 = 4'h4 < realFlowNum_0 ? _GEN_39053 : _GEN_35212; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_43279 = 4'h4 < realFlowNum_0 ? _GEN_39054 : _GEN_35213; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_43280 = 4'h4 < realFlowNum_0 ? _GEN_39055 : _GEN_35214; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_43281 = 4'h4 < realFlowNum_0 ? _GEN_39056 : _GEN_35215; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_43282 = 4'h4 < realFlowNum_0 ? _GEN_39057 : _GEN_35216; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_43283 = 4'h4 < realFlowNum_0 ? _GEN_39058 : _GEN_35217; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_43284 = 4'h4 < realFlowNum_0 ? _GEN_39059 : _GEN_35218; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_43285 = 4'h4 < realFlowNum_0 ? _GEN_39060 : _GEN_35219; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_43286 = 4'h4 < realFlowNum_0 ? _GEN_39061 : _GEN_35220; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_43287 = 4'h4 < realFlowNum_0 ? _GEN_39062 : _GEN_35221; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_43288 = 4'h4 < realFlowNum_0 ? _GEN_39063 : _GEN_35222; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_43289 = 4'h4 < realFlowNum_0 ? _GEN_39064 : _GEN_35223; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_43290 = 4'h4 < realFlowNum_0 ? _GEN_39065 : _GEN_35224; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_43291 = 4'h4 < realFlowNum_0 ? _GEN_39066 : _GEN_35225; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_43292 = 4'h4 < realFlowNum_0 ? _GEN_39067 : _GEN_35226; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_43293 = 4'h4 < realFlowNum_0 ? _GEN_39068 : _GEN_35227; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_43294 = 4'h4 < realFlowNum_0 ? _GEN_39069 : _GEN_35228; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_43295 = 4'h4 < realFlowNum_0 ? _GEN_39070 : _GEN_35229; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_43296 = 4'h4 < realFlowNum_0 ? _GEN_39071 : _GEN_35230; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_43297 = 4'h4 < realFlowNum_0 ? _GEN_39072 : _GEN_35231; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_43298 = 4'h4 < realFlowNum_0 ? _GEN_39073 : _GEN_35232; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_43299 = 4'h4 < realFlowNum_0 ? _GEN_39074 : _GEN_35233; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_43300 = 4'h4 < realFlowNum_0 ? _GEN_39075 : _GEN_35234; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_43301 = 4'h4 < realFlowNum_0 ? _GEN_39076 : _GEN_35235; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_43302 = 4'h4 < realFlowNum_0 ? _GEN_39077 : _GEN_35236; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_43303 = 4'h4 < realFlowNum_0 ? _GEN_39078 : _GEN_35237; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_43304 = 4'h4 < realFlowNum_0 ? _GEN_39079 : _GEN_35238; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_43850 = 4'h4 < realFlowNum_0 ? _GEN_39624 : _GEN_35784; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_43851 = 4'h4 < realFlowNum_0 ? _GEN_39625 : _GEN_35785; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_43852 = 4'h4 < realFlowNum_0 ? _GEN_39626 : _GEN_35786; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_43853 = 4'h4 < realFlowNum_0 ? _GEN_39627 : _GEN_35787; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_43854 = 4'h4 < realFlowNum_0 ? _GEN_39628 : _GEN_35788; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_43855 = 4'h4 < realFlowNum_0 ? _GEN_39629 : _GEN_35789; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_43856 = 4'h4 < realFlowNum_0 ? _GEN_39630 : _GEN_35790; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_43857 = 4'h4 < realFlowNum_0 ? _GEN_39631 : _GEN_35791; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_43858 = 4'h4 < realFlowNum_0 ? _GEN_39632 : _GEN_35792; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_43859 = 4'h4 < realFlowNum_0 ? _GEN_39633 : _GEN_35793; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_43860 = 4'h4 < realFlowNum_0 ? _GEN_39634 : _GEN_35794; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_43861 = 4'h4 < realFlowNum_0 ? _GEN_39635 : _GEN_35795; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_43862 = 4'h4 < realFlowNum_0 ? _GEN_39636 : _GEN_35796; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_43863 = 4'h4 < realFlowNum_0 ? _GEN_39637 : _GEN_35797; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_43864 = 4'h4 < realFlowNum_0 ? _GEN_39638 : _GEN_35798; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_43865 = 4'h4 < realFlowNum_0 ? _GEN_39639 : _GEN_35799; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_43866 = 4'h4 < realFlowNum_0 ? _GEN_39640 : _GEN_35800; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_43867 = 4'h4 < realFlowNum_0 ? _GEN_39641 : _GEN_35801; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_43868 = 4'h4 < realFlowNum_0 ? _GEN_39642 : _GEN_35802; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_43869 = 4'h4 < realFlowNum_0 ? _GEN_39643 : _GEN_35803; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_43870 = 4'h4 < realFlowNum_0 ? _GEN_39644 : _GEN_35804; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_43871 = 4'h4 < realFlowNum_0 ? _GEN_39645 : _GEN_35805; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_43872 = 4'h4 < realFlowNum_0 ? _GEN_39646 : _GEN_35806; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_43873 = 4'h4 < realFlowNum_0 ? _GEN_39647 : _GEN_35807; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_43874 = 4'h4 < realFlowNum_0 ? _GEN_39648 : _GEN_35808; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_43875 = 4'h4 < realFlowNum_0 ? _GEN_39649 : _GEN_35809; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_43876 = 4'h4 < realFlowNum_0 ? _GEN_39650 : _GEN_35810; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_43877 = 4'h4 < realFlowNum_0 ? _GEN_39651 : _GEN_35811; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_43878 = 4'h4 < realFlowNum_0 ? _GEN_39652 : _GEN_35812; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_43879 = 4'h4 < realFlowNum_0 ? _GEN_39653 : _GEN_35813; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_43880 = 4'h4 < realFlowNum_0 ? _GEN_39654 : _GEN_35814; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_43881 = 4'h4 < realFlowNum_0 ? _GEN_39655 : _GEN_35815; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_44138 = _GEN_161423 | _GEN_40297; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_44139 = _GEN_161424 | _GEN_40298; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_44140 = _GEN_161425 | _GEN_40299; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_44141 = _GEN_161426 | _GEN_40300; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_44142 = _GEN_161427 | _GEN_40301; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_44143 = _GEN_161428 | _GEN_40302; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_44144 = _GEN_161429 | _GEN_40303; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_44145 = _GEN_161430 | _GEN_40304; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_44146 = _GEN_161431 | _GEN_40305; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_44147 = _GEN_161432 | _GEN_40306; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_44148 = _GEN_161433 | _GEN_40307; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_44149 = _GEN_161434 | _GEN_40308; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_44150 = _GEN_161435 | _GEN_40309; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_44151 = _GEN_161436 | _GEN_40310; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_44152 = _GEN_161437 | _GEN_40311; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_44153 = _GEN_161438 | _GEN_40312; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_44154 = _GEN_161439 | _GEN_40313; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_44155 = _GEN_161440 | _GEN_40314; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_44156 = _GEN_161441 | _GEN_40315; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_44157 = _GEN_161442 | _GEN_40316; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_44158 = _GEN_161443 | _GEN_40317; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_44159 = _GEN_161444 | _GEN_40318; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_44160 = _GEN_161445 | _GEN_40319; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_44161 = _GEN_161446 | _GEN_40320; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_44162 = _GEN_161447 | _GEN_40321; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_44163 = _GEN_161448 | _GEN_40322; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_44164 = _GEN_161449 | _GEN_40323; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_44165 = _GEN_161450 | _GEN_40324; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_44166 = _GEN_161451 | _GEN_40325; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_44167 = _GEN_161452 | _GEN_40326; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_44168 = _GEN_161453 | _GEN_40327; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_44169 = _GEN_161454 | _GEN_40328; // @[Vlflowqueue.scala 197:{51,51}]
  wire [4:0] _GEN_47114 = 5'h0 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_43273; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_47115 = 5'h1 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_43274; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_47116 = 5'h2 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_43275; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_47117 = 5'h3 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_43276; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_47118 = 5'h4 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_43277; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_47119 = 5'h5 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_43278; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_47120 = 5'h6 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_43279; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_47121 = 5'h7 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_43280; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_47122 = 5'h8 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_43281; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_47123 = 5'h9 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_43282; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_47124 = 5'ha == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_43283; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_47125 = 5'hb == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_43284; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_47126 = 5'hc == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_43285; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_47127 = 5'hd == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_43286; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_47128 = 5'he == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_43287; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_47129 = 5'hf == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_43288; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_47130 = 5'h10 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_43289; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_47131 = 5'h11 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_43290; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_47132 = 5'h12 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_43291; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_47133 = 5'h13 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_43292; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_47134 = 5'h14 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_43293; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_47135 = 5'h15 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_43294; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_47136 = 5'h16 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_43295; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_47137 = 5'h17 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_43296; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_47138 = 5'h18 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_43297; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_47139 = 5'h19 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_43298; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_47140 = 5'h1a == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_43299; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_47141 = 5'h1b == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_43300; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_47142 = 5'h1c == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_43301; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_47143 = 5'h1d == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_43302; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_47144 = 5'h1e == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_43303; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_47145 = 5'h1f == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_43304; // @[Vlflowqueue.scala 198:{51,51}]
  wire [38:0] _GEN_47690 = 5'h0 == index_0 ? vaddr_0 : _GEN_43850; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_47691 = 5'h1 == index_0 ? vaddr_0 : _GEN_43851; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_47692 = 5'h2 == index_0 ? vaddr_0 : _GEN_43852; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_47693 = 5'h3 == index_0 ? vaddr_0 : _GEN_43853; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_47694 = 5'h4 == index_0 ? vaddr_0 : _GEN_43854; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_47695 = 5'h5 == index_0 ? vaddr_0 : _GEN_43855; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_47696 = 5'h6 == index_0 ? vaddr_0 : _GEN_43856; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_47697 = 5'h7 == index_0 ? vaddr_0 : _GEN_43857; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_47698 = 5'h8 == index_0 ? vaddr_0 : _GEN_43858; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_47699 = 5'h9 == index_0 ? vaddr_0 : _GEN_43859; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_47700 = 5'ha == index_0 ? vaddr_0 : _GEN_43860; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_47701 = 5'hb == index_0 ? vaddr_0 : _GEN_43861; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_47702 = 5'hc == index_0 ? vaddr_0 : _GEN_43862; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_47703 = 5'hd == index_0 ? vaddr_0 : _GEN_43863; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_47704 = 5'he == index_0 ? vaddr_0 : _GEN_43864; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_47705 = 5'hf == index_0 ? vaddr_0 : _GEN_43865; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_47706 = 5'h10 == index_0 ? vaddr_0 : _GEN_43866; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_47707 = 5'h11 == index_0 ? vaddr_0 : _GEN_43867; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_47708 = 5'h12 == index_0 ? vaddr_0 : _GEN_43868; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_47709 = 5'h13 == index_0 ? vaddr_0 : _GEN_43869; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_47710 = 5'h14 == index_0 ? vaddr_0 : _GEN_43870; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_47711 = 5'h15 == index_0 ? vaddr_0 : _GEN_43871; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_47712 = 5'h16 == index_0 ? vaddr_0 : _GEN_43872; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_47713 = 5'h17 == index_0 ? vaddr_0 : _GEN_43873; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_47714 = 5'h18 == index_0 ? vaddr_0 : _GEN_43874; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_47715 = 5'h19 == index_0 ? vaddr_0 : _GEN_43875; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_47716 = 5'h1a == index_0 ? vaddr_0 : _GEN_43876; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_47717 = 5'h1b == index_0 ? vaddr_0 : _GEN_43877; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_47718 = 5'h1c == index_0 ? vaddr_0 : _GEN_43878; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_47719 = 5'h1d == index_0 ? vaddr_0 : _GEN_43879; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_47720 = 5'h1e == index_0 ? vaddr_0 : _GEN_43880; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_47721 = 5'h1f == index_0 ? vaddr_0 : _GEN_43881; // @[Vlflowqueue.scala 203:{51,51}]
  wire  _GEN_48363 = 4'h5 < realFlowNum_0 ? _GEN_44138 : _GEN_40297; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_48364 = 4'h5 < realFlowNum_0 ? _GEN_44139 : _GEN_40298; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_48365 = 4'h5 < realFlowNum_0 ? _GEN_44140 : _GEN_40299; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_48366 = 4'h5 < realFlowNum_0 ? _GEN_44141 : _GEN_40300; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_48367 = 4'h5 < realFlowNum_0 ? _GEN_44142 : _GEN_40301; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_48368 = 4'h5 < realFlowNum_0 ? _GEN_44143 : _GEN_40302; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_48369 = 4'h5 < realFlowNum_0 ? _GEN_44144 : _GEN_40303; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_48370 = 4'h5 < realFlowNum_0 ? _GEN_44145 : _GEN_40304; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_48371 = 4'h5 < realFlowNum_0 ? _GEN_44146 : _GEN_40305; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_48372 = 4'h5 < realFlowNum_0 ? _GEN_44147 : _GEN_40306; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_48373 = 4'h5 < realFlowNum_0 ? _GEN_44148 : _GEN_40307; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_48374 = 4'h5 < realFlowNum_0 ? _GEN_44149 : _GEN_40308; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_48375 = 4'h5 < realFlowNum_0 ? _GEN_44150 : _GEN_40309; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_48376 = 4'h5 < realFlowNum_0 ? _GEN_44151 : _GEN_40310; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_48377 = 4'h5 < realFlowNum_0 ? _GEN_44152 : _GEN_40311; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_48378 = 4'h5 < realFlowNum_0 ? _GEN_44153 : _GEN_40312; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_48379 = 4'h5 < realFlowNum_0 ? _GEN_44154 : _GEN_40313; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_48380 = 4'h5 < realFlowNum_0 ? _GEN_44155 : _GEN_40314; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_48381 = 4'h5 < realFlowNum_0 ? _GEN_44156 : _GEN_40315; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_48382 = 4'h5 < realFlowNum_0 ? _GEN_44157 : _GEN_40316; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_48383 = 4'h5 < realFlowNum_0 ? _GEN_44158 : _GEN_40317; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_48384 = 4'h5 < realFlowNum_0 ? _GEN_44159 : _GEN_40318; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_48385 = 4'h5 < realFlowNum_0 ? _GEN_44160 : _GEN_40319; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_48386 = 4'h5 < realFlowNum_0 ? _GEN_44161 : _GEN_40320; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_48387 = 4'h5 < realFlowNum_0 ? _GEN_44162 : _GEN_40321; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_48388 = 4'h5 < realFlowNum_0 ? _GEN_44163 : _GEN_40322; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_48389 = 4'h5 < realFlowNum_0 ? _GEN_44164 : _GEN_40323; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_48390 = 4'h5 < realFlowNum_0 ? _GEN_44165 : _GEN_40324; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_48391 = 4'h5 < realFlowNum_0 ? _GEN_44166 : _GEN_40325; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_48392 = 4'h5 < realFlowNum_0 ? _GEN_44167 : _GEN_40326; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_48393 = 4'h5 < realFlowNum_0 ? _GEN_44168 : _GEN_40327; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_48394 = 4'h5 < realFlowNum_0 ? _GEN_44169 : _GEN_40328; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_51339 = 4'h5 < realFlowNum_0 ? _GEN_47114 : _GEN_43273; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_51340 = 4'h5 < realFlowNum_0 ? _GEN_47115 : _GEN_43274; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_51341 = 4'h5 < realFlowNum_0 ? _GEN_47116 : _GEN_43275; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_51342 = 4'h5 < realFlowNum_0 ? _GEN_47117 : _GEN_43276; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_51343 = 4'h5 < realFlowNum_0 ? _GEN_47118 : _GEN_43277; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_51344 = 4'h5 < realFlowNum_0 ? _GEN_47119 : _GEN_43278; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_51345 = 4'h5 < realFlowNum_0 ? _GEN_47120 : _GEN_43279; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_51346 = 4'h5 < realFlowNum_0 ? _GEN_47121 : _GEN_43280; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_51347 = 4'h5 < realFlowNum_0 ? _GEN_47122 : _GEN_43281; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_51348 = 4'h5 < realFlowNum_0 ? _GEN_47123 : _GEN_43282; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_51349 = 4'h5 < realFlowNum_0 ? _GEN_47124 : _GEN_43283; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_51350 = 4'h5 < realFlowNum_0 ? _GEN_47125 : _GEN_43284; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_51351 = 4'h5 < realFlowNum_0 ? _GEN_47126 : _GEN_43285; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_51352 = 4'h5 < realFlowNum_0 ? _GEN_47127 : _GEN_43286; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_51353 = 4'h5 < realFlowNum_0 ? _GEN_47128 : _GEN_43287; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_51354 = 4'h5 < realFlowNum_0 ? _GEN_47129 : _GEN_43288; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_51355 = 4'h5 < realFlowNum_0 ? _GEN_47130 : _GEN_43289; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_51356 = 4'h5 < realFlowNum_0 ? _GEN_47131 : _GEN_43290; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_51357 = 4'h5 < realFlowNum_0 ? _GEN_47132 : _GEN_43291; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_51358 = 4'h5 < realFlowNum_0 ? _GEN_47133 : _GEN_43292; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_51359 = 4'h5 < realFlowNum_0 ? _GEN_47134 : _GEN_43293; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_51360 = 4'h5 < realFlowNum_0 ? _GEN_47135 : _GEN_43294; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_51361 = 4'h5 < realFlowNum_0 ? _GEN_47136 : _GEN_43295; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_51362 = 4'h5 < realFlowNum_0 ? _GEN_47137 : _GEN_43296; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_51363 = 4'h5 < realFlowNum_0 ? _GEN_47138 : _GEN_43297; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_51364 = 4'h5 < realFlowNum_0 ? _GEN_47139 : _GEN_43298; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_51365 = 4'h5 < realFlowNum_0 ? _GEN_47140 : _GEN_43299; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_51366 = 4'h5 < realFlowNum_0 ? _GEN_47141 : _GEN_43300; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_51367 = 4'h5 < realFlowNum_0 ? _GEN_47142 : _GEN_43301; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_51368 = 4'h5 < realFlowNum_0 ? _GEN_47143 : _GEN_43302; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_51369 = 4'h5 < realFlowNum_0 ? _GEN_47144 : _GEN_43303; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_51370 = 4'h5 < realFlowNum_0 ? _GEN_47145 : _GEN_43304; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_51916 = 4'h5 < realFlowNum_0 ? _GEN_47690 : _GEN_43850; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_51917 = 4'h5 < realFlowNum_0 ? _GEN_47691 : _GEN_43851; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_51918 = 4'h5 < realFlowNum_0 ? _GEN_47692 : _GEN_43852; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_51919 = 4'h5 < realFlowNum_0 ? _GEN_47693 : _GEN_43853; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_51920 = 4'h5 < realFlowNum_0 ? _GEN_47694 : _GEN_43854; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_51921 = 4'h5 < realFlowNum_0 ? _GEN_47695 : _GEN_43855; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_51922 = 4'h5 < realFlowNum_0 ? _GEN_47696 : _GEN_43856; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_51923 = 4'h5 < realFlowNum_0 ? _GEN_47697 : _GEN_43857; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_51924 = 4'h5 < realFlowNum_0 ? _GEN_47698 : _GEN_43858; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_51925 = 4'h5 < realFlowNum_0 ? _GEN_47699 : _GEN_43859; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_51926 = 4'h5 < realFlowNum_0 ? _GEN_47700 : _GEN_43860; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_51927 = 4'h5 < realFlowNum_0 ? _GEN_47701 : _GEN_43861; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_51928 = 4'h5 < realFlowNum_0 ? _GEN_47702 : _GEN_43862; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_51929 = 4'h5 < realFlowNum_0 ? _GEN_47703 : _GEN_43863; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_51930 = 4'h5 < realFlowNum_0 ? _GEN_47704 : _GEN_43864; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_51931 = 4'h5 < realFlowNum_0 ? _GEN_47705 : _GEN_43865; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_51932 = 4'h5 < realFlowNum_0 ? _GEN_47706 : _GEN_43866; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_51933 = 4'h5 < realFlowNum_0 ? _GEN_47707 : _GEN_43867; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_51934 = 4'h5 < realFlowNum_0 ? _GEN_47708 : _GEN_43868; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_51935 = 4'h5 < realFlowNum_0 ? _GEN_47709 : _GEN_43869; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_51936 = 4'h5 < realFlowNum_0 ? _GEN_47710 : _GEN_43870; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_51937 = 4'h5 < realFlowNum_0 ? _GEN_47711 : _GEN_43871; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_51938 = 4'h5 < realFlowNum_0 ? _GEN_47712 : _GEN_43872; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_51939 = 4'h5 < realFlowNum_0 ? _GEN_47713 : _GEN_43873; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_51940 = 4'h5 < realFlowNum_0 ? _GEN_47714 : _GEN_43874; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_51941 = 4'h5 < realFlowNum_0 ? _GEN_47715 : _GEN_43875; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_51942 = 4'h5 < realFlowNum_0 ? _GEN_47716 : _GEN_43876; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_51943 = 4'h5 < realFlowNum_0 ? _GEN_47717 : _GEN_43877; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_51944 = 4'h5 < realFlowNum_0 ? _GEN_47718 : _GEN_43878; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_51945 = 4'h5 < realFlowNum_0 ? _GEN_47719 : _GEN_43879; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_51946 = 4'h5 < realFlowNum_0 ? _GEN_47720 : _GEN_43880; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_51947 = 4'h5 < realFlowNum_0 ? _GEN_47721 : _GEN_43881; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_52204 = _GEN_161423 | _GEN_48363; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_52205 = _GEN_161424 | _GEN_48364; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_52206 = _GEN_161425 | _GEN_48365; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_52207 = _GEN_161426 | _GEN_48366; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_52208 = _GEN_161427 | _GEN_48367; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_52209 = _GEN_161428 | _GEN_48368; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_52210 = _GEN_161429 | _GEN_48369; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_52211 = _GEN_161430 | _GEN_48370; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_52212 = _GEN_161431 | _GEN_48371; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_52213 = _GEN_161432 | _GEN_48372; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_52214 = _GEN_161433 | _GEN_48373; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_52215 = _GEN_161434 | _GEN_48374; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_52216 = _GEN_161435 | _GEN_48375; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_52217 = _GEN_161436 | _GEN_48376; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_52218 = _GEN_161437 | _GEN_48377; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_52219 = _GEN_161438 | _GEN_48378; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_52220 = _GEN_161439 | _GEN_48379; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_52221 = _GEN_161440 | _GEN_48380; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_52222 = _GEN_161441 | _GEN_48381; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_52223 = _GEN_161442 | _GEN_48382; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_52224 = _GEN_161443 | _GEN_48383; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_52225 = _GEN_161444 | _GEN_48384; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_52226 = _GEN_161445 | _GEN_48385; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_52227 = _GEN_161446 | _GEN_48386; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_52228 = _GEN_161447 | _GEN_48387; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_52229 = _GEN_161448 | _GEN_48388; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_52230 = _GEN_161449 | _GEN_48389; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_52231 = _GEN_161450 | _GEN_48390; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_52232 = _GEN_161451 | _GEN_48391; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_52233 = _GEN_161452 | _GEN_48392; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_52234 = _GEN_161453 | _GEN_48393; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_52235 = _GEN_161454 | _GEN_48394; // @[Vlflowqueue.scala 197:{51,51}]
  wire [4:0] _GEN_55180 = 5'h0 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_51339; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_55181 = 5'h1 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_51340; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_55182 = 5'h2 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_51341; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_55183 = 5'h3 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_51342; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_55184 = 5'h4 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_51343; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_55185 = 5'h5 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_51344; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_55186 = 5'h6 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_51345; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_55187 = 5'h7 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_51346; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_55188 = 5'h8 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_51347; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_55189 = 5'h9 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_51348; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_55190 = 5'ha == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_51349; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_55191 = 5'hb == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_51350; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_55192 = 5'hc == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_51351; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_55193 = 5'hd == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_51352; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_55194 = 5'he == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_51353; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_55195 = 5'hf == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_51354; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_55196 = 5'h10 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_51355; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_55197 = 5'h11 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_51356; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_55198 = 5'h12 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_51357; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_55199 = 5'h13 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_51358; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_55200 = 5'h14 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_51359; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_55201 = 5'h15 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_51360; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_55202 = 5'h16 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_51361; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_55203 = 5'h17 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_51362; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_55204 = 5'h18 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_51363; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_55205 = 5'h19 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_51364; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_55206 = 5'h1a == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_51365; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_55207 = 5'h1b == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_51366; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_55208 = 5'h1c == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_51367; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_55209 = 5'h1d == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_51368; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_55210 = 5'h1e == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_51369; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_55211 = 5'h1f == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_51370; // @[Vlflowqueue.scala 198:{51,51}]
  wire [38:0] _GEN_55756 = 5'h0 == index_0 ? vaddr_0 : _GEN_51916; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_55757 = 5'h1 == index_0 ? vaddr_0 : _GEN_51917; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_55758 = 5'h2 == index_0 ? vaddr_0 : _GEN_51918; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_55759 = 5'h3 == index_0 ? vaddr_0 : _GEN_51919; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_55760 = 5'h4 == index_0 ? vaddr_0 : _GEN_51920; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_55761 = 5'h5 == index_0 ? vaddr_0 : _GEN_51921; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_55762 = 5'h6 == index_0 ? vaddr_0 : _GEN_51922; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_55763 = 5'h7 == index_0 ? vaddr_0 : _GEN_51923; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_55764 = 5'h8 == index_0 ? vaddr_0 : _GEN_51924; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_55765 = 5'h9 == index_0 ? vaddr_0 : _GEN_51925; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_55766 = 5'ha == index_0 ? vaddr_0 : _GEN_51926; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_55767 = 5'hb == index_0 ? vaddr_0 : _GEN_51927; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_55768 = 5'hc == index_0 ? vaddr_0 : _GEN_51928; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_55769 = 5'hd == index_0 ? vaddr_0 : _GEN_51929; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_55770 = 5'he == index_0 ? vaddr_0 : _GEN_51930; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_55771 = 5'hf == index_0 ? vaddr_0 : _GEN_51931; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_55772 = 5'h10 == index_0 ? vaddr_0 : _GEN_51932; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_55773 = 5'h11 == index_0 ? vaddr_0 : _GEN_51933; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_55774 = 5'h12 == index_0 ? vaddr_0 : _GEN_51934; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_55775 = 5'h13 == index_0 ? vaddr_0 : _GEN_51935; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_55776 = 5'h14 == index_0 ? vaddr_0 : _GEN_51936; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_55777 = 5'h15 == index_0 ? vaddr_0 : _GEN_51937; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_55778 = 5'h16 == index_0 ? vaddr_0 : _GEN_51938; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_55779 = 5'h17 == index_0 ? vaddr_0 : _GEN_51939; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_55780 = 5'h18 == index_0 ? vaddr_0 : _GEN_51940; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_55781 = 5'h19 == index_0 ? vaddr_0 : _GEN_51941; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_55782 = 5'h1a == index_0 ? vaddr_0 : _GEN_51942; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_55783 = 5'h1b == index_0 ? vaddr_0 : _GEN_51943; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_55784 = 5'h1c == index_0 ? vaddr_0 : _GEN_51944; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_55785 = 5'h1d == index_0 ? vaddr_0 : _GEN_51945; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_55786 = 5'h1e == index_0 ? vaddr_0 : _GEN_51946; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_55787 = 5'h1f == index_0 ? vaddr_0 : _GEN_51947; // @[Vlflowqueue.scala 203:{51,51}]
  wire  _GEN_56429 = 4'h6 < realFlowNum_0 ? _GEN_52204 : _GEN_48363; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_56430 = 4'h6 < realFlowNum_0 ? _GEN_52205 : _GEN_48364; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_56431 = 4'h6 < realFlowNum_0 ? _GEN_52206 : _GEN_48365; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_56432 = 4'h6 < realFlowNum_0 ? _GEN_52207 : _GEN_48366; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_56433 = 4'h6 < realFlowNum_0 ? _GEN_52208 : _GEN_48367; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_56434 = 4'h6 < realFlowNum_0 ? _GEN_52209 : _GEN_48368; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_56435 = 4'h6 < realFlowNum_0 ? _GEN_52210 : _GEN_48369; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_56436 = 4'h6 < realFlowNum_0 ? _GEN_52211 : _GEN_48370; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_56437 = 4'h6 < realFlowNum_0 ? _GEN_52212 : _GEN_48371; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_56438 = 4'h6 < realFlowNum_0 ? _GEN_52213 : _GEN_48372; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_56439 = 4'h6 < realFlowNum_0 ? _GEN_52214 : _GEN_48373; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_56440 = 4'h6 < realFlowNum_0 ? _GEN_52215 : _GEN_48374; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_56441 = 4'h6 < realFlowNum_0 ? _GEN_52216 : _GEN_48375; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_56442 = 4'h6 < realFlowNum_0 ? _GEN_52217 : _GEN_48376; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_56443 = 4'h6 < realFlowNum_0 ? _GEN_52218 : _GEN_48377; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_56444 = 4'h6 < realFlowNum_0 ? _GEN_52219 : _GEN_48378; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_56445 = 4'h6 < realFlowNum_0 ? _GEN_52220 : _GEN_48379; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_56446 = 4'h6 < realFlowNum_0 ? _GEN_52221 : _GEN_48380; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_56447 = 4'h6 < realFlowNum_0 ? _GEN_52222 : _GEN_48381; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_56448 = 4'h6 < realFlowNum_0 ? _GEN_52223 : _GEN_48382; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_56449 = 4'h6 < realFlowNum_0 ? _GEN_52224 : _GEN_48383; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_56450 = 4'h6 < realFlowNum_0 ? _GEN_52225 : _GEN_48384; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_56451 = 4'h6 < realFlowNum_0 ? _GEN_52226 : _GEN_48385; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_56452 = 4'h6 < realFlowNum_0 ? _GEN_52227 : _GEN_48386; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_56453 = 4'h6 < realFlowNum_0 ? _GEN_52228 : _GEN_48387; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_56454 = 4'h6 < realFlowNum_0 ? _GEN_52229 : _GEN_48388; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_56455 = 4'h6 < realFlowNum_0 ? _GEN_52230 : _GEN_48389; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_56456 = 4'h6 < realFlowNum_0 ? _GEN_52231 : _GEN_48390; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_56457 = 4'h6 < realFlowNum_0 ? _GEN_52232 : _GEN_48391; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_56458 = 4'h6 < realFlowNum_0 ? _GEN_52233 : _GEN_48392; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_56459 = 4'h6 < realFlowNum_0 ? _GEN_52234 : _GEN_48393; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_56460 = 4'h6 < realFlowNum_0 ? _GEN_52235 : _GEN_48394; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_59405 = 4'h6 < realFlowNum_0 ? _GEN_55180 : _GEN_51339; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_59406 = 4'h6 < realFlowNum_0 ? _GEN_55181 : _GEN_51340; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_59407 = 4'h6 < realFlowNum_0 ? _GEN_55182 : _GEN_51341; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_59408 = 4'h6 < realFlowNum_0 ? _GEN_55183 : _GEN_51342; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_59409 = 4'h6 < realFlowNum_0 ? _GEN_55184 : _GEN_51343; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_59410 = 4'h6 < realFlowNum_0 ? _GEN_55185 : _GEN_51344; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_59411 = 4'h6 < realFlowNum_0 ? _GEN_55186 : _GEN_51345; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_59412 = 4'h6 < realFlowNum_0 ? _GEN_55187 : _GEN_51346; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_59413 = 4'h6 < realFlowNum_0 ? _GEN_55188 : _GEN_51347; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_59414 = 4'h6 < realFlowNum_0 ? _GEN_55189 : _GEN_51348; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_59415 = 4'h6 < realFlowNum_0 ? _GEN_55190 : _GEN_51349; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_59416 = 4'h6 < realFlowNum_0 ? _GEN_55191 : _GEN_51350; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_59417 = 4'h6 < realFlowNum_0 ? _GEN_55192 : _GEN_51351; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_59418 = 4'h6 < realFlowNum_0 ? _GEN_55193 : _GEN_51352; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_59419 = 4'h6 < realFlowNum_0 ? _GEN_55194 : _GEN_51353; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_59420 = 4'h6 < realFlowNum_0 ? _GEN_55195 : _GEN_51354; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_59421 = 4'h6 < realFlowNum_0 ? _GEN_55196 : _GEN_51355; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_59422 = 4'h6 < realFlowNum_0 ? _GEN_55197 : _GEN_51356; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_59423 = 4'h6 < realFlowNum_0 ? _GEN_55198 : _GEN_51357; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_59424 = 4'h6 < realFlowNum_0 ? _GEN_55199 : _GEN_51358; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_59425 = 4'h6 < realFlowNum_0 ? _GEN_55200 : _GEN_51359; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_59426 = 4'h6 < realFlowNum_0 ? _GEN_55201 : _GEN_51360; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_59427 = 4'h6 < realFlowNum_0 ? _GEN_55202 : _GEN_51361; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_59428 = 4'h6 < realFlowNum_0 ? _GEN_55203 : _GEN_51362; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_59429 = 4'h6 < realFlowNum_0 ? _GEN_55204 : _GEN_51363; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_59430 = 4'h6 < realFlowNum_0 ? _GEN_55205 : _GEN_51364; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_59431 = 4'h6 < realFlowNum_0 ? _GEN_55206 : _GEN_51365; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_59432 = 4'h6 < realFlowNum_0 ? _GEN_55207 : _GEN_51366; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_59433 = 4'h6 < realFlowNum_0 ? _GEN_55208 : _GEN_51367; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_59434 = 4'h6 < realFlowNum_0 ? _GEN_55209 : _GEN_51368; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_59435 = 4'h6 < realFlowNum_0 ? _GEN_55210 : _GEN_51369; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_59436 = 4'h6 < realFlowNum_0 ? _GEN_55211 : _GEN_51370; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_59982 = 4'h6 < realFlowNum_0 ? _GEN_55756 : _GEN_51916; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_59983 = 4'h6 < realFlowNum_0 ? _GEN_55757 : _GEN_51917; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_59984 = 4'h6 < realFlowNum_0 ? _GEN_55758 : _GEN_51918; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_59985 = 4'h6 < realFlowNum_0 ? _GEN_55759 : _GEN_51919; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_59986 = 4'h6 < realFlowNum_0 ? _GEN_55760 : _GEN_51920; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_59987 = 4'h6 < realFlowNum_0 ? _GEN_55761 : _GEN_51921; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_59988 = 4'h6 < realFlowNum_0 ? _GEN_55762 : _GEN_51922; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_59989 = 4'h6 < realFlowNum_0 ? _GEN_55763 : _GEN_51923; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_59990 = 4'h6 < realFlowNum_0 ? _GEN_55764 : _GEN_51924; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_59991 = 4'h6 < realFlowNum_0 ? _GEN_55765 : _GEN_51925; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_59992 = 4'h6 < realFlowNum_0 ? _GEN_55766 : _GEN_51926; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_59993 = 4'h6 < realFlowNum_0 ? _GEN_55767 : _GEN_51927; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_59994 = 4'h6 < realFlowNum_0 ? _GEN_55768 : _GEN_51928; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_59995 = 4'h6 < realFlowNum_0 ? _GEN_55769 : _GEN_51929; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_59996 = 4'h6 < realFlowNum_0 ? _GEN_55770 : _GEN_51930; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_59997 = 4'h6 < realFlowNum_0 ? _GEN_55771 : _GEN_51931; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_59998 = 4'h6 < realFlowNum_0 ? _GEN_55772 : _GEN_51932; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_59999 = 4'h6 < realFlowNum_0 ? _GEN_55773 : _GEN_51933; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_60000 = 4'h6 < realFlowNum_0 ? _GEN_55774 : _GEN_51934; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_60001 = 4'h6 < realFlowNum_0 ? _GEN_55775 : _GEN_51935; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_60002 = 4'h6 < realFlowNum_0 ? _GEN_55776 : _GEN_51936; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_60003 = 4'h6 < realFlowNum_0 ? _GEN_55777 : _GEN_51937; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_60004 = 4'h6 < realFlowNum_0 ? _GEN_55778 : _GEN_51938; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_60005 = 4'h6 < realFlowNum_0 ? _GEN_55779 : _GEN_51939; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_60006 = 4'h6 < realFlowNum_0 ? _GEN_55780 : _GEN_51940; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_60007 = 4'h6 < realFlowNum_0 ? _GEN_55781 : _GEN_51941; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_60008 = 4'h6 < realFlowNum_0 ? _GEN_55782 : _GEN_51942; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_60009 = 4'h6 < realFlowNum_0 ? _GEN_55783 : _GEN_51943; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_60010 = 4'h6 < realFlowNum_0 ? _GEN_55784 : _GEN_51944; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_60011 = 4'h6 < realFlowNum_0 ? _GEN_55785 : _GEN_51945; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_60012 = 4'h6 < realFlowNum_0 ? _GEN_55786 : _GEN_51946; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_60013 = 4'h6 < realFlowNum_0 ? _GEN_55787 : _GEN_51947; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_60270 = _GEN_161423 | _GEN_56429; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_60271 = _GEN_161424 | _GEN_56430; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_60272 = _GEN_161425 | _GEN_56431; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_60273 = _GEN_161426 | _GEN_56432; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_60274 = _GEN_161427 | _GEN_56433; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_60275 = _GEN_161428 | _GEN_56434; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_60276 = _GEN_161429 | _GEN_56435; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_60277 = _GEN_161430 | _GEN_56436; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_60278 = _GEN_161431 | _GEN_56437; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_60279 = _GEN_161432 | _GEN_56438; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_60280 = _GEN_161433 | _GEN_56439; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_60281 = _GEN_161434 | _GEN_56440; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_60282 = _GEN_161435 | _GEN_56441; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_60283 = _GEN_161436 | _GEN_56442; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_60284 = _GEN_161437 | _GEN_56443; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_60285 = _GEN_161438 | _GEN_56444; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_60286 = _GEN_161439 | _GEN_56445; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_60287 = _GEN_161440 | _GEN_56446; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_60288 = _GEN_161441 | _GEN_56447; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_60289 = _GEN_161442 | _GEN_56448; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_60290 = _GEN_161443 | _GEN_56449; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_60291 = _GEN_161444 | _GEN_56450; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_60292 = _GEN_161445 | _GEN_56451; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_60293 = _GEN_161446 | _GEN_56452; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_60294 = _GEN_161447 | _GEN_56453; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_60295 = _GEN_161448 | _GEN_56454; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_60296 = _GEN_161449 | _GEN_56455; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_60297 = _GEN_161450 | _GEN_56456; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_60298 = _GEN_161451 | _GEN_56457; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_60299 = _GEN_161452 | _GEN_56458; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_60300 = _GEN_161453 | _GEN_56459; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_60301 = _GEN_161454 | _GEN_56460; // @[Vlflowqueue.scala 197:{51,51}]
  wire [4:0] _GEN_63246 = 5'h0 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_59405; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_63247 = 5'h1 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_59406; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_63248 = 5'h2 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_59407; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_63249 = 5'h3 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_59408; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_63250 = 5'h4 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_59409; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_63251 = 5'h5 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_59410; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_63252 = 5'h6 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_59411; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_63253 = 5'h7 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_59412; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_63254 = 5'h8 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_59413; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_63255 = 5'h9 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_59414; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_63256 = 5'ha == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_59415; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_63257 = 5'hb == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_59416; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_63258 = 5'hc == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_59417; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_63259 = 5'hd == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_59418; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_63260 = 5'he == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_59419; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_63261 = 5'hf == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_59420; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_63262 = 5'h10 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_59421; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_63263 = 5'h11 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_59422; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_63264 = 5'h12 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_59423; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_63265 = 5'h13 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_59424; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_63266 = 5'h14 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_59425; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_63267 = 5'h15 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_59426; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_63268 = 5'h16 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_59427; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_63269 = 5'h17 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_59428; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_63270 = 5'h18 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_59429; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_63271 = 5'h19 == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_59430; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_63272 = 5'h1a == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_59431; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_63273 = 5'h1b == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_59432; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_63274 = 5'h1c == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_59433; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_63275 = 5'h1d == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_59434; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_63276 = 5'h1e == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_59435; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_63277 = 5'h1f == index_0 ? io_loadRegIn_0_bits_uop_robIdx_value : _GEN_59436; // @[Vlflowqueue.scala 198:{51,51}]
  wire [38:0] _GEN_63822 = 5'h0 == index_0 ? vaddr_0 : _GEN_59982; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_63823 = 5'h1 == index_0 ? vaddr_0 : _GEN_59983; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_63824 = 5'h2 == index_0 ? vaddr_0 : _GEN_59984; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_63825 = 5'h3 == index_0 ? vaddr_0 : _GEN_59985; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_63826 = 5'h4 == index_0 ? vaddr_0 : _GEN_59986; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_63827 = 5'h5 == index_0 ? vaddr_0 : _GEN_59987; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_63828 = 5'h6 == index_0 ? vaddr_0 : _GEN_59988; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_63829 = 5'h7 == index_0 ? vaddr_0 : _GEN_59989; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_63830 = 5'h8 == index_0 ? vaddr_0 : _GEN_59990; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_63831 = 5'h9 == index_0 ? vaddr_0 : _GEN_59991; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_63832 = 5'ha == index_0 ? vaddr_0 : _GEN_59992; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_63833 = 5'hb == index_0 ? vaddr_0 : _GEN_59993; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_63834 = 5'hc == index_0 ? vaddr_0 : _GEN_59994; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_63835 = 5'hd == index_0 ? vaddr_0 : _GEN_59995; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_63836 = 5'he == index_0 ? vaddr_0 : _GEN_59996; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_63837 = 5'hf == index_0 ? vaddr_0 : _GEN_59997; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_63838 = 5'h10 == index_0 ? vaddr_0 : _GEN_59998; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_63839 = 5'h11 == index_0 ? vaddr_0 : _GEN_59999; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_63840 = 5'h12 == index_0 ? vaddr_0 : _GEN_60000; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_63841 = 5'h13 == index_0 ? vaddr_0 : _GEN_60001; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_63842 = 5'h14 == index_0 ? vaddr_0 : _GEN_60002; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_63843 = 5'h15 == index_0 ? vaddr_0 : _GEN_60003; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_63844 = 5'h16 == index_0 ? vaddr_0 : _GEN_60004; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_63845 = 5'h17 == index_0 ? vaddr_0 : _GEN_60005; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_63846 = 5'h18 == index_0 ? vaddr_0 : _GEN_60006; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_63847 = 5'h19 == index_0 ? vaddr_0 : _GEN_60007; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_63848 = 5'h1a == index_0 ? vaddr_0 : _GEN_60008; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_63849 = 5'h1b == index_0 ? vaddr_0 : _GEN_60009; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_63850 = 5'h1c == index_0 ? vaddr_0 : _GEN_60010; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_63851 = 5'h1d == index_0 ? vaddr_0 : _GEN_60011; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_63852 = 5'h1e == index_0 ? vaddr_0 : _GEN_60012; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_63853 = 5'h1f == index_0 ? vaddr_0 : _GEN_60013; // @[Vlflowqueue.scala 203:{51,51}]
  wire  _GEN_64495 = 4'h7 < realFlowNum_0 ? _GEN_60270 : _GEN_56429; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_64496 = 4'h7 < realFlowNum_0 ? _GEN_60271 : _GEN_56430; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_64497 = 4'h7 < realFlowNum_0 ? _GEN_60272 : _GEN_56431; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_64498 = 4'h7 < realFlowNum_0 ? _GEN_60273 : _GEN_56432; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_64499 = 4'h7 < realFlowNum_0 ? _GEN_60274 : _GEN_56433; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_64500 = 4'h7 < realFlowNum_0 ? _GEN_60275 : _GEN_56434; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_64501 = 4'h7 < realFlowNum_0 ? _GEN_60276 : _GEN_56435; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_64502 = 4'h7 < realFlowNum_0 ? _GEN_60277 : _GEN_56436; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_64503 = 4'h7 < realFlowNum_0 ? _GEN_60278 : _GEN_56437; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_64504 = 4'h7 < realFlowNum_0 ? _GEN_60279 : _GEN_56438; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_64505 = 4'h7 < realFlowNum_0 ? _GEN_60280 : _GEN_56439; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_64506 = 4'h7 < realFlowNum_0 ? _GEN_60281 : _GEN_56440; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_64507 = 4'h7 < realFlowNum_0 ? _GEN_60282 : _GEN_56441; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_64508 = 4'h7 < realFlowNum_0 ? _GEN_60283 : _GEN_56442; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_64509 = 4'h7 < realFlowNum_0 ? _GEN_60284 : _GEN_56443; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_64510 = 4'h7 < realFlowNum_0 ? _GEN_60285 : _GEN_56444; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_64511 = 4'h7 < realFlowNum_0 ? _GEN_60286 : _GEN_56445; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_64512 = 4'h7 < realFlowNum_0 ? _GEN_60287 : _GEN_56446; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_64513 = 4'h7 < realFlowNum_0 ? _GEN_60288 : _GEN_56447; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_64514 = 4'h7 < realFlowNum_0 ? _GEN_60289 : _GEN_56448; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_64515 = 4'h7 < realFlowNum_0 ? _GEN_60290 : _GEN_56449; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_64516 = 4'h7 < realFlowNum_0 ? _GEN_60291 : _GEN_56450; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_64517 = 4'h7 < realFlowNum_0 ? _GEN_60292 : _GEN_56451; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_64518 = 4'h7 < realFlowNum_0 ? _GEN_60293 : _GEN_56452; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_64519 = 4'h7 < realFlowNum_0 ? _GEN_60294 : _GEN_56453; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_64520 = 4'h7 < realFlowNum_0 ? _GEN_60295 : _GEN_56454; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_64521 = 4'h7 < realFlowNum_0 ? _GEN_60296 : _GEN_56455; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_64522 = 4'h7 < realFlowNum_0 ? _GEN_60297 : _GEN_56456; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_64523 = 4'h7 < realFlowNum_0 ? _GEN_60298 : _GEN_56457; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_64524 = 4'h7 < realFlowNum_0 ? _GEN_60299 : _GEN_56458; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_64525 = 4'h7 < realFlowNum_0 ? _GEN_60300 : _GEN_56459; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_64526 = 4'h7 < realFlowNum_0 ? _GEN_60301 : _GEN_56460; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_67471 = 4'h7 < realFlowNum_0 ? _GEN_63246 : _GEN_59405; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_67472 = 4'h7 < realFlowNum_0 ? _GEN_63247 : _GEN_59406; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_67473 = 4'h7 < realFlowNum_0 ? _GEN_63248 : _GEN_59407; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_67474 = 4'h7 < realFlowNum_0 ? _GEN_63249 : _GEN_59408; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_67475 = 4'h7 < realFlowNum_0 ? _GEN_63250 : _GEN_59409; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_67476 = 4'h7 < realFlowNum_0 ? _GEN_63251 : _GEN_59410; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_67477 = 4'h7 < realFlowNum_0 ? _GEN_63252 : _GEN_59411; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_67478 = 4'h7 < realFlowNum_0 ? _GEN_63253 : _GEN_59412; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_67479 = 4'h7 < realFlowNum_0 ? _GEN_63254 : _GEN_59413; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_67480 = 4'h7 < realFlowNum_0 ? _GEN_63255 : _GEN_59414; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_67481 = 4'h7 < realFlowNum_0 ? _GEN_63256 : _GEN_59415; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_67482 = 4'h7 < realFlowNum_0 ? _GEN_63257 : _GEN_59416; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_67483 = 4'h7 < realFlowNum_0 ? _GEN_63258 : _GEN_59417; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_67484 = 4'h7 < realFlowNum_0 ? _GEN_63259 : _GEN_59418; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_67485 = 4'h7 < realFlowNum_0 ? _GEN_63260 : _GEN_59419; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_67486 = 4'h7 < realFlowNum_0 ? _GEN_63261 : _GEN_59420; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_67487 = 4'h7 < realFlowNum_0 ? _GEN_63262 : _GEN_59421; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_67488 = 4'h7 < realFlowNum_0 ? _GEN_63263 : _GEN_59422; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_67489 = 4'h7 < realFlowNum_0 ? _GEN_63264 : _GEN_59423; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_67490 = 4'h7 < realFlowNum_0 ? _GEN_63265 : _GEN_59424; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_67491 = 4'h7 < realFlowNum_0 ? _GEN_63266 : _GEN_59425; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_67492 = 4'h7 < realFlowNum_0 ? _GEN_63267 : _GEN_59426; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_67493 = 4'h7 < realFlowNum_0 ? _GEN_63268 : _GEN_59427; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_67494 = 4'h7 < realFlowNum_0 ? _GEN_63269 : _GEN_59428; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_67495 = 4'h7 < realFlowNum_0 ? _GEN_63270 : _GEN_59429; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_67496 = 4'h7 < realFlowNum_0 ? _GEN_63271 : _GEN_59430; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_67497 = 4'h7 < realFlowNum_0 ? _GEN_63272 : _GEN_59431; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_67498 = 4'h7 < realFlowNum_0 ? _GEN_63273 : _GEN_59432; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_67499 = 4'h7 < realFlowNum_0 ? _GEN_63274 : _GEN_59433; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_67500 = 4'h7 < realFlowNum_0 ? _GEN_63275 : _GEN_59434; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_67501 = 4'h7 < realFlowNum_0 ? _GEN_63276 : _GEN_59435; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_67502 = 4'h7 < realFlowNum_0 ? _GEN_63277 : _GEN_59436; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_68048 = 4'h7 < realFlowNum_0 ? _GEN_63822 : _GEN_59982; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_68049 = 4'h7 < realFlowNum_0 ? _GEN_63823 : _GEN_59983; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_68050 = 4'h7 < realFlowNum_0 ? _GEN_63824 : _GEN_59984; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_68051 = 4'h7 < realFlowNum_0 ? _GEN_63825 : _GEN_59985; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_68052 = 4'h7 < realFlowNum_0 ? _GEN_63826 : _GEN_59986; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_68053 = 4'h7 < realFlowNum_0 ? _GEN_63827 : _GEN_59987; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_68054 = 4'h7 < realFlowNum_0 ? _GEN_63828 : _GEN_59988; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_68055 = 4'h7 < realFlowNum_0 ? _GEN_63829 : _GEN_59989; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_68056 = 4'h7 < realFlowNum_0 ? _GEN_63830 : _GEN_59990; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_68057 = 4'h7 < realFlowNum_0 ? _GEN_63831 : _GEN_59991; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_68058 = 4'h7 < realFlowNum_0 ? _GEN_63832 : _GEN_59992; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_68059 = 4'h7 < realFlowNum_0 ? _GEN_63833 : _GEN_59993; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_68060 = 4'h7 < realFlowNum_0 ? _GEN_63834 : _GEN_59994; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_68061 = 4'h7 < realFlowNum_0 ? _GEN_63835 : _GEN_59995; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_68062 = 4'h7 < realFlowNum_0 ? _GEN_63836 : _GEN_59996; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_68063 = 4'h7 < realFlowNum_0 ? _GEN_63837 : _GEN_59997; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_68064 = 4'h7 < realFlowNum_0 ? _GEN_63838 : _GEN_59998; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_68065 = 4'h7 < realFlowNum_0 ? _GEN_63839 : _GEN_59999; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_68066 = 4'h7 < realFlowNum_0 ? _GEN_63840 : _GEN_60000; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_68067 = 4'h7 < realFlowNum_0 ? _GEN_63841 : _GEN_60001; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_68068 = 4'h7 < realFlowNum_0 ? _GEN_63842 : _GEN_60002; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_68069 = 4'h7 < realFlowNum_0 ? _GEN_63843 : _GEN_60003; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_68070 = 4'h7 < realFlowNum_0 ? _GEN_63844 : _GEN_60004; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_68071 = 4'h7 < realFlowNum_0 ? _GEN_63845 : _GEN_60005; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_68072 = 4'h7 < realFlowNum_0 ? _GEN_63846 : _GEN_60006; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_68073 = 4'h7 < realFlowNum_0 ? _GEN_63847 : _GEN_60007; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_68074 = 4'h7 < realFlowNum_0 ? _GEN_63848 : _GEN_60008; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_68075 = 4'h7 < realFlowNum_0 ? _GEN_63849 : _GEN_60009; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_68076 = 4'h7 < realFlowNum_0 ? _GEN_63850 : _GEN_60010; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_68077 = 4'h7 < realFlowNum_0 ? _GEN_63851 : _GEN_60011; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_68078 = 4'h7 < realFlowNum_0 ? _GEN_63852 : _GEN_60012; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_68079 = 4'h7 < realFlowNum_0 ? _GEN_63853 : _GEN_60013; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_68336 = _GEN_161423 | _GEN_64495; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_68337 = _GEN_161424 | _GEN_64496; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_68338 = _GEN_161425 | _GEN_64497; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_68339 = _GEN_161426 | _GEN_64498; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_68340 = _GEN_161427 | _GEN_64499; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_68341 = _GEN_161428 | _GEN_64500; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_68342 = _GEN_161429 | _GEN_64501; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_68343 = _GEN_161430 | _GEN_64502; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_68344 = _GEN_161431 | _GEN_64503; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_68345 = _GEN_161432 | _GEN_64504; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_68346 = _GEN_161433 | _GEN_64505; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_68347 = _GEN_161434 | _GEN_64506; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_68348 = _GEN_161435 | _GEN_64507; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_68349 = _GEN_161436 | _GEN_64508; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_68350 = _GEN_161437 | _GEN_64509; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_68351 = _GEN_161438 | _GEN_64510; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_68352 = _GEN_161439 | _GEN_64511; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_68353 = _GEN_161440 | _GEN_64512; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_68354 = _GEN_161441 | _GEN_64513; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_68355 = _GEN_161442 | _GEN_64514; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_68356 = _GEN_161443 | _GEN_64515; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_68357 = _GEN_161444 | _GEN_64516; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_68358 = _GEN_161445 | _GEN_64517; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_68359 = _GEN_161446 | _GEN_64518; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_68360 = _GEN_161447 | _GEN_64519; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_68361 = _GEN_161448 | _GEN_64520; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_68362 = _GEN_161449 | _GEN_64521; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_68363 = _GEN_161450 | _GEN_64522; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_68364 = _GEN_161451 | _GEN_64523; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_68365 = _GEN_161452 | _GEN_64524; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_68366 = _GEN_161453 | _GEN_64525; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_68367 = _GEN_161454 | _GEN_64526; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_72561 = 4'h8 < realFlowNum_0 ? _GEN_68336 : _GEN_64495; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_72562 = 4'h8 < realFlowNum_0 ? _GEN_68337 : _GEN_64496; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_72563 = 4'h8 < realFlowNum_0 ? _GEN_68338 : _GEN_64497; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_72564 = 4'h8 < realFlowNum_0 ? _GEN_68339 : _GEN_64498; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_72565 = 4'h8 < realFlowNum_0 ? _GEN_68340 : _GEN_64499; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_72566 = 4'h8 < realFlowNum_0 ? _GEN_68341 : _GEN_64500; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_72567 = 4'h8 < realFlowNum_0 ? _GEN_68342 : _GEN_64501; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_72568 = 4'h8 < realFlowNum_0 ? _GEN_68343 : _GEN_64502; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_72569 = 4'h8 < realFlowNum_0 ? _GEN_68344 : _GEN_64503; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_72570 = 4'h8 < realFlowNum_0 ? _GEN_68345 : _GEN_64504; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_72571 = 4'h8 < realFlowNum_0 ? _GEN_68346 : _GEN_64505; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_72572 = 4'h8 < realFlowNum_0 ? _GEN_68347 : _GEN_64506; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_72573 = 4'h8 < realFlowNum_0 ? _GEN_68348 : _GEN_64507; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_72574 = 4'h8 < realFlowNum_0 ? _GEN_68349 : _GEN_64508; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_72575 = 4'h8 < realFlowNum_0 ? _GEN_68350 : _GEN_64509; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_72576 = 4'h8 < realFlowNum_0 ? _GEN_68351 : _GEN_64510; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_72577 = 4'h8 < realFlowNum_0 ? _GEN_68352 : _GEN_64511; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_72578 = 4'h8 < realFlowNum_0 ? _GEN_68353 : _GEN_64512; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_72579 = 4'h8 < realFlowNum_0 ? _GEN_68354 : _GEN_64513; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_72580 = 4'h8 < realFlowNum_0 ? _GEN_68355 : _GEN_64514; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_72581 = 4'h8 < realFlowNum_0 ? _GEN_68356 : _GEN_64515; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_72582 = 4'h8 < realFlowNum_0 ? _GEN_68357 : _GEN_64516; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_72583 = 4'h8 < realFlowNum_0 ? _GEN_68358 : _GEN_64517; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_72584 = 4'h8 < realFlowNum_0 ? _GEN_68359 : _GEN_64518; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_72585 = 4'h8 < realFlowNum_0 ? _GEN_68360 : _GEN_64519; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_72586 = 4'h8 < realFlowNum_0 ? _GEN_68361 : _GEN_64520; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_72587 = 4'h8 < realFlowNum_0 ? _GEN_68362 : _GEN_64521; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_72588 = 4'h8 < realFlowNum_0 ? _GEN_68363 : _GEN_64522; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_72589 = 4'h8 < realFlowNum_0 ? _GEN_68364 : _GEN_64523; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_72590 = 4'h8 < realFlowNum_0 ? _GEN_68365 : _GEN_64524; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_72591 = 4'h8 < realFlowNum_0 ? _GEN_68366 : _GEN_64525; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_72592 = 4'h8 < realFlowNum_0 ? _GEN_68367 : _GEN_64526; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_76404 = needAlloc_0 ? _GEN_72561 : flow_entry_valid_0_0; // @[Vlflowqueue.scala 191:25 135:33]
  wire  _GEN_76405 = needAlloc_0 ? _GEN_72562 : flow_entry_valid_0_1; // @[Vlflowqueue.scala 191:25 135:33]
  wire  _GEN_76406 = needAlloc_0 ? _GEN_72563 : flow_entry_valid_0_2; // @[Vlflowqueue.scala 191:25 135:33]
  wire  _GEN_76407 = needAlloc_0 ? _GEN_72564 : flow_entry_valid_0_3; // @[Vlflowqueue.scala 191:25 135:33]
  wire  _GEN_76408 = needAlloc_0 ? _GEN_72565 : flow_entry_valid_0_4; // @[Vlflowqueue.scala 191:25 135:33]
  wire  _GEN_76409 = needAlloc_0 ? _GEN_72566 : flow_entry_valid_0_5; // @[Vlflowqueue.scala 191:25 135:33]
  wire  _GEN_76410 = needAlloc_0 ? _GEN_72567 : flow_entry_valid_0_6; // @[Vlflowqueue.scala 191:25 135:33]
  wire  _GEN_76411 = needAlloc_0 ? _GEN_72568 : flow_entry_valid_0_7; // @[Vlflowqueue.scala 191:25 135:33]
  wire  _GEN_76412 = needAlloc_0 ? _GEN_72569 : flow_entry_valid_0_8; // @[Vlflowqueue.scala 191:25 135:33]
  wire  _GEN_76413 = needAlloc_0 ? _GEN_72570 : flow_entry_valid_0_9; // @[Vlflowqueue.scala 191:25 135:33]
  wire  _GEN_76414 = needAlloc_0 ? _GEN_72571 : flow_entry_valid_0_10; // @[Vlflowqueue.scala 191:25 135:33]
  wire  _GEN_76415 = needAlloc_0 ? _GEN_72572 : flow_entry_valid_0_11; // @[Vlflowqueue.scala 191:25 135:33]
  wire  _GEN_76416 = needAlloc_0 ? _GEN_72573 : flow_entry_valid_0_12; // @[Vlflowqueue.scala 191:25 135:33]
  wire  _GEN_76417 = needAlloc_0 ? _GEN_72574 : flow_entry_valid_0_13; // @[Vlflowqueue.scala 191:25 135:33]
  wire  _GEN_76418 = needAlloc_0 ? _GEN_72575 : flow_entry_valid_0_14; // @[Vlflowqueue.scala 191:25 135:33]
  wire  _GEN_76419 = needAlloc_0 ? _GEN_72576 : flow_entry_valid_0_15; // @[Vlflowqueue.scala 191:25 135:33]
  wire  _GEN_76420 = needAlloc_0 ? _GEN_72577 : flow_entry_valid_0_16; // @[Vlflowqueue.scala 191:25 135:33]
  wire  _GEN_76421 = needAlloc_0 ? _GEN_72578 : flow_entry_valid_0_17; // @[Vlflowqueue.scala 191:25 135:33]
  wire  _GEN_76422 = needAlloc_0 ? _GEN_72579 : flow_entry_valid_0_18; // @[Vlflowqueue.scala 191:25 135:33]
  wire  _GEN_76423 = needAlloc_0 ? _GEN_72580 : flow_entry_valid_0_19; // @[Vlflowqueue.scala 191:25 135:33]
  wire  _GEN_76424 = needAlloc_0 ? _GEN_72581 : flow_entry_valid_0_20; // @[Vlflowqueue.scala 191:25 135:33]
  wire  _GEN_76425 = needAlloc_0 ? _GEN_72582 : flow_entry_valid_0_21; // @[Vlflowqueue.scala 191:25 135:33]
  wire  _GEN_76426 = needAlloc_0 ? _GEN_72583 : flow_entry_valid_0_22; // @[Vlflowqueue.scala 191:25 135:33]
  wire  _GEN_76427 = needAlloc_0 ? _GEN_72584 : flow_entry_valid_0_23; // @[Vlflowqueue.scala 191:25 135:33]
  wire  _GEN_76428 = needAlloc_0 ? _GEN_72585 : flow_entry_valid_0_24; // @[Vlflowqueue.scala 191:25 135:33]
  wire  _GEN_76429 = needAlloc_0 ? _GEN_72586 : flow_entry_valid_0_25; // @[Vlflowqueue.scala 191:25 135:33]
  wire  _GEN_76430 = needAlloc_0 ? _GEN_72587 : flow_entry_valid_0_26; // @[Vlflowqueue.scala 191:25 135:33]
  wire  _GEN_76431 = needAlloc_0 ? _GEN_72588 : flow_entry_valid_0_27; // @[Vlflowqueue.scala 191:25 135:33]
  wire  _GEN_76432 = needAlloc_0 ? _GEN_72589 : flow_entry_valid_0_28; // @[Vlflowqueue.scala 191:25 135:33]
  wire  _GEN_76433 = needAlloc_0 ? _GEN_72590 : flow_entry_valid_0_29; // @[Vlflowqueue.scala 191:25 135:33]
  wire  _GEN_76434 = needAlloc_0 ? _GEN_72591 : flow_entry_valid_0_30; // @[Vlflowqueue.scala 191:25 135:33]
  wire  _GEN_76435 = needAlloc_0 ? _GEN_72592 : flow_entry_valid_0_31; // @[Vlflowqueue.scala 191:25 135:33]
  wire [4:0] _index_1_T_17 = enqPtr_1_value + 5'h8; // @[Vlflowqueue.scala 195:39]
  wire [4:0] _index_1_T_15 = enqPtr_1_value + 5'h7; // @[Vlflowqueue.scala 195:39]
  wire [4:0] _index_1_T_13 = enqPtr_1_value + 5'h6; // @[Vlflowqueue.scala 195:39]
  wire [4:0] _index_1_T_11 = enqPtr_1_value + 5'h5; // @[Vlflowqueue.scala 195:39]
  wire [4:0] _index_1_T_9 = enqPtr_1_value + 5'h4; // @[Vlflowqueue.scala 195:39]
  wire [4:0] _index_1_T_7 = enqPtr_1_value + 5'h3; // @[Vlflowqueue.scala 195:39]
  wire [4:0] _index_1_T_5 = enqPtr_1_value + 5'h2; // @[Vlflowqueue.scala 195:39]
  wire [4:0] _index_1_T_3 = enqPtr_1_value + 5'h1; // @[Vlflowqueue.scala 195:39]
  wire [4:0] _GEN_96343 = 4'h1 < realFlowNum_1 ? _index_1_T_3 : _GEN_161420[4:0]; // @[Vlflowqueue.scala 194:37 195:20]
  wire [4:0] _GEN_104409 = 4'h2 < realFlowNum_1 ? _index_1_T_5 : _GEN_96343; // @[Vlflowqueue.scala 194:37 195:20]
  wire [4:0] _GEN_112475 = 4'h3 < realFlowNum_1 ? _index_1_T_7 : _GEN_104409; // @[Vlflowqueue.scala 194:37 195:20]
  wire [4:0] _GEN_120541 = 4'h4 < realFlowNum_1 ? _index_1_T_9 : _GEN_112475; // @[Vlflowqueue.scala 194:37 195:20]
  wire [4:0] _GEN_128607 = 4'h5 < realFlowNum_1 ? _index_1_T_11 : _GEN_120541; // @[Vlflowqueue.scala 194:37 195:20]
  wire [4:0] _GEN_136673 = 4'h6 < realFlowNum_1 ? _index_1_T_13 : _GEN_128607; // @[Vlflowqueue.scala 194:37 195:20]
  wire [4:0] _GEN_144739 = 4'h7 < realFlowNum_1 ? _index_1_T_15 : _GEN_136673; // @[Vlflowqueue.scala 194:37 195:20]
  wire [4:0] index_1 = 4'h8 < realFlowNum_1 ? _index_1_T_17 : _GEN_144739; // @[Vlflowqueue.scala 194:37 195:20]
  wire  _GEN_162068 = 5'h0 == index_1; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_84053 = 5'h0 == index_1 | flow_entry_valid_1_0; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_162069 = 5'h1 == index_1; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_84054 = 5'h1 == index_1 | flow_entry_valid_1_1; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_162070 = 5'h2 == index_1; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_84055 = 5'h2 == index_1 | flow_entry_valid_1_2; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_162071 = 5'h3 == index_1; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_84056 = 5'h3 == index_1 | flow_entry_valid_1_3; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_162072 = 5'h4 == index_1; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_84057 = 5'h4 == index_1 | flow_entry_valid_1_4; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_162073 = 5'h5 == index_1; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_84058 = 5'h5 == index_1 | flow_entry_valid_1_5; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_162074 = 5'h6 == index_1; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_84059 = 5'h6 == index_1 | flow_entry_valid_1_6; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_162075 = 5'h7 == index_1; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_84060 = 5'h7 == index_1 | flow_entry_valid_1_7; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_162076 = 5'h8 == index_1; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_84061 = 5'h8 == index_1 | flow_entry_valid_1_8; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_162077 = 5'h9 == index_1; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_84062 = 5'h9 == index_1 | flow_entry_valid_1_9; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_162078 = 5'ha == index_1; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_84063 = 5'ha == index_1 | flow_entry_valid_1_10; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_162079 = 5'hb == index_1; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_84064 = 5'hb == index_1 | flow_entry_valid_1_11; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_162080 = 5'hc == index_1; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_84065 = 5'hc == index_1 | flow_entry_valid_1_12; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_162081 = 5'hd == index_1; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_84066 = 5'hd == index_1 | flow_entry_valid_1_13; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_162082 = 5'he == index_1; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_84067 = 5'he == index_1 | flow_entry_valid_1_14; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_162083 = 5'hf == index_1; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_84068 = 5'hf == index_1 | flow_entry_valid_1_15; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_162084 = 5'h10 == index_1; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_84069 = 5'h10 == index_1 | flow_entry_valid_1_16; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_162085 = 5'h11 == index_1; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_84070 = 5'h11 == index_1 | flow_entry_valid_1_17; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_162086 = 5'h12 == index_1; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_84071 = 5'h12 == index_1 | flow_entry_valid_1_18; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_162087 = 5'h13 == index_1; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_84072 = 5'h13 == index_1 | flow_entry_valid_1_19; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_162088 = 5'h14 == index_1; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_84073 = 5'h14 == index_1 | flow_entry_valid_1_20; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_162089 = 5'h15 == index_1; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_84074 = 5'h15 == index_1 | flow_entry_valid_1_21; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_162090 = 5'h16 == index_1; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_84075 = 5'h16 == index_1 | flow_entry_valid_1_22; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_162091 = 5'h17 == index_1; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_84076 = 5'h17 == index_1 | flow_entry_valid_1_23; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_162092 = 5'h18 == index_1; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_84077 = 5'h18 == index_1 | flow_entry_valid_1_24; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_162093 = 5'h19 == index_1; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_84078 = 5'h19 == index_1 | flow_entry_valid_1_25; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_162094 = 5'h1a == index_1; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_84079 = 5'h1a == index_1 | flow_entry_valid_1_26; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_162095 = 5'h1b == index_1; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_84080 = 5'h1b == index_1 | flow_entry_valid_1_27; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_162096 = 5'h1c == index_1; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_84081 = 5'h1c == index_1 | flow_entry_valid_1_28; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_162097 = 5'h1d == index_1; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_84082 = 5'h1d == index_1 | flow_entry_valid_1_29; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_162098 = 5'h1e == index_1; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_84083 = 5'h1e == index_1 | flow_entry_valid_1_30; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_162099 = 5'h1f == index_1; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire  _GEN_84084 = 5'h1f == index_1 | flow_entry_valid_1_31; // @[Vlflowqueue.scala 135:33 197:{51,51}]
  wire [4:0] _GEN_87029 = 5'h0 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : flow_entry_1_0_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 198:{51,51}]
  wire [4:0] _GEN_87030 = 5'h1 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : flow_entry_1_1_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 198:{51,51}]
  wire [4:0] _GEN_87031 = 5'h2 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : flow_entry_1_2_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 198:{51,51}]
  wire [4:0] _GEN_87032 = 5'h3 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : flow_entry_1_3_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 198:{51,51}]
  wire [4:0] _GEN_87033 = 5'h4 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : flow_entry_1_4_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 198:{51,51}]
  wire [4:0] _GEN_87034 = 5'h5 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : flow_entry_1_5_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 198:{51,51}]
  wire [4:0] _GEN_87035 = 5'h6 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : flow_entry_1_6_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 198:{51,51}]
  wire [4:0] _GEN_87036 = 5'h7 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : flow_entry_1_7_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 198:{51,51}]
  wire [4:0] _GEN_87037 = 5'h8 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : flow_entry_1_8_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 198:{51,51}]
  wire [4:0] _GEN_87038 = 5'h9 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : flow_entry_1_9_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 198:{51,51}]
  wire [4:0] _GEN_87039 = 5'ha == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : flow_entry_1_10_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 198:{51,51}]
  wire [4:0] _GEN_87040 = 5'hb == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : flow_entry_1_11_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 198:{51,51}]
  wire [4:0] _GEN_87041 = 5'hc == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : flow_entry_1_12_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 198:{51,51}]
  wire [4:0] _GEN_87042 = 5'hd == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : flow_entry_1_13_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 198:{51,51}]
  wire [4:0] _GEN_87043 = 5'he == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : flow_entry_1_14_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 198:{51,51}]
  wire [4:0] _GEN_87044 = 5'hf == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : flow_entry_1_15_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 198:{51,51}]
  wire [4:0] _GEN_87045 = 5'h10 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : flow_entry_1_16_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 198:{51,51}]
  wire [4:0] _GEN_87046 = 5'h11 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : flow_entry_1_17_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 198:{51,51}]
  wire [4:0] _GEN_87047 = 5'h12 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : flow_entry_1_18_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 198:{51,51}]
  wire [4:0] _GEN_87048 = 5'h13 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : flow_entry_1_19_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 198:{51,51}]
  wire [4:0] _GEN_87049 = 5'h14 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : flow_entry_1_20_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 198:{51,51}]
  wire [4:0] _GEN_87050 = 5'h15 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : flow_entry_1_21_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 198:{51,51}]
  wire [4:0] _GEN_87051 = 5'h16 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : flow_entry_1_22_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 198:{51,51}]
  wire [4:0] _GEN_87052 = 5'h17 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : flow_entry_1_23_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 198:{51,51}]
  wire [4:0] _GEN_87053 = 5'h18 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : flow_entry_1_24_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 198:{51,51}]
  wire [4:0] _GEN_87054 = 5'h19 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : flow_entry_1_25_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 198:{51,51}]
  wire [4:0] _GEN_87055 = 5'h1a == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : flow_entry_1_26_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 198:{51,51}]
  wire [4:0] _GEN_87056 = 5'h1b == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : flow_entry_1_27_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 198:{51,51}]
  wire [4:0] _GEN_87057 = 5'h1c == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : flow_entry_1_28_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 198:{51,51}]
  wire [4:0] _GEN_87058 = 5'h1d == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : flow_entry_1_29_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 198:{51,51}]
  wire [4:0] _GEN_87059 = 5'h1e == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : flow_entry_1_30_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 198:{51,51}]
  wire [4:0] _GEN_87060 = 5'h1f == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : flow_entry_1_31_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 198:{51,51}]
  wire [39:0] _vaddr_1_T_1 = {{1'd0}, io_loadRegIn_1_bits_baseaddr}; // @[Vlflowqueue.scala 91:32]
  wire [38:0] _vaddr_1_T_162 = io_loadRegIn_1_bits_baseaddr + 39'h80; // @[Vlflowqueue.scala 91:32]
  wire [38:0] _vaddr_1_T_142 = io_loadRegIn_1_bits_baseaddr + 39'h70; // @[Vlflowqueue.scala 91:32]
  wire [38:0] _vaddr_1_T_122 = io_loadRegIn_1_bits_baseaddr + 39'h60; // @[Vlflowqueue.scala 91:32]
  wire [38:0] _vaddr_1_T_102 = io_loadRegIn_1_bits_baseaddr + 39'h50; // @[Vlflowqueue.scala 91:32]
  wire [38:0] _vaddr_1_T_82 = io_loadRegIn_1_bits_baseaddr + 39'h40; // @[Vlflowqueue.scala 91:32]
  wire [38:0] _vaddr_1_T_62 = io_loadRegIn_1_bits_baseaddr + 39'h30; // @[Vlflowqueue.scala 91:32]
  wire [38:0] _vaddr_1_T_42 = io_loadRegIn_1_bits_baseaddr + 39'h20; // @[Vlflowqueue.scala 91:32]
  wire [38:0] _vaddr_1_T_22 = io_loadRegIn_1_bits_baseaddr + 39'h10; // @[Vlflowqueue.scala 91:32]
  wire [38:0] _GEN_99864 = 4'h1 < realFlowNum_1 ? _vaddr_1_T_22 : _vaddr_1_T_1[38:0]; // @[Vlflowqueue.scala 194:37 201:51]
  wire [38:0] _GEN_107930 = 4'h2 < realFlowNum_1 ? _vaddr_1_T_42 : _GEN_99864; // @[Vlflowqueue.scala 194:37 201:51]
  wire [38:0] _GEN_115996 = 4'h3 < realFlowNum_1 ? _vaddr_1_T_62 : _GEN_107930; // @[Vlflowqueue.scala 194:37 201:51]
  wire [38:0] _GEN_124062 = 4'h4 < realFlowNum_1 ? _vaddr_1_T_82 : _GEN_115996; // @[Vlflowqueue.scala 194:37 201:51]
  wire [38:0] _GEN_132128 = 4'h5 < realFlowNum_1 ? _vaddr_1_T_102 : _GEN_124062; // @[Vlflowqueue.scala 194:37 201:51]
  wire [38:0] _GEN_140194 = 4'h6 < realFlowNum_1 ? _vaddr_1_T_122 : _GEN_132128; // @[Vlflowqueue.scala 194:37 201:51]
  wire [38:0] _GEN_148260 = 4'h7 < realFlowNum_1 ? _vaddr_1_T_142 : _GEN_140194; // @[Vlflowqueue.scala 194:37 201:51]
  wire [38:0] vaddr_1 = 4'h8 < realFlowNum_1 ? _vaddr_1_T_162 : _GEN_148260; // @[Vlflowqueue.scala 194:37 201:51]
  wire [38:0] _GEN_87605 = 5'h0 == index_1 ? vaddr_1 : flow_entry_1_0_vaddr; // @[Vlflowqueue.scala 134:29 203:{51,51}]
  wire [38:0] _GEN_87606 = 5'h1 == index_1 ? vaddr_1 : flow_entry_1_1_vaddr; // @[Vlflowqueue.scala 134:29 203:{51,51}]
  wire [38:0] _GEN_87607 = 5'h2 == index_1 ? vaddr_1 : flow_entry_1_2_vaddr; // @[Vlflowqueue.scala 134:29 203:{51,51}]
  wire [38:0] _GEN_87608 = 5'h3 == index_1 ? vaddr_1 : flow_entry_1_3_vaddr; // @[Vlflowqueue.scala 134:29 203:{51,51}]
  wire [38:0] _GEN_87609 = 5'h4 == index_1 ? vaddr_1 : flow_entry_1_4_vaddr; // @[Vlflowqueue.scala 134:29 203:{51,51}]
  wire [38:0] _GEN_87610 = 5'h5 == index_1 ? vaddr_1 : flow_entry_1_5_vaddr; // @[Vlflowqueue.scala 134:29 203:{51,51}]
  wire [38:0] _GEN_87611 = 5'h6 == index_1 ? vaddr_1 : flow_entry_1_6_vaddr; // @[Vlflowqueue.scala 134:29 203:{51,51}]
  wire [38:0] _GEN_87612 = 5'h7 == index_1 ? vaddr_1 : flow_entry_1_7_vaddr; // @[Vlflowqueue.scala 134:29 203:{51,51}]
  wire [38:0] _GEN_87613 = 5'h8 == index_1 ? vaddr_1 : flow_entry_1_8_vaddr; // @[Vlflowqueue.scala 134:29 203:{51,51}]
  wire [38:0] _GEN_87614 = 5'h9 == index_1 ? vaddr_1 : flow_entry_1_9_vaddr; // @[Vlflowqueue.scala 134:29 203:{51,51}]
  wire [38:0] _GEN_87615 = 5'ha == index_1 ? vaddr_1 : flow_entry_1_10_vaddr; // @[Vlflowqueue.scala 134:29 203:{51,51}]
  wire [38:0] _GEN_87616 = 5'hb == index_1 ? vaddr_1 : flow_entry_1_11_vaddr; // @[Vlflowqueue.scala 134:29 203:{51,51}]
  wire [38:0] _GEN_87617 = 5'hc == index_1 ? vaddr_1 : flow_entry_1_12_vaddr; // @[Vlflowqueue.scala 134:29 203:{51,51}]
  wire [38:0] _GEN_87618 = 5'hd == index_1 ? vaddr_1 : flow_entry_1_13_vaddr; // @[Vlflowqueue.scala 134:29 203:{51,51}]
  wire [38:0] _GEN_87619 = 5'he == index_1 ? vaddr_1 : flow_entry_1_14_vaddr; // @[Vlflowqueue.scala 134:29 203:{51,51}]
  wire [38:0] _GEN_87620 = 5'hf == index_1 ? vaddr_1 : flow_entry_1_15_vaddr; // @[Vlflowqueue.scala 134:29 203:{51,51}]
  wire [38:0] _GEN_87621 = 5'h10 == index_1 ? vaddr_1 : flow_entry_1_16_vaddr; // @[Vlflowqueue.scala 134:29 203:{51,51}]
  wire [38:0] _GEN_87622 = 5'h11 == index_1 ? vaddr_1 : flow_entry_1_17_vaddr; // @[Vlflowqueue.scala 134:29 203:{51,51}]
  wire [38:0] _GEN_87623 = 5'h12 == index_1 ? vaddr_1 : flow_entry_1_18_vaddr; // @[Vlflowqueue.scala 134:29 203:{51,51}]
  wire [38:0] _GEN_87624 = 5'h13 == index_1 ? vaddr_1 : flow_entry_1_19_vaddr; // @[Vlflowqueue.scala 134:29 203:{51,51}]
  wire [38:0] _GEN_87625 = 5'h14 == index_1 ? vaddr_1 : flow_entry_1_20_vaddr; // @[Vlflowqueue.scala 134:29 203:{51,51}]
  wire [38:0] _GEN_87626 = 5'h15 == index_1 ? vaddr_1 : flow_entry_1_21_vaddr; // @[Vlflowqueue.scala 134:29 203:{51,51}]
  wire [38:0] _GEN_87627 = 5'h16 == index_1 ? vaddr_1 : flow_entry_1_22_vaddr; // @[Vlflowqueue.scala 134:29 203:{51,51}]
  wire [38:0] _GEN_87628 = 5'h17 == index_1 ? vaddr_1 : flow_entry_1_23_vaddr; // @[Vlflowqueue.scala 134:29 203:{51,51}]
  wire [38:0] _GEN_87629 = 5'h18 == index_1 ? vaddr_1 : flow_entry_1_24_vaddr; // @[Vlflowqueue.scala 134:29 203:{51,51}]
  wire [38:0] _GEN_87630 = 5'h19 == index_1 ? vaddr_1 : flow_entry_1_25_vaddr; // @[Vlflowqueue.scala 134:29 203:{51,51}]
  wire [38:0] _GEN_87631 = 5'h1a == index_1 ? vaddr_1 : flow_entry_1_26_vaddr; // @[Vlflowqueue.scala 134:29 203:{51,51}]
  wire [38:0] _GEN_87632 = 5'h1b == index_1 ? vaddr_1 : flow_entry_1_27_vaddr; // @[Vlflowqueue.scala 134:29 203:{51,51}]
  wire [38:0] _GEN_87633 = 5'h1c == index_1 ? vaddr_1 : flow_entry_1_28_vaddr; // @[Vlflowqueue.scala 134:29 203:{51,51}]
  wire [38:0] _GEN_87634 = 5'h1d == index_1 ? vaddr_1 : flow_entry_1_29_vaddr; // @[Vlflowqueue.scala 134:29 203:{51,51}]
  wire [38:0] _GEN_87635 = 5'h1e == index_1 ? vaddr_1 : flow_entry_1_30_vaddr; // @[Vlflowqueue.scala 134:29 203:{51,51}]
  wire [38:0] _GEN_87636 = 5'h1f == index_1 ? vaddr_1 : flow_entry_1_31_vaddr; // @[Vlflowqueue.scala 134:29 203:{51,51}]
  wire  _GEN_88278 = 4'h0 < realFlowNum_1 ? _GEN_84053 : flow_entry_valid_1_0; // @[Vlflowqueue.scala 135:33 194:37]
  wire  _GEN_88279 = 4'h0 < realFlowNum_1 ? _GEN_84054 : flow_entry_valid_1_1; // @[Vlflowqueue.scala 135:33 194:37]
  wire  _GEN_88280 = 4'h0 < realFlowNum_1 ? _GEN_84055 : flow_entry_valid_1_2; // @[Vlflowqueue.scala 135:33 194:37]
  wire  _GEN_88281 = 4'h0 < realFlowNum_1 ? _GEN_84056 : flow_entry_valid_1_3; // @[Vlflowqueue.scala 135:33 194:37]
  wire  _GEN_88282 = 4'h0 < realFlowNum_1 ? _GEN_84057 : flow_entry_valid_1_4; // @[Vlflowqueue.scala 135:33 194:37]
  wire  _GEN_88283 = 4'h0 < realFlowNum_1 ? _GEN_84058 : flow_entry_valid_1_5; // @[Vlflowqueue.scala 135:33 194:37]
  wire  _GEN_88284 = 4'h0 < realFlowNum_1 ? _GEN_84059 : flow_entry_valid_1_6; // @[Vlflowqueue.scala 135:33 194:37]
  wire  _GEN_88285 = 4'h0 < realFlowNum_1 ? _GEN_84060 : flow_entry_valid_1_7; // @[Vlflowqueue.scala 135:33 194:37]
  wire  _GEN_88286 = 4'h0 < realFlowNum_1 ? _GEN_84061 : flow_entry_valid_1_8; // @[Vlflowqueue.scala 135:33 194:37]
  wire  _GEN_88287 = 4'h0 < realFlowNum_1 ? _GEN_84062 : flow_entry_valid_1_9; // @[Vlflowqueue.scala 135:33 194:37]
  wire  _GEN_88288 = 4'h0 < realFlowNum_1 ? _GEN_84063 : flow_entry_valid_1_10; // @[Vlflowqueue.scala 135:33 194:37]
  wire  _GEN_88289 = 4'h0 < realFlowNum_1 ? _GEN_84064 : flow_entry_valid_1_11; // @[Vlflowqueue.scala 135:33 194:37]
  wire  _GEN_88290 = 4'h0 < realFlowNum_1 ? _GEN_84065 : flow_entry_valid_1_12; // @[Vlflowqueue.scala 135:33 194:37]
  wire  _GEN_88291 = 4'h0 < realFlowNum_1 ? _GEN_84066 : flow_entry_valid_1_13; // @[Vlflowqueue.scala 135:33 194:37]
  wire  _GEN_88292 = 4'h0 < realFlowNum_1 ? _GEN_84067 : flow_entry_valid_1_14; // @[Vlflowqueue.scala 135:33 194:37]
  wire  _GEN_88293 = 4'h0 < realFlowNum_1 ? _GEN_84068 : flow_entry_valid_1_15; // @[Vlflowqueue.scala 135:33 194:37]
  wire  _GEN_88294 = 4'h0 < realFlowNum_1 ? _GEN_84069 : flow_entry_valid_1_16; // @[Vlflowqueue.scala 135:33 194:37]
  wire  _GEN_88295 = 4'h0 < realFlowNum_1 ? _GEN_84070 : flow_entry_valid_1_17; // @[Vlflowqueue.scala 135:33 194:37]
  wire  _GEN_88296 = 4'h0 < realFlowNum_1 ? _GEN_84071 : flow_entry_valid_1_18; // @[Vlflowqueue.scala 135:33 194:37]
  wire  _GEN_88297 = 4'h0 < realFlowNum_1 ? _GEN_84072 : flow_entry_valid_1_19; // @[Vlflowqueue.scala 135:33 194:37]
  wire  _GEN_88298 = 4'h0 < realFlowNum_1 ? _GEN_84073 : flow_entry_valid_1_20; // @[Vlflowqueue.scala 135:33 194:37]
  wire  _GEN_88299 = 4'h0 < realFlowNum_1 ? _GEN_84074 : flow_entry_valid_1_21; // @[Vlflowqueue.scala 135:33 194:37]
  wire  _GEN_88300 = 4'h0 < realFlowNum_1 ? _GEN_84075 : flow_entry_valid_1_22; // @[Vlflowqueue.scala 135:33 194:37]
  wire  _GEN_88301 = 4'h0 < realFlowNum_1 ? _GEN_84076 : flow_entry_valid_1_23; // @[Vlflowqueue.scala 135:33 194:37]
  wire  _GEN_88302 = 4'h0 < realFlowNum_1 ? _GEN_84077 : flow_entry_valid_1_24; // @[Vlflowqueue.scala 135:33 194:37]
  wire  _GEN_88303 = 4'h0 < realFlowNum_1 ? _GEN_84078 : flow_entry_valid_1_25; // @[Vlflowqueue.scala 135:33 194:37]
  wire  _GEN_88304 = 4'h0 < realFlowNum_1 ? _GEN_84079 : flow_entry_valid_1_26; // @[Vlflowqueue.scala 135:33 194:37]
  wire  _GEN_88305 = 4'h0 < realFlowNum_1 ? _GEN_84080 : flow_entry_valid_1_27; // @[Vlflowqueue.scala 135:33 194:37]
  wire  _GEN_88306 = 4'h0 < realFlowNum_1 ? _GEN_84081 : flow_entry_valid_1_28; // @[Vlflowqueue.scala 135:33 194:37]
  wire  _GEN_88307 = 4'h0 < realFlowNum_1 ? _GEN_84082 : flow_entry_valid_1_29; // @[Vlflowqueue.scala 135:33 194:37]
  wire  _GEN_88308 = 4'h0 < realFlowNum_1 ? _GEN_84083 : flow_entry_valid_1_30; // @[Vlflowqueue.scala 135:33 194:37]
  wire  _GEN_88309 = 4'h0 < realFlowNum_1 ? _GEN_84084 : flow_entry_valid_1_31; // @[Vlflowqueue.scala 135:33 194:37]
  wire [4:0] _GEN_91254 = 4'h0 < realFlowNum_1 ? _GEN_87029 : flow_entry_1_0_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 194:37]
  wire [4:0] _GEN_91255 = 4'h0 < realFlowNum_1 ? _GEN_87030 : flow_entry_1_1_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 194:37]
  wire [4:0] _GEN_91256 = 4'h0 < realFlowNum_1 ? _GEN_87031 : flow_entry_1_2_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 194:37]
  wire [4:0] _GEN_91257 = 4'h0 < realFlowNum_1 ? _GEN_87032 : flow_entry_1_3_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 194:37]
  wire [4:0] _GEN_91258 = 4'h0 < realFlowNum_1 ? _GEN_87033 : flow_entry_1_4_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 194:37]
  wire [4:0] _GEN_91259 = 4'h0 < realFlowNum_1 ? _GEN_87034 : flow_entry_1_5_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 194:37]
  wire [4:0] _GEN_91260 = 4'h0 < realFlowNum_1 ? _GEN_87035 : flow_entry_1_6_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 194:37]
  wire [4:0] _GEN_91261 = 4'h0 < realFlowNum_1 ? _GEN_87036 : flow_entry_1_7_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 194:37]
  wire [4:0] _GEN_91262 = 4'h0 < realFlowNum_1 ? _GEN_87037 : flow_entry_1_8_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 194:37]
  wire [4:0] _GEN_91263 = 4'h0 < realFlowNum_1 ? _GEN_87038 : flow_entry_1_9_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 194:37]
  wire [4:0] _GEN_91264 = 4'h0 < realFlowNum_1 ? _GEN_87039 : flow_entry_1_10_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 194:37]
  wire [4:0] _GEN_91265 = 4'h0 < realFlowNum_1 ? _GEN_87040 : flow_entry_1_11_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 194:37]
  wire [4:0] _GEN_91266 = 4'h0 < realFlowNum_1 ? _GEN_87041 : flow_entry_1_12_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 194:37]
  wire [4:0] _GEN_91267 = 4'h0 < realFlowNum_1 ? _GEN_87042 : flow_entry_1_13_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 194:37]
  wire [4:0] _GEN_91268 = 4'h0 < realFlowNum_1 ? _GEN_87043 : flow_entry_1_14_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 194:37]
  wire [4:0] _GEN_91269 = 4'h0 < realFlowNum_1 ? _GEN_87044 : flow_entry_1_15_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 194:37]
  wire [4:0] _GEN_91270 = 4'h0 < realFlowNum_1 ? _GEN_87045 : flow_entry_1_16_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 194:37]
  wire [4:0] _GEN_91271 = 4'h0 < realFlowNum_1 ? _GEN_87046 : flow_entry_1_17_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 194:37]
  wire [4:0] _GEN_91272 = 4'h0 < realFlowNum_1 ? _GEN_87047 : flow_entry_1_18_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 194:37]
  wire [4:0] _GEN_91273 = 4'h0 < realFlowNum_1 ? _GEN_87048 : flow_entry_1_19_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 194:37]
  wire [4:0] _GEN_91274 = 4'h0 < realFlowNum_1 ? _GEN_87049 : flow_entry_1_20_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 194:37]
  wire [4:0] _GEN_91275 = 4'h0 < realFlowNum_1 ? _GEN_87050 : flow_entry_1_21_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 194:37]
  wire [4:0] _GEN_91276 = 4'h0 < realFlowNum_1 ? _GEN_87051 : flow_entry_1_22_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 194:37]
  wire [4:0] _GEN_91277 = 4'h0 < realFlowNum_1 ? _GEN_87052 : flow_entry_1_23_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 194:37]
  wire [4:0] _GEN_91278 = 4'h0 < realFlowNum_1 ? _GEN_87053 : flow_entry_1_24_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 194:37]
  wire [4:0] _GEN_91279 = 4'h0 < realFlowNum_1 ? _GEN_87054 : flow_entry_1_25_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 194:37]
  wire [4:0] _GEN_91280 = 4'h0 < realFlowNum_1 ? _GEN_87055 : flow_entry_1_26_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 194:37]
  wire [4:0] _GEN_91281 = 4'h0 < realFlowNum_1 ? _GEN_87056 : flow_entry_1_27_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 194:37]
  wire [4:0] _GEN_91282 = 4'h0 < realFlowNum_1 ? _GEN_87057 : flow_entry_1_28_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 194:37]
  wire [4:0] _GEN_91283 = 4'h0 < realFlowNum_1 ? _GEN_87058 : flow_entry_1_29_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 194:37]
  wire [4:0] _GEN_91284 = 4'h0 < realFlowNum_1 ? _GEN_87059 : flow_entry_1_30_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 194:37]
  wire [4:0] _GEN_91285 = 4'h0 < realFlowNum_1 ? _GEN_87060 : flow_entry_1_31_uop_robIdx_value; // @[Vlflowqueue.scala 134:29 194:37]
  wire [38:0] _GEN_91831 = 4'h0 < realFlowNum_1 ? _GEN_87605 : flow_entry_1_0_vaddr; // @[Vlflowqueue.scala 134:29 194:37]
  wire [38:0] _GEN_91832 = 4'h0 < realFlowNum_1 ? _GEN_87606 : flow_entry_1_1_vaddr; // @[Vlflowqueue.scala 134:29 194:37]
  wire [38:0] _GEN_91833 = 4'h0 < realFlowNum_1 ? _GEN_87607 : flow_entry_1_2_vaddr; // @[Vlflowqueue.scala 134:29 194:37]
  wire [38:0] _GEN_91834 = 4'h0 < realFlowNum_1 ? _GEN_87608 : flow_entry_1_3_vaddr; // @[Vlflowqueue.scala 134:29 194:37]
  wire [38:0] _GEN_91835 = 4'h0 < realFlowNum_1 ? _GEN_87609 : flow_entry_1_4_vaddr; // @[Vlflowqueue.scala 134:29 194:37]
  wire [38:0] _GEN_91836 = 4'h0 < realFlowNum_1 ? _GEN_87610 : flow_entry_1_5_vaddr; // @[Vlflowqueue.scala 134:29 194:37]
  wire [38:0] _GEN_91837 = 4'h0 < realFlowNum_1 ? _GEN_87611 : flow_entry_1_6_vaddr; // @[Vlflowqueue.scala 134:29 194:37]
  wire [38:0] _GEN_91838 = 4'h0 < realFlowNum_1 ? _GEN_87612 : flow_entry_1_7_vaddr; // @[Vlflowqueue.scala 134:29 194:37]
  wire [38:0] _GEN_91839 = 4'h0 < realFlowNum_1 ? _GEN_87613 : flow_entry_1_8_vaddr; // @[Vlflowqueue.scala 134:29 194:37]
  wire [38:0] _GEN_91840 = 4'h0 < realFlowNum_1 ? _GEN_87614 : flow_entry_1_9_vaddr; // @[Vlflowqueue.scala 134:29 194:37]
  wire [38:0] _GEN_91841 = 4'h0 < realFlowNum_1 ? _GEN_87615 : flow_entry_1_10_vaddr; // @[Vlflowqueue.scala 134:29 194:37]
  wire [38:0] _GEN_91842 = 4'h0 < realFlowNum_1 ? _GEN_87616 : flow_entry_1_11_vaddr; // @[Vlflowqueue.scala 134:29 194:37]
  wire [38:0] _GEN_91843 = 4'h0 < realFlowNum_1 ? _GEN_87617 : flow_entry_1_12_vaddr; // @[Vlflowqueue.scala 134:29 194:37]
  wire [38:0] _GEN_91844 = 4'h0 < realFlowNum_1 ? _GEN_87618 : flow_entry_1_13_vaddr; // @[Vlflowqueue.scala 134:29 194:37]
  wire [38:0] _GEN_91845 = 4'h0 < realFlowNum_1 ? _GEN_87619 : flow_entry_1_14_vaddr; // @[Vlflowqueue.scala 134:29 194:37]
  wire [38:0] _GEN_91846 = 4'h0 < realFlowNum_1 ? _GEN_87620 : flow_entry_1_15_vaddr; // @[Vlflowqueue.scala 134:29 194:37]
  wire [38:0] _GEN_91847 = 4'h0 < realFlowNum_1 ? _GEN_87621 : flow_entry_1_16_vaddr; // @[Vlflowqueue.scala 134:29 194:37]
  wire [38:0] _GEN_91848 = 4'h0 < realFlowNum_1 ? _GEN_87622 : flow_entry_1_17_vaddr; // @[Vlflowqueue.scala 134:29 194:37]
  wire [38:0] _GEN_91849 = 4'h0 < realFlowNum_1 ? _GEN_87623 : flow_entry_1_18_vaddr; // @[Vlflowqueue.scala 134:29 194:37]
  wire [38:0] _GEN_91850 = 4'h0 < realFlowNum_1 ? _GEN_87624 : flow_entry_1_19_vaddr; // @[Vlflowqueue.scala 134:29 194:37]
  wire [38:0] _GEN_91851 = 4'h0 < realFlowNum_1 ? _GEN_87625 : flow_entry_1_20_vaddr; // @[Vlflowqueue.scala 134:29 194:37]
  wire [38:0] _GEN_91852 = 4'h0 < realFlowNum_1 ? _GEN_87626 : flow_entry_1_21_vaddr; // @[Vlflowqueue.scala 134:29 194:37]
  wire [38:0] _GEN_91853 = 4'h0 < realFlowNum_1 ? _GEN_87627 : flow_entry_1_22_vaddr; // @[Vlflowqueue.scala 134:29 194:37]
  wire [38:0] _GEN_91854 = 4'h0 < realFlowNum_1 ? _GEN_87628 : flow_entry_1_23_vaddr; // @[Vlflowqueue.scala 134:29 194:37]
  wire [38:0] _GEN_91855 = 4'h0 < realFlowNum_1 ? _GEN_87629 : flow_entry_1_24_vaddr; // @[Vlflowqueue.scala 134:29 194:37]
  wire [38:0] _GEN_91856 = 4'h0 < realFlowNum_1 ? _GEN_87630 : flow_entry_1_25_vaddr; // @[Vlflowqueue.scala 134:29 194:37]
  wire [38:0] _GEN_91857 = 4'h0 < realFlowNum_1 ? _GEN_87631 : flow_entry_1_26_vaddr; // @[Vlflowqueue.scala 134:29 194:37]
  wire [38:0] _GEN_91858 = 4'h0 < realFlowNum_1 ? _GEN_87632 : flow_entry_1_27_vaddr; // @[Vlflowqueue.scala 134:29 194:37]
  wire [38:0] _GEN_91859 = 4'h0 < realFlowNum_1 ? _GEN_87633 : flow_entry_1_28_vaddr; // @[Vlflowqueue.scala 134:29 194:37]
  wire [38:0] _GEN_91860 = 4'h0 < realFlowNum_1 ? _GEN_87634 : flow_entry_1_29_vaddr; // @[Vlflowqueue.scala 134:29 194:37]
  wire [38:0] _GEN_91861 = 4'h0 < realFlowNum_1 ? _GEN_87635 : flow_entry_1_30_vaddr; // @[Vlflowqueue.scala 134:29 194:37]
  wire [38:0] _GEN_91862 = 4'h0 < realFlowNum_1 ? _GEN_87636 : flow_entry_1_31_vaddr; // @[Vlflowqueue.scala 134:29 194:37]
  wire  _GEN_92119 = _GEN_162068 | _GEN_88278; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_92120 = _GEN_162069 | _GEN_88279; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_92121 = _GEN_162070 | _GEN_88280; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_92122 = _GEN_162071 | _GEN_88281; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_92123 = _GEN_162072 | _GEN_88282; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_92124 = _GEN_162073 | _GEN_88283; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_92125 = _GEN_162074 | _GEN_88284; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_92126 = _GEN_162075 | _GEN_88285; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_92127 = _GEN_162076 | _GEN_88286; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_92128 = _GEN_162077 | _GEN_88287; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_92129 = _GEN_162078 | _GEN_88288; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_92130 = _GEN_162079 | _GEN_88289; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_92131 = _GEN_162080 | _GEN_88290; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_92132 = _GEN_162081 | _GEN_88291; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_92133 = _GEN_162082 | _GEN_88292; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_92134 = _GEN_162083 | _GEN_88293; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_92135 = _GEN_162084 | _GEN_88294; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_92136 = _GEN_162085 | _GEN_88295; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_92137 = _GEN_162086 | _GEN_88296; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_92138 = _GEN_162087 | _GEN_88297; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_92139 = _GEN_162088 | _GEN_88298; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_92140 = _GEN_162089 | _GEN_88299; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_92141 = _GEN_162090 | _GEN_88300; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_92142 = _GEN_162091 | _GEN_88301; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_92143 = _GEN_162092 | _GEN_88302; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_92144 = _GEN_162093 | _GEN_88303; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_92145 = _GEN_162094 | _GEN_88304; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_92146 = _GEN_162095 | _GEN_88305; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_92147 = _GEN_162096 | _GEN_88306; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_92148 = _GEN_162097 | _GEN_88307; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_92149 = _GEN_162098 | _GEN_88308; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_92150 = _GEN_162099 | _GEN_88309; // @[Vlflowqueue.scala 197:{51,51}]
  wire [4:0] _GEN_95095 = 5'h0 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_91254; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_95096 = 5'h1 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_91255; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_95097 = 5'h2 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_91256; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_95098 = 5'h3 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_91257; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_95099 = 5'h4 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_91258; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_95100 = 5'h5 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_91259; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_95101 = 5'h6 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_91260; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_95102 = 5'h7 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_91261; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_95103 = 5'h8 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_91262; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_95104 = 5'h9 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_91263; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_95105 = 5'ha == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_91264; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_95106 = 5'hb == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_91265; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_95107 = 5'hc == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_91266; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_95108 = 5'hd == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_91267; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_95109 = 5'he == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_91268; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_95110 = 5'hf == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_91269; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_95111 = 5'h10 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_91270; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_95112 = 5'h11 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_91271; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_95113 = 5'h12 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_91272; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_95114 = 5'h13 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_91273; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_95115 = 5'h14 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_91274; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_95116 = 5'h15 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_91275; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_95117 = 5'h16 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_91276; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_95118 = 5'h17 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_91277; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_95119 = 5'h18 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_91278; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_95120 = 5'h19 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_91279; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_95121 = 5'h1a == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_91280; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_95122 = 5'h1b == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_91281; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_95123 = 5'h1c == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_91282; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_95124 = 5'h1d == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_91283; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_95125 = 5'h1e == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_91284; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_95126 = 5'h1f == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_91285; // @[Vlflowqueue.scala 198:{51,51}]
  wire [38:0] _GEN_95671 = 5'h0 == index_1 ? vaddr_1 : _GEN_91831; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_95672 = 5'h1 == index_1 ? vaddr_1 : _GEN_91832; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_95673 = 5'h2 == index_1 ? vaddr_1 : _GEN_91833; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_95674 = 5'h3 == index_1 ? vaddr_1 : _GEN_91834; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_95675 = 5'h4 == index_1 ? vaddr_1 : _GEN_91835; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_95676 = 5'h5 == index_1 ? vaddr_1 : _GEN_91836; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_95677 = 5'h6 == index_1 ? vaddr_1 : _GEN_91837; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_95678 = 5'h7 == index_1 ? vaddr_1 : _GEN_91838; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_95679 = 5'h8 == index_1 ? vaddr_1 : _GEN_91839; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_95680 = 5'h9 == index_1 ? vaddr_1 : _GEN_91840; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_95681 = 5'ha == index_1 ? vaddr_1 : _GEN_91841; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_95682 = 5'hb == index_1 ? vaddr_1 : _GEN_91842; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_95683 = 5'hc == index_1 ? vaddr_1 : _GEN_91843; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_95684 = 5'hd == index_1 ? vaddr_1 : _GEN_91844; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_95685 = 5'he == index_1 ? vaddr_1 : _GEN_91845; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_95686 = 5'hf == index_1 ? vaddr_1 : _GEN_91846; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_95687 = 5'h10 == index_1 ? vaddr_1 : _GEN_91847; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_95688 = 5'h11 == index_1 ? vaddr_1 : _GEN_91848; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_95689 = 5'h12 == index_1 ? vaddr_1 : _GEN_91849; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_95690 = 5'h13 == index_1 ? vaddr_1 : _GEN_91850; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_95691 = 5'h14 == index_1 ? vaddr_1 : _GEN_91851; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_95692 = 5'h15 == index_1 ? vaddr_1 : _GEN_91852; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_95693 = 5'h16 == index_1 ? vaddr_1 : _GEN_91853; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_95694 = 5'h17 == index_1 ? vaddr_1 : _GEN_91854; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_95695 = 5'h18 == index_1 ? vaddr_1 : _GEN_91855; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_95696 = 5'h19 == index_1 ? vaddr_1 : _GEN_91856; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_95697 = 5'h1a == index_1 ? vaddr_1 : _GEN_91857; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_95698 = 5'h1b == index_1 ? vaddr_1 : _GEN_91858; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_95699 = 5'h1c == index_1 ? vaddr_1 : _GEN_91859; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_95700 = 5'h1d == index_1 ? vaddr_1 : _GEN_91860; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_95701 = 5'h1e == index_1 ? vaddr_1 : _GEN_91861; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_95702 = 5'h1f == index_1 ? vaddr_1 : _GEN_91862; // @[Vlflowqueue.scala 203:{51,51}]
  wire  _GEN_96344 = 4'h1 < realFlowNum_1 ? _GEN_92119 : _GEN_88278; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_96345 = 4'h1 < realFlowNum_1 ? _GEN_92120 : _GEN_88279; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_96346 = 4'h1 < realFlowNum_1 ? _GEN_92121 : _GEN_88280; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_96347 = 4'h1 < realFlowNum_1 ? _GEN_92122 : _GEN_88281; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_96348 = 4'h1 < realFlowNum_1 ? _GEN_92123 : _GEN_88282; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_96349 = 4'h1 < realFlowNum_1 ? _GEN_92124 : _GEN_88283; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_96350 = 4'h1 < realFlowNum_1 ? _GEN_92125 : _GEN_88284; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_96351 = 4'h1 < realFlowNum_1 ? _GEN_92126 : _GEN_88285; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_96352 = 4'h1 < realFlowNum_1 ? _GEN_92127 : _GEN_88286; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_96353 = 4'h1 < realFlowNum_1 ? _GEN_92128 : _GEN_88287; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_96354 = 4'h1 < realFlowNum_1 ? _GEN_92129 : _GEN_88288; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_96355 = 4'h1 < realFlowNum_1 ? _GEN_92130 : _GEN_88289; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_96356 = 4'h1 < realFlowNum_1 ? _GEN_92131 : _GEN_88290; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_96357 = 4'h1 < realFlowNum_1 ? _GEN_92132 : _GEN_88291; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_96358 = 4'h1 < realFlowNum_1 ? _GEN_92133 : _GEN_88292; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_96359 = 4'h1 < realFlowNum_1 ? _GEN_92134 : _GEN_88293; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_96360 = 4'h1 < realFlowNum_1 ? _GEN_92135 : _GEN_88294; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_96361 = 4'h1 < realFlowNum_1 ? _GEN_92136 : _GEN_88295; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_96362 = 4'h1 < realFlowNum_1 ? _GEN_92137 : _GEN_88296; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_96363 = 4'h1 < realFlowNum_1 ? _GEN_92138 : _GEN_88297; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_96364 = 4'h1 < realFlowNum_1 ? _GEN_92139 : _GEN_88298; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_96365 = 4'h1 < realFlowNum_1 ? _GEN_92140 : _GEN_88299; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_96366 = 4'h1 < realFlowNum_1 ? _GEN_92141 : _GEN_88300; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_96367 = 4'h1 < realFlowNum_1 ? _GEN_92142 : _GEN_88301; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_96368 = 4'h1 < realFlowNum_1 ? _GEN_92143 : _GEN_88302; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_96369 = 4'h1 < realFlowNum_1 ? _GEN_92144 : _GEN_88303; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_96370 = 4'h1 < realFlowNum_1 ? _GEN_92145 : _GEN_88304; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_96371 = 4'h1 < realFlowNum_1 ? _GEN_92146 : _GEN_88305; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_96372 = 4'h1 < realFlowNum_1 ? _GEN_92147 : _GEN_88306; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_96373 = 4'h1 < realFlowNum_1 ? _GEN_92148 : _GEN_88307; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_96374 = 4'h1 < realFlowNum_1 ? _GEN_92149 : _GEN_88308; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_96375 = 4'h1 < realFlowNum_1 ? _GEN_92150 : _GEN_88309; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_99320 = 4'h1 < realFlowNum_1 ? _GEN_95095 : _GEN_91254; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_99321 = 4'h1 < realFlowNum_1 ? _GEN_95096 : _GEN_91255; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_99322 = 4'h1 < realFlowNum_1 ? _GEN_95097 : _GEN_91256; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_99323 = 4'h1 < realFlowNum_1 ? _GEN_95098 : _GEN_91257; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_99324 = 4'h1 < realFlowNum_1 ? _GEN_95099 : _GEN_91258; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_99325 = 4'h1 < realFlowNum_1 ? _GEN_95100 : _GEN_91259; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_99326 = 4'h1 < realFlowNum_1 ? _GEN_95101 : _GEN_91260; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_99327 = 4'h1 < realFlowNum_1 ? _GEN_95102 : _GEN_91261; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_99328 = 4'h1 < realFlowNum_1 ? _GEN_95103 : _GEN_91262; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_99329 = 4'h1 < realFlowNum_1 ? _GEN_95104 : _GEN_91263; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_99330 = 4'h1 < realFlowNum_1 ? _GEN_95105 : _GEN_91264; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_99331 = 4'h1 < realFlowNum_1 ? _GEN_95106 : _GEN_91265; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_99332 = 4'h1 < realFlowNum_1 ? _GEN_95107 : _GEN_91266; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_99333 = 4'h1 < realFlowNum_1 ? _GEN_95108 : _GEN_91267; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_99334 = 4'h1 < realFlowNum_1 ? _GEN_95109 : _GEN_91268; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_99335 = 4'h1 < realFlowNum_1 ? _GEN_95110 : _GEN_91269; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_99336 = 4'h1 < realFlowNum_1 ? _GEN_95111 : _GEN_91270; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_99337 = 4'h1 < realFlowNum_1 ? _GEN_95112 : _GEN_91271; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_99338 = 4'h1 < realFlowNum_1 ? _GEN_95113 : _GEN_91272; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_99339 = 4'h1 < realFlowNum_1 ? _GEN_95114 : _GEN_91273; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_99340 = 4'h1 < realFlowNum_1 ? _GEN_95115 : _GEN_91274; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_99341 = 4'h1 < realFlowNum_1 ? _GEN_95116 : _GEN_91275; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_99342 = 4'h1 < realFlowNum_1 ? _GEN_95117 : _GEN_91276; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_99343 = 4'h1 < realFlowNum_1 ? _GEN_95118 : _GEN_91277; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_99344 = 4'h1 < realFlowNum_1 ? _GEN_95119 : _GEN_91278; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_99345 = 4'h1 < realFlowNum_1 ? _GEN_95120 : _GEN_91279; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_99346 = 4'h1 < realFlowNum_1 ? _GEN_95121 : _GEN_91280; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_99347 = 4'h1 < realFlowNum_1 ? _GEN_95122 : _GEN_91281; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_99348 = 4'h1 < realFlowNum_1 ? _GEN_95123 : _GEN_91282; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_99349 = 4'h1 < realFlowNum_1 ? _GEN_95124 : _GEN_91283; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_99350 = 4'h1 < realFlowNum_1 ? _GEN_95125 : _GEN_91284; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_99351 = 4'h1 < realFlowNum_1 ? _GEN_95126 : _GEN_91285; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_99897 = 4'h1 < realFlowNum_1 ? _GEN_95671 : _GEN_91831; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_99898 = 4'h1 < realFlowNum_1 ? _GEN_95672 : _GEN_91832; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_99899 = 4'h1 < realFlowNum_1 ? _GEN_95673 : _GEN_91833; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_99900 = 4'h1 < realFlowNum_1 ? _GEN_95674 : _GEN_91834; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_99901 = 4'h1 < realFlowNum_1 ? _GEN_95675 : _GEN_91835; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_99902 = 4'h1 < realFlowNum_1 ? _GEN_95676 : _GEN_91836; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_99903 = 4'h1 < realFlowNum_1 ? _GEN_95677 : _GEN_91837; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_99904 = 4'h1 < realFlowNum_1 ? _GEN_95678 : _GEN_91838; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_99905 = 4'h1 < realFlowNum_1 ? _GEN_95679 : _GEN_91839; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_99906 = 4'h1 < realFlowNum_1 ? _GEN_95680 : _GEN_91840; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_99907 = 4'h1 < realFlowNum_1 ? _GEN_95681 : _GEN_91841; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_99908 = 4'h1 < realFlowNum_1 ? _GEN_95682 : _GEN_91842; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_99909 = 4'h1 < realFlowNum_1 ? _GEN_95683 : _GEN_91843; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_99910 = 4'h1 < realFlowNum_1 ? _GEN_95684 : _GEN_91844; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_99911 = 4'h1 < realFlowNum_1 ? _GEN_95685 : _GEN_91845; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_99912 = 4'h1 < realFlowNum_1 ? _GEN_95686 : _GEN_91846; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_99913 = 4'h1 < realFlowNum_1 ? _GEN_95687 : _GEN_91847; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_99914 = 4'h1 < realFlowNum_1 ? _GEN_95688 : _GEN_91848; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_99915 = 4'h1 < realFlowNum_1 ? _GEN_95689 : _GEN_91849; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_99916 = 4'h1 < realFlowNum_1 ? _GEN_95690 : _GEN_91850; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_99917 = 4'h1 < realFlowNum_1 ? _GEN_95691 : _GEN_91851; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_99918 = 4'h1 < realFlowNum_1 ? _GEN_95692 : _GEN_91852; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_99919 = 4'h1 < realFlowNum_1 ? _GEN_95693 : _GEN_91853; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_99920 = 4'h1 < realFlowNum_1 ? _GEN_95694 : _GEN_91854; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_99921 = 4'h1 < realFlowNum_1 ? _GEN_95695 : _GEN_91855; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_99922 = 4'h1 < realFlowNum_1 ? _GEN_95696 : _GEN_91856; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_99923 = 4'h1 < realFlowNum_1 ? _GEN_95697 : _GEN_91857; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_99924 = 4'h1 < realFlowNum_1 ? _GEN_95698 : _GEN_91858; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_99925 = 4'h1 < realFlowNum_1 ? _GEN_95699 : _GEN_91859; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_99926 = 4'h1 < realFlowNum_1 ? _GEN_95700 : _GEN_91860; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_99927 = 4'h1 < realFlowNum_1 ? _GEN_95701 : _GEN_91861; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_99928 = 4'h1 < realFlowNum_1 ? _GEN_95702 : _GEN_91862; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_100185 = _GEN_162068 | _GEN_96344; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_100186 = _GEN_162069 | _GEN_96345; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_100187 = _GEN_162070 | _GEN_96346; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_100188 = _GEN_162071 | _GEN_96347; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_100189 = _GEN_162072 | _GEN_96348; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_100190 = _GEN_162073 | _GEN_96349; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_100191 = _GEN_162074 | _GEN_96350; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_100192 = _GEN_162075 | _GEN_96351; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_100193 = _GEN_162076 | _GEN_96352; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_100194 = _GEN_162077 | _GEN_96353; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_100195 = _GEN_162078 | _GEN_96354; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_100196 = _GEN_162079 | _GEN_96355; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_100197 = _GEN_162080 | _GEN_96356; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_100198 = _GEN_162081 | _GEN_96357; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_100199 = _GEN_162082 | _GEN_96358; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_100200 = _GEN_162083 | _GEN_96359; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_100201 = _GEN_162084 | _GEN_96360; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_100202 = _GEN_162085 | _GEN_96361; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_100203 = _GEN_162086 | _GEN_96362; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_100204 = _GEN_162087 | _GEN_96363; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_100205 = _GEN_162088 | _GEN_96364; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_100206 = _GEN_162089 | _GEN_96365; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_100207 = _GEN_162090 | _GEN_96366; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_100208 = _GEN_162091 | _GEN_96367; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_100209 = _GEN_162092 | _GEN_96368; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_100210 = _GEN_162093 | _GEN_96369; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_100211 = _GEN_162094 | _GEN_96370; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_100212 = _GEN_162095 | _GEN_96371; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_100213 = _GEN_162096 | _GEN_96372; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_100214 = _GEN_162097 | _GEN_96373; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_100215 = _GEN_162098 | _GEN_96374; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_100216 = _GEN_162099 | _GEN_96375; // @[Vlflowqueue.scala 197:{51,51}]
  wire [4:0] _GEN_103161 = 5'h0 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_99320; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_103162 = 5'h1 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_99321; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_103163 = 5'h2 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_99322; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_103164 = 5'h3 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_99323; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_103165 = 5'h4 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_99324; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_103166 = 5'h5 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_99325; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_103167 = 5'h6 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_99326; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_103168 = 5'h7 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_99327; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_103169 = 5'h8 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_99328; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_103170 = 5'h9 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_99329; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_103171 = 5'ha == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_99330; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_103172 = 5'hb == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_99331; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_103173 = 5'hc == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_99332; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_103174 = 5'hd == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_99333; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_103175 = 5'he == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_99334; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_103176 = 5'hf == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_99335; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_103177 = 5'h10 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_99336; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_103178 = 5'h11 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_99337; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_103179 = 5'h12 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_99338; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_103180 = 5'h13 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_99339; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_103181 = 5'h14 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_99340; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_103182 = 5'h15 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_99341; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_103183 = 5'h16 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_99342; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_103184 = 5'h17 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_99343; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_103185 = 5'h18 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_99344; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_103186 = 5'h19 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_99345; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_103187 = 5'h1a == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_99346; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_103188 = 5'h1b == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_99347; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_103189 = 5'h1c == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_99348; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_103190 = 5'h1d == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_99349; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_103191 = 5'h1e == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_99350; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_103192 = 5'h1f == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_99351; // @[Vlflowqueue.scala 198:{51,51}]
  wire [38:0] _GEN_103737 = 5'h0 == index_1 ? vaddr_1 : _GEN_99897; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_103738 = 5'h1 == index_1 ? vaddr_1 : _GEN_99898; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_103739 = 5'h2 == index_1 ? vaddr_1 : _GEN_99899; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_103740 = 5'h3 == index_1 ? vaddr_1 : _GEN_99900; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_103741 = 5'h4 == index_1 ? vaddr_1 : _GEN_99901; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_103742 = 5'h5 == index_1 ? vaddr_1 : _GEN_99902; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_103743 = 5'h6 == index_1 ? vaddr_1 : _GEN_99903; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_103744 = 5'h7 == index_1 ? vaddr_1 : _GEN_99904; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_103745 = 5'h8 == index_1 ? vaddr_1 : _GEN_99905; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_103746 = 5'h9 == index_1 ? vaddr_1 : _GEN_99906; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_103747 = 5'ha == index_1 ? vaddr_1 : _GEN_99907; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_103748 = 5'hb == index_1 ? vaddr_1 : _GEN_99908; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_103749 = 5'hc == index_1 ? vaddr_1 : _GEN_99909; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_103750 = 5'hd == index_1 ? vaddr_1 : _GEN_99910; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_103751 = 5'he == index_1 ? vaddr_1 : _GEN_99911; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_103752 = 5'hf == index_1 ? vaddr_1 : _GEN_99912; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_103753 = 5'h10 == index_1 ? vaddr_1 : _GEN_99913; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_103754 = 5'h11 == index_1 ? vaddr_1 : _GEN_99914; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_103755 = 5'h12 == index_1 ? vaddr_1 : _GEN_99915; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_103756 = 5'h13 == index_1 ? vaddr_1 : _GEN_99916; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_103757 = 5'h14 == index_1 ? vaddr_1 : _GEN_99917; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_103758 = 5'h15 == index_1 ? vaddr_1 : _GEN_99918; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_103759 = 5'h16 == index_1 ? vaddr_1 : _GEN_99919; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_103760 = 5'h17 == index_1 ? vaddr_1 : _GEN_99920; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_103761 = 5'h18 == index_1 ? vaddr_1 : _GEN_99921; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_103762 = 5'h19 == index_1 ? vaddr_1 : _GEN_99922; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_103763 = 5'h1a == index_1 ? vaddr_1 : _GEN_99923; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_103764 = 5'h1b == index_1 ? vaddr_1 : _GEN_99924; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_103765 = 5'h1c == index_1 ? vaddr_1 : _GEN_99925; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_103766 = 5'h1d == index_1 ? vaddr_1 : _GEN_99926; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_103767 = 5'h1e == index_1 ? vaddr_1 : _GEN_99927; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_103768 = 5'h1f == index_1 ? vaddr_1 : _GEN_99928; // @[Vlflowqueue.scala 203:{51,51}]
  wire  _GEN_104410 = 4'h2 < realFlowNum_1 ? _GEN_100185 : _GEN_96344; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_104411 = 4'h2 < realFlowNum_1 ? _GEN_100186 : _GEN_96345; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_104412 = 4'h2 < realFlowNum_1 ? _GEN_100187 : _GEN_96346; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_104413 = 4'h2 < realFlowNum_1 ? _GEN_100188 : _GEN_96347; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_104414 = 4'h2 < realFlowNum_1 ? _GEN_100189 : _GEN_96348; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_104415 = 4'h2 < realFlowNum_1 ? _GEN_100190 : _GEN_96349; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_104416 = 4'h2 < realFlowNum_1 ? _GEN_100191 : _GEN_96350; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_104417 = 4'h2 < realFlowNum_1 ? _GEN_100192 : _GEN_96351; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_104418 = 4'h2 < realFlowNum_1 ? _GEN_100193 : _GEN_96352; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_104419 = 4'h2 < realFlowNum_1 ? _GEN_100194 : _GEN_96353; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_104420 = 4'h2 < realFlowNum_1 ? _GEN_100195 : _GEN_96354; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_104421 = 4'h2 < realFlowNum_1 ? _GEN_100196 : _GEN_96355; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_104422 = 4'h2 < realFlowNum_1 ? _GEN_100197 : _GEN_96356; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_104423 = 4'h2 < realFlowNum_1 ? _GEN_100198 : _GEN_96357; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_104424 = 4'h2 < realFlowNum_1 ? _GEN_100199 : _GEN_96358; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_104425 = 4'h2 < realFlowNum_1 ? _GEN_100200 : _GEN_96359; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_104426 = 4'h2 < realFlowNum_1 ? _GEN_100201 : _GEN_96360; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_104427 = 4'h2 < realFlowNum_1 ? _GEN_100202 : _GEN_96361; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_104428 = 4'h2 < realFlowNum_1 ? _GEN_100203 : _GEN_96362; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_104429 = 4'h2 < realFlowNum_1 ? _GEN_100204 : _GEN_96363; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_104430 = 4'h2 < realFlowNum_1 ? _GEN_100205 : _GEN_96364; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_104431 = 4'h2 < realFlowNum_1 ? _GEN_100206 : _GEN_96365; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_104432 = 4'h2 < realFlowNum_1 ? _GEN_100207 : _GEN_96366; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_104433 = 4'h2 < realFlowNum_1 ? _GEN_100208 : _GEN_96367; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_104434 = 4'h2 < realFlowNum_1 ? _GEN_100209 : _GEN_96368; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_104435 = 4'h2 < realFlowNum_1 ? _GEN_100210 : _GEN_96369; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_104436 = 4'h2 < realFlowNum_1 ? _GEN_100211 : _GEN_96370; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_104437 = 4'h2 < realFlowNum_1 ? _GEN_100212 : _GEN_96371; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_104438 = 4'h2 < realFlowNum_1 ? _GEN_100213 : _GEN_96372; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_104439 = 4'h2 < realFlowNum_1 ? _GEN_100214 : _GEN_96373; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_104440 = 4'h2 < realFlowNum_1 ? _GEN_100215 : _GEN_96374; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_104441 = 4'h2 < realFlowNum_1 ? _GEN_100216 : _GEN_96375; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_107386 = 4'h2 < realFlowNum_1 ? _GEN_103161 : _GEN_99320; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_107387 = 4'h2 < realFlowNum_1 ? _GEN_103162 : _GEN_99321; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_107388 = 4'h2 < realFlowNum_1 ? _GEN_103163 : _GEN_99322; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_107389 = 4'h2 < realFlowNum_1 ? _GEN_103164 : _GEN_99323; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_107390 = 4'h2 < realFlowNum_1 ? _GEN_103165 : _GEN_99324; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_107391 = 4'h2 < realFlowNum_1 ? _GEN_103166 : _GEN_99325; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_107392 = 4'h2 < realFlowNum_1 ? _GEN_103167 : _GEN_99326; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_107393 = 4'h2 < realFlowNum_1 ? _GEN_103168 : _GEN_99327; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_107394 = 4'h2 < realFlowNum_1 ? _GEN_103169 : _GEN_99328; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_107395 = 4'h2 < realFlowNum_1 ? _GEN_103170 : _GEN_99329; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_107396 = 4'h2 < realFlowNum_1 ? _GEN_103171 : _GEN_99330; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_107397 = 4'h2 < realFlowNum_1 ? _GEN_103172 : _GEN_99331; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_107398 = 4'h2 < realFlowNum_1 ? _GEN_103173 : _GEN_99332; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_107399 = 4'h2 < realFlowNum_1 ? _GEN_103174 : _GEN_99333; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_107400 = 4'h2 < realFlowNum_1 ? _GEN_103175 : _GEN_99334; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_107401 = 4'h2 < realFlowNum_1 ? _GEN_103176 : _GEN_99335; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_107402 = 4'h2 < realFlowNum_1 ? _GEN_103177 : _GEN_99336; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_107403 = 4'h2 < realFlowNum_1 ? _GEN_103178 : _GEN_99337; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_107404 = 4'h2 < realFlowNum_1 ? _GEN_103179 : _GEN_99338; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_107405 = 4'h2 < realFlowNum_1 ? _GEN_103180 : _GEN_99339; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_107406 = 4'h2 < realFlowNum_1 ? _GEN_103181 : _GEN_99340; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_107407 = 4'h2 < realFlowNum_1 ? _GEN_103182 : _GEN_99341; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_107408 = 4'h2 < realFlowNum_1 ? _GEN_103183 : _GEN_99342; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_107409 = 4'h2 < realFlowNum_1 ? _GEN_103184 : _GEN_99343; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_107410 = 4'h2 < realFlowNum_1 ? _GEN_103185 : _GEN_99344; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_107411 = 4'h2 < realFlowNum_1 ? _GEN_103186 : _GEN_99345; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_107412 = 4'h2 < realFlowNum_1 ? _GEN_103187 : _GEN_99346; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_107413 = 4'h2 < realFlowNum_1 ? _GEN_103188 : _GEN_99347; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_107414 = 4'h2 < realFlowNum_1 ? _GEN_103189 : _GEN_99348; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_107415 = 4'h2 < realFlowNum_1 ? _GEN_103190 : _GEN_99349; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_107416 = 4'h2 < realFlowNum_1 ? _GEN_103191 : _GEN_99350; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_107417 = 4'h2 < realFlowNum_1 ? _GEN_103192 : _GEN_99351; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_107963 = 4'h2 < realFlowNum_1 ? _GEN_103737 : _GEN_99897; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_107964 = 4'h2 < realFlowNum_1 ? _GEN_103738 : _GEN_99898; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_107965 = 4'h2 < realFlowNum_1 ? _GEN_103739 : _GEN_99899; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_107966 = 4'h2 < realFlowNum_1 ? _GEN_103740 : _GEN_99900; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_107967 = 4'h2 < realFlowNum_1 ? _GEN_103741 : _GEN_99901; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_107968 = 4'h2 < realFlowNum_1 ? _GEN_103742 : _GEN_99902; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_107969 = 4'h2 < realFlowNum_1 ? _GEN_103743 : _GEN_99903; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_107970 = 4'h2 < realFlowNum_1 ? _GEN_103744 : _GEN_99904; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_107971 = 4'h2 < realFlowNum_1 ? _GEN_103745 : _GEN_99905; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_107972 = 4'h2 < realFlowNum_1 ? _GEN_103746 : _GEN_99906; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_107973 = 4'h2 < realFlowNum_1 ? _GEN_103747 : _GEN_99907; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_107974 = 4'h2 < realFlowNum_1 ? _GEN_103748 : _GEN_99908; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_107975 = 4'h2 < realFlowNum_1 ? _GEN_103749 : _GEN_99909; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_107976 = 4'h2 < realFlowNum_1 ? _GEN_103750 : _GEN_99910; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_107977 = 4'h2 < realFlowNum_1 ? _GEN_103751 : _GEN_99911; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_107978 = 4'h2 < realFlowNum_1 ? _GEN_103752 : _GEN_99912; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_107979 = 4'h2 < realFlowNum_1 ? _GEN_103753 : _GEN_99913; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_107980 = 4'h2 < realFlowNum_1 ? _GEN_103754 : _GEN_99914; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_107981 = 4'h2 < realFlowNum_1 ? _GEN_103755 : _GEN_99915; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_107982 = 4'h2 < realFlowNum_1 ? _GEN_103756 : _GEN_99916; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_107983 = 4'h2 < realFlowNum_1 ? _GEN_103757 : _GEN_99917; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_107984 = 4'h2 < realFlowNum_1 ? _GEN_103758 : _GEN_99918; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_107985 = 4'h2 < realFlowNum_1 ? _GEN_103759 : _GEN_99919; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_107986 = 4'h2 < realFlowNum_1 ? _GEN_103760 : _GEN_99920; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_107987 = 4'h2 < realFlowNum_1 ? _GEN_103761 : _GEN_99921; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_107988 = 4'h2 < realFlowNum_1 ? _GEN_103762 : _GEN_99922; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_107989 = 4'h2 < realFlowNum_1 ? _GEN_103763 : _GEN_99923; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_107990 = 4'h2 < realFlowNum_1 ? _GEN_103764 : _GEN_99924; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_107991 = 4'h2 < realFlowNum_1 ? _GEN_103765 : _GEN_99925; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_107992 = 4'h2 < realFlowNum_1 ? _GEN_103766 : _GEN_99926; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_107993 = 4'h2 < realFlowNum_1 ? _GEN_103767 : _GEN_99927; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_107994 = 4'h2 < realFlowNum_1 ? _GEN_103768 : _GEN_99928; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_108251 = _GEN_162068 | _GEN_104410; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_108252 = _GEN_162069 | _GEN_104411; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_108253 = _GEN_162070 | _GEN_104412; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_108254 = _GEN_162071 | _GEN_104413; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_108255 = _GEN_162072 | _GEN_104414; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_108256 = _GEN_162073 | _GEN_104415; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_108257 = _GEN_162074 | _GEN_104416; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_108258 = _GEN_162075 | _GEN_104417; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_108259 = _GEN_162076 | _GEN_104418; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_108260 = _GEN_162077 | _GEN_104419; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_108261 = _GEN_162078 | _GEN_104420; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_108262 = _GEN_162079 | _GEN_104421; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_108263 = _GEN_162080 | _GEN_104422; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_108264 = _GEN_162081 | _GEN_104423; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_108265 = _GEN_162082 | _GEN_104424; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_108266 = _GEN_162083 | _GEN_104425; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_108267 = _GEN_162084 | _GEN_104426; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_108268 = _GEN_162085 | _GEN_104427; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_108269 = _GEN_162086 | _GEN_104428; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_108270 = _GEN_162087 | _GEN_104429; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_108271 = _GEN_162088 | _GEN_104430; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_108272 = _GEN_162089 | _GEN_104431; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_108273 = _GEN_162090 | _GEN_104432; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_108274 = _GEN_162091 | _GEN_104433; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_108275 = _GEN_162092 | _GEN_104434; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_108276 = _GEN_162093 | _GEN_104435; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_108277 = _GEN_162094 | _GEN_104436; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_108278 = _GEN_162095 | _GEN_104437; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_108279 = _GEN_162096 | _GEN_104438; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_108280 = _GEN_162097 | _GEN_104439; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_108281 = _GEN_162098 | _GEN_104440; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_108282 = _GEN_162099 | _GEN_104441; // @[Vlflowqueue.scala 197:{51,51}]
  wire [4:0] _GEN_111227 = 5'h0 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_107386; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_111228 = 5'h1 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_107387; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_111229 = 5'h2 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_107388; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_111230 = 5'h3 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_107389; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_111231 = 5'h4 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_107390; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_111232 = 5'h5 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_107391; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_111233 = 5'h6 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_107392; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_111234 = 5'h7 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_107393; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_111235 = 5'h8 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_107394; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_111236 = 5'h9 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_107395; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_111237 = 5'ha == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_107396; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_111238 = 5'hb == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_107397; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_111239 = 5'hc == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_107398; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_111240 = 5'hd == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_107399; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_111241 = 5'he == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_107400; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_111242 = 5'hf == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_107401; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_111243 = 5'h10 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_107402; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_111244 = 5'h11 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_107403; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_111245 = 5'h12 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_107404; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_111246 = 5'h13 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_107405; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_111247 = 5'h14 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_107406; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_111248 = 5'h15 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_107407; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_111249 = 5'h16 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_107408; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_111250 = 5'h17 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_107409; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_111251 = 5'h18 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_107410; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_111252 = 5'h19 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_107411; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_111253 = 5'h1a == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_107412; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_111254 = 5'h1b == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_107413; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_111255 = 5'h1c == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_107414; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_111256 = 5'h1d == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_107415; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_111257 = 5'h1e == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_107416; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_111258 = 5'h1f == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_107417; // @[Vlflowqueue.scala 198:{51,51}]
  wire [38:0] _GEN_111803 = 5'h0 == index_1 ? vaddr_1 : _GEN_107963; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_111804 = 5'h1 == index_1 ? vaddr_1 : _GEN_107964; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_111805 = 5'h2 == index_1 ? vaddr_1 : _GEN_107965; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_111806 = 5'h3 == index_1 ? vaddr_1 : _GEN_107966; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_111807 = 5'h4 == index_1 ? vaddr_1 : _GEN_107967; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_111808 = 5'h5 == index_1 ? vaddr_1 : _GEN_107968; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_111809 = 5'h6 == index_1 ? vaddr_1 : _GEN_107969; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_111810 = 5'h7 == index_1 ? vaddr_1 : _GEN_107970; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_111811 = 5'h8 == index_1 ? vaddr_1 : _GEN_107971; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_111812 = 5'h9 == index_1 ? vaddr_1 : _GEN_107972; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_111813 = 5'ha == index_1 ? vaddr_1 : _GEN_107973; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_111814 = 5'hb == index_1 ? vaddr_1 : _GEN_107974; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_111815 = 5'hc == index_1 ? vaddr_1 : _GEN_107975; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_111816 = 5'hd == index_1 ? vaddr_1 : _GEN_107976; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_111817 = 5'he == index_1 ? vaddr_1 : _GEN_107977; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_111818 = 5'hf == index_1 ? vaddr_1 : _GEN_107978; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_111819 = 5'h10 == index_1 ? vaddr_1 : _GEN_107979; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_111820 = 5'h11 == index_1 ? vaddr_1 : _GEN_107980; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_111821 = 5'h12 == index_1 ? vaddr_1 : _GEN_107981; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_111822 = 5'h13 == index_1 ? vaddr_1 : _GEN_107982; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_111823 = 5'h14 == index_1 ? vaddr_1 : _GEN_107983; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_111824 = 5'h15 == index_1 ? vaddr_1 : _GEN_107984; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_111825 = 5'h16 == index_1 ? vaddr_1 : _GEN_107985; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_111826 = 5'h17 == index_1 ? vaddr_1 : _GEN_107986; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_111827 = 5'h18 == index_1 ? vaddr_1 : _GEN_107987; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_111828 = 5'h19 == index_1 ? vaddr_1 : _GEN_107988; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_111829 = 5'h1a == index_1 ? vaddr_1 : _GEN_107989; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_111830 = 5'h1b == index_1 ? vaddr_1 : _GEN_107990; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_111831 = 5'h1c == index_1 ? vaddr_1 : _GEN_107991; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_111832 = 5'h1d == index_1 ? vaddr_1 : _GEN_107992; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_111833 = 5'h1e == index_1 ? vaddr_1 : _GEN_107993; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_111834 = 5'h1f == index_1 ? vaddr_1 : _GEN_107994; // @[Vlflowqueue.scala 203:{51,51}]
  wire  _GEN_112476 = 4'h3 < realFlowNum_1 ? _GEN_108251 : _GEN_104410; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_112477 = 4'h3 < realFlowNum_1 ? _GEN_108252 : _GEN_104411; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_112478 = 4'h3 < realFlowNum_1 ? _GEN_108253 : _GEN_104412; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_112479 = 4'h3 < realFlowNum_1 ? _GEN_108254 : _GEN_104413; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_112480 = 4'h3 < realFlowNum_1 ? _GEN_108255 : _GEN_104414; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_112481 = 4'h3 < realFlowNum_1 ? _GEN_108256 : _GEN_104415; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_112482 = 4'h3 < realFlowNum_1 ? _GEN_108257 : _GEN_104416; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_112483 = 4'h3 < realFlowNum_1 ? _GEN_108258 : _GEN_104417; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_112484 = 4'h3 < realFlowNum_1 ? _GEN_108259 : _GEN_104418; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_112485 = 4'h3 < realFlowNum_1 ? _GEN_108260 : _GEN_104419; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_112486 = 4'h3 < realFlowNum_1 ? _GEN_108261 : _GEN_104420; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_112487 = 4'h3 < realFlowNum_1 ? _GEN_108262 : _GEN_104421; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_112488 = 4'h3 < realFlowNum_1 ? _GEN_108263 : _GEN_104422; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_112489 = 4'h3 < realFlowNum_1 ? _GEN_108264 : _GEN_104423; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_112490 = 4'h3 < realFlowNum_1 ? _GEN_108265 : _GEN_104424; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_112491 = 4'h3 < realFlowNum_1 ? _GEN_108266 : _GEN_104425; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_112492 = 4'h3 < realFlowNum_1 ? _GEN_108267 : _GEN_104426; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_112493 = 4'h3 < realFlowNum_1 ? _GEN_108268 : _GEN_104427; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_112494 = 4'h3 < realFlowNum_1 ? _GEN_108269 : _GEN_104428; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_112495 = 4'h3 < realFlowNum_1 ? _GEN_108270 : _GEN_104429; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_112496 = 4'h3 < realFlowNum_1 ? _GEN_108271 : _GEN_104430; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_112497 = 4'h3 < realFlowNum_1 ? _GEN_108272 : _GEN_104431; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_112498 = 4'h3 < realFlowNum_1 ? _GEN_108273 : _GEN_104432; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_112499 = 4'h3 < realFlowNum_1 ? _GEN_108274 : _GEN_104433; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_112500 = 4'h3 < realFlowNum_1 ? _GEN_108275 : _GEN_104434; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_112501 = 4'h3 < realFlowNum_1 ? _GEN_108276 : _GEN_104435; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_112502 = 4'h3 < realFlowNum_1 ? _GEN_108277 : _GEN_104436; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_112503 = 4'h3 < realFlowNum_1 ? _GEN_108278 : _GEN_104437; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_112504 = 4'h3 < realFlowNum_1 ? _GEN_108279 : _GEN_104438; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_112505 = 4'h3 < realFlowNum_1 ? _GEN_108280 : _GEN_104439; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_112506 = 4'h3 < realFlowNum_1 ? _GEN_108281 : _GEN_104440; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_112507 = 4'h3 < realFlowNum_1 ? _GEN_108282 : _GEN_104441; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_115452 = 4'h3 < realFlowNum_1 ? _GEN_111227 : _GEN_107386; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_115453 = 4'h3 < realFlowNum_1 ? _GEN_111228 : _GEN_107387; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_115454 = 4'h3 < realFlowNum_1 ? _GEN_111229 : _GEN_107388; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_115455 = 4'h3 < realFlowNum_1 ? _GEN_111230 : _GEN_107389; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_115456 = 4'h3 < realFlowNum_1 ? _GEN_111231 : _GEN_107390; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_115457 = 4'h3 < realFlowNum_1 ? _GEN_111232 : _GEN_107391; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_115458 = 4'h3 < realFlowNum_1 ? _GEN_111233 : _GEN_107392; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_115459 = 4'h3 < realFlowNum_1 ? _GEN_111234 : _GEN_107393; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_115460 = 4'h3 < realFlowNum_1 ? _GEN_111235 : _GEN_107394; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_115461 = 4'h3 < realFlowNum_1 ? _GEN_111236 : _GEN_107395; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_115462 = 4'h3 < realFlowNum_1 ? _GEN_111237 : _GEN_107396; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_115463 = 4'h3 < realFlowNum_1 ? _GEN_111238 : _GEN_107397; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_115464 = 4'h3 < realFlowNum_1 ? _GEN_111239 : _GEN_107398; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_115465 = 4'h3 < realFlowNum_1 ? _GEN_111240 : _GEN_107399; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_115466 = 4'h3 < realFlowNum_1 ? _GEN_111241 : _GEN_107400; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_115467 = 4'h3 < realFlowNum_1 ? _GEN_111242 : _GEN_107401; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_115468 = 4'h3 < realFlowNum_1 ? _GEN_111243 : _GEN_107402; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_115469 = 4'h3 < realFlowNum_1 ? _GEN_111244 : _GEN_107403; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_115470 = 4'h3 < realFlowNum_1 ? _GEN_111245 : _GEN_107404; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_115471 = 4'h3 < realFlowNum_1 ? _GEN_111246 : _GEN_107405; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_115472 = 4'h3 < realFlowNum_1 ? _GEN_111247 : _GEN_107406; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_115473 = 4'h3 < realFlowNum_1 ? _GEN_111248 : _GEN_107407; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_115474 = 4'h3 < realFlowNum_1 ? _GEN_111249 : _GEN_107408; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_115475 = 4'h3 < realFlowNum_1 ? _GEN_111250 : _GEN_107409; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_115476 = 4'h3 < realFlowNum_1 ? _GEN_111251 : _GEN_107410; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_115477 = 4'h3 < realFlowNum_1 ? _GEN_111252 : _GEN_107411; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_115478 = 4'h3 < realFlowNum_1 ? _GEN_111253 : _GEN_107412; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_115479 = 4'h3 < realFlowNum_1 ? _GEN_111254 : _GEN_107413; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_115480 = 4'h3 < realFlowNum_1 ? _GEN_111255 : _GEN_107414; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_115481 = 4'h3 < realFlowNum_1 ? _GEN_111256 : _GEN_107415; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_115482 = 4'h3 < realFlowNum_1 ? _GEN_111257 : _GEN_107416; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_115483 = 4'h3 < realFlowNum_1 ? _GEN_111258 : _GEN_107417; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_116029 = 4'h3 < realFlowNum_1 ? _GEN_111803 : _GEN_107963; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_116030 = 4'h3 < realFlowNum_1 ? _GEN_111804 : _GEN_107964; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_116031 = 4'h3 < realFlowNum_1 ? _GEN_111805 : _GEN_107965; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_116032 = 4'h3 < realFlowNum_1 ? _GEN_111806 : _GEN_107966; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_116033 = 4'h3 < realFlowNum_1 ? _GEN_111807 : _GEN_107967; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_116034 = 4'h3 < realFlowNum_1 ? _GEN_111808 : _GEN_107968; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_116035 = 4'h3 < realFlowNum_1 ? _GEN_111809 : _GEN_107969; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_116036 = 4'h3 < realFlowNum_1 ? _GEN_111810 : _GEN_107970; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_116037 = 4'h3 < realFlowNum_1 ? _GEN_111811 : _GEN_107971; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_116038 = 4'h3 < realFlowNum_1 ? _GEN_111812 : _GEN_107972; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_116039 = 4'h3 < realFlowNum_1 ? _GEN_111813 : _GEN_107973; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_116040 = 4'h3 < realFlowNum_1 ? _GEN_111814 : _GEN_107974; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_116041 = 4'h3 < realFlowNum_1 ? _GEN_111815 : _GEN_107975; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_116042 = 4'h3 < realFlowNum_1 ? _GEN_111816 : _GEN_107976; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_116043 = 4'h3 < realFlowNum_1 ? _GEN_111817 : _GEN_107977; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_116044 = 4'h3 < realFlowNum_1 ? _GEN_111818 : _GEN_107978; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_116045 = 4'h3 < realFlowNum_1 ? _GEN_111819 : _GEN_107979; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_116046 = 4'h3 < realFlowNum_1 ? _GEN_111820 : _GEN_107980; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_116047 = 4'h3 < realFlowNum_1 ? _GEN_111821 : _GEN_107981; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_116048 = 4'h3 < realFlowNum_1 ? _GEN_111822 : _GEN_107982; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_116049 = 4'h3 < realFlowNum_1 ? _GEN_111823 : _GEN_107983; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_116050 = 4'h3 < realFlowNum_1 ? _GEN_111824 : _GEN_107984; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_116051 = 4'h3 < realFlowNum_1 ? _GEN_111825 : _GEN_107985; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_116052 = 4'h3 < realFlowNum_1 ? _GEN_111826 : _GEN_107986; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_116053 = 4'h3 < realFlowNum_1 ? _GEN_111827 : _GEN_107987; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_116054 = 4'h3 < realFlowNum_1 ? _GEN_111828 : _GEN_107988; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_116055 = 4'h3 < realFlowNum_1 ? _GEN_111829 : _GEN_107989; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_116056 = 4'h3 < realFlowNum_1 ? _GEN_111830 : _GEN_107990; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_116057 = 4'h3 < realFlowNum_1 ? _GEN_111831 : _GEN_107991; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_116058 = 4'h3 < realFlowNum_1 ? _GEN_111832 : _GEN_107992; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_116059 = 4'h3 < realFlowNum_1 ? _GEN_111833 : _GEN_107993; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_116060 = 4'h3 < realFlowNum_1 ? _GEN_111834 : _GEN_107994; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_116317 = _GEN_162068 | _GEN_112476; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_116318 = _GEN_162069 | _GEN_112477; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_116319 = _GEN_162070 | _GEN_112478; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_116320 = _GEN_162071 | _GEN_112479; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_116321 = _GEN_162072 | _GEN_112480; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_116322 = _GEN_162073 | _GEN_112481; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_116323 = _GEN_162074 | _GEN_112482; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_116324 = _GEN_162075 | _GEN_112483; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_116325 = _GEN_162076 | _GEN_112484; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_116326 = _GEN_162077 | _GEN_112485; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_116327 = _GEN_162078 | _GEN_112486; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_116328 = _GEN_162079 | _GEN_112487; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_116329 = _GEN_162080 | _GEN_112488; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_116330 = _GEN_162081 | _GEN_112489; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_116331 = _GEN_162082 | _GEN_112490; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_116332 = _GEN_162083 | _GEN_112491; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_116333 = _GEN_162084 | _GEN_112492; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_116334 = _GEN_162085 | _GEN_112493; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_116335 = _GEN_162086 | _GEN_112494; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_116336 = _GEN_162087 | _GEN_112495; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_116337 = _GEN_162088 | _GEN_112496; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_116338 = _GEN_162089 | _GEN_112497; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_116339 = _GEN_162090 | _GEN_112498; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_116340 = _GEN_162091 | _GEN_112499; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_116341 = _GEN_162092 | _GEN_112500; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_116342 = _GEN_162093 | _GEN_112501; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_116343 = _GEN_162094 | _GEN_112502; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_116344 = _GEN_162095 | _GEN_112503; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_116345 = _GEN_162096 | _GEN_112504; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_116346 = _GEN_162097 | _GEN_112505; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_116347 = _GEN_162098 | _GEN_112506; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_116348 = _GEN_162099 | _GEN_112507; // @[Vlflowqueue.scala 197:{51,51}]
  wire [4:0] _GEN_119293 = 5'h0 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_115452; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_119294 = 5'h1 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_115453; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_119295 = 5'h2 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_115454; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_119296 = 5'h3 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_115455; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_119297 = 5'h4 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_115456; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_119298 = 5'h5 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_115457; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_119299 = 5'h6 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_115458; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_119300 = 5'h7 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_115459; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_119301 = 5'h8 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_115460; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_119302 = 5'h9 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_115461; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_119303 = 5'ha == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_115462; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_119304 = 5'hb == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_115463; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_119305 = 5'hc == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_115464; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_119306 = 5'hd == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_115465; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_119307 = 5'he == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_115466; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_119308 = 5'hf == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_115467; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_119309 = 5'h10 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_115468; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_119310 = 5'h11 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_115469; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_119311 = 5'h12 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_115470; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_119312 = 5'h13 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_115471; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_119313 = 5'h14 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_115472; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_119314 = 5'h15 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_115473; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_119315 = 5'h16 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_115474; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_119316 = 5'h17 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_115475; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_119317 = 5'h18 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_115476; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_119318 = 5'h19 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_115477; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_119319 = 5'h1a == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_115478; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_119320 = 5'h1b == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_115479; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_119321 = 5'h1c == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_115480; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_119322 = 5'h1d == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_115481; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_119323 = 5'h1e == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_115482; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_119324 = 5'h1f == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_115483; // @[Vlflowqueue.scala 198:{51,51}]
  wire [38:0] _GEN_119869 = 5'h0 == index_1 ? vaddr_1 : _GEN_116029; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_119870 = 5'h1 == index_1 ? vaddr_1 : _GEN_116030; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_119871 = 5'h2 == index_1 ? vaddr_1 : _GEN_116031; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_119872 = 5'h3 == index_1 ? vaddr_1 : _GEN_116032; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_119873 = 5'h4 == index_1 ? vaddr_1 : _GEN_116033; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_119874 = 5'h5 == index_1 ? vaddr_1 : _GEN_116034; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_119875 = 5'h6 == index_1 ? vaddr_1 : _GEN_116035; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_119876 = 5'h7 == index_1 ? vaddr_1 : _GEN_116036; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_119877 = 5'h8 == index_1 ? vaddr_1 : _GEN_116037; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_119878 = 5'h9 == index_1 ? vaddr_1 : _GEN_116038; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_119879 = 5'ha == index_1 ? vaddr_1 : _GEN_116039; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_119880 = 5'hb == index_1 ? vaddr_1 : _GEN_116040; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_119881 = 5'hc == index_1 ? vaddr_1 : _GEN_116041; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_119882 = 5'hd == index_1 ? vaddr_1 : _GEN_116042; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_119883 = 5'he == index_1 ? vaddr_1 : _GEN_116043; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_119884 = 5'hf == index_1 ? vaddr_1 : _GEN_116044; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_119885 = 5'h10 == index_1 ? vaddr_1 : _GEN_116045; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_119886 = 5'h11 == index_1 ? vaddr_1 : _GEN_116046; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_119887 = 5'h12 == index_1 ? vaddr_1 : _GEN_116047; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_119888 = 5'h13 == index_1 ? vaddr_1 : _GEN_116048; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_119889 = 5'h14 == index_1 ? vaddr_1 : _GEN_116049; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_119890 = 5'h15 == index_1 ? vaddr_1 : _GEN_116050; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_119891 = 5'h16 == index_1 ? vaddr_1 : _GEN_116051; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_119892 = 5'h17 == index_1 ? vaddr_1 : _GEN_116052; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_119893 = 5'h18 == index_1 ? vaddr_1 : _GEN_116053; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_119894 = 5'h19 == index_1 ? vaddr_1 : _GEN_116054; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_119895 = 5'h1a == index_1 ? vaddr_1 : _GEN_116055; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_119896 = 5'h1b == index_1 ? vaddr_1 : _GEN_116056; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_119897 = 5'h1c == index_1 ? vaddr_1 : _GEN_116057; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_119898 = 5'h1d == index_1 ? vaddr_1 : _GEN_116058; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_119899 = 5'h1e == index_1 ? vaddr_1 : _GEN_116059; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_119900 = 5'h1f == index_1 ? vaddr_1 : _GEN_116060; // @[Vlflowqueue.scala 203:{51,51}]
  wire  _GEN_120542 = 4'h4 < realFlowNum_1 ? _GEN_116317 : _GEN_112476; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_120543 = 4'h4 < realFlowNum_1 ? _GEN_116318 : _GEN_112477; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_120544 = 4'h4 < realFlowNum_1 ? _GEN_116319 : _GEN_112478; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_120545 = 4'h4 < realFlowNum_1 ? _GEN_116320 : _GEN_112479; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_120546 = 4'h4 < realFlowNum_1 ? _GEN_116321 : _GEN_112480; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_120547 = 4'h4 < realFlowNum_1 ? _GEN_116322 : _GEN_112481; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_120548 = 4'h4 < realFlowNum_1 ? _GEN_116323 : _GEN_112482; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_120549 = 4'h4 < realFlowNum_1 ? _GEN_116324 : _GEN_112483; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_120550 = 4'h4 < realFlowNum_1 ? _GEN_116325 : _GEN_112484; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_120551 = 4'h4 < realFlowNum_1 ? _GEN_116326 : _GEN_112485; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_120552 = 4'h4 < realFlowNum_1 ? _GEN_116327 : _GEN_112486; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_120553 = 4'h4 < realFlowNum_1 ? _GEN_116328 : _GEN_112487; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_120554 = 4'h4 < realFlowNum_1 ? _GEN_116329 : _GEN_112488; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_120555 = 4'h4 < realFlowNum_1 ? _GEN_116330 : _GEN_112489; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_120556 = 4'h4 < realFlowNum_1 ? _GEN_116331 : _GEN_112490; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_120557 = 4'h4 < realFlowNum_1 ? _GEN_116332 : _GEN_112491; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_120558 = 4'h4 < realFlowNum_1 ? _GEN_116333 : _GEN_112492; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_120559 = 4'h4 < realFlowNum_1 ? _GEN_116334 : _GEN_112493; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_120560 = 4'h4 < realFlowNum_1 ? _GEN_116335 : _GEN_112494; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_120561 = 4'h4 < realFlowNum_1 ? _GEN_116336 : _GEN_112495; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_120562 = 4'h4 < realFlowNum_1 ? _GEN_116337 : _GEN_112496; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_120563 = 4'h4 < realFlowNum_1 ? _GEN_116338 : _GEN_112497; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_120564 = 4'h4 < realFlowNum_1 ? _GEN_116339 : _GEN_112498; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_120565 = 4'h4 < realFlowNum_1 ? _GEN_116340 : _GEN_112499; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_120566 = 4'h4 < realFlowNum_1 ? _GEN_116341 : _GEN_112500; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_120567 = 4'h4 < realFlowNum_1 ? _GEN_116342 : _GEN_112501; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_120568 = 4'h4 < realFlowNum_1 ? _GEN_116343 : _GEN_112502; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_120569 = 4'h4 < realFlowNum_1 ? _GEN_116344 : _GEN_112503; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_120570 = 4'h4 < realFlowNum_1 ? _GEN_116345 : _GEN_112504; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_120571 = 4'h4 < realFlowNum_1 ? _GEN_116346 : _GEN_112505; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_120572 = 4'h4 < realFlowNum_1 ? _GEN_116347 : _GEN_112506; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_120573 = 4'h4 < realFlowNum_1 ? _GEN_116348 : _GEN_112507; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_123518 = 4'h4 < realFlowNum_1 ? _GEN_119293 : _GEN_115452; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_123519 = 4'h4 < realFlowNum_1 ? _GEN_119294 : _GEN_115453; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_123520 = 4'h4 < realFlowNum_1 ? _GEN_119295 : _GEN_115454; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_123521 = 4'h4 < realFlowNum_1 ? _GEN_119296 : _GEN_115455; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_123522 = 4'h4 < realFlowNum_1 ? _GEN_119297 : _GEN_115456; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_123523 = 4'h4 < realFlowNum_1 ? _GEN_119298 : _GEN_115457; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_123524 = 4'h4 < realFlowNum_1 ? _GEN_119299 : _GEN_115458; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_123525 = 4'h4 < realFlowNum_1 ? _GEN_119300 : _GEN_115459; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_123526 = 4'h4 < realFlowNum_1 ? _GEN_119301 : _GEN_115460; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_123527 = 4'h4 < realFlowNum_1 ? _GEN_119302 : _GEN_115461; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_123528 = 4'h4 < realFlowNum_1 ? _GEN_119303 : _GEN_115462; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_123529 = 4'h4 < realFlowNum_1 ? _GEN_119304 : _GEN_115463; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_123530 = 4'h4 < realFlowNum_1 ? _GEN_119305 : _GEN_115464; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_123531 = 4'h4 < realFlowNum_1 ? _GEN_119306 : _GEN_115465; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_123532 = 4'h4 < realFlowNum_1 ? _GEN_119307 : _GEN_115466; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_123533 = 4'h4 < realFlowNum_1 ? _GEN_119308 : _GEN_115467; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_123534 = 4'h4 < realFlowNum_1 ? _GEN_119309 : _GEN_115468; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_123535 = 4'h4 < realFlowNum_1 ? _GEN_119310 : _GEN_115469; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_123536 = 4'h4 < realFlowNum_1 ? _GEN_119311 : _GEN_115470; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_123537 = 4'h4 < realFlowNum_1 ? _GEN_119312 : _GEN_115471; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_123538 = 4'h4 < realFlowNum_1 ? _GEN_119313 : _GEN_115472; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_123539 = 4'h4 < realFlowNum_1 ? _GEN_119314 : _GEN_115473; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_123540 = 4'h4 < realFlowNum_1 ? _GEN_119315 : _GEN_115474; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_123541 = 4'h4 < realFlowNum_1 ? _GEN_119316 : _GEN_115475; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_123542 = 4'h4 < realFlowNum_1 ? _GEN_119317 : _GEN_115476; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_123543 = 4'h4 < realFlowNum_1 ? _GEN_119318 : _GEN_115477; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_123544 = 4'h4 < realFlowNum_1 ? _GEN_119319 : _GEN_115478; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_123545 = 4'h4 < realFlowNum_1 ? _GEN_119320 : _GEN_115479; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_123546 = 4'h4 < realFlowNum_1 ? _GEN_119321 : _GEN_115480; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_123547 = 4'h4 < realFlowNum_1 ? _GEN_119322 : _GEN_115481; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_123548 = 4'h4 < realFlowNum_1 ? _GEN_119323 : _GEN_115482; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_123549 = 4'h4 < realFlowNum_1 ? _GEN_119324 : _GEN_115483; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_124095 = 4'h4 < realFlowNum_1 ? _GEN_119869 : _GEN_116029; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_124096 = 4'h4 < realFlowNum_1 ? _GEN_119870 : _GEN_116030; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_124097 = 4'h4 < realFlowNum_1 ? _GEN_119871 : _GEN_116031; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_124098 = 4'h4 < realFlowNum_1 ? _GEN_119872 : _GEN_116032; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_124099 = 4'h4 < realFlowNum_1 ? _GEN_119873 : _GEN_116033; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_124100 = 4'h4 < realFlowNum_1 ? _GEN_119874 : _GEN_116034; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_124101 = 4'h4 < realFlowNum_1 ? _GEN_119875 : _GEN_116035; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_124102 = 4'h4 < realFlowNum_1 ? _GEN_119876 : _GEN_116036; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_124103 = 4'h4 < realFlowNum_1 ? _GEN_119877 : _GEN_116037; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_124104 = 4'h4 < realFlowNum_1 ? _GEN_119878 : _GEN_116038; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_124105 = 4'h4 < realFlowNum_1 ? _GEN_119879 : _GEN_116039; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_124106 = 4'h4 < realFlowNum_1 ? _GEN_119880 : _GEN_116040; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_124107 = 4'h4 < realFlowNum_1 ? _GEN_119881 : _GEN_116041; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_124108 = 4'h4 < realFlowNum_1 ? _GEN_119882 : _GEN_116042; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_124109 = 4'h4 < realFlowNum_1 ? _GEN_119883 : _GEN_116043; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_124110 = 4'h4 < realFlowNum_1 ? _GEN_119884 : _GEN_116044; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_124111 = 4'h4 < realFlowNum_1 ? _GEN_119885 : _GEN_116045; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_124112 = 4'h4 < realFlowNum_1 ? _GEN_119886 : _GEN_116046; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_124113 = 4'h4 < realFlowNum_1 ? _GEN_119887 : _GEN_116047; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_124114 = 4'h4 < realFlowNum_1 ? _GEN_119888 : _GEN_116048; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_124115 = 4'h4 < realFlowNum_1 ? _GEN_119889 : _GEN_116049; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_124116 = 4'h4 < realFlowNum_1 ? _GEN_119890 : _GEN_116050; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_124117 = 4'h4 < realFlowNum_1 ? _GEN_119891 : _GEN_116051; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_124118 = 4'h4 < realFlowNum_1 ? _GEN_119892 : _GEN_116052; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_124119 = 4'h4 < realFlowNum_1 ? _GEN_119893 : _GEN_116053; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_124120 = 4'h4 < realFlowNum_1 ? _GEN_119894 : _GEN_116054; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_124121 = 4'h4 < realFlowNum_1 ? _GEN_119895 : _GEN_116055; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_124122 = 4'h4 < realFlowNum_1 ? _GEN_119896 : _GEN_116056; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_124123 = 4'h4 < realFlowNum_1 ? _GEN_119897 : _GEN_116057; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_124124 = 4'h4 < realFlowNum_1 ? _GEN_119898 : _GEN_116058; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_124125 = 4'h4 < realFlowNum_1 ? _GEN_119899 : _GEN_116059; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_124126 = 4'h4 < realFlowNum_1 ? _GEN_119900 : _GEN_116060; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_124383 = _GEN_162068 | _GEN_120542; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_124384 = _GEN_162069 | _GEN_120543; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_124385 = _GEN_162070 | _GEN_120544; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_124386 = _GEN_162071 | _GEN_120545; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_124387 = _GEN_162072 | _GEN_120546; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_124388 = _GEN_162073 | _GEN_120547; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_124389 = _GEN_162074 | _GEN_120548; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_124390 = _GEN_162075 | _GEN_120549; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_124391 = _GEN_162076 | _GEN_120550; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_124392 = _GEN_162077 | _GEN_120551; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_124393 = _GEN_162078 | _GEN_120552; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_124394 = _GEN_162079 | _GEN_120553; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_124395 = _GEN_162080 | _GEN_120554; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_124396 = _GEN_162081 | _GEN_120555; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_124397 = _GEN_162082 | _GEN_120556; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_124398 = _GEN_162083 | _GEN_120557; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_124399 = _GEN_162084 | _GEN_120558; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_124400 = _GEN_162085 | _GEN_120559; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_124401 = _GEN_162086 | _GEN_120560; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_124402 = _GEN_162087 | _GEN_120561; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_124403 = _GEN_162088 | _GEN_120562; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_124404 = _GEN_162089 | _GEN_120563; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_124405 = _GEN_162090 | _GEN_120564; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_124406 = _GEN_162091 | _GEN_120565; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_124407 = _GEN_162092 | _GEN_120566; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_124408 = _GEN_162093 | _GEN_120567; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_124409 = _GEN_162094 | _GEN_120568; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_124410 = _GEN_162095 | _GEN_120569; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_124411 = _GEN_162096 | _GEN_120570; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_124412 = _GEN_162097 | _GEN_120571; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_124413 = _GEN_162098 | _GEN_120572; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_124414 = _GEN_162099 | _GEN_120573; // @[Vlflowqueue.scala 197:{51,51}]
  wire [4:0] _GEN_127359 = 5'h0 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_123518; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_127360 = 5'h1 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_123519; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_127361 = 5'h2 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_123520; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_127362 = 5'h3 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_123521; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_127363 = 5'h4 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_123522; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_127364 = 5'h5 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_123523; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_127365 = 5'h6 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_123524; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_127366 = 5'h7 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_123525; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_127367 = 5'h8 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_123526; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_127368 = 5'h9 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_123527; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_127369 = 5'ha == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_123528; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_127370 = 5'hb == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_123529; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_127371 = 5'hc == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_123530; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_127372 = 5'hd == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_123531; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_127373 = 5'he == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_123532; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_127374 = 5'hf == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_123533; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_127375 = 5'h10 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_123534; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_127376 = 5'h11 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_123535; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_127377 = 5'h12 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_123536; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_127378 = 5'h13 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_123537; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_127379 = 5'h14 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_123538; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_127380 = 5'h15 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_123539; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_127381 = 5'h16 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_123540; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_127382 = 5'h17 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_123541; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_127383 = 5'h18 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_123542; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_127384 = 5'h19 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_123543; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_127385 = 5'h1a == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_123544; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_127386 = 5'h1b == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_123545; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_127387 = 5'h1c == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_123546; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_127388 = 5'h1d == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_123547; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_127389 = 5'h1e == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_123548; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_127390 = 5'h1f == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_123549; // @[Vlflowqueue.scala 198:{51,51}]
  wire [38:0] _GEN_127935 = 5'h0 == index_1 ? vaddr_1 : _GEN_124095; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_127936 = 5'h1 == index_1 ? vaddr_1 : _GEN_124096; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_127937 = 5'h2 == index_1 ? vaddr_1 : _GEN_124097; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_127938 = 5'h3 == index_1 ? vaddr_1 : _GEN_124098; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_127939 = 5'h4 == index_1 ? vaddr_1 : _GEN_124099; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_127940 = 5'h5 == index_1 ? vaddr_1 : _GEN_124100; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_127941 = 5'h6 == index_1 ? vaddr_1 : _GEN_124101; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_127942 = 5'h7 == index_1 ? vaddr_1 : _GEN_124102; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_127943 = 5'h8 == index_1 ? vaddr_1 : _GEN_124103; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_127944 = 5'h9 == index_1 ? vaddr_1 : _GEN_124104; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_127945 = 5'ha == index_1 ? vaddr_1 : _GEN_124105; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_127946 = 5'hb == index_1 ? vaddr_1 : _GEN_124106; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_127947 = 5'hc == index_1 ? vaddr_1 : _GEN_124107; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_127948 = 5'hd == index_1 ? vaddr_1 : _GEN_124108; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_127949 = 5'he == index_1 ? vaddr_1 : _GEN_124109; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_127950 = 5'hf == index_1 ? vaddr_1 : _GEN_124110; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_127951 = 5'h10 == index_1 ? vaddr_1 : _GEN_124111; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_127952 = 5'h11 == index_1 ? vaddr_1 : _GEN_124112; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_127953 = 5'h12 == index_1 ? vaddr_1 : _GEN_124113; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_127954 = 5'h13 == index_1 ? vaddr_1 : _GEN_124114; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_127955 = 5'h14 == index_1 ? vaddr_1 : _GEN_124115; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_127956 = 5'h15 == index_1 ? vaddr_1 : _GEN_124116; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_127957 = 5'h16 == index_1 ? vaddr_1 : _GEN_124117; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_127958 = 5'h17 == index_1 ? vaddr_1 : _GEN_124118; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_127959 = 5'h18 == index_1 ? vaddr_1 : _GEN_124119; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_127960 = 5'h19 == index_1 ? vaddr_1 : _GEN_124120; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_127961 = 5'h1a == index_1 ? vaddr_1 : _GEN_124121; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_127962 = 5'h1b == index_1 ? vaddr_1 : _GEN_124122; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_127963 = 5'h1c == index_1 ? vaddr_1 : _GEN_124123; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_127964 = 5'h1d == index_1 ? vaddr_1 : _GEN_124124; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_127965 = 5'h1e == index_1 ? vaddr_1 : _GEN_124125; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_127966 = 5'h1f == index_1 ? vaddr_1 : _GEN_124126; // @[Vlflowqueue.scala 203:{51,51}]
  wire  _GEN_128608 = 4'h5 < realFlowNum_1 ? _GEN_124383 : _GEN_120542; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_128609 = 4'h5 < realFlowNum_1 ? _GEN_124384 : _GEN_120543; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_128610 = 4'h5 < realFlowNum_1 ? _GEN_124385 : _GEN_120544; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_128611 = 4'h5 < realFlowNum_1 ? _GEN_124386 : _GEN_120545; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_128612 = 4'h5 < realFlowNum_1 ? _GEN_124387 : _GEN_120546; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_128613 = 4'h5 < realFlowNum_1 ? _GEN_124388 : _GEN_120547; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_128614 = 4'h5 < realFlowNum_1 ? _GEN_124389 : _GEN_120548; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_128615 = 4'h5 < realFlowNum_1 ? _GEN_124390 : _GEN_120549; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_128616 = 4'h5 < realFlowNum_1 ? _GEN_124391 : _GEN_120550; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_128617 = 4'h5 < realFlowNum_1 ? _GEN_124392 : _GEN_120551; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_128618 = 4'h5 < realFlowNum_1 ? _GEN_124393 : _GEN_120552; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_128619 = 4'h5 < realFlowNum_1 ? _GEN_124394 : _GEN_120553; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_128620 = 4'h5 < realFlowNum_1 ? _GEN_124395 : _GEN_120554; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_128621 = 4'h5 < realFlowNum_1 ? _GEN_124396 : _GEN_120555; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_128622 = 4'h5 < realFlowNum_1 ? _GEN_124397 : _GEN_120556; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_128623 = 4'h5 < realFlowNum_1 ? _GEN_124398 : _GEN_120557; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_128624 = 4'h5 < realFlowNum_1 ? _GEN_124399 : _GEN_120558; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_128625 = 4'h5 < realFlowNum_1 ? _GEN_124400 : _GEN_120559; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_128626 = 4'h5 < realFlowNum_1 ? _GEN_124401 : _GEN_120560; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_128627 = 4'h5 < realFlowNum_1 ? _GEN_124402 : _GEN_120561; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_128628 = 4'h5 < realFlowNum_1 ? _GEN_124403 : _GEN_120562; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_128629 = 4'h5 < realFlowNum_1 ? _GEN_124404 : _GEN_120563; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_128630 = 4'h5 < realFlowNum_1 ? _GEN_124405 : _GEN_120564; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_128631 = 4'h5 < realFlowNum_1 ? _GEN_124406 : _GEN_120565; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_128632 = 4'h5 < realFlowNum_1 ? _GEN_124407 : _GEN_120566; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_128633 = 4'h5 < realFlowNum_1 ? _GEN_124408 : _GEN_120567; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_128634 = 4'h5 < realFlowNum_1 ? _GEN_124409 : _GEN_120568; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_128635 = 4'h5 < realFlowNum_1 ? _GEN_124410 : _GEN_120569; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_128636 = 4'h5 < realFlowNum_1 ? _GEN_124411 : _GEN_120570; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_128637 = 4'h5 < realFlowNum_1 ? _GEN_124412 : _GEN_120571; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_128638 = 4'h5 < realFlowNum_1 ? _GEN_124413 : _GEN_120572; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_128639 = 4'h5 < realFlowNum_1 ? _GEN_124414 : _GEN_120573; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_131584 = 4'h5 < realFlowNum_1 ? _GEN_127359 : _GEN_123518; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_131585 = 4'h5 < realFlowNum_1 ? _GEN_127360 : _GEN_123519; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_131586 = 4'h5 < realFlowNum_1 ? _GEN_127361 : _GEN_123520; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_131587 = 4'h5 < realFlowNum_1 ? _GEN_127362 : _GEN_123521; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_131588 = 4'h5 < realFlowNum_1 ? _GEN_127363 : _GEN_123522; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_131589 = 4'h5 < realFlowNum_1 ? _GEN_127364 : _GEN_123523; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_131590 = 4'h5 < realFlowNum_1 ? _GEN_127365 : _GEN_123524; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_131591 = 4'h5 < realFlowNum_1 ? _GEN_127366 : _GEN_123525; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_131592 = 4'h5 < realFlowNum_1 ? _GEN_127367 : _GEN_123526; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_131593 = 4'h5 < realFlowNum_1 ? _GEN_127368 : _GEN_123527; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_131594 = 4'h5 < realFlowNum_1 ? _GEN_127369 : _GEN_123528; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_131595 = 4'h5 < realFlowNum_1 ? _GEN_127370 : _GEN_123529; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_131596 = 4'h5 < realFlowNum_1 ? _GEN_127371 : _GEN_123530; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_131597 = 4'h5 < realFlowNum_1 ? _GEN_127372 : _GEN_123531; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_131598 = 4'h5 < realFlowNum_1 ? _GEN_127373 : _GEN_123532; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_131599 = 4'h5 < realFlowNum_1 ? _GEN_127374 : _GEN_123533; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_131600 = 4'h5 < realFlowNum_1 ? _GEN_127375 : _GEN_123534; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_131601 = 4'h5 < realFlowNum_1 ? _GEN_127376 : _GEN_123535; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_131602 = 4'h5 < realFlowNum_1 ? _GEN_127377 : _GEN_123536; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_131603 = 4'h5 < realFlowNum_1 ? _GEN_127378 : _GEN_123537; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_131604 = 4'h5 < realFlowNum_1 ? _GEN_127379 : _GEN_123538; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_131605 = 4'h5 < realFlowNum_1 ? _GEN_127380 : _GEN_123539; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_131606 = 4'h5 < realFlowNum_1 ? _GEN_127381 : _GEN_123540; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_131607 = 4'h5 < realFlowNum_1 ? _GEN_127382 : _GEN_123541; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_131608 = 4'h5 < realFlowNum_1 ? _GEN_127383 : _GEN_123542; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_131609 = 4'h5 < realFlowNum_1 ? _GEN_127384 : _GEN_123543; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_131610 = 4'h5 < realFlowNum_1 ? _GEN_127385 : _GEN_123544; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_131611 = 4'h5 < realFlowNum_1 ? _GEN_127386 : _GEN_123545; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_131612 = 4'h5 < realFlowNum_1 ? _GEN_127387 : _GEN_123546; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_131613 = 4'h5 < realFlowNum_1 ? _GEN_127388 : _GEN_123547; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_131614 = 4'h5 < realFlowNum_1 ? _GEN_127389 : _GEN_123548; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_131615 = 4'h5 < realFlowNum_1 ? _GEN_127390 : _GEN_123549; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_132161 = 4'h5 < realFlowNum_1 ? _GEN_127935 : _GEN_124095; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_132162 = 4'h5 < realFlowNum_1 ? _GEN_127936 : _GEN_124096; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_132163 = 4'h5 < realFlowNum_1 ? _GEN_127937 : _GEN_124097; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_132164 = 4'h5 < realFlowNum_1 ? _GEN_127938 : _GEN_124098; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_132165 = 4'h5 < realFlowNum_1 ? _GEN_127939 : _GEN_124099; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_132166 = 4'h5 < realFlowNum_1 ? _GEN_127940 : _GEN_124100; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_132167 = 4'h5 < realFlowNum_1 ? _GEN_127941 : _GEN_124101; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_132168 = 4'h5 < realFlowNum_1 ? _GEN_127942 : _GEN_124102; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_132169 = 4'h5 < realFlowNum_1 ? _GEN_127943 : _GEN_124103; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_132170 = 4'h5 < realFlowNum_1 ? _GEN_127944 : _GEN_124104; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_132171 = 4'h5 < realFlowNum_1 ? _GEN_127945 : _GEN_124105; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_132172 = 4'h5 < realFlowNum_1 ? _GEN_127946 : _GEN_124106; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_132173 = 4'h5 < realFlowNum_1 ? _GEN_127947 : _GEN_124107; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_132174 = 4'h5 < realFlowNum_1 ? _GEN_127948 : _GEN_124108; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_132175 = 4'h5 < realFlowNum_1 ? _GEN_127949 : _GEN_124109; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_132176 = 4'h5 < realFlowNum_1 ? _GEN_127950 : _GEN_124110; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_132177 = 4'h5 < realFlowNum_1 ? _GEN_127951 : _GEN_124111; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_132178 = 4'h5 < realFlowNum_1 ? _GEN_127952 : _GEN_124112; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_132179 = 4'h5 < realFlowNum_1 ? _GEN_127953 : _GEN_124113; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_132180 = 4'h5 < realFlowNum_1 ? _GEN_127954 : _GEN_124114; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_132181 = 4'h5 < realFlowNum_1 ? _GEN_127955 : _GEN_124115; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_132182 = 4'h5 < realFlowNum_1 ? _GEN_127956 : _GEN_124116; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_132183 = 4'h5 < realFlowNum_1 ? _GEN_127957 : _GEN_124117; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_132184 = 4'h5 < realFlowNum_1 ? _GEN_127958 : _GEN_124118; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_132185 = 4'h5 < realFlowNum_1 ? _GEN_127959 : _GEN_124119; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_132186 = 4'h5 < realFlowNum_1 ? _GEN_127960 : _GEN_124120; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_132187 = 4'h5 < realFlowNum_1 ? _GEN_127961 : _GEN_124121; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_132188 = 4'h5 < realFlowNum_1 ? _GEN_127962 : _GEN_124122; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_132189 = 4'h5 < realFlowNum_1 ? _GEN_127963 : _GEN_124123; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_132190 = 4'h5 < realFlowNum_1 ? _GEN_127964 : _GEN_124124; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_132191 = 4'h5 < realFlowNum_1 ? _GEN_127965 : _GEN_124125; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_132192 = 4'h5 < realFlowNum_1 ? _GEN_127966 : _GEN_124126; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_132449 = _GEN_162068 | _GEN_128608; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_132450 = _GEN_162069 | _GEN_128609; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_132451 = _GEN_162070 | _GEN_128610; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_132452 = _GEN_162071 | _GEN_128611; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_132453 = _GEN_162072 | _GEN_128612; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_132454 = _GEN_162073 | _GEN_128613; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_132455 = _GEN_162074 | _GEN_128614; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_132456 = _GEN_162075 | _GEN_128615; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_132457 = _GEN_162076 | _GEN_128616; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_132458 = _GEN_162077 | _GEN_128617; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_132459 = _GEN_162078 | _GEN_128618; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_132460 = _GEN_162079 | _GEN_128619; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_132461 = _GEN_162080 | _GEN_128620; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_132462 = _GEN_162081 | _GEN_128621; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_132463 = _GEN_162082 | _GEN_128622; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_132464 = _GEN_162083 | _GEN_128623; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_132465 = _GEN_162084 | _GEN_128624; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_132466 = _GEN_162085 | _GEN_128625; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_132467 = _GEN_162086 | _GEN_128626; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_132468 = _GEN_162087 | _GEN_128627; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_132469 = _GEN_162088 | _GEN_128628; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_132470 = _GEN_162089 | _GEN_128629; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_132471 = _GEN_162090 | _GEN_128630; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_132472 = _GEN_162091 | _GEN_128631; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_132473 = _GEN_162092 | _GEN_128632; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_132474 = _GEN_162093 | _GEN_128633; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_132475 = _GEN_162094 | _GEN_128634; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_132476 = _GEN_162095 | _GEN_128635; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_132477 = _GEN_162096 | _GEN_128636; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_132478 = _GEN_162097 | _GEN_128637; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_132479 = _GEN_162098 | _GEN_128638; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_132480 = _GEN_162099 | _GEN_128639; // @[Vlflowqueue.scala 197:{51,51}]
  wire [4:0] _GEN_135425 = 5'h0 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_131584; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_135426 = 5'h1 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_131585; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_135427 = 5'h2 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_131586; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_135428 = 5'h3 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_131587; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_135429 = 5'h4 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_131588; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_135430 = 5'h5 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_131589; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_135431 = 5'h6 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_131590; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_135432 = 5'h7 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_131591; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_135433 = 5'h8 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_131592; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_135434 = 5'h9 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_131593; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_135435 = 5'ha == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_131594; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_135436 = 5'hb == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_131595; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_135437 = 5'hc == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_131596; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_135438 = 5'hd == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_131597; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_135439 = 5'he == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_131598; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_135440 = 5'hf == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_131599; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_135441 = 5'h10 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_131600; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_135442 = 5'h11 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_131601; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_135443 = 5'h12 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_131602; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_135444 = 5'h13 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_131603; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_135445 = 5'h14 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_131604; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_135446 = 5'h15 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_131605; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_135447 = 5'h16 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_131606; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_135448 = 5'h17 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_131607; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_135449 = 5'h18 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_131608; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_135450 = 5'h19 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_131609; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_135451 = 5'h1a == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_131610; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_135452 = 5'h1b == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_131611; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_135453 = 5'h1c == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_131612; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_135454 = 5'h1d == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_131613; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_135455 = 5'h1e == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_131614; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_135456 = 5'h1f == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_131615; // @[Vlflowqueue.scala 198:{51,51}]
  wire [38:0] _GEN_136001 = 5'h0 == index_1 ? vaddr_1 : _GEN_132161; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_136002 = 5'h1 == index_1 ? vaddr_1 : _GEN_132162; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_136003 = 5'h2 == index_1 ? vaddr_1 : _GEN_132163; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_136004 = 5'h3 == index_1 ? vaddr_1 : _GEN_132164; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_136005 = 5'h4 == index_1 ? vaddr_1 : _GEN_132165; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_136006 = 5'h5 == index_1 ? vaddr_1 : _GEN_132166; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_136007 = 5'h6 == index_1 ? vaddr_1 : _GEN_132167; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_136008 = 5'h7 == index_1 ? vaddr_1 : _GEN_132168; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_136009 = 5'h8 == index_1 ? vaddr_1 : _GEN_132169; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_136010 = 5'h9 == index_1 ? vaddr_1 : _GEN_132170; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_136011 = 5'ha == index_1 ? vaddr_1 : _GEN_132171; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_136012 = 5'hb == index_1 ? vaddr_1 : _GEN_132172; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_136013 = 5'hc == index_1 ? vaddr_1 : _GEN_132173; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_136014 = 5'hd == index_1 ? vaddr_1 : _GEN_132174; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_136015 = 5'he == index_1 ? vaddr_1 : _GEN_132175; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_136016 = 5'hf == index_1 ? vaddr_1 : _GEN_132176; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_136017 = 5'h10 == index_1 ? vaddr_1 : _GEN_132177; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_136018 = 5'h11 == index_1 ? vaddr_1 : _GEN_132178; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_136019 = 5'h12 == index_1 ? vaddr_1 : _GEN_132179; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_136020 = 5'h13 == index_1 ? vaddr_1 : _GEN_132180; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_136021 = 5'h14 == index_1 ? vaddr_1 : _GEN_132181; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_136022 = 5'h15 == index_1 ? vaddr_1 : _GEN_132182; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_136023 = 5'h16 == index_1 ? vaddr_1 : _GEN_132183; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_136024 = 5'h17 == index_1 ? vaddr_1 : _GEN_132184; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_136025 = 5'h18 == index_1 ? vaddr_1 : _GEN_132185; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_136026 = 5'h19 == index_1 ? vaddr_1 : _GEN_132186; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_136027 = 5'h1a == index_1 ? vaddr_1 : _GEN_132187; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_136028 = 5'h1b == index_1 ? vaddr_1 : _GEN_132188; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_136029 = 5'h1c == index_1 ? vaddr_1 : _GEN_132189; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_136030 = 5'h1d == index_1 ? vaddr_1 : _GEN_132190; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_136031 = 5'h1e == index_1 ? vaddr_1 : _GEN_132191; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_136032 = 5'h1f == index_1 ? vaddr_1 : _GEN_132192; // @[Vlflowqueue.scala 203:{51,51}]
  wire  _GEN_136674 = 4'h6 < realFlowNum_1 ? _GEN_132449 : _GEN_128608; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_136675 = 4'h6 < realFlowNum_1 ? _GEN_132450 : _GEN_128609; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_136676 = 4'h6 < realFlowNum_1 ? _GEN_132451 : _GEN_128610; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_136677 = 4'h6 < realFlowNum_1 ? _GEN_132452 : _GEN_128611; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_136678 = 4'h6 < realFlowNum_1 ? _GEN_132453 : _GEN_128612; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_136679 = 4'h6 < realFlowNum_1 ? _GEN_132454 : _GEN_128613; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_136680 = 4'h6 < realFlowNum_1 ? _GEN_132455 : _GEN_128614; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_136681 = 4'h6 < realFlowNum_1 ? _GEN_132456 : _GEN_128615; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_136682 = 4'h6 < realFlowNum_1 ? _GEN_132457 : _GEN_128616; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_136683 = 4'h6 < realFlowNum_1 ? _GEN_132458 : _GEN_128617; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_136684 = 4'h6 < realFlowNum_1 ? _GEN_132459 : _GEN_128618; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_136685 = 4'h6 < realFlowNum_1 ? _GEN_132460 : _GEN_128619; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_136686 = 4'h6 < realFlowNum_1 ? _GEN_132461 : _GEN_128620; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_136687 = 4'h6 < realFlowNum_1 ? _GEN_132462 : _GEN_128621; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_136688 = 4'h6 < realFlowNum_1 ? _GEN_132463 : _GEN_128622; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_136689 = 4'h6 < realFlowNum_1 ? _GEN_132464 : _GEN_128623; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_136690 = 4'h6 < realFlowNum_1 ? _GEN_132465 : _GEN_128624; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_136691 = 4'h6 < realFlowNum_1 ? _GEN_132466 : _GEN_128625; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_136692 = 4'h6 < realFlowNum_1 ? _GEN_132467 : _GEN_128626; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_136693 = 4'h6 < realFlowNum_1 ? _GEN_132468 : _GEN_128627; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_136694 = 4'h6 < realFlowNum_1 ? _GEN_132469 : _GEN_128628; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_136695 = 4'h6 < realFlowNum_1 ? _GEN_132470 : _GEN_128629; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_136696 = 4'h6 < realFlowNum_1 ? _GEN_132471 : _GEN_128630; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_136697 = 4'h6 < realFlowNum_1 ? _GEN_132472 : _GEN_128631; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_136698 = 4'h6 < realFlowNum_1 ? _GEN_132473 : _GEN_128632; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_136699 = 4'h6 < realFlowNum_1 ? _GEN_132474 : _GEN_128633; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_136700 = 4'h6 < realFlowNum_1 ? _GEN_132475 : _GEN_128634; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_136701 = 4'h6 < realFlowNum_1 ? _GEN_132476 : _GEN_128635; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_136702 = 4'h6 < realFlowNum_1 ? _GEN_132477 : _GEN_128636; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_136703 = 4'h6 < realFlowNum_1 ? _GEN_132478 : _GEN_128637; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_136704 = 4'h6 < realFlowNum_1 ? _GEN_132479 : _GEN_128638; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_136705 = 4'h6 < realFlowNum_1 ? _GEN_132480 : _GEN_128639; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_139650 = 4'h6 < realFlowNum_1 ? _GEN_135425 : _GEN_131584; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_139651 = 4'h6 < realFlowNum_1 ? _GEN_135426 : _GEN_131585; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_139652 = 4'h6 < realFlowNum_1 ? _GEN_135427 : _GEN_131586; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_139653 = 4'h6 < realFlowNum_1 ? _GEN_135428 : _GEN_131587; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_139654 = 4'h6 < realFlowNum_1 ? _GEN_135429 : _GEN_131588; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_139655 = 4'h6 < realFlowNum_1 ? _GEN_135430 : _GEN_131589; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_139656 = 4'h6 < realFlowNum_1 ? _GEN_135431 : _GEN_131590; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_139657 = 4'h6 < realFlowNum_1 ? _GEN_135432 : _GEN_131591; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_139658 = 4'h6 < realFlowNum_1 ? _GEN_135433 : _GEN_131592; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_139659 = 4'h6 < realFlowNum_1 ? _GEN_135434 : _GEN_131593; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_139660 = 4'h6 < realFlowNum_1 ? _GEN_135435 : _GEN_131594; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_139661 = 4'h6 < realFlowNum_1 ? _GEN_135436 : _GEN_131595; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_139662 = 4'h6 < realFlowNum_1 ? _GEN_135437 : _GEN_131596; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_139663 = 4'h6 < realFlowNum_1 ? _GEN_135438 : _GEN_131597; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_139664 = 4'h6 < realFlowNum_1 ? _GEN_135439 : _GEN_131598; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_139665 = 4'h6 < realFlowNum_1 ? _GEN_135440 : _GEN_131599; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_139666 = 4'h6 < realFlowNum_1 ? _GEN_135441 : _GEN_131600; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_139667 = 4'h6 < realFlowNum_1 ? _GEN_135442 : _GEN_131601; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_139668 = 4'h6 < realFlowNum_1 ? _GEN_135443 : _GEN_131602; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_139669 = 4'h6 < realFlowNum_1 ? _GEN_135444 : _GEN_131603; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_139670 = 4'h6 < realFlowNum_1 ? _GEN_135445 : _GEN_131604; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_139671 = 4'h6 < realFlowNum_1 ? _GEN_135446 : _GEN_131605; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_139672 = 4'h6 < realFlowNum_1 ? _GEN_135447 : _GEN_131606; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_139673 = 4'h6 < realFlowNum_1 ? _GEN_135448 : _GEN_131607; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_139674 = 4'h6 < realFlowNum_1 ? _GEN_135449 : _GEN_131608; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_139675 = 4'h6 < realFlowNum_1 ? _GEN_135450 : _GEN_131609; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_139676 = 4'h6 < realFlowNum_1 ? _GEN_135451 : _GEN_131610; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_139677 = 4'h6 < realFlowNum_1 ? _GEN_135452 : _GEN_131611; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_139678 = 4'h6 < realFlowNum_1 ? _GEN_135453 : _GEN_131612; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_139679 = 4'h6 < realFlowNum_1 ? _GEN_135454 : _GEN_131613; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_139680 = 4'h6 < realFlowNum_1 ? _GEN_135455 : _GEN_131614; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_139681 = 4'h6 < realFlowNum_1 ? _GEN_135456 : _GEN_131615; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_140227 = 4'h6 < realFlowNum_1 ? _GEN_136001 : _GEN_132161; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_140228 = 4'h6 < realFlowNum_1 ? _GEN_136002 : _GEN_132162; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_140229 = 4'h6 < realFlowNum_1 ? _GEN_136003 : _GEN_132163; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_140230 = 4'h6 < realFlowNum_1 ? _GEN_136004 : _GEN_132164; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_140231 = 4'h6 < realFlowNum_1 ? _GEN_136005 : _GEN_132165; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_140232 = 4'h6 < realFlowNum_1 ? _GEN_136006 : _GEN_132166; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_140233 = 4'h6 < realFlowNum_1 ? _GEN_136007 : _GEN_132167; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_140234 = 4'h6 < realFlowNum_1 ? _GEN_136008 : _GEN_132168; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_140235 = 4'h6 < realFlowNum_1 ? _GEN_136009 : _GEN_132169; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_140236 = 4'h6 < realFlowNum_1 ? _GEN_136010 : _GEN_132170; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_140237 = 4'h6 < realFlowNum_1 ? _GEN_136011 : _GEN_132171; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_140238 = 4'h6 < realFlowNum_1 ? _GEN_136012 : _GEN_132172; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_140239 = 4'h6 < realFlowNum_1 ? _GEN_136013 : _GEN_132173; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_140240 = 4'h6 < realFlowNum_1 ? _GEN_136014 : _GEN_132174; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_140241 = 4'h6 < realFlowNum_1 ? _GEN_136015 : _GEN_132175; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_140242 = 4'h6 < realFlowNum_1 ? _GEN_136016 : _GEN_132176; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_140243 = 4'h6 < realFlowNum_1 ? _GEN_136017 : _GEN_132177; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_140244 = 4'h6 < realFlowNum_1 ? _GEN_136018 : _GEN_132178; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_140245 = 4'h6 < realFlowNum_1 ? _GEN_136019 : _GEN_132179; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_140246 = 4'h6 < realFlowNum_1 ? _GEN_136020 : _GEN_132180; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_140247 = 4'h6 < realFlowNum_1 ? _GEN_136021 : _GEN_132181; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_140248 = 4'h6 < realFlowNum_1 ? _GEN_136022 : _GEN_132182; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_140249 = 4'h6 < realFlowNum_1 ? _GEN_136023 : _GEN_132183; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_140250 = 4'h6 < realFlowNum_1 ? _GEN_136024 : _GEN_132184; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_140251 = 4'h6 < realFlowNum_1 ? _GEN_136025 : _GEN_132185; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_140252 = 4'h6 < realFlowNum_1 ? _GEN_136026 : _GEN_132186; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_140253 = 4'h6 < realFlowNum_1 ? _GEN_136027 : _GEN_132187; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_140254 = 4'h6 < realFlowNum_1 ? _GEN_136028 : _GEN_132188; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_140255 = 4'h6 < realFlowNum_1 ? _GEN_136029 : _GEN_132189; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_140256 = 4'h6 < realFlowNum_1 ? _GEN_136030 : _GEN_132190; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_140257 = 4'h6 < realFlowNum_1 ? _GEN_136031 : _GEN_132191; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_140258 = 4'h6 < realFlowNum_1 ? _GEN_136032 : _GEN_132192; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_140515 = _GEN_162068 | _GEN_136674; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_140516 = _GEN_162069 | _GEN_136675; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_140517 = _GEN_162070 | _GEN_136676; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_140518 = _GEN_162071 | _GEN_136677; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_140519 = _GEN_162072 | _GEN_136678; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_140520 = _GEN_162073 | _GEN_136679; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_140521 = _GEN_162074 | _GEN_136680; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_140522 = _GEN_162075 | _GEN_136681; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_140523 = _GEN_162076 | _GEN_136682; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_140524 = _GEN_162077 | _GEN_136683; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_140525 = _GEN_162078 | _GEN_136684; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_140526 = _GEN_162079 | _GEN_136685; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_140527 = _GEN_162080 | _GEN_136686; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_140528 = _GEN_162081 | _GEN_136687; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_140529 = _GEN_162082 | _GEN_136688; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_140530 = _GEN_162083 | _GEN_136689; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_140531 = _GEN_162084 | _GEN_136690; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_140532 = _GEN_162085 | _GEN_136691; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_140533 = _GEN_162086 | _GEN_136692; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_140534 = _GEN_162087 | _GEN_136693; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_140535 = _GEN_162088 | _GEN_136694; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_140536 = _GEN_162089 | _GEN_136695; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_140537 = _GEN_162090 | _GEN_136696; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_140538 = _GEN_162091 | _GEN_136697; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_140539 = _GEN_162092 | _GEN_136698; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_140540 = _GEN_162093 | _GEN_136699; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_140541 = _GEN_162094 | _GEN_136700; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_140542 = _GEN_162095 | _GEN_136701; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_140543 = _GEN_162096 | _GEN_136702; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_140544 = _GEN_162097 | _GEN_136703; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_140545 = _GEN_162098 | _GEN_136704; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_140546 = _GEN_162099 | _GEN_136705; // @[Vlflowqueue.scala 197:{51,51}]
  wire [4:0] _GEN_143491 = 5'h0 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_139650; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_143492 = 5'h1 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_139651; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_143493 = 5'h2 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_139652; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_143494 = 5'h3 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_139653; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_143495 = 5'h4 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_139654; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_143496 = 5'h5 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_139655; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_143497 = 5'h6 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_139656; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_143498 = 5'h7 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_139657; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_143499 = 5'h8 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_139658; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_143500 = 5'h9 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_139659; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_143501 = 5'ha == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_139660; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_143502 = 5'hb == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_139661; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_143503 = 5'hc == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_139662; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_143504 = 5'hd == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_139663; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_143505 = 5'he == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_139664; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_143506 = 5'hf == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_139665; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_143507 = 5'h10 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_139666; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_143508 = 5'h11 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_139667; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_143509 = 5'h12 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_139668; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_143510 = 5'h13 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_139669; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_143511 = 5'h14 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_139670; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_143512 = 5'h15 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_139671; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_143513 = 5'h16 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_139672; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_143514 = 5'h17 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_139673; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_143515 = 5'h18 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_139674; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_143516 = 5'h19 == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_139675; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_143517 = 5'h1a == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_139676; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_143518 = 5'h1b == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_139677; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_143519 = 5'h1c == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_139678; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_143520 = 5'h1d == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_139679; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_143521 = 5'h1e == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_139680; // @[Vlflowqueue.scala 198:{51,51}]
  wire [4:0] _GEN_143522 = 5'h1f == index_1 ? io_loadRegIn_1_bits_uop_robIdx_value : _GEN_139681; // @[Vlflowqueue.scala 198:{51,51}]
  wire [38:0] _GEN_144067 = 5'h0 == index_1 ? vaddr_1 : _GEN_140227; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_144068 = 5'h1 == index_1 ? vaddr_1 : _GEN_140228; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_144069 = 5'h2 == index_1 ? vaddr_1 : _GEN_140229; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_144070 = 5'h3 == index_1 ? vaddr_1 : _GEN_140230; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_144071 = 5'h4 == index_1 ? vaddr_1 : _GEN_140231; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_144072 = 5'h5 == index_1 ? vaddr_1 : _GEN_140232; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_144073 = 5'h6 == index_1 ? vaddr_1 : _GEN_140233; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_144074 = 5'h7 == index_1 ? vaddr_1 : _GEN_140234; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_144075 = 5'h8 == index_1 ? vaddr_1 : _GEN_140235; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_144076 = 5'h9 == index_1 ? vaddr_1 : _GEN_140236; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_144077 = 5'ha == index_1 ? vaddr_1 : _GEN_140237; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_144078 = 5'hb == index_1 ? vaddr_1 : _GEN_140238; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_144079 = 5'hc == index_1 ? vaddr_1 : _GEN_140239; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_144080 = 5'hd == index_1 ? vaddr_1 : _GEN_140240; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_144081 = 5'he == index_1 ? vaddr_1 : _GEN_140241; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_144082 = 5'hf == index_1 ? vaddr_1 : _GEN_140242; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_144083 = 5'h10 == index_1 ? vaddr_1 : _GEN_140243; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_144084 = 5'h11 == index_1 ? vaddr_1 : _GEN_140244; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_144085 = 5'h12 == index_1 ? vaddr_1 : _GEN_140245; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_144086 = 5'h13 == index_1 ? vaddr_1 : _GEN_140246; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_144087 = 5'h14 == index_1 ? vaddr_1 : _GEN_140247; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_144088 = 5'h15 == index_1 ? vaddr_1 : _GEN_140248; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_144089 = 5'h16 == index_1 ? vaddr_1 : _GEN_140249; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_144090 = 5'h17 == index_1 ? vaddr_1 : _GEN_140250; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_144091 = 5'h18 == index_1 ? vaddr_1 : _GEN_140251; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_144092 = 5'h19 == index_1 ? vaddr_1 : _GEN_140252; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_144093 = 5'h1a == index_1 ? vaddr_1 : _GEN_140253; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_144094 = 5'h1b == index_1 ? vaddr_1 : _GEN_140254; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_144095 = 5'h1c == index_1 ? vaddr_1 : _GEN_140255; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_144096 = 5'h1d == index_1 ? vaddr_1 : _GEN_140256; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_144097 = 5'h1e == index_1 ? vaddr_1 : _GEN_140257; // @[Vlflowqueue.scala 203:{51,51}]
  wire [38:0] _GEN_144098 = 5'h1f == index_1 ? vaddr_1 : _GEN_140258; // @[Vlflowqueue.scala 203:{51,51}]
  wire  _GEN_144740 = 4'h7 < realFlowNum_1 ? _GEN_140515 : _GEN_136674; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_144741 = 4'h7 < realFlowNum_1 ? _GEN_140516 : _GEN_136675; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_144742 = 4'h7 < realFlowNum_1 ? _GEN_140517 : _GEN_136676; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_144743 = 4'h7 < realFlowNum_1 ? _GEN_140518 : _GEN_136677; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_144744 = 4'h7 < realFlowNum_1 ? _GEN_140519 : _GEN_136678; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_144745 = 4'h7 < realFlowNum_1 ? _GEN_140520 : _GEN_136679; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_144746 = 4'h7 < realFlowNum_1 ? _GEN_140521 : _GEN_136680; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_144747 = 4'h7 < realFlowNum_1 ? _GEN_140522 : _GEN_136681; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_144748 = 4'h7 < realFlowNum_1 ? _GEN_140523 : _GEN_136682; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_144749 = 4'h7 < realFlowNum_1 ? _GEN_140524 : _GEN_136683; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_144750 = 4'h7 < realFlowNum_1 ? _GEN_140525 : _GEN_136684; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_144751 = 4'h7 < realFlowNum_1 ? _GEN_140526 : _GEN_136685; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_144752 = 4'h7 < realFlowNum_1 ? _GEN_140527 : _GEN_136686; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_144753 = 4'h7 < realFlowNum_1 ? _GEN_140528 : _GEN_136687; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_144754 = 4'h7 < realFlowNum_1 ? _GEN_140529 : _GEN_136688; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_144755 = 4'h7 < realFlowNum_1 ? _GEN_140530 : _GEN_136689; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_144756 = 4'h7 < realFlowNum_1 ? _GEN_140531 : _GEN_136690; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_144757 = 4'h7 < realFlowNum_1 ? _GEN_140532 : _GEN_136691; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_144758 = 4'h7 < realFlowNum_1 ? _GEN_140533 : _GEN_136692; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_144759 = 4'h7 < realFlowNum_1 ? _GEN_140534 : _GEN_136693; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_144760 = 4'h7 < realFlowNum_1 ? _GEN_140535 : _GEN_136694; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_144761 = 4'h7 < realFlowNum_1 ? _GEN_140536 : _GEN_136695; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_144762 = 4'h7 < realFlowNum_1 ? _GEN_140537 : _GEN_136696; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_144763 = 4'h7 < realFlowNum_1 ? _GEN_140538 : _GEN_136697; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_144764 = 4'h7 < realFlowNum_1 ? _GEN_140539 : _GEN_136698; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_144765 = 4'h7 < realFlowNum_1 ? _GEN_140540 : _GEN_136699; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_144766 = 4'h7 < realFlowNum_1 ? _GEN_140541 : _GEN_136700; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_144767 = 4'h7 < realFlowNum_1 ? _GEN_140542 : _GEN_136701; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_144768 = 4'h7 < realFlowNum_1 ? _GEN_140543 : _GEN_136702; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_144769 = 4'h7 < realFlowNum_1 ? _GEN_140544 : _GEN_136703; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_144770 = 4'h7 < realFlowNum_1 ? _GEN_140545 : _GEN_136704; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_144771 = 4'h7 < realFlowNum_1 ? _GEN_140546 : _GEN_136705; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_147716 = 4'h7 < realFlowNum_1 ? _GEN_143491 : _GEN_139650; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_147717 = 4'h7 < realFlowNum_1 ? _GEN_143492 : _GEN_139651; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_147718 = 4'h7 < realFlowNum_1 ? _GEN_143493 : _GEN_139652; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_147719 = 4'h7 < realFlowNum_1 ? _GEN_143494 : _GEN_139653; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_147720 = 4'h7 < realFlowNum_1 ? _GEN_143495 : _GEN_139654; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_147721 = 4'h7 < realFlowNum_1 ? _GEN_143496 : _GEN_139655; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_147722 = 4'h7 < realFlowNum_1 ? _GEN_143497 : _GEN_139656; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_147723 = 4'h7 < realFlowNum_1 ? _GEN_143498 : _GEN_139657; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_147724 = 4'h7 < realFlowNum_1 ? _GEN_143499 : _GEN_139658; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_147725 = 4'h7 < realFlowNum_1 ? _GEN_143500 : _GEN_139659; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_147726 = 4'h7 < realFlowNum_1 ? _GEN_143501 : _GEN_139660; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_147727 = 4'h7 < realFlowNum_1 ? _GEN_143502 : _GEN_139661; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_147728 = 4'h7 < realFlowNum_1 ? _GEN_143503 : _GEN_139662; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_147729 = 4'h7 < realFlowNum_1 ? _GEN_143504 : _GEN_139663; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_147730 = 4'h7 < realFlowNum_1 ? _GEN_143505 : _GEN_139664; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_147731 = 4'h7 < realFlowNum_1 ? _GEN_143506 : _GEN_139665; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_147732 = 4'h7 < realFlowNum_1 ? _GEN_143507 : _GEN_139666; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_147733 = 4'h7 < realFlowNum_1 ? _GEN_143508 : _GEN_139667; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_147734 = 4'h7 < realFlowNum_1 ? _GEN_143509 : _GEN_139668; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_147735 = 4'h7 < realFlowNum_1 ? _GEN_143510 : _GEN_139669; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_147736 = 4'h7 < realFlowNum_1 ? _GEN_143511 : _GEN_139670; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_147737 = 4'h7 < realFlowNum_1 ? _GEN_143512 : _GEN_139671; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_147738 = 4'h7 < realFlowNum_1 ? _GEN_143513 : _GEN_139672; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_147739 = 4'h7 < realFlowNum_1 ? _GEN_143514 : _GEN_139673; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_147740 = 4'h7 < realFlowNum_1 ? _GEN_143515 : _GEN_139674; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_147741 = 4'h7 < realFlowNum_1 ? _GEN_143516 : _GEN_139675; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_147742 = 4'h7 < realFlowNum_1 ? _GEN_143517 : _GEN_139676; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_147743 = 4'h7 < realFlowNum_1 ? _GEN_143518 : _GEN_139677; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_147744 = 4'h7 < realFlowNum_1 ? _GEN_143519 : _GEN_139678; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_147745 = 4'h7 < realFlowNum_1 ? _GEN_143520 : _GEN_139679; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_147746 = 4'h7 < realFlowNum_1 ? _GEN_143521 : _GEN_139680; // @[Vlflowqueue.scala 194:37]
  wire [4:0] _GEN_147747 = 4'h7 < realFlowNum_1 ? _GEN_143522 : _GEN_139681; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_148293 = 4'h7 < realFlowNum_1 ? _GEN_144067 : _GEN_140227; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_148294 = 4'h7 < realFlowNum_1 ? _GEN_144068 : _GEN_140228; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_148295 = 4'h7 < realFlowNum_1 ? _GEN_144069 : _GEN_140229; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_148296 = 4'h7 < realFlowNum_1 ? _GEN_144070 : _GEN_140230; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_148297 = 4'h7 < realFlowNum_1 ? _GEN_144071 : _GEN_140231; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_148298 = 4'h7 < realFlowNum_1 ? _GEN_144072 : _GEN_140232; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_148299 = 4'h7 < realFlowNum_1 ? _GEN_144073 : _GEN_140233; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_148300 = 4'h7 < realFlowNum_1 ? _GEN_144074 : _GEN_140234; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_148301 = 4'h7 < realFlowNum_1 ? _GEN_144075 : _GEN_140235; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_148302 = 4'h7 < realFlowNum_1 ? _GEN_144076 : _GEN_140236; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_148303 = 4'h7 < realFlowNum_1 ? _GEN_144077 : _GEN_140237; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_148304 = 4'h7 < realFlowNum_1 ? _GEN_144078 : _GEN_140238; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_148305 = 4'h7 < realFlowNum_1 ? _GEN_144079 : _GEN_140239; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_148306 = 4'h7 < realFlowNum_1 ? _GEN_144080 : _GEN_140240; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_148307 = 4'h7 < realFlowNum_1 ? _GEN_144081 : _GEN_140241; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_148308 = 4'h7 < realFlowNum_1 ? _GEN_144082 : _GEN_140242; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_148309 = 4'h7 < realFlowNum_1 ? _GEN_144083 : _GEN_140243; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_148310 = 4'h7 < realFlowNum_1 ? _GEN_144084 : _GEN_140244; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_148311 = 4'h7 < realFlowNum_1 ? _GEN_144085 : _GEN_140245; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_148312 = 4'h7 < realFlowNum_1 ? _GEN_144086 : _GEN_140246; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_148313 = 4'h7 < realFlowNum_1 ? _GEN_144087 : _GEN_140247; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_148314 = 4'h7 < realFlowNum_1 ? _GEN_144088 : _GEN_140248; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_148315 = 4'h7 < realFlowNum_1 ? _GEN_144089 : _GEN_140249; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_148316 = 4'h7 < realFlowNum_1 ? _GEN_144090 : _GEN_140250; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_148317 = 4'h7 < realFlowNum_1 ? _GEN_144091 : _GEN_140251; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_148318 = 4'h7 < realFlowNum_1 ? _GEN_144092 : _GEN_140252; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_148319 = 4'h7 < realFlowNum_1 ? _GEN_144093 : _GEN_140253; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_148320 = 4'h7 < realFlowNum_1 ? _GEN_144094 : _GEN_140254; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_148321 = 4'h7 < realFlowNum_1 ? _GEN_144095 : _GEN_140255; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_148322 = 4'h7 < realFlowNum_1 ? _GEN_144096 : _GEN_140256; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_148323 = 4'h7 < realFlowNum_1 ? _GEN_144097 : _GEN_140257; // @[Vlflowqueue.scala 194:37]
  wire [38:0] _GEN_148324 = 4'h7 < realFlowNum_1 ? _GEN_144098 : _GEN_140258; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_148581 = _GEN_162068 | _GEN_144740; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_148582 = _GEN_162069 | _GEN_144741; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_148583 = _GEN_162070 | _GEN_144742; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_148584 = _GEN_162071 | _GEN_144743; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_148585 = _GEN_162072 | _GEN_144744; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_148586 = _GEN_162073 | _GEN_144745; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_148587 = _GEN_162074 | _GEN_144746; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_148588 = _GEN_162075 | _GEN_144747; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_148589 = _GEN_162076 | _GEN_144748; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_148590 = _GEN_162077 | _GEN_144749; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_148591 = _GEN_162078 | _GEN_144750; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_148592 = _GEN_162079 | _GEN_144751; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_148593 = _GEN_162080 | _GEN_144752; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_148594 = _GEN_162081 | _GEN_144753; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_148595 = _GEN_162082 | _GEN_144754; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_148596 = _GEN_162083 | _GEN_144755; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_148597 = _GEN_162084 | _GEN_144756; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_148598 = _GEN_162085 | _GEN_144757; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_148599 = _GEN_162086 | _GEN_144758; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_148600 = _GEN_162087 | _GEN_144759; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_148601 = _GEN_162088 | _GEN_144760; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_148602 = _GEN_162089 | _GEN_144761; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_148603 = _GEN_162090 | _GEN_144762; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_148604 = _GEN_162091 | _GEN_144763; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_148605 = _GEN_162092 | _GEN_144764; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_148606 = _GEN_162093 | _GEN_144765; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_148607 = _GEN_162094 | _GEN_144766; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_148608 = _GEN_162095 | _GEN_144767; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_148609 = _GEN_162096 | _GEN_144768; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_148610 = _GEN_162097 | _GEN_144769; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_148611 = _GEN_162098 | _GEN_144770; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_148612 = _GEN_162099 | _GEN_144771; // @[Vlflowqueue.scala 197:{51,51}]
  wire  _GEN_152806 = 4'h8 < realFlowNum_1 ? _GEN_148581 : _GEN_144740; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_152807 = 4'h8 < realFlowNum_1 ? _GEN_148582 : _GEN_144741; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_152808 = 4'h8 < realFlowNum_1 ? _GEN_148583 : _GEN_144742; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_152809 = 4'h8 < realFlowNum_1 ? _GEN_148584 : _GEN_144743; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_152810 = 4'h8 < realFlowNum_1 ? _GEN_148585 : _GEN_144744; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_152811 = 4'h8 < realFlowNum_1 ? _GEN_148586 : _GEN_144745; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_152812 = 4'h8 < realFlowNum_1 ? _GEN_148587 : _GEN_144746; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_152813 = 4'h8 < realFlowNum_1 ? _GEN_148588 : _GEN_144747; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_152814 = 4'h8 < realFlowNum_1 ? _GEN_148589 : _GEN_144748; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_152815 = 4'h8 < realFlowNum_1 ? _GEN_148590 : _GEN_144749; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_152816 = 4'h8 < realFlowNum_1 ? _GEN_148591 : _GEN_144750; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_152817 = 4'h8 < realFlowNum_1 ? _GEN_148592 : _GEN_144751; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_152818 = 4'h8 < realFlowNum_1 ? _GEN_148593 : _GEN_144752; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_152819 = 4'h8 < realFlowNum_1 ? _GEN_148594 : _GEN_144753; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_152820 = 4'h8 < realFlowNum_1 ? _GEN_148595 : _GEN_144754; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_152821 = 4'h8 < realFlowNum_1 ? _GEN_148596 : _GEN_144755; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_152822 = 4'h8 < realFlowNum_1 ? _GEN_148597 : _GEN_144756; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_152823 = 4'h8 < realFlowNum_1 ? _GEN_148598 : _GEN_144757; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_152824 = 4'h8 < realFlowNum_1 ? _GEN_148599 : _GEN_144758; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_152825 = 4'h8 < realFlowNum_1 ? _GEN_148600 : _GEN_144759; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_152826 = 4'h8 < realFlowNum_1 ? _GEN_148601 : _GEN_144760; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_152827 = 4'h8 < realFlowNum_1 ? _GEN_148602 : _GEN_144761; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_152828 = 4'h8 < realFlowNum_1 ? _GEN_148603 : _GEN_144762; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_152829 = 4'h8 < realFlowNum_1 ? _GEN_148604 : _GEN_144763; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_152830 = 4'h8 < realFlowNum_1 ? _GEN_148605 : _GEN_144764; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_152831 = 4'h8 < realFlowNum_1 ? _GEN_148606 : _GEN_144765; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_152832 = 4'h8 < realFlowNum_1 ? _GEN_148607 : _GEN_144766; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_152833 = 4'h8 < realFlowNum_1 ? _GEN_148608 : _GEN_144767; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_152834 = 4'h8 < realFlowNum_1 ? _GEN_148609 : _GEN_144768; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_152835 = 4'h8 < realFlowNum_1 ? _GEN_148610 : _GEN_144769; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_152836 = 4'h8 < realFlowNum_1 ? _GEN_148611 : _GEN_144770; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_152837 = 4'h8 < realFlowNum_1 ? _GEN_148612 : _GEN_144771; // @[Vlflowqueue.scala 194:37]
  wire  _GEN_156649 = needAlloc_1 ? _GEN_152806 : flow_entry_valid_1_0; // @[Vlflowqueue.scala 191:25 135:33]
  wire  _GEN_156650 = needAlloc_1 ? _GEN_152807 : flow_entry_valid_1_1; // @[Vlflowqueue.scala 191:25 135:33]
  wire  _GEN_156651 = needAlloc_1 ? _GEN_152808 : flow_entry_valid_1_2; // @[Vlflowqueue.scala 191:25 135:33]
  wire  _GEN_156652 = needAlloc_1 ? _GEN_152809 : flow_entry_valid_1_3; // @[Vlflowqueue.scala 191:25 135:33]
  wire  _GEN_156653 = needAlloc_1 ? _GEN_152810 : flow_entry_valid_1_4; // @[Vlflowqueue.scala 191:25 135:33]
  wire  _GEN_156654 = needAlloc_1 ? _GEN_152811 : flow_entry_valid_1_5; // @[Vlflowqueue.scala 191:25 135:33]
  wire  _GEN_156655 = needAlloc_1 ? _GEN_152812 : flow_entry_valid_1_6; // @[Vlflowqueue.scala 191:25 135:33]
  wire  _GEN_156656 = needAlloc_1 ? _GEN_152813 : flow_entry_valid_1_7; // @[Vlflowqueue.scala 191:25 135:33]
  wire  _GEN_156657 = needAlloc_1 ? _GEN_152814 : flow_entry_valid_1_8; // @[Vlflowqueue.scala 191:25 135:33]
  wire  _GEN_156658 = needAlloc_1 ? _GEN_152815 : flow_entry_valid_1_9; // @[Vlflowqueue.scala 191:25 135:33]
  wire  _GEN_156659 = needAlloc_1 ? _GEN_152816 : flow_entry_valid_1_10; // @[Vlflowqueue.scala 191:25 135:33]
  wire  _GEN_156660 = needAlloc_1 ? _GEN_152817 : flow_entry_valid_1_11; // @[Vlflowqueue.scala 191:25 135:33]
  wire  _GEN_156661 = needAlloc_1 ? _GEN_152818 : flow_entry_valid_1_12; // @[Vlflowqueue.scala 191:25 135:33]
  wire  _GEN_156662 = needAlloc_1 ? _GEN_152819 : flow_entry_valid_1_13; // @[Vlflowqueue.scala 191:25 135:33]
  wire  _GEN_156663 = needAlloc_1 ? _GEN_152820 : flow_entry_valid_1_14; // @[Vlflowqueue.scala 191:25 135:33]
  wire  _GEN_156664 = needAlloc_1 ? _GEN_152821 : flow_entry_valid_1_15; // @[Vlflowqueue.scala 191:25 135:33]
  wire  _GEN_156665 = needAlloc_1 ? _GEN_152822 : flow_entry_valid_1_16; // @[Vlflowqueue.scala 191:25 135:33]
  wire  _GEN_156666 = needAlloc_1 ? _GEN_152823 : flow_entry_valid_1_17; // @[Vlflowqueue.scala 191:25 135:33]
  wire  _GEN_156667 = needAlloc_1 ? _GEN_152824 : flow_entry_valid_1_18; // @[Vlflowqueue.scala 191:25 135:33]
  wire  _GEN_156668 = needAlloc_1 ? _GEN_152825 : flow_entry_valid_1_19; // @[Vlflowqueue.scala 191:25 135:33]
  wire  _GEN_156669 = needAlloc_1 ? _GEN_152826 : flow_entry_valid_1_20; // @[Vlflowqueue.scala 191:25 135:33]
  wire  _GEN_156670 = needAlloc_1 ? _GEN_152827 : flow_entry_valid_1_21; // @[Vlflowqueue.scala 191:25 135:33]
  wire  _GEN_156671 = needAlloc_1 ? _GEN_152828 : flow_entry_valid_1_22; // @[Vlflowqueue.scala 191:25 135:33]
  wire  _GEN_156672 = needAlloc_1 ? _GEN_152829 : flow_entry_valid_1_23; // @[Vlflowqueue.scala 191:25 135:33]
  wire  _GEN_156673 = needAlloc_1 ? _GEN_152830 : flow_entry_valid_1_24; // @[Vlflowqueue.scala 191:25 135:33]
  wire  _GEN_156674 = needAlloc_1 ? _GEN_152831 : flow_entry_valid_1_25; // @[Vlflowqueue.scala 191:25 135:33]
  wire  _GEN_156675 = needAlloc_1 ? _GEN_152832 : flow_entry_valid_1_26; // @[Vlflowqueue.scala 191:25 135:33]
  wire  _GEN_156676 = needAlloc_1 ? _GEN_152833 : flow_entry_valid_1_27; // @[Vlflowqueue.scala 191:25 135:33]
  wire  _GEN_156677 = needAlloc_1 ? _GEN_152834 : flow_entry_valid_1_28; // @[Vlflowqueue.scala 191:25 135:33]
  wire  _GEN_156678 = needAlloc_1 ? _GEN_152835 : flow_entry_valid_1_29; // @[Vlflowqueue.scala 191:25 135:33]
  wire  _GEN_156679 = needAlloc_1 ? _GEN_152836 : flow_entry_valid_1_30; // @[Vlflowqueue.scala 191:25 135:33]
  wire  _GEN_156680 = needAlloc_1 ? _GEN_152837 : flow_entry_valid_1_31; // @[Vlflowqueue.scala 191:25 135:33]
  wire  _GEN_160491 = 5'h1 == deqPtr_0_value ? flow_entry_valid_0_1 : flow_entry_valid_0_0; // @[Vlflowqueue.scala 236:{48,48}]
  wire  _GEN_160492 = 5'h2 == deqPtr_0_value ? flow_entry_valid_0_2 : _GEN_160491; // @[Vlflowqueue.scala 236:{48,48}]
  wire  _GEN_160493 = 5'h3 == deqPtr_0_value ? flow_entry_valid_0_3 : _GEN_160492; // @[Vlflowqueue.scala 236:{48,48}]
  wire  _GEN_160494 = 5'h4 == deqPtr_0_value ? flow_entry_valid_0_4 : _GEN_160493; // @[Vlflowqueue.scala 236:{48,48}]
  wire  _GEN_160495 = 5'h5 == deqPtr_0_value ? flow_entry_valid_0_5 : _GEN_160494; // @[Vlflowqueue.scala 236:{48,48}]
  wire  _GEN_160496 = 5'h6 == deqPtr_0_value ? flow_entry_valid_0_6 : _GEN_160495; // @[Vlflowqueue.scala 236:{48,48}]
  wire  _GEN_160497 = 5'h7 == deqPtr_0_value ? flow_entry_valid_0_7 : _GEN_160496; // @[Vlflowqueue.scala 236:{48,48}]
  wire  _GEN_160498 = 5'h8 == deqPtr_0_value ? flow_entry_valid_0_8 : _GEN_160497; // @[Vlflowqueue.scala 236:{48,48}]
  wire  _GEN_160499 = 5'h9 == deqPtr_0_value ? flow_entry_valid_0_9 : _GEN_160498; // @[Vlflowqueue.scala 236:{48,48}]
  wire  _GEN_160500 = 5'ha == deqPtr_0_value ? flow_entry_valid_0_10 : _GEN_160499; // @[Vlflowqueue.scala 236:{48,48}]
  wire  _GEN_160501 = 5'hb == deqPtr_0_value ? flow_entry_valid_0_11 : _GEN_160500; // @[Vlflowqueue.scala 236:{48,48}]
  wire  _GEN_160502 = 5'hc == deqPtr_0_value ? flow_entry_valid_0_12 : _GEN_160501; // @[Vlflowqueue.scala 236:{48,48}]
  wire  _GEN_160503 = 5'hd == deqPtr_0_value ? flow_entry_valid_0_13 : _GEN_160502; // @[Vlflowqueue.scala 236:{48,48}]
  wire  _GEN_160504 = 5'he == deqPtr_0_value ? flow_entry_valid_0_14 : _GEN_160503; // @[Vlflowqueue.scala 236:{48,48}]
  wire  _GEN_160505 = 5'hf == deqPtr_0_value ? flow_entry_valid_0_15 : _GEN_160504; // @[Vlflowqueue.scala 236:{48,48}]
  wire  _GEN_160506 = 5'h10 == deqPtr_0_value ? flow_entry_valid_0_16 : _GEN_160505; // @[Vlflowqueue.scala 236:{48,48}]
  wire  _GEN_160507 = 5'h11 == deqPtr_0_value ? flow_entry_valid_0_17 : _GEN_160506; // @[Vlflowqueue.scala 236:{48,48}]
  wire  _GEN_160508 = 5'h12 == deqPtr_0_value ? flow_entry_valid_0_18 : _GEN_160507; // @[Vlflowqueue.scala 236:{48,48}]
  wire  _GEN_160509 = 5'h13 == deqPtr_0_value ? flow_entry_valid_0_19 : _GEN_160508; // @[Vlflowqueue.scala 236:{48,48}]
  wire  _GEN_160510 = 5'h14 == deqPtr_0_value ? flow_entry_valid_0_20 : _GEN_160509; // @[Vlflowqueue.scala 236:{48,48}]
  wire  _GEN_160511 = 5'h15 == deqPtr_0_value ? flow_entry_valid_0_21 : _GEN_160510; // @[Vlflowqueue.scala 236:{48,48}]
  wire  _GEN_160512 = 5'h16 == deqPtr_0_value ? flow_entry_valid_0_22 : _GEN_160511; // @[Vlflowqueue.scala 236:{48,48}]
  wire  _GEN_160513 = 5'h17 == deqPtr_0_value ? flow_entry_valid_0_23 : _GEN_160512; // @[Vlflowqueue.scala 236:{48,48}]
  wire  _GEN_160514 = 5'h18 == deqPtr_0_value ? flow_entry_valid_0_24 : _GEN_160513; // @[Vlflowqueue.scala 236:{48,48}]
  wire  _GEN_160515 = 5'h19 == deqPtr_0_value ? flow_entry_valid_0_25 : _GEN_160514; // @[Vlflowqueue.scala 236:{48,48}]
  wire  _GEN_160516 = 5'h1a == deqPtr_0_value ? flow_entry_valid_0_26 : _GEN_160515; // @[Vlflowqueue.scala 236:{48,48}]
  wire  _GEN_160517 = 5'h1b == deqPtr_0_value ? flow_entry_valid_0_27 : _GEN_160516; // @[Vlflowqueue.scala 236:{48,48}]
  wire  _GEN_160518 = 5'h1c == deqPtr_0_value ? flow_entry_valid_0_28 : _GEN_160517; // @[Vlflowqueue.scala 236:{48,48}]
  wire  _GEN_160519 = 5'h1d == deqPtr_0_value ? flow_entry_valid_0_29 : _GEN_160518; // @[Vlflowqueue.scala 236:{48,48}]
  wire  _GEN_160520 = 5'h1e == deqPtr_0_value ? flow_entry_valid_0_30 : _GEN_160519; // @[Vlflowqueue.scala 236:{48,48}]
  wire [38:0] _GEN_160555 = 5'h1 == deqPtr_0_value ? flow_entry_0_1_vaddr : flow_entry_0_0_vaddr; // @[Vlflowqueue.scala 239:{50,50}]
  wire [38:0] _GEN_160556 = 5'h2 == deqPtr_0_value ? flow_entry_0_2_vaddr : _GEN_160555; // @[Vlflowqueue.scala 239:{50,50}]
  wire [38:0] _GEN_160557 = 5'h3 == deqPtr_0_value ? flow_entry_0_3_vaddr : _GEN_160556; // @[Vlflowqueue.scala 239:{50,50}]
  wire [38:0] _GEN_160558 = 5'h4 == deqPtr_0_value ? flow_entry_0_4_vaddr : _GEN_160557; // @[Vlflowqueue.scala 239:{50,50}]
  wire [38:0] _GEN_160559 = 5'h5 == deqPtr_0_value ? flow_entry_0_5_vaddr : _GEN_160558; // @[Vlflowqueue.scala 239:{50,50}]
  wire [38:0] _GEN_160560 = 5'h6 == deqPtr_0_value ? flow_entry_0_6_vaddr : _GEN_160559; // @[Vlflowqueue.scala 239:{50,50}]
  wire [38:0] _GEN_160561 = 5'h7 == deqPtr_0_value ? flow_entry_0_7_vaddr : _GEN_160560; // @[Vlflowqueue.scala 239:{50,50}]
  wire [38:0] _GEN_160562 = 5'h8 == deqPtr_0_value ? flow_entry_0_8_vaddr : _GEN_160561; // @[Vlflowqueue.scala 239:{50,50}]
  wire [38:0] _GEN_160563 = 5'h9 == deqPtr_0_value ? flow_entry_0_9_vaddr : _GEN_160562; // @[Vlflowqueue.scala 239:{50,50}]
  wire [38:0] _GEN_160564 = 5'ha == deqPtr_0_value ? flow_entry_0_10_vaddr : _GEN_160563; // @[Vlflowqueue.scala 239:{50,50}]
  wire [38:0] _GEN_160565 = 5'hb == deqPtr_0_value ? flow_entry_0_11_vaddr : _GEN_160564; // @[Vlflowqueue.scala 239:{50,50}]
  wire [38:0] _GEN_160566 = 5'hc == deqPtr_0_value ? flow_entry_0_12_vaddr : _GEN_160565; // @[Vlflowqueue.scala 239:{50,50}]
  wire [38:0] _GEN_160567 = 5'hd == deqPtr_0_value ? flow_entry_0_13_vaddr : _GEN_160566; // @[Vlflowqueue.scala 239:{50,50}]
  wire [38:0] _GEN_160568 = 5'he == deqPtr_0_value ? flow_entry_0_14_vaddr : _GEN_160567; // @[Vlflowqueue.scala 239:{50,50}]
  wire [38:0] _GEN_160569 = 5'hf == deqPtr_0_value ? flow_entry_0_15_vaddr : _GEN_160568; // @[Vlflowqueue.scala 239:{50,50}]
  wire [38:0] _GEN_160570 = 5'h10 == deqPtr_0_value ? flow_entry_0_16_vaddr : _GEN_160569; // @[Vlflowqueue.scala 239:{50,50}]
  wire [38:0] _GEN_160571 = 5'h11 == deqPtr_0_value ? flow_entry_0_17_vaddr : _GEN_160570; // @[Vlflowqueue.scala 239:{50,50}]
  wire [38:0] _GEN_160572 = 5'h12 == deqPtr_0_value ? flow_entry_0_18_vaddr : _GEN_160571; // @[Vlflowqueue.scala 239:{50,50}]
  wire [38:0] _GEN_160573 = 5'h13 == deqPtr_0_value ? flow_entry_0_19_vaddr : _GEN_160572; // @[Vlflowqueue.scala 239:{50,50}]
  wire [38:0] _GEN_160574 = 5'h14 == deqPtr_0_value ? flow_entry_0_20_vaddr : _GEN_160573; // @[Vlflowqueue.scala 239:{50,50}]
  wire [38:0] _GEN_160575 = 5'h15 == deqPtr_0_value ? flow_entry_0_21_vaddr : _GEN_160574; // @[Vlflowqueue.scala 239:{50,50}]
  wire [38:0] _GEN_160576 = 5'h16 == deqPtr_0_value ? flow_entry_0_22_vaddr : _GEN_160575; // @[Vlflowqueue.scala 239:{50,50}]
  wire [38:0] _GEN_160577 = 5'h17 == deqPtr_0_value ? flow_entry_0_23_vaddr : _GEN_160576; // @[Vlflowqueue.scala 239:{50,50}]
  wire [38:0] _GEN_160578 = 5'h18 == deqPtr_0_value ? flow_entry_0_24_vaddr : _GEN_160577; // @[Vlflowqueue.scala 239:{50,50}]
  wire [38:0] _GEN_160579 = 5'h19 == deqPtr_0_value ? flow_entry_0_25_vaddr : _GEN_160578; // @[Vlflowqueue.scala 239:{50,50}]
  wire [38:0] _GEN_160580 = 5'h1a == deqPtr_0_value ? flow_entry_0_26_vaddr : _GEN_160579; // @[Vlflowqueue.scala 239:{50,50}]
  wire [38:0] _GEN_160581 = 5'h1b == deqPtr_0_value ? flow_entry_0_27_vaddr : _GEN_160580; // @[Vlflowqueue.scala 239:{50,50}]
  wire [38:0] _GEN_160582 = 5'h1c == deqPtr_0_value ? flow_entry_0_28_vaddr : _GEN_160581; // @[Vlflowqueue.scala 239:{50,50}]
  wire [38:0] _GEN_160583 = 5'h1d == deqPtr_0_value ? flow_entry_0_29_vaddr : _GEN_160582; // @[Vlflowqueue.scala 239:{50,50}]
  wire [38:0] _GEN_160584 = 5'h1e == deqPtr_0_value ? flow_entry_0_30_vaddr : _GEN_160583; // @[Vlflowqueue.scala 239:{50,50}]
  wire  _GEN_160887 = 5'h1 == deqPtr_1_value ? flow_entry_valid_1_1 : flow_entry_valid_1_0; // @[Vlflowqueue.scala 236:{48,48}]
  wire  _GEN_160888 = 5'h2 == deqPtr_1_value ? flow_entry_valid_1_2 : _GEN_160887; // @[Vlflowqueue.scala 236:{48,48}]
  wire  _GEN_160889 = 5'h3 == deqPtr_1_value ? flow_entry_valid_1_3 : _GEN_160888; // @[Vlflowqueue.scala 236:{48,48}]
  wire  _GEN_160890 = 5'h4 == deqPtr_1_value ? flow_entry_valid_1_4 : _GEN_160889; // @[Vlflowqueue.scala 236:{48,48}]
  wire  _GEN_160891 = 5'h5 == deqPtr_1_value ? flow_entry_valid_1_5 : _GEN_160890; // @[Vlflowqueue.scala 236:{48,48}]
  wire  _GEN_160892 = 5'h6 == deqPtr_1_value ? flow_entry_valid_1_6 : _GEN_160891; // @[Vlflowqueue.scala 236:{48,48}]
  wire  _GEN_160893 = 5'h7 == deqPtr_1_value ? flow_entry_valid_1_7 : _GEN_160892; // @[Vlflowqueue.scala 236:{48,48}]
  wire  _GEN_160894 = 5'h8 == deqPtr_1_value ? flow_entry_valid_1_8 : _GEN_160893; // @[Vlflowqueue.scala 236:{48,48}]
  wire  _GEN_160895 = 5'h9 == deqPtr_1_value ? flow_entry_valid_1_9 : _GEN_160894; // @[Vlflowqueue.scala 236:{48,48}]
  wire  _GEN_160896 = 5'ha == deqPtr_1_value ? flow_entry_valid_1_10 : _GEN_160895; // @[Vlflowqueue.scala 236:{48,48}]
  wire  _GEN_160897 = 5'hb == deqPtr_1_value ? flow_entry_valid_1_11 : _GEN_160896; // @[Vlflowqueue.scala 236:{48,48}]
  wire  _GEN_160898 = 5'hc == deqPtr_1_value ? flow_entry_valid_1_12 : _GEN_160897; // @[Vlflowqueue.scala 236:{48,48}]
  wire  _GEN_160899 = 5'hd == deqPtr_1_value ? flow_entry_valid_1_13 : _GEN_160898; // @[Vlflowqueue.scala 236:{48,48}]
  wire  _GEN_160900 = 5'he == deqPtr_1_value ? flow_entry_valid_1_14 : _GEN_160899; // @[Vlflowqueue.scala 236:{48,48}]
  wire  _GEN_160901 = 5'hf == deqPtr_1_value ? flow_entry_valid_1_15 : _GEN_160900; // @[Vlflowqueue.scala 236:{48,48}]
  wire  _GEN_160902 = 5'h10 == deqPtr_1_value ? flow_entry_valid_1_16 : _GEN_160901; // @[Vlflowqueue.scala 236:{48,48}]
  wire  _GEN_160903 = 5'h11 == deqPtr_1_value ? flow_entry_valid_1_17 : _GEN_160902; // @[Vlflowqueue.scala 236:{48,48}]
  wire  _GEN_160904 = 5'h12 == deqPtr_1_value ? flow_entry_valid_1_18 : _GEN_160903; // @[Vlflowqueue.scala 236:{48,48}]
  wire  _GEN_160905 = 5'h13 == deqPtr_1_value ? flow_entry_valid_1_19 : _GEN_160904; // @[Vlflowqueue.scala 236:{48,48}]
  wire  _GEN_160906 = 5'h14 == deqPtr_1_value ? flow_entry_valid_1_20 : _GEN_160905; // @[Vlflowqueue.scala 236:{48,48}]
  wire  _GEN_160907 = 5'h15 == deqPtr_1_value ? flow_entry_valid_1_21 : _GEN_160906; // @[Vlflowqueue.scala 236:{48,48}]
  wire  _GEN_160908 = 5'h16 == deqPtr_1_value ? flow_entry_valid_1_22 : _GEN_160907; // @[Vlflowqueue.scala 236:{48,48}]
  wire  _GEN_160909 = 5'h17 == deqPtr_1_value ? flow_entry_valid_1_23 : _GEN_160908; // @[Vlflowqueue.scala 236:{48,48}]
  wire  _GEN_160910 = 5'h18 == deqPtr_1_value ? flow_entry_valid_1_24 : _GEN_160909; // @[Vlflowqueue.scala 236:{48,48}]
  wire  _GEN_160911 = 5'h19 == deqPtr_1_value ? flow_entry_valid_1_25 : _GEN_160910; // @[Vlflowqueue.scala 236:{48,48}]
  wire  _GEN_160912 = 5'h1a == deqPtr_1_value ? flow_entry_valid_1_26 : _GEN_160911; // @[Vlflowqueue.scala 236:{48,48}]
  wire  _GEN_160913 = 5'h1b == deqPtr_1_value ? flow_entry_valid_1_27 : _GEN_160912; // @[Vlflowqueue.scala 236:{48,48}]
  wire  _GEN_160914 = 5'h1c == deqPtr_1_value ? flow_entry_valid_1_28 : _GEN_160913; // @[Vlflowqueue.scala 236:{48,48}]
  wire  _GEN_160915 = 5'h1d == deqPtr_1_value ? flow_entry_valid_1_29 : _GEN_160914; // @[Vlflowqueue.scala 236:{48,48}]
  wire  _GEN_160916 = 5'h1e == deqPtr_1_value ? flow_entry_valid_1_30 : _GEN_160915; // @[Vlflowqueue.scala 236:{48,48}]
  wire [38:0] _GEN_160951 = 5'h1 == deqPtr_1_value ? flow_entry_1_1_vaddr : flow_entry_1_0_vaddr; // @[Vlflowqueue.scala 239:{50,50}]
  wire [38:0] _GEN_160952 = 5'h2 == deqPtr_1_value ? flow_entry_1_2_vaddr : _GEN_160951; // @[Vlflowqueue.scala 239:{50,50}]
  wire [38:0] _GEN_160953 = 5'h3 == deqPtr_1_value ? flow_entry_1_3_vaddr : _GEN_160952; // @[Vlflowqueue.scala 239:{50,50}]
  wire [38:0] _GEN_160954 = 5'h4 == deqPtr_1_value ? flow_entry_1_4_vaddr : _GEN_160953; // @[Vlflowqueue.scala 239:{50,50}]
  wire [38:0] _GEN_160955 = 5'h5 == deqPtr_1_value ? flow_entry_1_5_vaddr : _GEN_160954; // @[Vlflowqueue.scala 239:{50,50}]
  wire [38:0] _GEN_160956 = 5'h6 == deqPtr_1_value ? flow_entry_1_6_vaddr : _GEN_160955; // @[Vlflowqueue.scala 239:{50,50}]
  wire [38:0] _GEN_160957 = 5'h7 == deqPtr_1_value ? flow_entry_1_7_vaddr : _GEN_160956; // @[Vlflowqueue.scala 239:{50,50}]
  wire [38:0] _GEN_160958 = 5'h8 == deqPtr_1_value ? flow_entry_1_8_vaddr : _GEN_160957; // @[Vlflowqueue.scala 239:{50,50}]
  wire [38:0] _GEN_160959 = 5'h9 == deqPtr_1_value ? flow_entry_1_9_vaddr : _GEN_160958; // @[Vlflowqueue.scala 239:{50,50}]
  wire [38:0] _GEN_160960 = 5'ha == deqPtr_1_value ? flow_entry_1_10_vaddr : _GEN_160959; // @[Vlflowqueue.scala 239:{50,50}]
  wire [38:0] _GEN_160961 = 5'hb == deqPtr_1_value ? flow_entry_1_11_vaddr : _GEN_160960; // @[Vlflowqueue.scala 239:{50,50}]
  wire [38:0] _GEN_160962 = 5'hc == deqPtr_1_value ? flow_entry_1_12_vaddr : _GEN_160961; // @[Vlflowqueue.scala 239:{50,50}]
  wire [38:0] _GEN_160963 = 5'hd == deqPtr_1_value ? flow_entry_1_13_vaddr : _GEN_160962; // @[Vlflowqueue.scala 239:{50,50}]
  wire [38:0] _GEN_160964 = 5'he == deqPtr_1_value ? flow_entry_1_14_vaddr : _GEN_160963; // @[Vlflowqueue.scala 239:{50,50}]
  wire [38:0] _GEN_160965 = 5'hf == deqPtr_1_value ? flow_entry_1_15_vaddr : _GEN_160964; // @[Vlflowqueue.scala 239:{50,50}]
  wire [38:0] _GEN_160966 = 5'h10 == deqPtr_1_value ? flow_entry_1_16_vaddr : _GEN_160965; // @[Vlflowqueue.scala 239:{50,50}]
  wire [38:0] _GEN_160967 = 5'h11 == deqPtr_1_value ? flow_entry_1_17_vaddr : _GEN_160966; // @[Vlflowqueue.scala 239:{50,50}]
  wire [38:0] _GEN_160968 = 5'h12 == deqPtr_1_value ? flow_entry_1_18_vaddr : _GEN_160967; // @[Vlflowqueue.scala 239:{50,50}]
  wire [38:0] _GEN_160969 = 5'h13 == deqPtr_1_value ? flow_entry_1_19_vaddr : _GEN_160968; // @[Vlflowqueue.scala 239:{50,50}]
  wire [38:0] _GEN_160970 = 5'h14 == deqPtr_1_value ? flow_entry_1_20_vaddr : _GEN_160969; // @[Vlflowqueue.scala 239:{50,50}]
  wire [38:0] _GEN_160971 = 5'h15 == deqPtr_1_value ? flow_entry_1_21_vaddr : _GEN_160970; // @[Vlflowqueue.scala 239:{50,50}]
  wire [38:0] _GEN_160972 = 5'h16 == deqPtr_1_value ? flow_entry_1_22_vaddr : _GEN_160971; // @[Vlflowqueue.scala 239:{50,50}]
  wire [38:0] _GEN_160973 = 5'h17 == deqPtr_1_value ? flow_entry_1_23_vaddr : _GEN_160972; // @[Vlflowqueue.scala 239:{50,50}]
  wire [38:0] _GEN_160974 = 5'h18 == deqPtr_1_value ? flow_entry_1_24_vaddr : _GEN_160973; // @[Vlflowqueue.scala 239:{50,50}]
  wire [38:0] _GEN_160975 = 5'h19 == deqPtr_1_value ? flow_entry_1_25_vaddr : _GEN_160974; // @[Vlflowqueue.scala 239:{50,50}]
  wire [38:0] _GEN_160976 = 5'h1a == deqPtr_1_value ? flow_entry_1_26_vaddr : _GEN_160975; // @[Vlflowqueue.scala 239:{50,50}]
  wire [38:0] _GEN_160977 = 5'h1b == deqPtr_1_value ? flow_entry_1_27_vaddr : _GEN_160976; // @[Vlflowqueue.scala 239:{50,50}]
  wire [38:0] _GEN_160978 = 5'h1c == deqPtr_1_value ? flow_entry_1_28_vaddr : _GEN_160977; // @[Vlflowqueue.scala 239:{50,50}]
  wire [38:0] _GEN_160979 = 5'h1d == deqPtr_1_value ? flow_entry_1_29_vaddr : _GEN_160978; // @[Vlflowqueue.scala 239:{50,50}]
  wire [38:0] _GEN_160980 = 5'h1e == deqPtr_1_value ? flow_entry_1_30_vaddr : _GEN_160979; // @[Vlflowqueue.scala 239:{50,50}]
  wire  _T_90 = io_loadPipeOut_0_ready & io_loadPipeOut_0_valid; // @[Decoupled.scala 50:35]
  wire [5:0] _deqPtr_0_new_ptr_T = {deqPtr_0_flag,deqPtr_0_value}; // @[Cat.scala 31:58]
  wire [5:0] _deqPtr_0_new_ptr_T_2 = _deqPtr_0_new_ptr_T + 6'h1; // @[CircularQueuePtr.scala 39:46]
  wire [4:0] deqPtr_0_new_ptr_value = _deqPtr_0_new_ptr_T_2[4:0]; // @[CircularQueuePtr.scala 39:59]
  wire  deqPtr_0_new_ptr_flag = _deqPtr_0_new_ptr_T_2[5]; // @[CircularQueuePtr.scala 39:59]
  wire  _T_91 = io_loadPipeOut_1_ready & io_loadPipeOut_1_valid; // @[Decoupled.scala 50:35]
  wire [5:0] _deqPtr_1_new_ptr_T = {deqPtr_1_flag,deqPtr_1_value}; // @[Cat.scala 31:58]
  wire [5:0] _deqPtr_1_new_ptr_T_2 = _deqPtr_1_new_ptr_T + 6'h1; // @[CircularQueuePtr.scala 39:46]
  wire [4:0] deqPtr_1_new_ptr_value = _deqPtr_1_new_ptr_T_2[4:0]; // @[CircularQueuePtr.scala 39:59]
  wire  deqPtr_1_new_ptr_flag = _deqPtr_1_new_ptr_T_2[5]; // @[CircularQueuePtr.scala 39:59]
  assign io_loadPipeOut_0_valid = 5'h1f == deqPtr_0_value ? flow_entry_valid_0_31 : _GEN_160520; // @[Vlflowqueue.scala 236:{48,48}]
  assign io_loadPipeOut_0_bits_vaddr = 5'h1f == deqPtr_0_value ? flow_entry_0_31_vaddr : _GEN_160584; // @[Vlflowqueue.scala 239:{50,50}]
  assign io_loadPipeOut_1_valid = 5'h1f == deqPtr_1_value ? flow_entry_valid_1_31 : _GEN_160916; // @[Vlflowqueue.scala 236:{48,48}]
  assign io_loadPipeOut_1_bits_vaddr = 5'h1f == deqPtr_1_value ? flow_entry_1_31_vaddr : _GEN_160980; // @[Vlflowqueue.scala 239:{50,50}]
  always @(posedge clock) begin
    if (needAlloc_0) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
        if (5'h0 == index_0) begin // @[Vlflowqueue.scala 198:51]
          flow_entry_0_0_uop_robIdx_value <= io_loadRegIn_0_bits_uop_robIdx_value; // @[Vlflowqueue.scala 198:51]
        end else begin
          flow_entry_0_0_uop_robIdx_value <= _GEN_67471;
        end
      end else begin
        flow_entry_0_0_uop_robIdx_value <= _GEN_67471;
      end
    end
    if (needAlloc_0) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
        if (5'h0 == index_0) begin // @[Vlflowqueue.scala 203:51]
          if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
            flow_entry_0_0_vaddr <= _vaddr_0_T_162; // @[Vlflowqueue.scala 201:51]
          end else begin
            flow_entry_0_0_vaddr <= _GEN_68015;
          end
        end else begin
          flow_entry_0_0_vaddr <= _GEN_68048;
        end
      end else begin
        flow_entry_0_0_vaddr <= _GEN_68048;
      end
    end
    if (needAlloc_0) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
        if (5'h1 == index_0) begin // @[Vlflowqueue.scala 198:51]
          flow_entry_0_1_uop_robIdx_value <= io_loadRegIn_0_bits_uop_robIdx_value; // @[Vlflowqueue.scala 198:51]
        end else begin
          flow_entry_0_1_uop_robIdx_value <= _GEN_67472;
        end
      end else begin
        flow_entry_0_1_uop_robIdx_value <= _GEN_67472;
      end
    end
    if (needAlloc_0) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
        if (5'h1 == index_0) begin // @[Vlflowqueue.scala 203:51]
          if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
            flow_entry_0_1_vaddr <= _vaddr_0_T_162; // @[Vlflowqueue.scala 201:51]
          end else begin
            flow_entry_0_1_vaddr <= _GEN_68015;
          end
        end else begin
          flow_entry_0_1_vaddr <= _GEN_68049;
        end
      end else begin
        flow_entry_0_1_vaddr <= _GEN_68049;
      end
    end
    if (needAlloc_0) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
        if (5'h2 == index_0) begin // @[Vlflowqueue.scala 198:51]
          flow_entry_0_2_uop_robIdx_value <= io_loadRegIn_0_bits_uop_robIdx_value; // @[Vlflowqueue.scala 198:51]
        end else begin
          flow_entry_0_2_uop_robIdx_value <= _GEN_67473;
        end
      end else begin
        flow_entry_0_2_uop_robIdx_value <= _GEN_67473;
      end
    end
    if (needAlloc_0) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
        if (5'h2 == index_0) begin // @[Vlflowqueue.scala 203:51]
          if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
            flow_entry_0_2_vaddr <= _vaddr_0_T_162; // @[Vlflowqueue.scala 201:51]
          end else begin
            flow_entry_0_2_vaddr <= _GEN_68015;
          end
        end else begin
          flow_entry_0_2_vaddr <= _GEN_68050;
        end
      end else begin
        flow_entry_0_2_vaddr <= _GEN_68050;
      end
    end
    if (needAlloc_0) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
        if (5'h3 == index_0) begin // @[Vlflowqueue.scala 198:51]
          flow_entry_0_3_uop_robIdx_value <= io_loadRegIn_0_bits_uop_robIdx_value; // @[Vlflowqueue.scala 198:51]
        end else begin
          flow_entry_0_3_uop_robIdx_value <= _GEN_67474;
        end
      end else begin
        flow_entry_0_3_uop_robIdx_value <= _GEN_67474;
      end
    end
    if (needAlloc_0) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
        if (5'h3 == index_0) begin // @[Vlflowqueue.scala 203:51]
          if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
            flow_entry_0_3_vaddr <= _vaddr_0_T_162; // @[Vlflowqueue.scala 201:51]
          end else begin
            flow_entry_0_3_vaddr <= _GEN_68015;
          end
        end else begin
          flow_entry_0_3_vaddr <= _GEN_68051;
        end
      end else begin
        flow_entry_0_3_vaddr <= _GEN_68051;
      end
    end
    if (needAlloc_0) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
        if (5'h4 == index_0) begin // @[Vlflowqueue.scala 198:51]
          flow_entry_0_4_uop_robIdx_value <= io_loadRegIn_0_bits_uop_robIdx_value; // @[Vlflowqueue.scala 198:51]
        end else begin
          flow_entry_0_4_uop_robIdx_value <= _GEN_67475;
        end
      end else begin
        flow_entry_0_4_uop_robIdx_value <= _GEN_67475;
      end
    end
    if (needAlloc_0) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
        if (5'h4 == index_0) begin // @[Vlflowqueue.scala 203:51]
          if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
            flow_entry_0_4_vaddr <= _vaddr_0_T_162; // @[Vlflowqueue.scala 201:51]
          end else begin
            flow_entry_0_4_vaddr <= _GEN_68015;
          end
        end else begin
          flow_entry_0_4_vaddr <= _GEN_68052;
        end
      end else begin
        flow_entry_0_4_vaddr <= _GEN_68052;
      end
    end
    if (needAlloc_0) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
        if (5'h5 == index_0) begin // @[Vlflowqueue.scala 198:51]
          flow_entry_0_5_uop_robIdx_value <= io_loadRegIn_0_bits_uop_robIdx_value; // @[Vlflowqueue.scala 198:51]
        end else begin
          flow_entry_0_5_uop_robIdx_value <= _GEN_67476;
        end
      end else begin
        flow_entry_0_5_uop_robIdx_value <= _GEN_67476;
      end
    end
    if (needAlloc_0) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
        if (5'h5 == index_0) begin // @[Vlflowqueue.scala 203:51]
          if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
            flow_entry_0_5_vaddr <= _vaddr_0_T_162; // @[Vlflowqueue.scala 201:51]
          end else begin
            flow_entry_0_5_vaddr <= _GEN_68015;
          end
        end else begin
          flow_entry_0_5_vaddr <= _GEN_68053;
        end
      end else begin
        flow_entry_0_5_vaddr <= _GEN_68053;
      end
    end
    if (needAlloc_0) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
        if (5'h6 == index_0) begin // @[Vlflowqueue.scala 198:51]
          flow_entry_0_6_uop_robIdx_value <= io_loadRegIn_0_bits_uop_robIdx_value; // @[Vlflowqueue.scala 198:51]
        end else begin
          flow_entry_0_6_uop_robIdx_value <= _GEN_67477;
        end
      end else begin
        flow_entry_0_6_uop_robIdx_value <= _GEN_67477;
      end
    end
    if (needAlloc_0) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
        if (5'h6 == index_0) begin // @[Vlflowqueue.scala 203:51]
          if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
            flow_entry_0_6_vaddr <= _vaddr_0_T_162; // @[Vlflowqueue.scala 201:51]
          end else begin
            flow_entry_0_6_vaddr <= _GEN_68015;
          end
        end else begin
          flow_entry_0_6_vaddr <= _GEN_68054;
        end
      end else begin
        flow_entry_0_6_vaddr <= _GEN_68054;
      end
    end
    if (needAlloc_0) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
        if (5'h7 == index_0) begin // @[Vlflowqueue.scala 198:51]
          flow_entry_0_7_uop_robIdx_value <= io_loadRegIn_0_bits_uop_robIdx_value; // @[Vlflowqueue.scala 198:51]
        end else begin
          flow_entry_0_7_uop_robIdx_value <= _GEN_67478;
        end
      end else begin
        flow_entry_0_7_uop_robIdx_value <= _GEN_67478;
      end
    end
    if (needAlloc_0) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
        if (5'h7 == index_0) begin // @[Vlflowqueue.scala 203:51]
          if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
            flow_entry_0_7_vaddr <= _vaddr_0_T_162; // @[Vlflowqueue.scala 201:51]
          end else begin
            flow_entry_0_7_vaddr <= _GEN_68015;
          end
        end else begin
          flow_entry_0_7_vaddr <= _GEN_68055;
        end
      end else begin
        flow_entry_0_7_vaddr <= _GEN_68055;
      end
    end
    if (needAlloc_0) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
        if (5'h8 == index_0) begin // @[Vlflowqueue.scala 198:51]
          flow_entry_0_8_uop_robIdx_value <= io_loadRegIn_0_bits_uop_robIdx_value; // @[Vlflowqueue.scala 198:51]
        end else begin
          flow_entry_0_8_uop_robIdx_value <= _GEN_67479;
        end
      end else begin
        flow_entry_0_8_uop_robIdx_value <= _GEN_67479;
      end
    end
    if (needAlloc_0) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
        if (5'h8 == index_0) begin // @[Vlflowqueue.scala 203:51]
          if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
            flow_entry_0_8_vaddr <= _vaddr_0_T_162; // @[Vlflowqueue.scala 201:51]
          end else begin
            flow_entry_0_8_vaddr <= _GEN_68015;
          end
        end else begin
          flow_entry_0_8_vaddr <= _GEN_68056;
        end
      end else begin
        flow_entry_0_8_vaddr <= _GEN_68056;
      end
    end
    if (needAlloc_0) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
        if (5'h9 == index_0) begin // @[Vlflowqueue.scala 198:51]
          flow_entry_0_9_uop_robIdx_value <= io_loadRegIn_0_bits_uop_robIdx_value; // @[Vlflowqueue.scala 198:51]
        end else begin
          flow_entry_0_9_uop_robIdx_value <= _GEN_67480;
        end
      end else begin
        flow_entry_0_9_uop_robIdx_value <= _GEN_67480;
      end
    end
    if (needAlloc_0) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
        if (5'h9 == index_0) begin // @[Vlflowqueue.scala 203:51]
          if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
            flow_entry_0_9_vaddr <= _vaddr_0_T_162; // @[Vlflowqueue.scala 201:51]
          end else begin
            flow_entry_0_9_vaddr <= _GEN_68015;
          end
        end else begin
          flow_entry_0_9_vaddr <= _GEN_68057;
        end
      end else begin
        flow_entry_0_9_vaddr <= _GEN_68057;
      end
    end
    if (needAlloc_0) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
        if (5'ha == index_0) begin // @[Vlflowqueue.scala 198:51]
          flow_entry_0_10_uop_robIdx_value <= io_loadRegIn_0_bits_uop_robIdx_value; // @[Vlflowqueue.scala 198:51]
        end else begin
          flow_entry_0_10_uop_robIdx_value <= _GEN_67481;
        end
      end else begin
        flow_entry_0_10_uop_robIdx_value <= _GEN_67481;
      end
    end
    if (needAlloc_0) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
        if (5'ha == index_0) begin // @[Vlflowqueue.scala 203:51]
          if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
            flow_entry_0_10_vaddr <= _vaddr_0_T_162; // @[Vlflowqueue.scala 201:51]
          end else begin
            flow_entry_0_10_vaddr <= _GEN_68015;
          end
        end else begin
          flow_entry_0_10_vaddr <= _GEN_68058;
        end
      end else begin
        flow_entry_0_10_vaddr <= _GEN_68058;
      end
    end
    if (needAlloc_0) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
        if (5'hb == index_0) begin // @[Vlflowqueue.scala 198:51]
          flow_entry_0_11_uop_robIdx_value <= io_loadRegIn_0_bits_uop_robIdx_value; // @[Vlflowqueue.scala 198:51]
        end else begin
          flow_entry_0_11_uop_robIdx_value <= _GEN_67482;
        end
      end else begin
        flow_entry_0_11_uop_robIdx_value <= _GEN_67482;
      end
    end
    if (needAlloc_0) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
        if (5'hb == index_0) begin // @[Vlflowqueue.scala 203:51]
          if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
            flow_entry_0_11_vaddr <= _vaddr_0_T_162; // @[Vlflowqueue.scala 201:51]
          end else begin
            flow_entry_0_11_vaddr <= _GEN_68015;
          end
        end else begin
          flow_entry_0_11_vaddr <= _GEN_68059;
        end
      end else begin
        flow_entry_0_11_vaddr <= _GEN_68059;
      end
    end
    if (needAlloc_0) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
        if (5'hc == index_0) begin // @[Vlflowqueue.scala 198:51]
          flow_entry_0_12_uop_robIdx_value <= io_loadRegIn_0_bits_uop_robIdx_value; // @[Vlflowqueue.scala 198:51]
        end else begin
          flow_entry_0_12_uop_robIdx_value <= _GEN_67483;
        end
      end else begin
        flow_entry_0_12_uop_robIdx_value <= _GEN_67483;
      end
    end
    if (needAlloc_0) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
        if (5'hc == index_0) begin // @[Vlflowqueue.scala 203:51]
          if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
            flow_entry_0_12_vaddr <= _vaddr_0_T_162; // @[Vlflowqueue.scala 201:51]
          end else begin
            flow_entry_0_12_vaddr <= _GEN_68015;
          end
        end else begin
          flow_entry_0_12_vaddr <= _GEN_68060;
        end
      end else begin
        flow_entry_0_12_vaddr <= _GEN_68060;
      end
    end
    if (needAlloc_0) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
        if (5'hd == index_0) begin // @[Vlflowqueue.scala 198:51]
          flow_entry_0_13_uop_robIdx_value <= io_loadRegIn_0_bits_uop_robIdx_value; // @[Vlflowqueue.scala 198:51]
        end else begin
          flow_entry_0_13_uop_robIdx_value <= _GEN_67484;
        end
      end else begin
        flow_entry_0_13_uop_robIdx_value <= _GEN_67484;
      end
    end
    if (needAlloc_0) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
        if (5'hd == index_0) begin // @[Vlflowqueue.scala 203:51]
          if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
            flow_entry_0_13_vaddr <= _vaddr_0_T_162; // @[Vlflowqueue.scala 201:51]
          end else begin
            flow_entry_0_13_vaddr <= _GEN_68015;
          end
        end else begin
          flow_entry_0_13_vaddr <= _GEN_68061;
        end
      end else begin
        flow_entry_0_13_vaddr <= _GEN_68061;
      end
    end
    if (needAlloc_0) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
        if (5'he == index_0) begin // @[Vlflowqueue.scala 198:51]
          flow_entry_0_14_uop_robIdx_value <= io_loadRegIn_0_bits_uop_robIdx_value; // @[Vlflowqueue.scala 198:51]
        end else begin
          flow_entry_0_14_uop_robIdx_value <= _GEN_67485;
        end
      end else begin
        flow_entry_0_14_uop_robIdx_value <= _GEN_67485;
      end
    end
    if (needAlloc_0) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
        if (5'he == index_0) begin // @[Vlflowqueue.scala 203:51]
          if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
            flow_entry_0_14_vaddr <= _vaddr_0_T_162; // @[Vlflowqueue.scala 201:51]
          end else begin
            flow_entry_0_14_vaddr <= _GEN_68015;
          end
        end else begin
          flow_entry_0_14_vaddr <= _GEN_68062;
        end
      end else begin
        flow_entry_0_14_vaddr <= _GEN_68062;
      end
    end
    if (needAlloc_0) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
        if (5'hf == index_0) begin // @[Vlflowqueue.scala 198:51]
          flow_entry_0_15_uop_robIdx_value <= io_loadRegIn_0_bits_uop_robIdx_value; // @[Vlflowqueue.scala 198:51]
        end else begin
          flow_entry_0_15_uop_robIdx_value <= _GEN_67486;
        end
      end else begin
        flow_entry_0_15_uop_robIdx_value <= _GEN_67486;
      end
    end
    if (needAlloc_0) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
        if (5'hf == index_0) begin // @[Vlflowqueue.scala 203:51]
          if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
            flow_entry_0_15_vaddr <= _vaddr_0_T_162; // @[Vlflowqueue.scala 201:51]
          end else begin
            flow_entry_0_15_vaddr <= _GEN_68015;
          end
        end else begin
          flow_entry_0_15_vaddr <= _GEN_68063;
        end
      end else begin
        flow_entry_0_15_vaddr <= _GEN_68063;
      end
    end
    if (needAlloc_0) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
        if (5'h10 == index_0) begin // @[Vlflowqueue.scala 198:51]
          flow_entry_0_16_uop_robIdx_value <= io_loadRegIn_0_bits_uop_robIdx_value; // @[Vlflowqueue.scala 198:51]
        end else begin
          flow_entry_0_16_uop_robIdx_value <= _GEN_67487;
        end
      end else begin
        flow_entry_0_16_uop_robIdx_value <= _GEN_67487;
      end
    end
    if (needAlloc_0) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
        if (5'h10 == index_0) begin // @[Vlflowqueue.scala 203:51]
          if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
            flow_entry_0_16_vaddr <= _vaddr_0_T_162; // @[Vlflowqueue.scala 201:51]
          end else begin
            flow_entry_0_16_vaddr <= _GEN_68015;
          end
        end else begin
          flow_entry_0_16_vaddr <= _GEN_68064;
        end
      end else begin
        flow_entry_0_16_vaddr <= _GEN_68064;
      end
    end
    if (needAlloc_0) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
        if (5'h11 == index_0) begin // @[Vlflowqueue.scala 198:51]
          flow_entry_0_17_uop_robIdx_value <= io_loadRegIn_0_bits_uop_robIdx_value; // @[Vlflowqueue.scala 198:51]
        end else begin
          flow_entry_0_17_uop_robIdx_value <= _GEN_67488;
        end
      end else begin
        flow_entry_0_17_uop_robIdx_value <= _GEN_67488;
      end
    end
    if (needAlloc_0) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
        if (5'h11 == index_0) begin // @[Vlflowqueue.scala 203:51]
          if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
            flow_entry_0_17_vaddr <= _vaddr_0_T_162; // @[Vlflowqueue.scala 201:51]
          end else begin
            flow_entry_0_17_vaddr <= _GEN_68015;
          end
        end else begin
          flow_entry_0_17_vaddr <= _GEN_68065;
        end
      end else begin
        flow_entry_0_17_vaddr <= _GEN_68065;
      end
    end
    if (needAlloc_0) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
        if (5'h12 == index_0) begin // @[Vlflowqueue.scala 198:51]
          flow_entry_0_18_uop_robIdx_value <= io_loadRegIn_0_bits_uop_robIdx_value; // @[Vlflowqueue.scala 198:51]
        end else begin
          flow_entry_0_18_uop_robIdx_value <= _GEN_67489;
        end
      end else begin
        flow_entry_0_18_uop_robIdx_value <= _GEN_67489;
      end
    end
    if (needAlloc_0) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
        if (5'h12 == index_0) begin // @[Vlflowqueue.scala 203:51]
          if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
            flow_entry_0_18_vaddr <= _vaddr_0_T_162; // @[Vlflowqueue.scala 201:51]
          end else begin
            flow_entry_0_18_vaddr <= _GEN_68015;
          end
        end else begin
          flow_entry_0_18_vaddr <= _GEN_68066;
        end
      end else begin
        flow_entry_0_18_vaddr <= _GEN_68066;
      end
    end
    if (needAlloc_0) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
        if (5'h13 == index_0) begin // @[Vlflowqueue.scala 198:51]
          flow_entry_0_19_uop_robIdx_value <= io_loadRegIn_0_bits_uop_robIdx_value; // @[Vlflowqueue.scala 198:51]
        end else begin
          flow_entry_0_19_uop_robIdx_value <= _GEN_67490;
        end
      end else begin
        flow_entry_0_19_uop_robIdx_value <= _GEN_67490;
      end
    end
    if (needAlloc_0) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
        if (5'h13 == index_0) begin // @[Vlflowqueue.scala 203:51]
          if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
            flow_entry_0_19_vaddr <= _vaddr_0_T_162; // @[Vlflowqueue.scala 201:51]
          end else begin
            flow_entry_0_19_vaddr <= _GEN_68015;
          end
        end else begin
          flow_entry_0_19_vaddr <= _GEN_68067;
        end
      end else begin
        flow_entry_0_19_vaddr <= _GEN_68067;
      end
    end
    if (needAlloc_0) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
        if (5'h14 == index_0) begin // @[Vlflowqueue.scala 198:51]
          flow_entry_0_20_uop_robIdx_value <= io_loadRegIn_0_bits_uop_robIdx_value; // @[Vlflowqueue.scala 198:51]
        end else begin
          flow_entry_0_20_uop_robIdx_value <= _GEN_67491;
        end
      end else begin
        flow_entry_0_20_uop_robIdx_value <= _GEN_67491;
      end
    end
    if (needAlloc_0) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
        if (5'h14 == index_0) begin // @[Vlflowqueue.scala 203:51]
          if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
            flow_entry_0_20_vaddr <= _vaddr_0_T_162; // @[Vlflowqueue.scala 201:51]
          end else begin
            flow_entry_0_20_vaddr <= _GEN_68015;
          end
        end else begin
          flow_entry_0_20_vaddr <= _GEN_68068;
        end
      end else begin
        flow_entry_0_20_vaddr <= _GEN_68068;
      end
    end
    if (needAlloc_0) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
        if (5'h15 == index_0) begin // @[Vlflowqueue.scala 198:51]
          flow_entry_0_21_uop_robIdx_value <= io_loadRegIn_0_bits_uop_robIdx_value; // @[Vlflowqueue.scala 198:51]
        end else begin
          flow_entry_0_21_uop_robIdx_value <= _GEN_67492;
        end
      end else begin
        flow_entry_0_21_uop_robIdx_value <= _GEN_67492;
      end
    end
    if (needAlloc_0) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
        if (5'h15 == index_0) begin // @[Vlflowqueue.scala 203:51]
          if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
            flow_entry_0_21_vaddr <= _vaddr_0_T_162; // @[Vlflowqueue.scala 201:51]
          end else begin
            flow_entry_0_21_vaddr <= _GEN_68015;
          end
        end else begin
          flow_entry_0_21_vaddr <= _GEN_68069;
        end
      end else begin
        flow_entry_0_21_vaddr <= _GEN_68069;
      end
    end
    if (needAlloc_0) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
        if (5'h16 == index_0) begin // @[Vlflowqueue.scala 198:51]
          flow_entry_0_22_uop_robIdx_value <= io_loadRegIn_0_bits_uop_robIdx_value; // @[Vlflowqueue.scala 198:51]
        end else begin
          flow_entry_0_22_uop_robIdx_value <= _GEN_67493;
        end
      end else begin
        flow_entry_0_22_uop_robIdx_value <= _GEN_67493;
      end
    end
    if (needAlloc_0) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
        if (5'h16 == index_0) begin // @[Vlflowqueue.scala 203:51]
          if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
            flow_entry_0_22_vaddr <= _vaddr_0_T_162; // @[Vlflowqueue.scala 201:51]
          end else begin
            flow_entry_0_22_vaddr <= _GEN_68015;
          end
        end else begin
          flow_entry_0_22_vaddr <= _GEN_68070;
        end
      end else begin
        flow_entry_0_22_vaddr <= _GEN_68070;
      end
    end
    if (needAlloc_0) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
        if (5'h17 == index_0) begin // @[Vlflowqueue.scala 198:51]
          flow_entry_0_23_uop_robIdx_value <= io_loadRegIn_0_bits_uop_robIdx_value; // @[Vlflowqueue.scala 198:51]
        end else begin
          flow_entry_0_23_uop_robIdx_value <= _GEN_67494;
        end
      end else begin
        flow_entry_0_23_uop_robIdx_value <= _GEN_67494;
      end
    end
    if (needAlloc_0) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
        if (5'h17 == index_0) begin // @[Vlflowqueue.scala 203:51]
          if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
            flow_entry_0_23_vaddr <= _vaddr_0_T_162; // @[Vlflowqueue.scala 201:51]
          end else begin
            flow_entry_0_23_vaddr <= _GEN_68015;
          end
        end else begin
          flow_entry_0_23_vaddr <= _GEN_68071;
        end
      end else begin
        flow_entry_0_23_vaddr <= _GEN_68071;
      end
    end
    if (needAlloc_0) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
        if (5'h18 == index_0) begin // @[Vlflowqueue.scala 198:51]
          flow_entry_0_24_uop_robIdx_value <= io_loadRegIn_0_bits_uop_robIdx_value; // @[Vlflowqueue.scala 198:51]
        end else begin
          flow_entry_0_24_uop_robIdx_value <= _GEN_67495;
        end
      end else begin
        flow_entry_0_24_uop_robIdx_value <= _GEN_67495;
      end
    end
    if (needAlloc_0) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
        if (5'h18 == index_0) begin // @[Vlflowqueue.scala 203:51]
          if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
            flow_entry_0_24_vaddr <= _vaddr_0_T_162; // @[Vlflowqueue.scala 201:51]
          end else begin
            flow_entry_0_24_vaddr <= _GEN_68015;
          end
        end else begin
          flow_entry_0_24_vaddr <= _GEN_68072;
        end
      end else begin
        flow_entry_0_24_vaddr <= _GEN_68072;
      end
    end
    if (needAlloc_0) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
        if (5'h19 == index_0) begin // @[Vlflowqueue.scala 198:51]
          flow_entry_0_25_uop_robIdx_value <= io_loadRegIn_0_bits_uop_robIdx_value; // @[Vlflowqueue.scala 198:51]
        end else begin
          flow_entry_0_25_uop_robIdx_value <= _GEN_67496;
        end
      end else begin
        flow_entry_0_25_uop_robIdx_value <= _GEN_67496;
      end
    end
    if (needAlloc_0) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
        if (5'h19 == index_0) begin // @[Vlflowqueue.scala 203:51]
          if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
            flow_entry_0_25_vaddr <= _vaddr_0_T_162; // @[Vlflowqueue.scala 201:51]
          end else begin
            flow_entry_0_25_vaddr <= _GEN_68015;
          end
        end else begin
          flow_entry_0_25_vaddr <= _GEN_68073;
        end
      end else begin
        flow_entry_0_25_vaddr <= _GEN_68073;
      end
    end
    if (needAlloc_0) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
        if (5'h1a == index_0) begin // @[Vlflowqueue.scala 198:51]
          flow_entry_0_26_uop_robIdx_value <= io_loadRegIn_0_bits_uop_robIdx_value; // @[Vlflowqueue.scala 198:51]
        end else begin
          flow_entry_0_26_uop_robIdx_value <= _GEN_67497;
        end
      end else begin
        flow_entry_0_26_uop_robIdx_value <= _GEN_67497;
      end
    end
    if (needAlloc_0) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
        if (5'h1a == index_0) begin // @[Vlflowqueue.scala 203:51]
          if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
            flow_entry_0_26_vaddr <= _vaddr_0_T_162; // @[Vlflowqueue.scala 201:51]
          end else begin
            flow_entry_0_26_vaddr <= _GEN_68015;
          end
        end else begin
          flow_entry_0_26_vaddr <= _GEN_68074;
        end
      end else begin
        flow_entry_0_26_vaddr <= _GEN_68074;
      end
    end
    if (needAlloc_0) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
        if (5'h1b == index_0) begin // @[Vlflowqueue.scala 198:51]
          flow_entry_0_27_uop_robIdx_value <= io_loadRegIn_0_bits_uop_robIdx_value; // @[Vlflowqueue.scala 198:51]
        end else begin
          flow_entry_0_27_uop_robIdx_value <= _GEN_67498;
        end
      end else begin
        flow_entry_0_27_uop_robIdx_value <= _GEN_67498;
      end
    end
    if (needAlloc_0) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
        if (5'h1b == index_0) begin // @[Vlflowqueue.scala 203:51]
          if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
            flow_entry_0_27_vaddr <= _vaddr_0_T_162; // @[Vlflowqueue.scala 201:51]
          end else begin
            flow_entry_0_27_vaddr <= _GEN_68015;
          end
        end else begin
          flow_entry_0_27_vaddr <= _GEN_68075;
        end
      end else begin
        flow_entry_0_27_vaddr <= _GEN_68075;
      end
    end
    if (needAlloc_0) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
        if (5'h1c == index_0) begin // @[Vlflowqueue.scala 198:51]
          flow_entry_0_28_uop_robIdx_value <= io_loadRegIn_0_bits_uop_robIdx_value; // @[Vlflowqueue.scala 198:51]
        end else begin
          flow_entry_0_28_uop_robIdx_value <= _GEN_67499;
        end
      end else begin
        flow_entry_0_28_uop_robIdx_value <= _GEN_67499;
      end
    end
    if (needAlloc_0) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
        if (5'h1c == index_0) begin // @[Vlflowqueue.scala 203:51]
          if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
            flow_entry_0_28_vaddr <= _vaddr_0_T_162; // @[Vlflowqueue.scala 201:51]
          end else begin
            flow_entry_0_28_vaddr <= _GEN_68015;
          end
        end else begin
          flow_entry_0_28_vaddr <= _GEN_68076;
        end
      end else begin
        flow_entry_0_28_vaddr <= _GEN_68076;
      end
    end
    if (needAlloc_0) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
        if (5'h1d == index_0) begin // @[Vlflowqueue.scala 198:51]
          flow_entry_0_29_uop_robIdx_value <= io_loadRegIn_0_bits_uop_robIdx_value; // @[Vlflowqueue.scala 198:51]
        end else begin
          flow_entry_0_29_uop_robIdx_value <= _GEN_67500;
        end
      end else begin
        flow_entry_0_29_uop_robIdx_value <= _GEN_67500;
      end
    end
    if (needAlloc_0) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
        if (5'h1d == index_0) begin // @[Vlflowqueue.scala 203:51]
          if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
            flow_entry_0_29_vaddr <= _vaddr_0_T_162; // @[Vlflowqueue.scala 201:51]
          end else begin
            flow_entry_0_29_vaddr <= _GEN_68015;
          end
        end else begin
          flow_entry_0_29_vaddr <= _GEN_68077;
        end
      end else begin
        flow_entry_0_29_vaddr <= _GEN_68077;
      end
    end
    if (needAlloc_0) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
        if (5'h1e == index_0) begin // @[Vlflowqueue.scala 198:51]
          flow_entry_0_30_uop_robIdx_value <= io_loadRegIn_0_bits_uop_robIdx_value; // @[Vlflowqueue.scala 198:51]
        end else begin
          flow_entry_0_30_uop_robIdx_value <= _GEN_67501;
        end
      end else begin
        flow_entry_0_30_uop_robIdx_value <= _GEN_67501;
      end
    end
    if (needAlloc_0) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
        if (5'h1e == index_0) begin // @[Vlflowqueue.scala 203:51]
          if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
            flow_entry_0_30_vaddr <= _vaddr_0_T_162; // @[Vlflowqueue.scala 201:51]
          end else begin
            flow_entry_0_30_vaddr <= _GEN_68015;
          end
        end else begin
          flow_entry_0_30_vaddr <= _GEN_68078;
        end
      end else begin
        flow_entry_0_30_vaddr <= _GEN_68078;
      end
    end
    if (needAlloc_0) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
        if (5'h1f == index_0) begin // @[Vlflowqueue.scala 198:51]
          flow_entry_0_31_uop_robIdx_value <= io_loadRegIn_0_bits_uop_robIdx_value; // @[Vlflowqueue.scala 198:51]
        end else begin
          flow_entry_0_31_uop_robIdx_value <= _GEN_67502;
        end
      end else begin
        flow_entry_0_31_uop_robIdx_value <= _GEN_67502;
      end
    end
    if (needAlloc_0) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
        if (5'h1f == index_0) begin // @[Vlflowqueue.scala 203:51]
          if (4'h8 < realFlowNum_0) begin // @[Vlflowqueue.scala 194:37]
            flow_entry_0_31_vaddr <= _vaddr_0_T_162; // @[Vlflowqueue.scala 201:51]
          end else begin
            flow_entry_0_31_vaddr <= _GEN_68015;
          end
        end else begin
          flow_entry_0_31_vaddr <= _GEN_68079;
        end
      end else begin
        flow_entry_0_31_vaddr <= _GEN_68079;
      end
    end
    if (needAlloc_1) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
        if (5'h0 == index_1) begin // @[Vlflowqueue.scala 198:51]
          flow_entry_1_0_uop_robIdx_value <= io_loadRegIn_1_bits_uop_robIdx_value; // @[Vlflowqueue.scala 198:51]
        end else begin
          flow_entry_1_0_uop_robIdx_value <= _GEN_147716;
        end
      end else begin
        flow_entry_1_0_uop_robIdx_value <= _GEN_147716;
      end
    end
    if (needAlloc_1) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
        if (5'h0 == index_1) begin // @[Vlflowqueue.scala 203:51]
          if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
            flow_entry_1_0_vaddr <= _vaddr_1_T_162; // @[Vlflowqueue.scala 201:51]
          end else begin
            flow_entry_1_0_vaddr <= _GEN_148260;
          end
        end else begin
          flow_entry_1_0_vaddr <= _GEN_148293;
        end
      end else begin
        flow_entry_1_0_vaddr <= _GEN_148293;
      end
    end
    if (needAlloc_1) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
        if (5'h1 == index_1) begin // @[Vlflowqueue.scala 198:51]
          flow_entry_1_1_uop_robIdx_value <= io_loadRegIn_1_bits_uop_robIdx_value; // @[Vlflowqueue.scala 198:51]
        end else begin
          flow_entry_1_1_uop_robIdx_value <= _GEN_147717;
        end
      end else begin
        flow_entry_1_1_uop_robIdx_value <= _GEN_147717;
      end
    end
    if (needAlloc_1) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
        if (5'h1 == index_1) begin // @[Vlflowqueue.scala 203:51]
          if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
            flow_entry_1_1_vaddr <= _vaddr_1_T_162; // @[Vlflowqueue.scala 201:51]
          end else begin
            flow_entry_1_1_vaddr <= _GEN_148260;
          end
        end else begin
          flow_entry_1_1_vaddr <= _GEN_148294;
        end
      end else begin
        flow_entry_1_1_vaddr <= _GEN_148294;
      end
    end
    if (needAlloc_1) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
        if (5'h2 == index_1) begin // @[Vlflowqueue.scala 198:51]
          flow_entry_1_2_uop_robIdx_value <= io_loadRegIn_1_bits_uop_robIdx_value; // @[Vlflowqueue.scala 198:51]
        end else begin
          flow_entry_1_2_uop_robIdx_value <= _GEN_147718;
        end
      end else begin
        flow_entry_1_2_uop_robIdx_value <= _GEN_147718;
      end
    end
    if (needAlloc_1) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
        if (5'h2 == index_1) begin // @[Vlflowqueue.scala 203:51]
          if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
            flow_entry_1_2_vaddr <= _vaddr_1_T_162; // @[Vlflowqueue.scala 201:51]
          end else begin
            flow_entry_1_2_vaddr <= _GEN_148260;
          end
        end else begin
          flow_entry_1_2_vaddr <= _GEN_148295;
        end
      end else begin
        flow_entry_1_2_vaddr <= _GEN_148295;
      end
    end
    if (needAlloc_1) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
        if (5'h3 == index_1) begin // @[Vlflowqueue.scala 198:51]
          flow_entry_1_3_uop_robIdx_value <= io_loadRegIn_1_bits_uop_robIdx_value; // @[Vlflowqueue.scala 198:51]
        end else begin
          flow_entry_1_3_uop_robIdx_value <= _GEN_147719;
        end
      end else begin
        flow_entry_1_3_uop_robIdx_value <= _GEN_147719;
      end
    end
    if (needAlloc_1) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
        if (5'h3 == index_1) begin // @[Vlflowqueue.scala 203:51]
          if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
            flow_entry_1_3_vaddr <= _vaddr_1_T_162; // @[Vlflowqueue.scala 201:51]
          end else begin
            flow_entry_1_3_vaddr <= _GEN_148260;
          end
        end else begin
          flow_entry_1_3_vaddr <= _GEN_148296;
        end
      end else begin
        flow_entry_1_3_vaddr <= _GEN_148296;
      end
    end
    if (needAlloc_1) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
        if (5'h4 == index_1) begin // @[Vlflowqueue.scala 198:51]
          flow_entry_1_4_uop_robIdx_value <= io_loadRegIn_1_bits_uop_robIdx_value; // @[Vlflowqueue.scala 198:51]
        end else begin
          flow_entry_1_4_uop_robIdx_value <= _GEN_147720;
        end
      end else begin
        flow_entry_1_4_uop_robIdx_value <= _GEN_147720;
      end
    end
    if (needAlloc_1) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
        if (5'h4 == index_1) begin // @[Vlflowqueue.scala 203:51]
          if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
            flow_entry_1_4_vaddr <= _vaddr_1_T_162; // @[Vlflowqueue.scala 201:51]
          end else begin
            flow_entry_1_4_vaddr <= _GEN_148260;
          end
        end else begin
          flow_entry_1_4_vaddr <= _GEN_148297;
        end
      end else begin
        flow_entry_1_4_vaddr <= _GEN_148297;
      end
    end
    if (needAlloc_1) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
        if (5'h5 == index_1) begin // @[Vlflowqueue.scala 198:51]
          flow_entry_1_5_uop_robIdx_value <= io_loadRegIn_1_bits_uop_robIdx_value; // @[Vlflowqueue.scala 198:51]
        end else begin
          flow_entry_1_5_uop_robIdx_value <= _GEN_147721;
        end
      end else begin
        flow_entry_1_5_uop_robIdx_value <= _GEN_147721;
      end
    end
    if (needAlloc_1) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
        if (5'h5 == index_1) begin // @[Vlflowqueue.scala 203:51]
          if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
            flow_entry_1_5_vaddr <= _vaddr_1_T_162; // @[Vlflowqueue.scala 201:51]
          end else begin
            flow_entry_1_5_vaddr <= _GEN_148260;
          end
        end else begin
          flow_entry_1_5_vaddr <= _GEN_148298;
        end
      end else begin
        flow_entry_1_5_vaddr <= _GEN_148298;
      end
    end
    if (needAlloc_1) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
        if (5'h6 == index_1) begin // @[Vlflowqueue.scala 198:51]
          flow_entry_1_6_uop_robIdx_value <= io_loadRegIn_1_bits_uop_robIdx_value; // @[Vlflowqueue.scala 198:51]
        end else begin
          flow_entry_1_6_uop_robIdx_value <= _GEN_147722;
        end
      end else begin
        flow_entry_1_6_uop_robIdx_value <= _GEN_147722;
      end
    end
    if (needAlloc_1) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
        if (5'h6 == index_1) begin // @[Vlflowqueue.scala 203:51]
          if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
            flow_entry_1_6_vaddr <= _vaddr_1_T_162; // @[Vlflowqueue.scala 201:51]
          end else begin
            flow_entry_1_6_vaddr <= _GEN_148260;
          end
        end else begin
          flow_entry_1_6_vaddr <= _GEN_148299;
        end
      end else begin
        flow_entry_1_6_vaddr <= _GEN_148299;
      end
    end
    if (needAlloc_1) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
        if (5'h7 == index_1) begin // @[Vlflowqueue.scala 198:51]
          flow_entry_1_7_uop_robIdx_value <= io_loadRegIn_1_bits_uop_robIdx_value; // @[Vlflowqueue.scala 198:51]
        end else begin
          flow_entry_1_7_uop_robIdx_value <= _GEN_147723;
        end
      end else begin
        flow_entry_1_7_uop_robIdx_value <= _GEN_147723;
      end
    end
    if (needAlloc_1) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
        if (5'h7 == index_1) begin // @[Vlflowqueue.scala 203:51]
          if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
            flow_entry_1_7_vaddr <= _vaddr_1_T_162; // @[Vlflowqueue.scala 201:51]
          end else begin
            flow_entry_1_7_vaddr <= _GEN_148260;
          end
        end else begin
          flow_entry_1_7_vaddr <= _GEN_148300;
        end
      end else begin
        flow_entry_1_7_vaddr <= _GEN_148300;
      end
    end
    if (needAlloc_1) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
        if (5'h8 == index_1) begin // @[Vlflowqueue.scala 198:51]
          flow_entry_1_8_uop_robIdx_value <= io_loadRegIn_1_bits_uop_robIdx_value; // @[Vlflowqueue.scala 198:51]
        end else begin
          flow_entry_1_8_uop_robIdx_value <= _GEN_147724;
        end
      end else begin
        flow_entry_1_8_uop_robIdx_value <= _GEN_147724;
      end
    end
    if (needAlloc_1) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
        if (5'h8 == index_1) begin // @[Vlflowqueue.scala 203:51]
          if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
            flow_entry_1_8_vaddr <= _vaddr_1_T_162; // @[Vlflowqueue.scala 201:51]
          end else begin
            flow_entry_1_8_vaddr <= _GEN_148260;
          end
        end else begin
          flow_entry_1_8_vaddr <= _GEN_148301;
        end
      end else begin
        flow_entry_1_8_vaddr <= _GEN_148301;
      end
    end
    if (needAlloc_1) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
        if (5'h9 == index_1) begin // @[Vlflowqueue.scala 198:51]
          flow_entry_1_9_uop_robIdx_value <= io_loadRegIn_1_bits_uop_robIdx_value; // @[Vlflowqueue.scala 198:51]
        end else begin
          flow_entry_1_9_uop_robIdx_value <= _GEN_147725;
        end
      end else begin
        flow_entry_1_9_uop_robIdx_value <= _GEN_147725;
      end
    end
    if (needAlloc_1) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
        if (5'h9 == index_1) begin // @[Vlflowqueue.scala 203:51]
          if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
            flow_entry_1_9_vaddr <= _vaddr_1_T_162; // @[Vlflowqueue.scala 201:51]
          end else begin
            flow_entry_1_9_vaddr <= _GEN_148260;
          end
        end else begin
          flow_entry_1_9_vaddr <= _GEN_148302;
        end
      end else begin
        flow_entry_1_9_vaddr <= _GEN_148302;
      end
    end
    if (needAlloc_1) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
        if (5'ha == index_1) begin // @[Vlflowqueue.scala 198:51]
          flow_entry_1_10_uop_robIdx_value <= io_loadRegIn_1_bits_uop_robIdx_value; // @[Vlflowqueue.scala 198:51]
        end else begin
          flow_entry_1_10_uop_robIdx_value <= _GEN_147726;
        end
      end else begin
        flow_entry_1_10_uop_robIdx_value <= _GEN_147726;
      end
    end
    if (needAlloc_1) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
        if (5'ha == index_1) begin // @[Vlflowqueue.scala 203:51]
          if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
            flow_entry_1_10_vaddr <= _vaddr_1_T_162; // @[Vlflowqueue.scala 201:51]
          end else begin
            flow_entry_1_10_vaddr <= _GEN_148260;
          end
        end else begin
          flow_entry_1_10_vaddr <= _GEN_148303;
        end
      end else begin
        flow_entry_1_10_vaddr <= _GEN_148303;
      end
    end
    if (needAlloc_1) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
        if (5'hb == index_1) begin // @[Vlflowqueue.scala 198:51]
          flow_entry_1_11_uop_robIdx_value <= io_loadRegIn_1_bits_uop_robIdx_value; // @[Vlflowqueue.scala 198:51]
        end else begin
          flow_entry_1_11_uop_robIdx_value <= _GEN_147727;
        end
      end else begin
        flow_entry_1_11_uop_robIdx_value <= _GEN_147727;
      end
    end
    if (needAlloc_1) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
        if (5'hb == index_1) begin // @[Vlflowqueue.scala 203:51]
          if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
            flow_entry_1_11_vaddr <= _vaddr_1_T_162; // @[Vlflowqueue.scala 201:51]
          end else begin
            flow_entry_1_11_vaddr <= _GEN_148260;
          end
        end else begin
          flow_entry_1_11_vaddr <= _GEN_148304;
        end
      end else begin
        flow_entry_1_11_vaddr <= _GEN_148304;
      end
    end
    if (needAlloc_1) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
        if (5'hc == index_1) begin // @[Vlflowqueue.scala 198:51]
          flow_entry_1_12_uop_robIdx_value <= io_loadRegIn_1_bits_uop_robIdx_value; // @[Vlflowqueue.scala 198:51]
        end else begin
          flow_entry_1_12_uop_robIdx_value <= _GEN_147728;
        end
      end else begin
        flow_entry_1_12_uop_robIdx_value <= _GEN_147728;
      end
    end
    if (needAlloc_1) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
        if (5'hc == index_1) begin // @[Vlflowqueue.scala 203:51]
          if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
            flow_entry_1_12_vaddr <= _vaddr_1_T_162; // @[Vlflowqueue.scala 201:51]
          end else begin
            flow_entry_1_12_vaddr <= _GEN_148260;
          end
        end else begin
          flow_entry_1_12_vaddr <= _GEN_148305;
        end
      end else begin
        flow_entry_1_12_vaddr <= _GEN_148305;
      end
    end
    if (needAlloc_1) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
        if (5'hd == index_1) begin // @[Vlflowqueue.scala 198:51]
          flow_entry_1_13_uop_robIdx_value <= io_loadRegIn_1_bits_uop_robIdx_value; // @[Vlflowqueue.scala 198:51]
        end else begin
          flow_entry_1_13_uop_robIdx_value <= _GEN_147729;
        end
      end else begin
        flow_entry_1_13_uop_robIdx_value <= _GEN_147729;
      end
    end
    if (needAlloc_1) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
        if (5'hd == index_1) begin // @[Vlflowqueue.scala 203:51]
          if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
            flow_entry_1_13_vaddr <= _vaddr_1_T_162; // @[Vlflowqueue.scala 201:51]
          end else begin
            flow_entry_1_13_vaddr <= _GEN_148260;
          end
        end else begin
          flow_entry_1_13_vaddr <= _GEN_148306;
        end
      end else begin
        flow_entry_1_13_vaddr <= _GEN_148306;
      end
    end
    if (needAlloc_1) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
        if (5'he == index_1) begin // @[Vlflowqueue.scala 198:51]
          flow_entry_1_14_uop_robIdx_value <= io_loadRegIn_1_bits_uop_robIdx_value; // @[Vlflowqueue.scala 198:51]
        end else begin
          flow_entry_1_14_uop_robIdx_value <= _GEN_147730;
        end
      end else begin
        flow_entry_1_14_uop_robIdx_value <= _GEN_147730;
      end
    end
    if (needAlloc_1) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
        if (5'he == index_1) begin // @[Vlflowqueue.scala 203:51]
          if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
            flow_entry_1_14_vaddr <= _vaddr_1_T_162; // @[Vlflowqueue.scala 201:51]
          end else begin
            flow_entry_1_14_vaddr <= _GEN_148260;
          end
        end else begin
          flow_entry_1_14_vaddr <= _GEN_148307;
        end
      end else begin
        flow_entry_1_14_vaddr <= _GEN_148307;
      end
    end
    if (needAlloc_1) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
        if (5'hf == index_1) begin // @[Vlflowqueue.scala 198:51]
          flow_entry_1_15_uop_robIdx_value <= io_loadRegIn_1_bits_uop_robIdx_value; // @[Vlflowqueue.scala 198:51]
        end else begin
          flow_entry_1_15_uop_robIdx_value <= _GEN_147731;
        end
      end else begin
        flow_entry_1_15_uop_robIdx_value <= _GEN_147731;
      end
    end
    if (needAlloc_1) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
        if (5'hf == index_1) begin // @[Vlflowqueue.scala 203:51]
          if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
            flow_entry_1_15_vaddr <= _vaddr_1_T_162; // @[Vlflowqueue.scala 201:51]
          end else begin
            flow_entry_1_15_vaddr <= _GEN_148260;
          end
        end else begin
          flow_entry_1_15_vaddr <= _GEN_148308;
        end
      end else begin
        flow_entry_1_15_vaddr <= _GEN_148308;
      end
    end
    if (needAlloc_1) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
        if (5'h10 == index_1) begin // @[Vlflowqueue.scala 198:51]
          flow_entry_1_16_uop_robIdx_value <= io_loadRegIn_1_bits_uop_robIdx_value; // @[Vlflowqueue.scala 198:51]
        end else begin
          flow_entry_1_16_uop_robIdx_value <= _GEN_147732;
        end
      end else begin
        flow_entry_1_16_uop_robIdx_value <= _GEN_147732;
      end
    end
    if (needAlloc_1) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
        if (5'h10 == index_1) begin // @[Vlflowqueue.scala 203:51]
          if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
            flow_entry_1_16_vaddr <= _vaddr_1_T_162; // @[Vlflowqueue.scala 201:51]
          end else begin
            flow_entry_1_16_vaddr <= _GEN_148260;
          end
        end else begin
          flow_entry_1_16_vaddr <= _GEN_148309;
        end
      end else begin
        flow_entry_1_16_vaddr <= _GEN_148309;
      end
    end
    if (needAlloc_1) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
        if (5'h11 == index_1) begin // @[Vlflowqueue.scala 198:51]
          flow_entry_1_17_uop_robIdx_value <= io_loadRegIn_1_bits_uop_robIdx_value; // @[Vlflowqueue.scala 198:51]
        end else begin
          flow_entry_1_17_uop_robIdx_value <= _GEN_147733;
        end
      end else begin
        flow_entry_1_17_uop_robIdx_value <= _GEN_147733;
      end
    end
    if (needAlloc_1) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
        if (5'h11 == index_1) begin // @[Vlflowqueue.scala 203:51]
          if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
            flow_entry_1_17_vaddr <= _vaddr_1_T_162; // @[Vlflowqueue.scala 201:51]
          end else begin
            flow_entry_1_17_vaddr <= _GEN_148260;
          end
        end else begin
          flow_entry_1_17_vaddr <= _GEN_148310;
        end
      end else begin
        flow_entry_1_17_vaddr <= _GEN_148310;
      end
    end
    if (needAlloc_1) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
        if (5'h12 == index_1) begin // @[Vlflowqueue.scala 198:51]
          flow_entry_1_18_uop_robIdx_value <= io_loadRegIn_1_bits_uop_robIdx_value; // @[Vlflowqueue.scala 198:51]
        end else begin
          flow_entry_1_18_uop_robIdx_value <= _GEN_147734;
        end
      end else begin
        flow_entry_1_18_uop_robIdx_value <= _GEN_147734;
      end
    end
    if (needAlloc_1) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
        if (5'h12 == index_1) begin // @[Vlflowqueue.scala 203:51]
          if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
            flow_entry_1_18_vaddr <= _vaddr_1_T_162; // @[Vlflowqueue.scala 201:51]
          end else begin
            flow_entry_1_18_vaddr <= _GEN_148260;
          end
        end else begin
          flow_entry_1_18_vaddr <= _GEN_148311;
        end
      end else begin
        flow_entry_1_18_vaddr <= _GEN_148311;
      end
    end
    if (needAlloc_1) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
        if (5'h13 == index_1) begin // @[Vlflowqueue.scala 198:51]
          flow_entry_1_19_uop_robIdx_value <= io_loadRegIn_1_bits_uop_robIdx_value; // @[Vlflowqueue.scala 198:51]
        end else begin
          flow_entry_1_19_uop_robIdx_value <= _GEN_147735;
        end
      end else begin
        flow_entry_1_19_uop_robIdx_value <= _GEN_147735;
      end
    end
    if (needAlloc_1) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
        if (5'h13 == index_1) begin // @[Vlflowqueue.scala 203:51]
          if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
            flow_entry_1_19_vaddr <= _vaddr_1_T_162; // @[Vlflowqueue.scala 201:51]
          end else begin
            flow_entry_1_19_vaddr <= _GEN_148260;
          end
        end else begin
          flow_entry_1_19_vaddr <= _GEN_148312;
        end
      end else begin
        flow_entry_1_19_vaddr <= _GEN_148312;
      end
    end
    if (needAlloc_1) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
        if (5'h14 == index_1) begin // @[Vlflowqueue.scala 198:51]
          flow_entry_1_20_uop_robIdx_value <= io_loadRegIn_1_bits_uop_robIdx_value; // @[Vlflowqueue.scala 198:51]
        end else begin
          flow_entry_1_20_uop_robIdx_value <= _GEN_147736;
        end
      end else begin
        flow_entry_1_20_uop_robIdx_value <= _GEN_147736;
      end
    end
    if (needAlloc_1) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
        if (5'h14 == index_1) begin // @[Vlflowqueue.scala 203:51]
          if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
            flow_entry_1_20_vaddr <= _vaddr_1_T_162; // @[Vlflowqueue.scala 201:51]
          end else begin
            flow_entry_1_20_vaddr <= _GEN_148260;
          end
        end else begin
          flow_entry_1_20_vaddr <= _GEN_148313;
        end
      end else begin
        flow_entry_1_20_vaddr <= _GEN_148313;
      end
    end
    if (needAlloc_1) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
        if (5'h15 == index_1) begin // @[Vlflowqueue.scala 198:51]
          flow_entry_1_21_uop_robIdx_value <= io_loadRegIn_1_bits_uop_robIdx_value; // @[Vlflowqueue.scala 198:51]
        end else begin
          flow_entry_1_21_uop_robIdx_value <= _GEN_147737;
        end
      end else begin
        flow_entry_1_21_uop_robIdx_value <= _GEN_147737;
      end
    end
    if (needAlloc_1) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
        if (5'h15 == index_1) begin // @[Vlflowqueue.scala 203:51]
          if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
            flow_entry_1_21_vaddr <= _vaddr_1_T_162; // @[Vlflowqueue.scala 201:51]
          end else begin
            flow_entry_1_21_vaddr <= _GEN_148260;
          end
        end else begin
          flow_entry_1_21_vaddr <= _GEN_148314;
        end
      end else begin
        flow_entry_1_21_vaddr <= _GEN_148314;
      end
    end
    if (needAlloc_1) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
        if (5'h16 == index_1) begin // @[Vlflowqueue.scala 198:51]
          flow_entry_1_22_uop_robIdx_value <= io_loadRegIn_1_bits_uop_robIdx_value; // @[Vlflowqueue.scala 198:51]
        end else begin
          flow_entry_1_22_uop_robIdx_value <= _GEN_147738;
        end
      end else begin
        flow_entry_1_22_uop_robIdx_value <= _GEN_147738;
      end
    end
    if (needAlloc_1) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
        if (5'h16 == index_1) begin // @[Vlflowqueue.scala 203:51]
          if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
            flow_entry_1_22_vaddr <= _vaddr_1_T_162; // @[Vlflowqueue.scala 201:51]
          end else begin
            flow_entry_1_22_vaddr <= _GEN_148260;
          end
        end else begin
          flow_entry_1_22_vaddr <= _GEN_148315;
        end
      end else begin
        flow_entry_1_22_vaddr <= _GEN_148315;
      end
    end
    if (needAlloc_1) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
        if (5'h17 == index_1) begin // @[Vlflowqueue.scala 198:51]
          flow_entry_1_23_uop_robIdx_value <= io_loadRegIn_1_bits_uop_robIdx_value; // @[Vlflowqueue.scala 198:51]
        end else begin
          flow_entry_1_23_uop_robIdx_value <= _GEN_147739;
        end
      end else begin
        flow_entry_1_23_uop_robIdx_value <= _GEN_147739;
      end
    end
    if (needAlloc_1) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
        if (5'h17 == index_1) begin // @[Vlflowqueue.scala 203:51]
          if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
            flow_entry_1_23_vaddr <= _vaddr_1_T_162; // @[Vlflowqueue.scala 201:51]
          end else begin
            flow_entry_1_23_vaddr <= _GEN_148260;
          end
        end else begin
          flow_entry_1_23_vaddr <= _GEN_148316;
        end
      end else begin
        flow_entry_1_23_vaddr <= _GEN_148316;
      end
    end
    if (needAlloc_1) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
        if (5'h18 == index_1) begin // @[Vlflowqueue.scala 198:51]
          flow_entry_1_24_uop_robIdx_value <= io_loadRegIn_1_bits_uop_robIdx_value; // @[Vlflowqueue.scala 198:51]
        end else begin
          flow_entry_1_24_uop_robIdx_value <= _GEN_147740;
        end
      end else begin
        flow_entry_1_24_uop_robIdx_value <= _GEN_147740;
      end
    end
    if (needAlloc_1) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
        if (5'h18 == index_1) begin // @[Vlflowqueue.scala 203:51]
          if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
            flow_entry_1_24_vaddr <= _vaddr_1_T_162; // @[Vlflowqueue.scala 201:51]
          end else begin
            flow_entry_1_24_vaddr <= _GEN_148260;
          end
        end else begin
          flow_entry_1_24_vaddr <= _GEN_148317;
        end
      end else begin
        flow_entry_1_24_vaddr <= _GEN_148317;
      end
    end
    if (needAlloc_1) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
        if (5'h19 == index_1) begin // @[Vlflowqueue.scala 198:51]
          flow_entry_1_25_uop_robIdx_value <= io_loadRegIn_1_bits_uop_robIdx_value; // @[Vlflowqueue.scala 198:51]
        end else begin
          flow_entry_1_25_uop_robIdx_value <= _GEN_147741;
        end
      end else begin
        flow_entry_1_25_uop_robIdx_value <= _GEN_147741;
      end
    end
    if (needAlloc_1) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
        if (5'h19 == index_1) begin // @[Vlflowqueue.scala 203:51]
          if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
            flow_entry_1_25_vaddr <= _vaddr_1_T_162; // @[Vlflowqueue.scala 201:51]
          end else begin
            flow_entry_1_25_vaddr <= _GEN_148260;
          end
        end else begin
          flow_entry_1_25_vaddr <= _GEN_148318;
        end
      end else begin
        flow_entry_1_25_vaddr <= _GEN_148318;
      end
    end
    if (needAlloc_1) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
        if (5'h1a == index_1) begin // @[Vlflowqueue.scala 198:51]
          flow_entry_1_26_uop_robIdx_value <= io_loadRegIn_1_bits_uop_robIdx_value; // @[Vlflowqueue.scala 198:51]
        end else begin
          flow_entry_1_26_uop_robIdx_value <= _GEN_147742;
        end
      end else begin
        flow_entry_1_26_uop_robIdx_value <= _GEN_147742;
      end
    end
    if (needAlloc_1) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
        if (5'h1a == index_1) begin // @[Vlflowqueue.scala 203:51]
          if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
            flow_entry_1_26_vaddr <= _vaddr_1_T_162; // @[Vlflowqueue.scala 201:51]
          end else begin
            flow_entry_1_26_vaddr <= _GEN_148260;
          end
        end else begin
          flow_entry_1_26_vaddr <= _GEN_148319;
        end
      end else begin
        flow_entry_1_26_vaddr <= _GEN_148319;
      end
    end
    if (needAlloc_1) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
        if (5'h1b == index_1) begin // @[Vlflowqueue.scala 198:51]
          flow_entry_1_27_uop_robIdx_value <= io_loadRegIn_1_bits_uop_robIdx_value; // @[Vlflowqueue.scala 198:51]
        end else begin
          flow_entry_1_27_uop_robIdx_value <= _GEN_147743;
        end
      end else begin
        flow_entry_1_27_uop_robIdx_value <= _GEN_147743;
      end
    end
    if (needAlloc_1) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
        if (5'h1b == index_1) begin // @[Vlflowqueue.scala 203:51]
          if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
            flow_entry_1_27_vaddr <= _vaddr_1_T_162; // @[Vlflowqueue.scala 201:51]
          end else begin
            flow_entry_1_27_vaddr <= _GEN_148260;
          end
        end else begin
          flow_entry_1_27_vaddr <= _GEN_148320;
        end
      end else begin
        flow_entry_1_27_vaddr <= _GEN_148320;
      end
    end
    if (needAlloc_1) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
        if (5'h1c == index_1) begin // @[Vlflowqueue.scala 198:51]
          flow_entry_1_28_uop_robIdx_value <= io_loadRegIn_1_bits_uop_robIdx_value; // @[Vlflowqueue.scala 198:51]
        end else begin
          flow_entry_1_28_uop_robIdx_value <= _GEN_147744;
        end
      end else begin
        flow_entry_1_28_uop_robIdx_value <= _GEN_147744;
      end
    end
    if (needAlloc_1) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
        if (5'h1c == index_1) begin // @[Vlflowqueue.scala 203:51]
          if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
            flow_entry_1_28_vaddr <= _vaddr_1_T_162; // @[Vlflowqueue.scala 201:51]
          end else begin
            flow_entry_1_28_vaddr <= _GEN_148260;
          end
        end else begin
          flow_entry_1_28_vaddr <= _GEN_148321;
        end
      end else begin
        flow_entry_1_28_vaddr <= _GEN_148321;
      end
    end
    if (needAlloc_1) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
        if (5'h1d == index_1) begin // @[Vlflowqueue.scala 198:51]
          flow_entry_1_29_uop_robIdx_value <= io_loadRegIn_1_bits_uop_robIdx_value; // @[Vlflowqueue.scala 198:51]
        end else begin
          flow_entry_1_29_uop_robIdx_value <= _GEN_147745;
        end
      end else begin
        flow_entry_1_29_uop_robIdx_value <= _GEN_147745;
      end
    end
    if (needAlloc_1) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
        if (5'h1d == index_1) begin // @[Vlflowqueue.scala 203:51]
          if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
            flow_entry_1_29_vaddr <= _vaddr_1_T_162; // @[Vlflowqueue.scala 201:51]
          end else begin
            flow_entry_1_29_vaddr <= _GEN_148260;
          end
        end else begin
          flow_entry_1_29_vaddr <= _GEN_148322;
        end
      end else begin
        flow_entry_1_29_vaddr <= _GEN_148322;
      end
    end
    if (needAlloc_1) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
        if (5'h1e == index_1) begin // @[Vlflowqueue.scala 198:51]
          flow_entry_1_30_uop_robIdx_value <= io_loadRegIn_1_bits_uop_robIdx_value; // @[Vlflowqueue.scala 198:51]
        end else begin
          flow_entry_1_30_uop_robIdx_value <= _GEN_147746;
        end
      end else begin
        flow_entry_1_30_uop_robIdx_value <= _GEN_147746;
      end
    end
    if (needAlloc_1) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
        if (5'h1e == index_1) begin // @[Vlflowqueue.scala 203:51]
          if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
            flow_entry_1_30_vaddr <= _vaddr_1_T_162; // @[Vlflowqueue.scala 201:51]
          end else begin
            flow_entry_1_30_vaddr <= _GEN_148260;
          end
        end else begin
          flow_entry_1_30_vaddr <= _GEN_148323;
        end
      end else begin
        flow_entry_1_30_vaddr <= _GEN_148323;
      end
    end
    if (needAlloc_1) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
        if (5'h1f == index_1) begin // @[Vlflowqueue.scala 198:51]
          flow_entry_1_31_uop_robIdx_value <= io_loadRegIn_1_bits_uop_robIdx_value; // @[Vlflowqueue.scala 198:51]
        end else begin
          flow_entry_1_31_uop_robIdx_value <= _GEN_147747;
        end
      end else begin
        flow_entry_1_31_uop_robIdx_value <= _GEN_147747;
      end
    end
    if (needAlloc_1) begin // @[Vlflowqueue.scala 191:25]
      if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
        if (5'h1f == index_1) begin // @[Vlflowqueue.scala 203:51]
          if (4'h8 < realFlowNum_1) begin // @[Vlflowqueue.scala 194:37]
            flow_entry_1_31_vaddr <= _vaddr_1_T_162; // @[Vlflowqueue.scala 201:51]
          end else begin
            flow_entry_1_31_vaddr <= _GEN_148260;
          end
        end else begin
          flow_entry_1_31_vaddr <= _GEN_148324;
        end
      end else begin
        flow_entry_1_31_vaddr <= _GEN_148324;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Vlflowqueue.scala 250:35]
      flow_entry_valid_0_0 <= 1'h0; // @[Vlflowqueue.scala 251:{44,44}]
    end else if (_T_90) begin
      if (5'h0 == deqPtr_0_value) begin
        flow_entry_valid_0_0 <= 1'h0;
      end else begin
        flow_entry_valid_0_0 <= _GEN_76404;
      end
    end else begin
      flow_entry_valid_0_0 <= _GEN_76404;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Vlflowqueue.scala 250:35]
      flow_entry_valid_0_1 <= 1'h0; // @[Vlflowqueue.scala 251:{44,44}]
    end else if (_T_90) begin
      if (5'h1 == deqPtr_0_value) begin
        flow_entry_valid_0_1 <= 1'h0;
      end else begin
        flow_entry_valid_0_1 <= _GEN_76405;
      end
    end else begin
      flow_entry_valid_0_1 <= _GEN_76405;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Vlflowqueue.scala 250:35]
      flow_entry_valid_0_2 <= 1'h0; // @[Vlflowqueue.scala 251:{44,44}]
    end else if (_T_90) begin
      if (5'h2 == deqPtr_0_value) begin
        flow_entry_valid_0_2 <= 1'h0;
      end else begin
        flow_entry_valid_0_2 <= _GEN_76406;
      end
    end else begin
      flow_entry_valid_0_2 <= _GEN_76406;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Vlflowqueue.scala 250:35]
      flow_entry_valid_0_3 <= 1'h0; // @[Vlflowqueue.scala 251:{44,44}]
    end else if (_T_90) begin
      if (5'h3 == deqPtr_0_value) begin
        flow_entry_valid_0_3 <= 1'h0;
      end else begin
        flow_entry_valid_0_3 <= _GEN_76407;
      end
    end else begin
      flow_entry_valid_0_3 <= _GEN_76407;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Vlflowqueue.scala 250:35]
      flow_entry_valid_0_4 <= 1'h0; // @[Vlflowqueue.scala 251:{44,44}]
    end else if (_T_90) begin
      if (5'h4 == deqPtr_0_value) begin
        flow_entry_valid_0_4 <= 1'h0;
      end else begin
        flow_entry_valid_0_4 <= _GEN_76408;
      end
    end else begin
      flow_entry_valid_0_4 <= _GEN_76408;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Vlflowqueue.scala 250:35]
      flow_entry_valid_0_5 <= 1'h0; // @[Vlflowqueue.scala 251:{44,44}]
    end else if (_T_90) begin
      if (5'h5 == deqPtr_0_value) begin
        flow_entry_valid_0_5 <= 1'h0;
      end else begin
        flow_entry_valid_0_5 <= _GEN_76409;
      end
    end else begin
      flow_entry_valid_0_5 <= _GEN_76409;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Vlflowqueue.scala 250:35]
      flow_entry_valid_0_6 <= 1'h0; // @[Vlflowqueue.scala 251:{44,44}]
    end else if (_T_90) begin
      if (5'h6 == deqPtr_0_value) begin
        flow_entry_valid_0_6 <= 1'h0;
      end else begin
        flow_entry_valid_0_6 <= _GEN_76410;
      end
    end else begin
      flow_entry_valid_0_6 <= _GEN_76410;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Vlflowqueue.scala 250:35]
      flow_entry_valid_0_7 <= 1'h0; // @[Vlflowqueue.scala 251:{44,44}]
    end else if (_T_90) begin
      if (5'h7 == deqPtr_0_value) begin
        flow_entry_valid_0_7 <= 1'h0;
      end else begin
        flow_entry_valid_0_7 <= _GEN_76411;
      end
    end else begin
      flow_entry_valid_0_7 <= _GEN_76411;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Vlflowqueue.scala 250:35]
      flow_entry_valid_0_8 <= 1'h0; // @[Vlflowqueue.scala 251:{44,44}]
    end else if (_T_90) begin
      if (5'h8 == deqPtr_0_value) begin
        flow_entry_valid_0_8 <= 1'h0;
      end else begin
        flow_entry_valid_0_8 <= _GEN_76412;
      end
    end else begin
      flow_entry_valid_0_8 <= _GEN_76412;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Vlflowqueue.scala 250:35]
      flow_entry_valid_0_9 <= 1'h0; // @[Vlflowqueue.scala 251:{44,44}]
    end else if (_T_90) begin
      if (5'h9 == deqPtr_0_value) begin
        flow_entry_valid_0_9 <= 1'h0;
      end else begin
        flow_entry_valid_0_9 <= _GEN_76413;
      end
    end else begin
      flow_entry_valid_0_9 <= _GEN_76413;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Vlflowqueue.scala 250:35]
      flow_entry_valid_0_10 <= 1'h0; // @[Vlflowqueue.scala 251:{44,44}]
    end else if (_T_90) begin
      if (5'ha == deqPtr_0_value) begin
        flow_entry_valid_0_10 <= 1'h0;
      end else begin
        flow_entry_valid_0_10 <= _GEN_76414;
      end
    end else begin
      flow_entry_valid_0_10 <= _GEN_76414;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Vlflowqueue.scala 250:35]
      flow_entry_valid_0_11 <= 1'h0; // @[Vlflowqueue.scala 251:{44,44}]
    end else if (_T_90) begin
      if (5'hb == deqPtr_0_value) begin
        flow_entry_valid_0_11 <= 1'h0;
      end else begin
        flow_entry_valid_0_11 <= _GEN_76415;
      end
    end else begin
      flow_entry_valid_0_11 <= _GEN_76415;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Vlflowqueue.scala 250:35]
      flow_entry_valid_0_12 <= 1'h0; // @[Vlflowqueue.scala 251:{44,44}]
    end else if (_T_90) begin
      if (5'hc == deqPtr_0_value) begin
        flow_entry_valid_0_12 <= 1'h0;
      end else begin
        flow_entry_valid_0_12 <= _GEN_76416;
      end
    end else begin
      flow_entry_valid_0_12 <= _GEN_76416;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Vlflowqueue.scala 250:35]
      flow_entry_valid_0_13 <= 1'h0; // @[Vlflowqueue.scala 251:{44,44}]
    end else if (_T_90) begin
      if (5'hd == deqPtr_0_value) begin
        flow_entry_valid_0_13 <= 1'h0;
      end else begin
        flow_entry_valid_0_13 <= _GEN_76417;
      end
    end else begin
      flow_entry_valid_0_13 <= _GEN_76417;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Vlflowqueue.scala 250:35]
      flow_entry_valid_0_14 <= 1'h0; // @[Vlflowqueue.scala 251:{44,44}]
    end else if (_T_90) begin
      if (5'he == deqPtr_0_value) begin
        flow_entry_valid_0_14 <= 1'h0;
      end else begin
        flow_entry_valid_0_14 <= _GEN_76418;
      end
    end else begin
      flow_entry_valid_0_14 <= _GEN_76418;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Vlflowqueue.scala 250:35]
      flow_entry_valid_0_15 <= 1'h0; // @[Vlflowqueue.scala 251:{44,44}]
    end else if (_T_90) begin
      if (5'hf == deqPtr_0_value) begin
        flow_entry_valid_0_15 <= 1'h0;
      end else begin
        flow_entry_valid_0_15 <= _GEN_76419;
      end
    end else begin
      flow_entry_valid_0_15 <= _GEN_76419;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Vlflowqueue.scala 250:35]
      flow_entry_valid_0_16 <= 1'h0; // @[Vlflowqueue.scala 251:{44,44}]
    end else if (_T_90) begin
      if (5'h10 == deqPtr_0_value) begin
        flow_entry_valid_0_16 <= 1'h0;
      end else begin
        flow_entry_valid_0_16 <= _GEN_76420;
      end
    end else begin
      flow_entry_valid_0_16 <= _GEN_76420;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Vlflowqueue.scala 250:35]
      flow_entry_valid_0_17 <= 1'h0; // @[Vlflowqueue.scala 251:{44,44}]
    end else if (_T_90) begin
      if (5'h11 == deqPtr_0_value) begin
        flow_entry_valid_0_17 <= 1'h0;
      end else begin
        flow_entry_valid_0_17 <= _GEN_76421;
      end
    end else begin
      flow_entry_valid_0_17 <= _GEN_76421;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Vlflowqueue.scala 250:35]
      flow_entry_valid_0_18 <= 1'h0; // @[Vlflowqueue.scala 251:{44,44}]
    end else if (_T_90) begin
      if (5'h12 == deqPtr_0_value) begin
        flow_entry_valid_0_18 <= 1'h0;
      end else begin
        flow_entry_valid_0_18 <= _GEN_76422;
      end
    end else begin
      flow_entry_valid_0_18 <= _GEN_76422;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Vlflowqueue.scala 250:35]
      flow_entry_valid_0_19 <= 1'h0; // @[Vlflowqueue.scala 251:{44,44}]
    end else if (_T_90) begin
      if (5'h13 == deqPtr_0_value) begin
        flow_entry_valid_0_19 <= 1'h0;
      end else begin
        flow_entry_valid_0_19 <= _GEN_76423;
      end
    end else begin
      flow_entry_valid_0_19 <= _GEN_76423;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Vlflowqueue.scala 250:35]
      flow_entry_valid_0_20 <= 1'h0; // @[Vlflowqueue.scala 251:{44,44}]
    end else if (_T_90) begin
      if (5'h14 == deqPtr_0_value) begin
        flow_entry_valid_0_20 <= 1'h0;
      end else begin
        flow_entry_valid_0_20 <= _GEN_76424;
      end
    end else begin
      flow_entry_valid_0_20 <= _GEN_76424;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Vlflowqueue.scala 250:35]
      flow_entry_valid_0_21 <= 1'h0; // @[Vlflowqueue.scala 251:{44,44}]
    end else if (_T_90) begin
      if (5'h15 == deqPtr_0_value) begin
        flow_entry_valid_0_21 <= 1'h0;
      end else begin
        flow_entry_valid_0_21 <= _GEN_76425;
      end
    end else begin
      flow_entry_valid_0_21 <= _GEN_76425;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Vlflowqueue.scala 250:35]
      flow_entry_valid_0_22 <= 1'h0; // @[Vlflowqueue.scala 251:{44,44}]
    end else if (_T_90) begin
      if (5'h16 == deqPtr_0_value) begin
        flow_entry_valid_0_22 <= 1'h0;
      end else begin
        flow_entry_valid_0_22 <= _GEN_76426;
      end
    end else begin
      flow_entry_valid_0_22 <= _GEN_76426;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Vlflowqueue.scala 250:35]
      flow_entry_valid_0_23 <= 1'h0; // @[Vlflowqueue.scala 251:{44,44}]
    end else if (_T_90) begin
      if (5'h17 == deqPtr_0_value) begin
        flow_entry_valid_0_23 <= 1'h0;
      end else begin
        flow_entry_valid_0_23 <= _GEN_76427;
      end
    end else begin
      flow_entry_valid_0_23 <= _GEN_76427;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Vlflowqueue.scala 250:35]
      flow_entry_valid_0_24 <= 1'h0; // @[Vlflowqueue.scala 251:{44,44}]
    end else if (_T_90) begin
      if (5'h18 == deqPtr_0_value) begin
        flow_entry_valid_0_24 <= 1'h0;
      end else begin
        flow_entry_valid_0_24 <= _GEN_76428;
      end
    end else begin
      flow_entry_valid_0_24 <= _GEN_76428;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Vlflowqueue.scala 250:35]
      flow_entry_valid_0_25 <= 1'h0; // @[Vlflowqueue.scala 251:{44,44}]
    end else if (_T_90) begin
      if (5'h19 == deqPtr_0_value) begin
        flow_entry_valid_0_25 <= 1'h0;
      end else begin
        flow_entry_valid_0_25 <= _GEN_76429;
      end
    end else begin
      flow_entry_valid_0_25 <= _GEN_76429;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Vlflowqueue.scala 250:35]
      flow_entry_valid_0_26 <= 1'h0; // @[Vlflowqueue.scala 251:{44,44}]
    end else if (_T_90) begin
      if (5'h1a == deqPtr_0_value) begin
        flow_entry_valid_0_26 <= 1'h0;
      end else begin
        flow_entry_valid_0_26 <= _GEN_76430;
      end
    end else begin
      flow_entry_valid_0_26 <= _GEN_76430;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Vlflowqueue.scala 250:35]
      flow_entry_valid_0_27 <= 1'h0; // @[Vlflowqueue.scala 251:{44,44}]
    end else if (_T_90) begin
      if (5'h1b == deqPtr_0_value) begin
        flow_entry_valid_0_27 <= 1'h0;
      end else begin
        flow_entry_valid_0_27 <= _GEN_76431;
      end
    end else begin
      flow_entry_valid_0_27 <= _GEN_76431;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Vlflowqueue.scala 250:35]
      flow_entry_valid_0_28 <= 1'h0; // @[Vlflowqueue.scala 251:{44,44}]
    end else if (_T_90) begin
      if (5'h1c == deqPtr_0_value) begin
        flow_entry_valid_0_28 <= 1'h0;
      end else begin
        flow_entry_valid_0_28 <= _GEN_76432;
      end
    end else begin
      flow_entry_valid_0_28 <= _GEN_76432;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Vlflowqueue.scala 250:35]
      flow_entry_valid_0_29 <= 1'h0; // @[Vlflowqueue.scala 251:{44,44}]
    end else if (_T_90) begin
      if (5'h1d == deqPtr_0_value) begin
        flow_entry_valid_0_29 <= 1'h0;
      end else begin
        flow_entry_valid_0_29 <= _GEN_76433;
      end
    end else begin
      flow_entry_valid_0_29 <= _GEN_76433;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Vlflowqueue.scala 250:35]
      flow_entry_valid_0_30 <= 1'h0; // @[Vlflowqueue.scala 251:{44,44}]
    end else if (_T_90) begin
      if (5'h1e == deqPtr_0_value) begin
        flow_entry_valid_0_30 <= 1'h0;
      end else begin
        flow_entry_valid_0_30 <= _GEN_76434;
      end
    end else begin
      flow_entry_valid_0_30 <= _GEN_76434;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Vlflowqueue.scala 250:35]
      flow_entry_valid_0_31 <= 1'h0; // @[Vlflowqueue.scala 251:{44,44}]
    end else if (_T_90) begin
      if (5'h1f == deqPtr_0_value) begin
        flow_entry_valid_0_31 <= 1'h0;
      end else begin
        flow_entry_valid_0_31 <= _GEN_76435;
      end
    end else begin
      flow_entry_valid_0_31 <= _GEN_76435;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Vlflowqueue.scala 250:35]
      flow_entry_valid_1_0 <= 1'h0; // @[Vlflowqueue.scala 251:{44,44}]
    end else if (_T_91) begin
      if (5'h0 == deqPtr_1_value) begin
        flow_entry_valid_1_0 <= 1'h0;
      end else begin
        flow_entry_valid_1_0 <= _GEN_156649;
      end
    end else begin
      flow_entry_valid_1_0 <= _GEN_156649;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Vlflowqueue.scala 250:35]
      flow_entry_valid_1_1 <= 1'h0; // @[Vlflowqueue.scala 251:{44,44}]
    end else if (_T_91) begin
      if (5'h1 == deqPtr_1_value) begin
        flow_entry_valid_1_1 <= 1'h0;
      end else begin
        flow_entry_valid_1_1 <= _GEN_156650;
      end
    end else begin
      flow_entry_valid_1_1 <= _GEN_156650;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Vlflowqueue.scala 250:35]
      flow_entry_valid_1_2 <= 1'h0; // @[Vlflowqueue.scala 251:{44,44}]
    end else if (_T_91) begin
      if (5'h2 == deqPtr_1_value) begin
        flow_entry_valid_1_2 <= 1'h0;
      end else begin
        flow_entry_valid_1_2 <= _GEN_156651;
      end
    end else begin
      flow_entry_valid_1_2 <= _GEN_156651;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Vlflowqueue.scala 250:35]
      flow_entry_valid_1_3 <= 1'h0; // @[Vlflowqueue.scala 251:{44,44}]
    end else if (_T_91) begin
      if (5'h3 == deqPtr_1_value) begin
        flow_entry_valid_1_3 <= 1'h0;
      end else begin
        flow_entry_valid_1_3 <= _GEN_156652;
      end
    end else begin
      flow_entry_valid_1_3 <= _GEN_156652;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Vlflowqueue.scala 250:35]
      flow_entry_valid_1_4 <= 1'h0; // @[Vlflowqueue.scala 251:{44,44}]
    end else if (_T_91) begin
      if (5'h4 == deqPtr_1_value) begin
        flow_entry_valid_1_4 <= 1'h0;
      end else begin
        flow_entry_valid_1_4 <= _GEN_156653;
      end
    end else begin
      flow_entry_valid_1_4 <= _GEN_156653;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Vlflowqueue.scala 250:35]
      flow_entry_valid_1_5 <= 1'h0; // @[Vlflowqueue.scala 251:{44,44}]
    end else if (_T_91) begin
      if (5'h5 == deqPtr_1_value) begin
        flow_entry_valid_1_5 <= 1'h0;
      end else begin
        flow_entry_valid_1_5 <= _GEN_156654;
      end
    end else begin
      flow_entry_valid_1_5 <= _GEN_156654;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Vlflowqueue.scala 250:35]
      flow_entry_valid_1_6 <= 1'h0; // @[Vlflowqueue.scala 251:{44,44}]
    end else if (_T_91) begin
      if (5'h6 == deqPtr_1_value) begin
        flow_entry_valid_1_6 <= 1'h0;
      end else begin
        flow_entry_valid_1_6 <= _GEN_156655;
      end
    end else begin
      flow_entry_valid_1_6 <= _GEN_156655;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Vlflowqueue.scala 250:35]
      flow_entry_valid_1_7 <= 1'h0; // @[Vlflowqueue.scala 251:{44,44}]
    end else if (_T_91) begin
      if (5'h7 == deqPtr_1_value) begin
        flow_entry_valid_1_7 <= 1'h0;
      end else begin
        flow_entry_valid_1_7 <= _GEN_156656;
      end
    end else begin
      flow_entry_valid_1_7 <= _GEN_156656;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Vlflowqueue.scala 250:35]
      flow_entry_valid_1_8 <= 1'h0; // @[Vlflowqueue.scala 251:{44,44}]
    end else if (_T_91) begin
      if (5'h8 == deqPtr_1_value) begin
        flow_entry_valid_1_8 <= 1'h0;
      end else begin
        flow_entry_valid_1_8 <= _GEN_156657;
      end
    end else begin
      flow_entry_valid_1_8 <= _GEN_156657;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Vlflowqueue.scala 250:35]
      flow_entry_valid_1_9 <= 1'h0; // @[Vlflowqueue.scala 251:{44,44}]
    end else if (_T_91) begin
      if (5'h9 == deqPtr_1_value) begin
        flow_entry_valid_1_9 <= 1'h0;
      end else begin
        flow_entry_valid_1_9 <= _GEN_156658;
      end
    end else begin
      flow_entry_valid_1_9 <= _GEN_156658;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Vlflowqueue.scala 250:35]
      flow_entry_valid_1_10 <= 1'h0; // @[Vlflowqueue.scala 251:{44,44}]
    end else if (_T_91) begin
      if (5'ha == deqPtr_1_value) begin
        flow_entry_valid_1_10 <= 1'h0;
      end else begin
        flow_entry_valid_1_10 <= _GEN_156659;
      end
    end else begin
      flow_entry_valid_1_10 <= _GEN_156659;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Vlflowqueue.scala 250:35]
      flow_entry_valid_1_11 <= 1'h0; // @[Vlflowqueue.scala 251:{44,44}]
    end else if (_T_91) begin
      if (5'hb == deqPtr_1_value) begin
        flow_entry_valid_1_11 <= 1'h0;
      end else begin
        flow_entry_valid_1_11 <= _GEN_156660;
      end
    end else begin
      flow_entry_valid_1_11 <= _GEN_156660;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Vlflowqueue.scala 250:35]
      flow_entry_valid_1_12 <= 1'h0; // @[Vlflowqueue.scala 251:{44,44}]
    end else if (_T_91) begin
      if (5'hc == deqPtr_1_value) begin
        flow_entry_valid_1_12 <= 1'h0;
      end else begin
        flow_entry_valid_1_12 <= _GEN_156661;
      end
    end else begin
      flow_entry_valid_1_12 <= _GEN_156661;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Vlflowqueue.scala 250:35]
      flow_entry_valid_1_13 <= 1'h0; // @[Vlflowqueue.scala 251:{44,44}]
    end else if (_T_91) begin
      if (5'hd == deqPtr_1_value) begin
        flow_entry_valid_1_13 <= 1'h0;
      end else begin
        flow_entry_valid_1_13 <= _GEN_156662;
      end
    end else begin
      flow_entry_valid_1_13 <= _GEN_156662;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Vlflowqueue.scala 250:35]
      flow_entry_valid_1_14 <= 1'h0; // @[Vlflowqueue.scala 251:{44,44}]
    end else if (_T_91) begin
      if (5'he == deqPtr_1_value) begin
        flow_entry_valid_1_14 <= 1'h0;
      end else begin
        flow_entry_valid_1_14 <= _GEN_156663;
      end
    end else begin
      flow_entry_valid_1_14 <= _GEN_156663;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Vlflowqueue.scala 250:35]
      flow_entry_valid_1_15 <= 1'h0; // @[Vlflowqueue.scala 251:{44,44}]
    end else if (_T_91) begin
      if (5'hf == deqPtr_1_value) begin
        flow_entry_valid_1_15 <= 1'h0;
      end else begin
        flow_entry_valid_1_15 <= _GEN_156664;
      end
    end else begin
      flow_entry_valid_1_15 <= _GEN_156664;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Vlflowqueue.scala 250:35]
      flow_entry_valid_1_16 <= 1'h0; // @[Vlflowqueue.scala 251:{44,44}]
    end else if (_T_91) begin
      if (5'h10 == deqPtr_1_value) begin
        flow_entry_valid_1_16 <= 1'h0;
      end else begin
        flow_entry_valid_1_16 <= _GEN_156665;
      end
    end else begin
      flow_entry_valid_1_16 <= _GEN_156665;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Vlflowqueue.scala 250:35]
      flow_entry_valid_1_17 <= 1'h0; // @[Vlflowqueue.scala 251:{44,44}]
    end else if (_T_91) begin
      if (5'h11 == deqPtr_1_value) begin
        flow_entry_valid_1_17 <= 1'h0;
      end else begin
        flow_entry_valid_1_17 <= _GEN_156666;
      end
    end else begin
      flow_entry_valid_1_17 <= _GEN_156666;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Vlflowqueue.scala 250:35]
      flow_entry_valid_1_18 <= 1'h0; // @[Vlflowqueue.scala 251:{44,44}]
    end else if (_T_91) begin
      if (5'h12 == deqPtr_1_value) begin
        flow_entry_valid_1_18 <= 1'h0;
      end else begin
        flow_entry_valid_1_18 <= _GEN_156667;
      end
    end else begin
      flow_entry_valid_1_18 <= _GEN_156667;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Vlflowqueue.scala 250:35]
      flow_entry_valid_1_19 <= 1'h0; // @[Vlflowqueue.scala 251:{44,44}]
    end else if (_T_91) begin
      if (5'h13 == deqPtr_1_value) begin
        flow_entry_valid_1_19 <= 1'h0;
      end else begin
        flow_entry_valid_1_19 <= _GEN_156668;
      end
    end else begin
      flow_entry_valid_1_19 <= _GEN_156668;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Vlflowqueue.scala 250:35]
      flow_entry_valid_1_20 <= 1'h0; // @[Vlflowqueue.scala 251:{44,44}]
    end else if (_T_91) begin
      if (5'h14 == deqPtr_1_value) begin
        flow_entry_valid_1_20 <= 1'h0;
      end else begin
        flow_entry_valid_1_20 <= _GEN_156669;
      end
    end else begin
      flow_entry_valid_1_20 <= _GEN_156669;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Vlflowqueue.scala 250:35]
      flow_entry_valid_1_21 <= 1'h0; // @[Vlflowqueue.scala 251:{44,44}]
    end else if (_T_91) begin
      if (5'h15 == deqPtr_1_value) begin
        flow_entry_valid_1_21 <= 1'h0;
      end else begin
        flow_entry_valid_1_21 <= _GEN_156670;
      end
    end else begin
      flow_entry_valid_1_21 <= _GEN_156670;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Vlflowqueue.scala 250:35]
      flow_entry_valid_1_22 <= 1'h0; // @[Vlflowqueue.scala 251:{44,44}]
    end else if (_T_91) begin
      if (5'h16 == deqPtr_1_value) begin
        flow_entry_valid_1_22 <= 1'h0;
      end else begin
        flow_entry_valid_1_22 <= _GEN_156671;
      end
    end else begin
      flow_entry_valid_1_22 <= _GEN_156671;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Vlflowqueue.scala 250:35]
      flow_entry_valid_1_23 <= 1'h0; // @[Vlflowqueue.scala 251:{44,44}]
    end else if (_T_91) begin
      if (5'h17 == deqPtr_1_value) begin
        flow_entry_valid_1_23 <= 1'h0;
      end else begin
        flow_entry_valid_1_23 <= _GEN_156672;
      end
    end else begin
      flow_entry_valid_1_23 <= _GEN_156672;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Vlflowqueue.scala 250:35]
      flow_entry_valid_1_24 <= 1'h0; // @[Vlflowqueue.scala 251:{44,44}]
    end else if (_T_91) begin
      if (5'h18 == deqPtr_1_value) begin
        flow_entry_valid_1_24 <= 1'h0;
      end else begin
        flow_entry_valid_1_24 <= _GEN_156673;
      end
    end else begin
      flow_entry_valid_1_24 <= _GEN_156673;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Vlflowqueue.scala 250:35]
      flow_entry_valid_1_25 <= 1'h0; // @[Vlflowqueue.scala 251:{44,44}]
    end else if (_T_91) begin
      if (5'h19 == deqPtr_1_value) begin
        flow_entry_valid_1_25 <= 1'h0;
      end else begin
        flow_entry_valid_1_25 <= _GEN_156674;
      end
    end else begin
      flow_entry_valid_1_25 <= _GEN_156674;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Vlflowqueue.scala 250:35]
      flow_entry_valid_1_26 <= 1'h0; // @[Vlflowqueue.scala 251:{44,44}]
    end else if (_T_91) begin
      if (5'h1a == deqPtr_1_value) begin
        flow_entry_valid_1_26 <= 1'h0;
      end else begin
        flow_entry_valid_1_26 <= _GEN_156675;
      end
    end else begin
      flow_entry_valid_1_26 <= _GEN_156675;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Vlflowqueue.scala 250:35]
      flow_entry_valid_1_27 <= 1'h0; // @[Vlflowqueue.scala 251:{44,44}]
    end else if (_T_91) begin
      if (5'h1b == deqPtr_1_value) begin
        flow_entry_valid_1_27 <= 1'h0;
      end else begin
        flow_entry_valid_1_27 <= _GEN_156676;
      end
    end else begin
      flow_entry_valid_1_27 <= _GEN_156676;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Vlflowqueue.scala 250:35]
      flow_entry_valid_1_28 <= 1'h0; // @[Vlflowqueue.scala 251:{44,44}]
    end else if (_T_91) begin
      if (5'h1c == deqPtr_1_value) begin
        flow_entry_valid_1_28 <= 1'h0;
      end else begin
        flow_entry_valid_1_28 <= _GEN_156677;
      end
    end else begin
      flow_entry_valid_1_28 <= _GEN_156677;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Vlflowqueue.scala 250:35]
      flow_entry_valid_1_29 <= 1'h0; // @[Vlflowqueue.scala 251:{44,44}]
    end else if (_T_91) begin
      if (5'h1d == deqPtr_1_value) begin
        flow_entry_valid_1_29 <= 1'h0;
      end else begin
        flow_entry_valid_1_29 <= _GEN_156678;
      end
    end else begin
      flow_entry_valid_1_29 <= _GEN_156678;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Vlflowqueue.scala 250:35]
      flow_entry_valid_1_30 <= 1'h0; // @[Vlflowqueue.scala 251:{44,44}]
    end else if (_T_91) begin
      if (5'h1e == deqPtr_1_value) begin
        flow_entry_valid_1_30 <= 1'h0;
      end else begin
        flow_entry_valid_1_30 <= _GEN_156679;
      end
    end else begin
      flow_entry_valid_1_30 <= _GEN_156679;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Vlflowqueue.scala 250:35]
      flow_entry_valid_1_31 <= 1'h0; // @[Vlflowqueue.scala 251:{44,44}]
    end else if (_T_91) begin
      if (5'h1f == deqPtr_1_value) begin
        flow_entry_valid_1_31 <= 1'h0;
      end else begin
        flow_entry_valid_1_31 <= _GEN_156680;
      end
    end else begin
      flow_entry_valid_1_31 <= _GEN_156680;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Vlflowqueue.scala 178:40]
      enqPtr_0_value <= 5'h0;
    end else begin
      enqPtr_0_value <= enqPtr_0_value + _GEN_161415;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Vlflowqueue.scala 178:40]
      enqPtr_1_value <= 5'h0;
    end else begin
      enqPtr_1_value <= enqPtr_1_value + _GEN_161417;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Vlflowqueue.scala 250:35]
      deqPtr_0_flag <= 1'h0; // @[Vlflowqueue.scala 252:17]
    end else if (_T_90) begin // @[Vlflowqueue.scala 172:23]
      deqPtr_0_flag <= deqPtr_0_new_ptr_flag;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Vlflowqueue.scala 250:35]
      deqPtr_0_value <= 5'h0; // @[Vlflowqueue.scala 252:17]
    end else if (_T_90) begin // @[Vlflowqueue.scala 172:23]
      deqPtr_0_value <= deqPtr_0_new_ptr_value;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Vlflowqueue.scala 250:35]
      deqPtr_1_flag <= 1'h0; // @[Vlflowqueue.scala 252:17]
    end else if (_T_91) begin // @[Vlflowqueue.scala 172:23]
      deqPtr_1_flag <= deqPtr_1_new_ptr_flag;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Vlflowqueue.scala 250:35]
      deqPtr_1_value <= 5'h0; // @[Vlflowqueue.scala 252:17]
    end else if (_T_91) begin // @[Vlflowqueue.scala 172:23]
      deqPtr_1_value <= deqPtr_1_new_ptr_value;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  flow_entry_0_0_uop_robIdx_value = _RAND_0[4:0];
  _RAND_1 = {2{`RANDOM}};
  flow_entry_0_0_vaddr = _RAND_1[38:0];
  _RAND_2 = {1{`RANDOM}};
  flow_entry_0_1_uop_robIdx_value = _RAND_2[4:0];
  _RAND_3 = {2{`RANDOM}};
  flow_entry_0_1_vaddr = _RAND_3[38:0];
  _RAND_4 = {1{`RANDOM}};
  flow_entry_0_2_uop_robIdx_value = _RAND_4[4:0];
  _RAND_5 = {2{`RANDOM}};
  flow_entry_0_2_vaddr = _RAND_5[38:0];
  _RAND_6 = {1{`RANDOM}};
  flow_entry_0_3_uop_robIdx_value = _RAND_6[4:0];
  _RAND_7 = {2{`RANDOM}};
  flow_entry_0_3_vaddr = _RAND_7[38:0];
  _RAND_8 = {1{`RANDOM}};
  flow_entry_0_4_uop_robIdx_value = _RAND_8[4:0];
  _RAND_9 = {2{`RANDOM}};
  flow_entry_0_4_vaddr = _RAND_9[38:0];
  _RAND_10 = {1{`RANDOM}};
  flow_entry_0_5_uop_robIdx_value = _RAND_10[4:0];
  _RAND_11 = {2{`RANDOM}};
  flow_entry_0_5_vaddr = _RAND_11[38:0];
  _RAND_12 = {1{`RANDOM}};
  flow_entry_0_6_uop_robIdx_value = _RAND_12[4:0];
  _RAND_13 = {2{`RANDOM}};
  flow_entry_0_6_vaddr = _RAND_13[38:0];
  _RAND_14 = {1{`RANDOM}};
  flow_entry_0_7_uop_robIdx_value = _RAND_14[4:0];
  _RAND_15 = {2{`RANDOM}};
  flow_entry_0_7_vaddr = _RAND_15[38:0];
  _RAND_16 = {1{`RANDOM}};
  flow_entry_0_8_uop_robIdx_value = _RAND_16[4:0];
  _RAND_17 = {2{`RANDOM}};
  flow_entry_0_8_vaddr = _RAND_17[38:0];
  _RAND_18 = {1{`RANDOM}};
  flow_entry_0_9_uop_robIdx_value = _RAND_18[4:0];
  _RAND_19 = {2{`RANDOM}};
  flow_entry_0_9_vaddr = _RAND_19[38:0];
  _RAND_20 = {1{`RANDOM}};
  flow_entry_0_10_uop_robIdx_value = _RAND_20[4:0];
  _RAND_21 = {2{`RANDOM}};
  flow_entry_0_10_vaddr = _RAND_21[38:0];
  _RAND_22 = {1{`RANDOM}};
  flow_entry_0_11_uop_robIdx_value = _RAND_22[4:0];
  _RAND_23 = {2{`RANDOM}};
  flow_entry_0_11_vaddr = _RAND_23[38:0];
  _RAND_24 = {1{`RANDOM}};
  flow_entry_0_12_uop_robIdx_value = _RAND_24[4:0];
  _RAND_25 = {2{`RANDOM}};
  flow_entry_0_12_vaddr = _RAND_25[38:0];
  _RAND_26 = {1{`RANDOM}};
  flow_entry_0_13_uop_robIdx_value = _RAND_26[4:0];
  _RAND_27 = {2{`RANDOM}};
  flow_entry_0_13_vaddr = _RAND_27[38:0];
  _RAND_28 = {1{`RANDOM}};
  flow_entry_0_14_uop_robIdx_value = _RAND_28[4:0];
  _RAND_29 = {2{`RANDOM}};
  flow_entry_0_14_vaddr = _RAND_29[38:0];
  _RAND_30 = {1{`RANDOM}};
  flow_entry_0_15_uop_robIdx_value = _RAND_30[4:0];
  _RAND_31 = {2{`RANDOM}};
  flow_entry_0_15_vaddr = _RAND_31[38:0];
  _RAND_32 = {1{`RANDOM}};
  flow_entry_0_16_uop_robIdx_value = _RAND_32[4:0];
  _RAND_33 = {2{`RANDOM}};
  flow_entry_0_16_vaddr = _RAND_33[38:0];
  _RAND_34 = {1{`RANDOM}};
  flow_entry_0_17_uop_robIdx_value = _RAND_34[4:0];
  _RAND_35 = {2{`RANDOM}};
  flow_entry_0_17_vaddr = _RAND_35[38:0];
  _RAND_36 = {1{`RANDOM}};
  flow_entry_0_18_uop_robIdx_value = _RAND_36[4:0];
  _RAND_37 = {2{`RANDOM}};
  flow_entry_0_18_vaddr = _RAND_37[38:0];
  _RAND_38 = {1{`RANDOM}};
  flow_entry_0_19_uop_robIdx_value = _RAND_38[4:0];
  _RAND_39 = {2{`RANDOM}};
  flow_entry_0_19_vaddr = _RAND_39[38:0];
  _RAND_40 = {1{`RANDOM}};
  flow_entry_0_20_uop_robIdx_value = _RAND_40[4:0];
  _RAND_41 = {2{`RANDOM}};
  flow_entry_0_20_vaddr = _RAND_41[38:0];
  _RAND_42 = {1{`RANDOM}};
  flow_entry_0_21_uop_robIdx_value = _RAND_42[4:0];
  _RAND_43 = {2{`RANDOM}};
  flow_entry_0_21_vaddr = _RAND_43[38:0];
  _RAND_44 = {1{`RANDOM}};
  flow_entry_0_22_uop_robIdx_value = _RAND_44[4:0];
  _RAND_45 = {2{`RANDOM}};
  flow_entry_0_22_vaddr = _RAND_45[38:0];
  _RAND_46 = {1{`RANDOM}};
  flow_entry_0_23_uop_robIdx_value = _RAND_46[4:0];
  _RAND_47 = {2{`RANDOM}};
  flow_entry_0_23_vaddr = _RAND_47[38:0];
  _RAND_48 = {1{`RANDOM}};
  flow_entry_0_24_uop_robIdx_value = _RAND_48[4:0];
  _RAND_49 = {2{`RANDOM}};
  flow_entry_0_24_vaddr = _RAND_49[38:0];
  _RAND_50 = {1{`RANDOM}};
  flow_entry_0_25_uop_robIdx_value = _RAND_50[4:0];
  _RAND_51 = {2{`RANDOM}};
  flow_entry_0_25_vaddr = _RAND_51[38:0];
  _RAND_52 = {1{`RANDOM}};
  flow_entry_0_26_uop_robIdx_value = _RAND_52[4:0];
  _RAND_53 = {2{`RANDOM}};
  flow_entry_0_26_vaddr = _RAND_53[38:0];
  _RAND_54 = {1{`RANDOM}};
  flow_entry_0_27_uop_robIdx_value = _RAND_54[4:0];
  _RAND_55 = {2{`RANDOM}};
  flow_entry_0_27_vaddr = _RAND_55[38:0];
  _RAND_56 = {1{`RANDOM}};
  flow_entry_0_28_uop_robIdx_value = _RAND_56[4:0];
  _RAND_57 = {2{`RANDOM}};
  flow_entry_0_28_vaddr = _RAND_57[38:0];
  _RAND_58 = {1{`RANDOM}};
  flow_entry_0_29_uop_robIdx_value = _RAND_58[4:0];
  _RAND_59 = {2{`RANDOM}};
  flow_entry_0_29_vaddr = _RAND_59[38:0];
  _RAND_60 = {1{`RANDOM}};
  flow_entry_0_30_uop_robIdx_value = _RAND_60[4:0];
  _RAND_61 = {2{`RANDOM}};
  flow_entry_0_30_vaddr = _RAND_61[38:0];
  _RAND_62 = {1{`RANDOM}};
  flow_entry_0_31_uop_robIdx_value = _RAND_62[4:0];
  _RAND_63 = {2{`RANDOM}};
  flow_entry_0_31_vaddr = _RAND_63[38:0];
  _RAND_64 = {1{`RANDOM}};
  flow_entry_1_0_uop_robIdx_value = _RAND_64[4:0];
  _RAND_65 = {2{`RANDOM}};
  flow_entry_1_0_vaddr = _RAND_65[38:0];
  _RAND_66 = {1{`RANDOM}};
  flow_entry_1_1_uop_robIdx_value = _RAND_66[4:0];
  _RAND_67 = {2{`RANDOM}};
  flow_entry_1_1_vaddr = _RAND_67[38:0];
  _RAND_68 = {1{`RANDOM}};
  flow_entry_1_2_uop_robIdx_value = _RAND_68[4:0];
  _RAND_69 = {2{`RANDOM}};
  flow_entry_1_2_vaddr = _RAND_69[38:0];
  _RAND_70 = {1{`RANDOM}};
  flow_entry_1_3_uop_robIdx_value = _RAND_70[4:0];
  _RAND_71 = {2{`RANDOM}};
  flow_entry_1_3_vaddr = _RAND_71[38:0];
  _RAND_72 = {1{`RANDOM}};
  flow_entry_1_4_uop_robIdx_value = _RAND_72[4:0];
  _RAND_73 = {2{`RANDOM}};
  flow_entry_1_4_vaddr = _RAND_73[38:0];
  _RAND_74 = {1{`RANDOM}};
  flow_entry_1_5_uop_robIdx_value = _RAND_74[4:0];
  _RAND_75 = {2{`RANDOM}};
  flow_entry_1_5_vaddr = _RAND_75[38:0];
  _RAND_76 = {1{`RANDOM}};
  flow_entry_1_6_uop_robIdx_value = _RAND_76[4:0];
  _RAND_77 = {2{`RANDOM}};
  flow_entry_1_6_vaddr = _RAND_77[38:0];
  _RAND_78 = {1{`RANDOM}};
  flow_entry_1_7_uop_robIdx_value = _RAND_78[4:0];
  _RAND_79 = {2{`RANDOM}};
  flow_entry_1_7_vaddr = _RAND_79[38:0];
  _RAND_80 = {1{`RANDOM}};
  flow_entry_1_8_uop_robIdx_value = _RAND_80[4:0];
  _RAND_81 = {2{`RANDOM}};
  flow_entry_1_8_vaddr = _RAND_81[38:0];
  _RAND_82 = {1{`RANDOM}};
  flow_entry_1_9_uop_robIdx_value = _RAND_82[4:0];
  _RAND_83 = {2{`RANDOM}};
  flow_entry_1_9_vaddr = _RAND_83[38:0];
  _RAND_84 = {1{`RANDOM}};
  flow_entry_1_10_uop_robIdx_value = _RAND_84[4:0];
  _RAND_85 = {2{`RANDOM}};
  flow_entry_1_10_vaddr = _RAND_85[38:0];
  _RAND_86 = {1{`RANDOM}};
  flow_entry_1_11_uop_robIdx_value = _RAND_86[4:0];
  _RAND_87 = {2{`RANDOM}};
  flow_entry_1_11_vaddr = _RAND_87[38:0];
  _RAND_88 = {1{`RANDOM}};
  flow_entry_1_12_uop_robIdx_value = _RAND_88[4:0];
  _RAND_89 = {2{`RANDOM}};
  flow_entry_1_12_vaddr = _RAND_89[38:0];
  _RAND_90 = {1{`RANDOM}};
  flow_entry_1_13_uop_robIdx_value = _RAND_90[4:0];
  _RAND_91 = {2{`RANDOM}};
  flow_entry_1_13_vaddr = _RAND_91[38:0];
  _RAND_92 = {1{`RANDOM}};
  flow_entry_1_14_uop_robIdx_value = _RAND_92[4:0];
  _RAND_93 = {2{`RANDOM}};
  flow_entry_1_14_vaddr = _RAND_93[38:0];
  _RAND_94 = {1{`RANDOM}};
  flow_entry_1_15_uop_robIdx_value = _RAND_94[4:0];
  _RAND_95 = {2{`RANDOM}};
  flow_entry_1_15_vaddr = _RAND_95[38:0];
  _RAND_96 = {1{`RANDOM}};
  flow_entry_1_16_uop_robIdx_value = _RAND_96[4:0];
  _RAND_97 = {2{`RANDOM}};
  flow_entry_1_16_vaddr = _RAND_97[38:0];
  _RAND_98 = {1{`RANDOM}};
  flow_entry_1_17_uop_robIdx_value = _RAND_98[4:0];
  _RAND_99 = {2{`RANDOM}};
  flow_entry_1_17_vaddr = _RAND_99[38:0];
  _RAND_100 = {1{`RANDOM}};
  flow_entry_1_18_uop_robIdx_value = _RAND_100[4:0];
  _RAND_101 = {2{`RANDOM}};
  flow_entry_1_18_vaddr = _RAND_101[38:0];
  _RAND_102 = {1{`RANDOM}};
  flow_entry_1_19_uop_robIdx_value = _RAND_102[4:0];
  _RAND_103 = {2{`RANDOM}};
  flow_entry_1_19_vaddr = _RAND_103[38:0];
  _RAND_104 = {1{`RANDOM}};
  flow_entry_1_20_uop_robIdx_value = _RAND_104[4:0];
  _RAND_105 = {2{`RANDOM}};
  flow_entry_1_20_vaddr = _RAND_105[38:0];
  _RAND_106 = {1{`RANDOM}};
  flow_entry_1_21_uop_robIdx_value = _RAND_106[4:0];
  _RAND_107 = {2{`RANDOM}};
  flow_entry_1_21_vaddr = _RAND_107[38:0];
  _RAND_108 = {1{`RANDOM}};
  flow_entry_1_22_uop_robIdx_value = _RAND_108[4:0];
  _RAND_109 = {2{`RANDOM}};
  flow_entry_1_22_vaddr = _RAND_109[38:0];
  _RAND_110 = {1{`RANDOM}};
  flow_entry_1_23_uop_robIdx_value = _RAND_110[4:0];
  _RAND_111 = {2{`RANDOM}};
  flow_entry_1_23_vaddr = _RAND_111[38:0];
  _RAND_112 = {1{`RANDOM}};
  flow_entry_1_24_uop_robIdx_value = _RAND_112[4:0];
  _RAND_113 = {2{`RANDOM}};
  flow_entry_1_24_vaddr = _RAND_113[38:0];
  _RAND_114 = {1{`RANDOM}};
  flow_entry_1_25_uop_robIdx_value = _RAND_114[4:0];
  _RAND_115 = {2{`RANDOM}};
  flow_entry_1_25_vaddr = _RAND_115[38:0];
  _RAND_116 = {1{`RANDOM}};
  flow_entry_1_26_uop_robIdx_value = _RAND_116[4:0];
  _RAND_117 = {2{`RANDOM}};
  flow_entry_1_26_vaddr = _RAND_117[38:0];
  _RAND_118 = {1{`RANDOM}};
  flow_entry_1_27_uop_robIdx_value = _RAND_118[4:0];
  _RAND_119 = {2{`RANDOM}};
  flow_entry_1_27_vaddr = _RAND_119[38:0];
  _RAND_120 = {1{`RANDOM}};
  flow_entry_1_28_uop_robIdx_value = _RAND_120[4:0];
  _RAND_121 = {2{`RANDOM}};
  flow_entry_1_28_vaddr = _RAND_121[38:0];
  _RAND_122 = {1{`RANDOM}};
  flow_entry_1_29_uop_robIdx_value = _RAND_122[4:0];
  _RAND_123 = {2{`RANDOM}};
  flow_entry_1_29_vaddr = _RAND_123[38:0];
  _RAND_124 = {1{`RANDOM}};
  flow_entry_1_30_uop_robIdx_value = _RAND_124[4:0];
  _RAND_125 = {2{`RANDOM}};
  flow_entry_1_30_vaddr = _RAND_125[38:0];
  _RAND_126 = {1{`RANDOM}};
  flow_entry_1_31_uop_robIdx_value = _RAND_126[4:0];
  _RAND_127 = {2{`RANDOM}};
  flow_entry_1_31_vaddr = _RAND_127[38:0];
  _RAND_128 = {1{`RANDOM}};
  flow_entry_valid_0_0 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  flow_entry_valid_0_1 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  flow_entry_valid_0_2 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  flow_entry_valid_0_3 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  flow_entry_valid_0_4 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  flow_entry_valid_0_5 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  flow_entry_valid_0_6 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  flow_entry_valid_0_7 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  flow_entry_valid_0_8 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  flow_entry_valid_0_9 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  flow_entry_valid_0_10 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  flow_entry_valid_0_11 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  flow_entry_valid_0_12 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  flow_entry_valid_0_13 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  flow_entry_valid_0_14 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  flow_entry_valid_0_15 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  flow_entry_valid_0_16 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  flow_entry_valid_0_17 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  flow_entry_valid_0_18 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  flow_entry_valid_0_19 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  flow_entry_valid_0_20 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  flow_entry_valid_0_21 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  flow_entry_valid_0_22 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  flow_entry_valid_0_23 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  flow_entry_valid_0_24 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  flow_entry_valid_0_25 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  flow_entry_valid_0_26 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  flow_entry_valid_0_27 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  flow_entry_valid_0_28 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  flow_entry_valid_0_29 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  flow_entry_valid_0_30 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  flow_entry_valid_0_31 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  flow_entry_valid_1_0 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  flow_entry_valid_1_1 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  flow_entry_valid_1_2 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  flow_entry_valid_1_3 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  flow_entry_valid_1_4 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  flow_entry_valid_1_5 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  flow_entry_valid_1_6 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  flow_entry_valid_1_7 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  flow_entry_valid_1_8 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  flow_entry_valid_1_9 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  flow_entry_valid_1_10 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  flow_entry_valid_1_11 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  flow_entry_valid_1_12 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  flow_entry_valid_1_13 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  flow_entry_valid_1_14 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  flow_entry_valid_1_15 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  flow_entry_valid_1_16 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  flow_entry_valid_1_17 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  flow_entry_valid_1_18 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  flow_entry_valid_1_19 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  flow_entry_valid_1_20 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  flow_entry_valid_1_21 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  flow_entry_valid_1_22 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  flow_entry_valid_1_23 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  flow_entry_valid_1_24 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  flow_entry_valid_1_25 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  flow_entry_valid_1_26 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  flow_entry_valid_1_27 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  flow_entry_valid_1_28 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  flow_entry_valid_1_29 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  flow_entry_valid_1_30 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  flow_entry_valid_1_31 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  enqPtr_0_value = _RAND_192[4:0];
  _RAND_193 = {1{`RANDOM}};
  enqPtr_1_value = _RAND_193[4:0];
  _RAND_194 = {1{`RANDOM}};
  deqPtr_0_flag = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  deqPtr_0_value = _RAND_195[4:0];
  _RAND_196 = {1{`RANDOM}};
  deqPtr_1_flag = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  deqPtr_1_value = _RAND_197[4:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    flow_entry_valid_0_0 = 1'h0;
  end
  if (reset) begin
    flow_entry_valid_0_1 = 1'h0;
  end
  if (reset) begin
    flow_entry_valid_0_2 = 1'h0;
  end
  if (reset) begin
    flow_entry_valid_0_3 = 1'h0;
  end
  if (reset) begin
    flow_entry_valid_0_4 = 1'h0;
  end
  if (reset) begin
    flow_entry_valid_0_5 = 1'h0;
  end
  if (reset) begin
    flow_entry_valid_0_6 = 1'h0;
  end
  if (reset) begin
    flow_entry_valid_0_7 = 1'h0;
  end
  if (reset) begin
    flow_entry_valid_0_8 = 1'h0;
  end
  if (reset) begin
    flow_entry_valid_0_9 = 1'h0;
  end
  if (reset) begin
    flow_entry_valid_0_10 = 1'h0;
  end
  if (reset) begin
    flow_entry_valid_0_11 = 1'h0;
  end
  if (reset) begin
    flow_entry_valid_0_12 = 1'h0;
  end
  if (reset) begin
    flow_entry_valid_0_13 = 1'h0;
  end
  if (reset) begin
    flow_entry_valid_0_14 = 1'h0;
  end
  if (reset) begin
    flow_entry_valid_0_15 = 1'h0;
  end
  if (reset) begin
    flow_entry_valid_0_16 = 1'h0;
  end
  if (reset) begin
    flow_entry_valid_0_17 = 1'h0;
  end
  if (reset) begin
    flow_entry_valid_0_18 = 1'h0;
  end
  if (reset) begin
    flow_entry_valid_0_19 = 1'h0;
  end
  if (reset) begin
    flow_entry_valid_0_20 = 1'h0;
  end
  if (reset) begin
    flow_entry_valid_0_21 = 1'h0;
  end
  if (reset) begin
    flow_entry_valid_0_22 = 1'h0;
  end
  if (reset) begin
    flow_entry_valid_0_23 = 1'h0;
  end
  if (reset) begin
    flow_entry_valid_0_24 = 1'h0;
  end
  if (reset) begin
    flow_entry_valid_0_25 = 1'h0;
  end
  if (reset) begin
    flow_entry_valid_0_26 = 1'h0;
  end
  if (reset) begin
    flow_entry_valid_0_27 = 1'h0;
  end
  if (reset) begin
    flow_entry_valid_0_28 = 1'h0;
  end
  if (reset) begin
    flow_entry_valid_0_29 = 1'h0;
  end
  if (reset) begin
    flow_entry_valid_0_30 = 1'h0;
  end
  if (reset) begin
    flow_entry_valid_0_31 = 1'h0;
  end
  if (reset) begin
    flow_entry_valid_1_0 = 1'h0;
  end
  if (reset) begin
    flow_entry_valid_1_1 = 1'h0;
  end
  if (reset) begin
    flow_entry_valid_1_2 = 1'h0;
  end
  if (reset) begin
    flow_entry_valid_1_3 = 1'h0;
  end
  if (reset) begin
    flow_entry_valid_1_4 = 1'h0;
  end
  if (reset) begin
    flow_entry_valid_1_5 = 1'h0;
  end
  if (reset) begin
    flow_entry_valid_1_6 = 1'h0;
  end
  if (reset) begin
    flow_entry_valid_1_7 = 1'h0;
  end
  if (reset) begin
    flow_entry_valid_1_8 = 1'h0;
  end
  if (reset) begin
    flow_entry_valid_1_9 = 1'h0;
  end
  if (reset) begin
    flow_entry_valid_1_10 = 1'h0;
  end
  if (reset) begin
    flow_entry_valid_1_11 = 1'h0;
  end
  if (reset) begin
    flow_entry_valid_1_12 = 1'h0;
  end
  if (reset) begin
    flow_entry_valid_1_13 = 1'h0;
  end
  if (reset) begin
    flow_entry_valid_1_14 = 1'h0;
  end
  if (reset) begin
    flow_entry_valid_1_15 = 1'h0;
  end
  if (reset) begin
    flow_entry_valid_1_16 = 1'h0;
  end
  if (reset) begin
    flow_entry_valid_1_17 = 1'h0;
  end
  if (reset) begin
    flow_entry_valid_1_18 = 1'h0;
  end
  if (reset) begin
    flow_entry_valid_1_19 = 1'h0;
  end
  if (reset) begin
    flow_entry_valid_1_20 = 1'h0;
  end
  if (reset) begin
    flow_entry_valid_1_21 = 1'h0;
  end
  if (reset) begin
    flow_entry_valid_1_22 = 1'h0;
  end
  if (reset) begin
    flow_entry_valid_1_23 = 1'h0;
  end
  if (reset) begin
    flow_entry_valid_1_24 = 1'h0;
  end
  if (reset) begin
    flow_entry_valid_1_25 = 1'h0;
  end
  if (reset) begin
    flow_entry_valid_1_26 = 1'h0;
  end
  if (reset) begin
    flow_entry_valid_1_27 = 1'h0;
  end
  if (reset) begin
    flow_entry_valid_1_28 = 1'h0;
  end
  if (reset) begin
    flow_entry_valid_1_29 = 1'h0;
  end
  if (reset) begin
    flow_entry_valid_1_30 = 1'h0;
  end
  if (reset) begin
    flow_entry_valid_1_31 = 1'h0;
  end
  if (reset) begin
    enqPtr_0_value = 5'h0;
  end
  if (reset) begin
    enqPtr_1_value = 5'h0;
  end
  if (reset) begin
    deqPtr_0_flag = 1'h0;
  end
  if (reset) begin
    deqPtr_0_value = 5'h0;
  end
  if (reset) begin
    deqPtr_1_flag = 1'h0;
  end
  if (reset) begin
    deqPtr_1_value = 5'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule

