module Dispatch2Rs_5(
  output  io_in_0_ready,
  input   io_out_0_ready
);
  assign io_in_0_ready = io_out_0_ready; // @[Dispatch2Rs.scala 122:15 135:31 136:17]
endmodule

