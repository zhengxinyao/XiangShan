module L2TLB(
  input          clock,
  input          reset,
  input          auto_out_a_ready,
  output         auto_out_a_valid,
  output [2:0]   auto_out_a_bits_source,
  output [35:0]  auto_out_a_bits_address,
  input          auto_out_d_valid,
  input  [2:0]   auto_out_d_bits_opcode,
  input  [2:0]   auto_out_d_bits_size,
  input  [2:0]   auto_out_d_bits_source,
  input  [255:0] auto_out_d_bits_data,
  output         io_tlb_0_req_0_ready,
  input          io_tlb_0_req_0_valid,
  input  [26:0]  io_tlb_0_req_0_bits_vpn,
  input          io_tlb_0_resp_ready,
  output         io_tlb_0_resp_valid,
  output [26:0]  io_tlb_0_resp_bits_entry_tag,
  output [15:0]  io_tlb_0_resp_bits_entry_asid,
  output [23:0]  io_tlb_0_resp_bits_entry_ppn,
  output         io_tlb_0_resp_bits_entry_perm_d,
  output         io_tlb_0_resp_bits_entry_perm_a,
  output         io_tlb_0_resp_bits_entry_perm_g,
  output         io_tlb_0_resp_bits_entry_perm_u,
  output         io_tlb_0_resp_bits_entry_perm_x,
  output         io_tlb_0_resp_bits_entry_perm_w,
  output         io_tlb_0_resp_bits_entry_perm_r,
  output [1:0]   io_tlb_0_resp_bits_entry_level,
  output         io_tlb_0_resp_bits_pf,
  output         io_tlb_0_resp_bits_af,
  output         io_tlb_1_req_0_ready,
  input          io_tlb_1_req_0_valid,
  input  [26:0]  io_tlb_1_req_0_bits_vpn,
  input          io_tlb_1_resp_ready,
  output         io_tlb_1_resp_valid,
  output [26:0]  io_tlb_1_resp_bits_entry_tag,
  output [15:0]  io_tlb_1_resp_bits_entry_asid,
  output [23:0]  io_tlb_1_resp_bits_entry_ppn,
  output         io_tlb_1_resp_bits_entry_perm_d,
  output         io_tlb_1_resp_bits_entry_perm_a,
  output         io_tlb_1_resp_bits_entry_perm_g,
  output         io_tlb_1_resp_bits_entry_perm_u,
  output         io_tlb_1_resp_bits_entry_perm_x,
  output         io_tlb_1_resp_bits_entry_perm_w,
  output         io_tlb_1_resp_bits_entry_perm_r,
  output [1:0]   io_tlb_1_resp_bits_entry_level,
  output         io_tlb_1_resp_bits_pf,
  output         io_tlb_1_resp_bits_af,
  input          io_sfence_valid,
  input          io_sfence_bits_rs1,
  input          io_sfence_bits_rs2,
  input  [38:0]  io_sfence_bits_addr,
  input  [15:0]  io_sfence_bits_asid,
  input  [15:0]  io_csr_tlb_satp_asid,
  input  [43:0]  io_csr_tlb_satp_ppn,
  input          io_csr_tlb_satp_changed,
  input          io_csr_distribute_csr_wvalid,
  input  [11:0]  io_csr_distribute_csr_waddr,
  input  [63:0]  io_csr_distribute_csr_wdata,
  output [5:0]   io_perf_0_value,
  output [5:0]   io_perf_1_value,
  output [5:0]   io_perf_2_value,
  output [5:0]   io_perf_3_value,
  output [5:0]   io_perf_4_value,
  output [5:0]   io_perf_5_value,
  output [5:0]   io_perf_6_value,
  output [5:0]   io_perf_7_value,
  output [5:0]   io_perf_8_value,
  output [5:0]   io_perf_9_value,
  output [5:0]   io_perf_10_value,
  output [5:0]   io_perf_11_value,
  output [5:0]   io_perf_12_value,
  output [5:0]   io_perf_13_value,
  output [5:0]   io_perf_14_value,
  output [5:0]   io_perf_15_value,
  output [5:0]   io_perf_16_value,
  output [5:0]   io_perf_17_value,
  output [5:0]   io_perf_18_value
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [255:0] _RAND_49;
  reg [255:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [63:0] _RAND_52;
  reg [63:0] _RAND_53;
  reg [63:0] _RAND_54;
  reg [63:0] _RAND_55;
  reg [63:0] _RAND_56;
  reg [63:0] _RAND_57;
  reg [63:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [63:0] _RAND_75;
  reg [63:0] _RAND_76;
  reg [63:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [63:0] _RAND_116;
  reg [63:0] _RAND_117;
  reg [63:0] _RAND_118;
  reg [63:0] _RAND_119;
  reg [63:0] _RAND_120;
  reg [63:0] _RAND_121;
  reg [63:0] _RAND_122;
  reg [63:0] _RAND_123;
  reg [63:0] _RAND_124;
  reg [63:0] _RAND_125;
  reg [63:0] _RAND_126;
`endif // RANDOMIZE_REG_INIT
  wire  sfence_tmp_delay_clock; // @[Hold.scala 97:23]
  wire  sfence_tmp_delay_io_in_valid; // @[Hold.scala 97:23]
  wire  sfence_tmp_delay_io_in_bits_rs1; // @[Hold.scala 97:23]
  wire  sfence_tmp_delay_io_in_bits_rs2; // @[Hold.scala 97:23]
  wire [38:0] sfence_tmp_delay_io_in_bits_addr; // @[Hold.scala 97:23]
  wire [15:0] sfence_tmp_delay_io_in_bits_asid; // @[Hold.scala 97:23]
  wire  sfence_tmp_delay_io_out_valid; // @[Hold.scala 97:23]
  wire  sfence_tmp_delay_io_out_bits_rs1; // @[Hold.scala 97:23]
  wire  sfence_tmp_delay_io_out_bits_rs2; // @[Hold.scala 97:23]
  wire [38:0] sfence_tmp_delay_io_out_bits_addr; // @[Hold.scala 97:23]
  wire [15:0] sfence_tmp_delay_io_out_bits_asid; // @[Hold.scala 97:23]
  wire  csr_tmp_delay_clock; // @[Hold.scala 97:23]
  wire [15:0] csr_tmp_delay_io_in_satp_asid; // @[Hold.scala 97:23]
  wire [43:0] csr_tmp_delay_io_in_satp_ppn; // @[Hold.scala 97:23]
  wire  csr_tmp_delay_io_in_satp_changed; // @[Hold.scala 97:23]
  wire [15:0] csr_tmp_delay_io_out_satp_asid; // @[Hold.scala 97:23]
  wire [43:0] csr_tmp_delay_io_out_satp_ppn; // @[Hold.scala 97:23]
  wire  csr_tmp_delay_io_out_satp_changed; // @[Hold.scala 97:23]
  wire  pmp_clock; // @[L2TLB.scala 88:19]
  wire  pmp_reset; // @[L2TLB.scala 88:19]
  wire  pmp_io_distribute_csr_wvalid; // @[L2TLB.scala 88:19]
  wire [11:0] pmp_io_distribute_csr_waddr; // @[L2TLB.scala 88:19]
  wire [63:0] pmp_io_distribute_csr_wdata; // @[L2TLB.scala 88:19]
  wire  pmp_io_pmp_0_cfg_l; // @[L2TLB.scala 88:19]
  wire [1:0] pmp_io_pmp_0_cfg_a; // @[L2TLB.scala 88:19]
  wire  pmp_io_pmp_0_cfg_x; // @[L2TLB.scala 88:19]
  wire  pmp_io_pmp_0_cfg_w; // @[L2TLB.scala 88:19]
  wire  pmp_io_pmp_0_cfg_r; // @[L2TLB.scala 88:19]
  wire [33:0] pmp_io_pmp_0_addr; // @[L2TLB.scala 88:19]
  wire [35:0] pmp_io_pmp_0_mask; // @[L2TLB.scala 88:19]
  wire  pmp_io_pmp_1_cfg_l; // @[L2TLB.scala 88:19]
  wire [1:0] pmp_io_pmp_1_cfg_a; // @[L2TLB.scala 88:19]
  wire  pmp_io_pmp_1_cfg_x; // @[L2TLB.scala 88:19]
  wire  pmp_io_pmp_1_cfg_w; // @[L2TLB.scala 88:19]
  wire  pmp_io_pmp_1_cfg_r; // @[L2TLB.scala 88:19]
  wire [33:0] pmp_io_pmp_1_addr; // @[L2TLB.scala 88:19]
  wire [35:0] pmp_io_pmp_1_mask; // @[L2TLB.scala 88:19]
  wire  pmp_io_pmp_2_cfg_l; // @[L2TLB.scala 88:19]
  wire [1:0] pmp_io_pmp_2_cfg_a; // @[L2TLB.scala 88:19]
  wire  pmp_io_pmp_2_cfg_x; // @[L2TLB.scala 88:19]
  wire  pmp_io_pmp_2_cfg_w; // @[L2TLB.scala 88:19]
  wire  pmp_io_pmp_2_cfg_r; // @[L2TLB.scala 88:19]
  wire [33:0] pmp_io_pmp_2_addr; // @[L2TLB.scala 88:19]
  wire [35:0] pmp_io_pmp_2_mask; // @[L2TLB.scala 88:19]
  wire  pmp_io_pmp_3_cfg_l; // @[L2TLB.scala 88:19]
  wire [1:0] pmp_io_pmp_3_cfg_a; // @[L2TLB.scala 88:19]
  wire  pmp_io_pmp_3_cfg_x; // @[L2TLB.scala 88:19]
  wire  pmp_io_pmp_3_cfg_w; // @[L2TLB.scala 88:19]
  wire  pmp_io_pmp_3_cfg_r; // @[L2TLB.scala 88:19]
  wire [33:0] pmp_io_pmp_3_addr; // @[L2TLB.scala 88:19]
  wire [35:0] pmp_io_pmp_3_mask; // @[L2TLB.scala 88:19]
  wire  pmp_io_pmp_4_cfg_l; // @[L2TLB.scala 88:19]
  wire [1:0] pmp_io_pmp_4_cfg_a; // @[L2TLB.scala 88:19]
  wire  pmp_io_pmp_4_cfg_x; // @[L2TLB.scala 88:19]
  wire  pmp_io_pmp_4_cfg_w; // @[L2TLB.scala 88:19]
  wire  pmp_io_pmp_4_cfg_r; // @[L2TLB.scala 88:19]
  wire [33:0] pmp_io_pmp_4_addr; // @[L2TLB.scala 88:19]
  wire [35:0] pmp_io_pmp_4_mask; // @[L2TLB.scala 88:19]
  wire  pmp_io_pmp_5_cfg_l; // @[L2TLB.scala 88:19]
  wire [1:0] pmp_io_pmp_5_cfg_a; // @[L2TLB.scala 88:19]
  wire  pmp_io_pmp_5_cfg_x; // @[L2TLB.scala 88:19]
  wire  pmp_io_pmp_5_cfg_w; // @[L2TLB.scala 88:19]
  wire  pmp_io_pmp_5_cfg_r; // @[L2TLB.scala 88:19]
  wire [33:0] pmp_io_pmp_5_addr; // @[L2TLB.scala 88:19]
  wire [35:0] pmp_io_pmp_5_mask; // @[L2TLB.scala 88:19]
  wire  pmp_io_pmp_6_cfg_l; // @[L2TLB.scala 88:19]
  wire [1:0] pmp_io_pmp_6_cfg_a; // @[L2TLB.scala 88:19]
  wire  pmp_io_pmp_6_cfg_x; // @[L2TLB.scala 88:19]
  wire  pmp_io_pmp_6_cfg_w; // @[L2TLB.scala 88:19]
  wire  pmp_io_pmp_6_cfg_r; // @[L2TLB.scala 88:19]
  wire [33:0] pmp_io_pmp_6_addr; // @[L2TLB.scala 88:19]
  wire [35:0] pmp_io_pmp_6_mask; // @[L2TLB.scala 88:19]
  wire  pmp_io_pmp_7_cfg_l; // @[L2TLB.scala 88:19]
  wire [1:0] pmp_io_pmp_7_cfg_a; // @[L2TLB.scala 88:19]
  wire  pmp_io_pmp_7_cfg_x; // @[L2TLB.scala 88:19]
  wire  pmp_io_pmp_7_cfg_w; // @[L2TLB.scala 88:19]
  wire  pmp_io_pmp_7_cfg_r; // @[L2TLB.scala 88:19]
  wire [33:0] pmp_io_pmp_7_addr; // @[L2TLB.scala 88:19]
  wire [35:0] pmp_io_pmp_7_mask; // @[L2TLB.scala 88:19]
  wire  pmp_io_pmp_8_cfg_l; // @[L2TLB.scala 88:19]
  wire [1:0] pmp_io_pmp_8_cfg_a; // @[L2TLB.scala 88:19]
  wire  pmp_io_pmp_8_cfg_x; // @[L2TLB.scala 88:19]
  wire  pmp_io_pmp_8_cfg_w; // @[L2TLB.scala 88:19]
  wire  pmp_io_pmp_8_cfg_r; // @[L2TLB.scala 88:19]
  wire [33:0] pmp_io_pmp_8_addr; // @[L2TLB.scala 88:19]
  wire [35:0] pmp_io_pmp_8_mask; // @[L2TLB.scala 88:19]
  wire  pmp_io_pmp_9_cfg_l; // @[L2TLB.scala 88:19]
  wire [1:0] pmp_io_pmp_9_cfg_a; // @[L2TLB.scala 88:19]
  wire  pmp_io_pmp_9_cfg_x; // @[L2TLB.scala 88:19]
  wire  pmp_io_pmp_9_cfg_w; // @[L2TLB.scala 88:19]
  wire  pmp_io_pmp_9_cfg_r; // @[L2TLB.scala 88:19]
  wire [33:0] pmp_io_pmp_9_addr; // @[L2TLB.scala 88:19]
  wire [35:0] pmp_io_pmp_9_mask; // @[L2TLB.scala 88:19]
  wire  pmp_io_pmp_10_cfg_l; // @[L2TLB.scala 88:19]
  wire [1:0] pmp_io_pmp_10_cfg_a; // @[L2TLB.scala 88:19]
  wire  pmp_io_pmp_10_cfg_x; // @[L2TLB.scala 88:19]
  wire  pmp_io_pmp_10_cfg_w; // @[L2TLB.scala 88:19]
  wire  pmp_io_pmp_10_cfg_r; // @[L2TLB.scala 88:19]
  wire [33:0] pmp_io_pmp_10_addr; // @[L2TLB.scala 88:19]
  wire [35:0] pmp_io_pmp_10_mask; // @[L2TLB.scala 88:19]
  wire  pmp_io_pmp_11_cfg_l; // @[L2TLB.scala 88:19]
  wire [1:0] pmp_io_pmp_11_cfg_a; // @[L2TLB.scala 88:19]
  wire  pmp_io_pmp_11_cfg_x; // @[L2TLB.scala 88:19]
  wire  pmp_io_pmp_11_cfg_w; // @[L2TLB.scala 88:19]
  wire  pmp_io_pmp_11_cfg_r; // @[L2TLB.scala 88:19]
  wire [33:0] pmp_io_pmp_11_addr; // @[L2TLB.scala 88:19]
  wire [35:0] pmp_io_pmp_11_mask; // @[L2TLB.scala 88:19]
  wire  pmp_io_pmp_12_cfg_l; // @[L2TLB.scala 88:19]
  wire [1:0] pmp_io_pmp_12_cfg_a; // @[L2TLB.scala 88:19]
  wire  pmp_io_pmp_12_cfg_x; // @[L2TLB.scala 88:19]
  wire  pmp_io_pmp_12_cfg_w; // @[L2TLB.scala 88:19]
  wire  pmp_io_pmp_12_cfg_r; // @[L2TLB.scala 88:19]
  wire [33:0] pmp_io_pmp_12_addr; // @[L2TLB.scala 88:19]
  wire [35:0] pmp_io_pmp_12_mask; // @[L2TLB.scala 88:19]
  wire  pmp_io_pmp_13_cfg_l; // @[L2TLB.scala 88:19]
  wire [1:0] pmp_io_pmp_13_cfg_a; // @[L2TLB.scala 88:19]
  wire  pmp_io_pmp_13_cfg_x; // @[L2TLB.scala 88:19]
  wire  pmp_io_pmp_13_cfg_w; // @[L2TLB.scala 88:19]
  wire  pmp_io_pmp_13_cfg_r; // @[L2TLB.scala 88:19]
  wire [33:0] pmp_io_pmp_13_addr; // @[L2TLB.scala 88:19]
  wire [35:0] pmp_io_pmp_13_mask; // @[L2TLB.scala 88:19]
  wire  pmp_io_pmp_14_cfg_l; // @[L2TLB.scala 88:19]
  wire [1:0] pmp_io_pmp_14_cfg_a; // @[L2TLB.scala 88:19]
  wire  pmp_io_pmp_14_cfg_x; // @[L2TLB.scala 88:19]
  wire  pmp_io_pmp_14_cfg_w; // @[L2TLB.scala 88:19]
  wire  pmp_io_pmp_14_cfg_r; // @[L2TLB.scala 88:19]
  wire [33:0] pmp_io_pmp_14_addr; // @[L2TLB.scala 88:19]
  wire [35:0] pmp_io_pmp_14_mask; // @[L2TLB.scala 88:19]
  wire  pmp_io_pmp_15_cfg_l; // @[L2TLB.scala 88:19]
  wire [1:0] pmp_io_pmp_15_cfg_a; // @[L2TLB.scala 88:19]
  wire  pmp_io_pmp_15_cfg_x; // @[L2TLB.scala 88:19]
  wire  pmp_io_pmp_15_cfg_w; // @[L2TLB.scala 88:19]
  wire  pmp_io_pmp_15_cfg_r; // @[L2TLB.scala 88:19]
  wire [33:0] pmp_io_pmp_15_addr; // @[L2TLB.scala 88:19]
  wire [35:0] pmp_io_pmp_15_mask; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_0_cfg_c; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_0_cfg_atomic; // @[L2TLB.scala 88:19]
  wire [1:0] pmp_io_pma_0_cfg_a; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_0_cfg_x; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_0_cfg_w; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_0_cfg_r; // @[L2TLB.scala 88:19]
  wire [33:0] pmp_io_pma_0_addr; // @[L2TLB.scala 88:19]
  wire [35:0] pmp_io_pma_0_mask; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_1_cfg_c; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_1_cfg_atomic; // @[L2TLB.scala 88:19]
  wire [1:0] pmp_io_pma_1_cfg_a; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_1_cfg_x; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_1_cfg_w; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_1_cfg_r; // @[L2TLB.scala 88:19]
  wire [33:0] pmp_io_pma_1_addr; // @[L2TLB.scala 88:19]
  wire [35:0] pmp_io_pma_1_mask; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_2_cfg_c; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_2_cfg_atomic; // @[L2TLB.scala 88:19]
  wire [1:0] pmp_io_pma_2_cfg_a; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_2_cfg_x; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_2_cfg_w; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_2_cfg_r; // @[L2TLB.scala 88:19]
  wire [33:0] pmp_io_pma_2_addr; // @[L2TLB.scala 88:19]
  wire [35:0] pmp_io_pma_2_mask; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_3_cfg_c; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_3_cfg_atomic; // @[L2TLB.scala 88:19]
  wire [1:0] pmp_io_pma_3_cfg_a; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_3_cfg_x; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_3_cfg_w; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_3_cfg_r; // @[L2TLB.scala 88:19]
  wire [33:0] pmp_io_pma_3_addr; // @[L2TLB.scala 88:19]
  wire [35:0] pmp_io_pma_3_mask; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_4_cfg_c; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_4_cfg_atomic; // @[L2TLB.scala 88:19]
  wire [1:0] pmp_io_pma_4_cfg_a; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_4_cfg_x; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_4_cfg_w; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_4_cfg_r; // @[L2TLB.scala 88:19]
  wire [33:0] pmp_io_pma_4_addr; // @[L2TLB.scala 88:19]
  wire [35:0] pmp_io_pma_4_mask; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_5_cfg_c; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_5_cfg_atomic; // @[L2TLB.scala 88:19]
  wire [1:0] pmp_io_pma_5_cfg_a; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_5_cfg_x; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_5_cfg_w; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_5_cfg_r; // @[L2TLB.scala 88:19]
  wire [33:0] pmp_io_pma_5_addr; // @[L2TLB.scala 88:19]
  wire [35:0] pmp_io_pma_5_mask; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_6_cfg_c; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_6_cfg_atomic; // @[L2TLB.scala 88:19]
  wire [1:0] pmp_io_pma_6_cfg_a; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_6_cfg_x; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_6_cfg_w; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_6_cfg_r; // @[L2TLB.scala 88:19]
  wire [33:0] pmp_io_pma_6_addr; // @[L2TLB.scala 88:19]
  wire [35:0] pmp_io_pma_6_mask; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_7_cfg_c; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_7_cfg_atomic; // @[L2TLB.scala 88:19]
  wire [1:0] pmp_io_pma_7_cfg_a; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_7_cfg_x; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_7_cfg_w; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_7_cfg_r; // @[L2TLB.scala 88:19]
  wire [33:0] pmp_io_pma_7_addr; // @[L2TLB.scala 88:19]
  wire [35:0] pmp_io_pma_7_mask; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_8_cfg_c; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_8_cfg_atomic; // @[L2TLB.scala 88:19]
  wire [1:0] pmp_io_pma_8_cfg_a; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_8_cfg_x; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_8_cfg_w; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_8_cfg_r; // @[L2TLB.scala 88:19]
  wire [33:0] pmp_io_pma_8_addr; // @[L2TLB.scala 88:19]
  wire [35:0] pmp_io_pma_8_mask; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_9_cfg_c; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_9_cfg_atomic; // @[L2TLB.scala 88:19]
  wire [1:0] pmp_io_pma_9_cfg_a; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_9_cfg_x; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_9_cfg_w; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_9_cfg_r; // @[L2TLB.scala 88:19]
  wire [33:0] pmp_io_pma_9_addr; // @[L2TLB.scala 88:19]
  wire [35:0] pmp_io_pma_9_mask; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_10_cfg_c; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_10_cfg_atomic; // @[L2TLB.scala 88:19]
  wire [1:0] pmp_io_pma_10_cfg_a; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_10_cfg_x; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_10_cfg_w; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_10_cfg_r; // @[L2TLB.scala 88:19]
  wire [33:0] pmp_io_pma_10_addr; // @[L2TLB.scala 88:19]
  wire [35:0] pmp_io_pma_10_mask; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_11_cfg_c; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_11_cfg_atomic; // @[L2TLB.scala 88:19]
  wire [1:0] pmp_io_pma_11_cfg_a; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_11_cfg_x; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_11_cfg_w; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_11_cfg_r; // @[L2TLB.scala 88:19]
  wire [33:0] pmp_io_pma_11_addr; // @[L2TLB.scala 88:19]
  wire [35:0] pmp_io_pma_11_mask; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_12_cfg_c; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_12_cfg_atomic; // @[L2TLB.scala 88:19]
  wire [1:0] pmp_io_pma_12_cfg_a; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_12_cfg_x; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_12_cfg_w; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_12_cfg_r; // @[L2TLB.scala 88:19]
  wire [33:0] pmp_io_pma_12_addr; // @[L2TLB.scala 88:19]
  wire [35:0] pmp_io_pma_12_mask; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_13_cfg_c; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_13_cfg_atomic; // @[L2TLB.scala 88:19]
  wire [1:0] pmp_io_pma_13_cfg_a; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_13_cfg_x; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_13_cfg_w; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_13_cfg_r; // @[L2TLB.scala 88:19]
  wire [33:0] pmp_io_pma_13_addr; // @[L2TLB.scala 88:19]
  wire [35:0] pmp_io_pma_13_mask; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_14_cfg_c; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_14_cfg_atomic; // @[L2TLB.scala 88:19]
  wire [1:0] pmp_io_pma_14_cfg_a; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_14_cfg_x; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_14_cfg_w; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_14_cfg_r; // @[L2TLB.scala 88:19]
  wire [33:0] pmp_io_pma_14_addr; // @[L2TLB.scala 88:19]
  wire [35:0] pmp_io_pma_14_mask; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_15_cfg_c; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_15_cfg_atomic; // @[L2TLB.scala 88:19]
  wire [1:0] pmp_io_pma_15_cfg_a; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_15_cfg_x; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_15_cfg_w; // @[L2TLB.scala 88:19]
  wire  pmp_io_pma_15_cfg_r; // @[L2TLB.scala 88:19]
  wire [33:0] pmp_io_pma_15_addr; // @[L2TLB.scala 88:19]
  wire [35:0] pmp_io_pma_15_mask; // @[L2TLB.scala 88:19]
  wire [1:0] PMPChecker_io_check_env_mode; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pmp_0_cfg_l; // @[L2TLB.scala 89:45]
  wire [1:0] PMPChecker_io_check_env_pmp_0_cfg_a; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pmp_0_cfg_x; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pmp_0_cfg_w; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pmp_0_cfg_r; // @[L2TLB.scala 89:45]
  wire [33:0] PMPChecker_io_check_env_pmp_0_addr; // @[L2TLB.scala 89:45]
  wire [35:0] PMPChecker_io_check_env_pmp_0_mask; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pmp_1_cfg_l; // @[L2TLB.scala 89:45]
  wire [1:0] PMPChecker_io_check_env_pmp_1_cfg_a; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pmp_1_cfg_x; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pmp_1_cfg_w; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pmp_1_cfg_r; // @[L2TLB.scala 89:45]
  wire [33:0] PMPChecker_io_check_env_pmp_1_addr; // @[L2TLB.scala 89:45]
  wire [35:0] PMPChecker_io_check_env_pmp_1_mask; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pmp_2_cfg_l; // @[L2TLB.scala 89:45]
  wire [1:0] PMPChecker_io_check_env_pmp_2_cfg_a; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pmp_2_cfg_x; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pmp_2_cfg_w; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pmp_2_cfg_r; // @[L2TLB.scala 89:45]
  wire [33:0] PMPChecker_io_check_env_pmp_2_addr; // @[L2TLB.scala 89:45]
  wire [35:0] PMPChecker_io_check_env_pmp_2_mask; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pmp_3_cfg_l; // @[L2TLB.scala 89:45]
  wire [1:0] PMPChecker_io_check_env_pmp_3_cfg_a; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pmp_3_cfg_x; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pmp_3_cfg_w; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pmp_3_cfg_r; // @[L2TLB.scala 89:45]
  wire [33:0] PMPChecker_io_check_env_pmp_3_addr; // @[L2TLB.scala 89:45]
  wire [35:0] PMPChecker_io_check_env_pmp_3_mask; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pmp_4_cfg_l; // @[L2TLB.scala 89:45]
  wire [1:0] PMPChecker_io_check_env_pmp_4_cfg_a; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pmp_4_cfg_x; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pmp_4_cfg_w; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pmp_4_cfg_r; // @[L2TLB.scala 89:45]
  wire [33:0] PMPChecker_io_check_env_pmp_4_addr; // @[L2TLB.scala 89:45]
  wire [35:0] PMPChecker_io_check_env_pmp_4_mask; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pmp_5_cfg_l; // @[L2TLB.scala 89:45]
  wire [1:0] PMPChecker_io_check_env_pmp_5_cfg_a; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pmp_5_cfg_x; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pmp_5_cfg_w; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pmp_5_cfg_r; // @[L2TLB.scala 89:45]
  wire [33:0] PMPChecker_io_check_env_pmp_5_addr; // @[L2TLB.scala 89:45]
  wire [35:0] PMPChecker_io_check_env_pmp_5_mask; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pmp_6_cfg_l; // @[L2TLB.scala 89:45]
  wire [1:0] PMPChecker_io_check_env_pmp_6_cfg_a; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pmp_6_cfg_x; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pmp_6_cfg_w; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pmp_6_cfg_r; // @[L2TLB.scala 89:45]
  wire [33:0] PMPChecker_io_check_env_pmp_6_addr; // @[L2TLB.scala 89:45]
  wire [35:0] PMPChecker_io_check_env_pmp_6_mask; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pmp_7_cfg_l; // @[L2TLB.scala 89:45]
  wire [1:0] PMPChecker_io_check_env_pmp_7_cfg_a; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pmp_7_cfg_x; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pmp_7_cfg_w; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pmp_7_cfg_r; // @[L2TLB.scala 89:45]
  wire [33:0] PMPChecker_io_check_env_pmp_7_addr; // @[L2TLB.scala 89:45]
  wire [35:0] PMPChecker_io_check_env_pmp_7_mask; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pmp_8_cfg_l; // @[L2TLB.scala 89:45]
  wire [1:0] PMPChecker_io_check_env_pmp_8_cfg_a; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pmp_8_cfg_x; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pmp_8_cfg_w; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pmp_8_cfg_r; // @[L2TLB.scala 89:45]
  wire [33:0] PMPChecker_io_check_env_pmp_8_addr; // @[L2TLB.scala 89:45]
  wire [35:0] PMPChecker_io_check_env_pmp_8_mask; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pmp_9_cfg_l; // @[L2TLB.scala 89:45]
  wire [1:0] PMPChecker_io_check_env_pmp_9_cfg_a; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pmp_9_cfg_x; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pmp_9_cfg_w; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pmp_9_cfg_r; // @[L2TLB.scala 89:45]
  wire [33:0] PMPChecker_io_check_env_pmp_9_addr; // @[L2TLB.scala 89:45]
  wire [35:0] PMPChecker_io_check_env_pmp_9_mask; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pmp_10_cfg_l; // @[L2TLB.scala 89:45]
  wire [1:0] PMPChecker_io_check_env_pmp_10_cfg_a; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pmp_10_cfg_x; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pmp_10_cfg_w; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pmp_10_cfg_r; // @[L2TLB.scala 89:45]
  wire [33:0] PMPChecker_io_check_env_pmp_10_addr; // @[L2TLB.scala 89:45]
  wire [35:0] PMPChecker_io_check_env_pmp_10_mask; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pmp_11_cfg_l; // @[L2TLB.scala 89:45]
  wire [1:0] PMPChecker_io_check_env_pmp_11_cfg_a; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pmp_11_cfg_x; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pmp_11_cfg_w; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pmp_11_cfg_r; // @[L2TLB.scala 89:45]
  wire [33:0] PMPChecker_io_check_env_pmp_11_addr; // @[L2TLB.scala 89:45]
  wire [35:0] PMPChecker_io_check_env_pmp_11_mask; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pmp_12_cfg_l; // @[L2TLB.scala 89:45]
  wire [1:0] PMPChecker_io_check_env_pmp_12_cfg_a; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pmp_12_cfg_x; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pmp_12_cfg_w; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pmp_12_cfg_r; // @[L2TLB.scala 89:45]
  wire [33:0] PMPChecker_io_check_env_pmp_12_addr; // @[L2TLB.scala 89:45]
  wire [35:0] PMPChecker_io_check_env_pmp_12_mask; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pmp_13_cfg_l; // @[L2TLB.scala 89:45]
  wire [1:0] PMPChecker_io_check_env_pmp_13_cfg_a; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pmp_13_cfg_x; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pmp_13_cfg_w; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pmp_13_cfg_r; // @[L2TLB.scala 89:45]
  wire [33:0] PMPChecker_io_check_env_pmp_13_addr; // @[L2TLB.scala 89:45]
  wire [35:0] PMPChecker_io_check_env_pmp_13_mask; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pmp_14_cfg_l; // @[L2TLB.scala 89:45]
  wire [1:0] PMPChecker_io_check_env_pmp_14_cfg_a; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pmp_14_cfg_x; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pmp_14_cfg_w; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pmp_14_cfg_r; // @[L2TLB.scala 89:45]
  wire [33:0] PMPChecker_io_check_env_pmp_14_addr; // @[L2TLB.scala 89:45]
  wire [35:0] PMPChecker_io_check_env_pmp_14_mask; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pmp_15_cfg_l; // @[L2TLB.scala 89:45]
  wire [1:0] PMPChecker_io_check_env_pmp_15_cfg_a; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pmp_15_cfg_x; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pmp_15_cfg_w; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pmp_15_cfg_r; // @[L2TLB.scala 89:45]
  wire [33:0] PMPChecker_io_check_env_pmp_15_addr; // @[L2TLB.scala 89:45]
  wire [35:0] PMPChecker_io_check_env_pmp_15_mask; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_0_cfg_c; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_0_cfg_atomic; // @[L2TLB.scala 89:45]
  wire [1:0] PMPChecker_io_check_env_pma_0_cfg_a; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_0_cfg_x; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_0_cfg_w; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_0_cfg_r; // @[L2TLB.scala 89:45]
  wire [33:0] PMPChecker_io_check_env_pma_0_addr; // @[L2TLB.scala 89:45]
  wire [35:0] PMPChecker_io_check_env_pma_0_mask; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_1_cfg_c; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_1_cfg_atomic; // @[L2TLB.scala 89:45]
  wire [1:0] PMPChecker_io_check_env_pma_1_cfg_a; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_1_cfg_x; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_1_cfg_w; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_1_cfg_r; // @[L2TLB.scala 89:45]
  wire [33:0] PMPChecker_io_check_env_pma_1_addr; // @[L2TLB.scala 89:45]
  wire [35:0] PMPChecker_io_check_env_pma_1_mask; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_2_cfg_c; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_2_cfg_atomic; // @[L2TLB.scala 89:45]
  wire [1:0] PMPChecker_io_check_env_pma_2_cfg_a; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_2_cfg_x; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_2_cfg_w; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_2_cfg_r; // @[L2TLB.scala 89:45]
  wire [33:0] PMPChecker_io_check_env_pma_2_addr; // @[L2TLB.scala 89:45]
  wire [35:0] PMPChecker_io_check_env_pma_2_mask; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_3_cfg_c; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_3_cfg_atomic; // @[L2TLB.scala 89:45]
  wire [1:0] PMPChecker_io_check_env_pma_3_cfg_a; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_3_cfg_x; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_3_cfg_w; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_3_cfg_r; // @[L2TLB.scala 89:45]
  wire [33:0] PMPChecker_io_check_env_pma_3_addr; // @[L2TLB.scala 89:45]
  wire [35:0] PMPChecker_io_check_env_pma_3_mask; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_4_cfg_c; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_4_cfg_atomic; // @[L2TLB.scala 89:45]
  wire [1:0] PMPChecker_io_check_env_pma_4_cfg_a; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_4_cfg_x; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_4_cfg_w; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_4_cfg_r; // @[L2TLB.scala 89:45]
  wire [33:0] PMPChecker_io_check_env_pma_4_addr; // @[L2TLB.scala 89:45]
  wire [35:0] PMPChecker_io_check_env_pma_4_mask; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_5_cfg_c; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_5_cfg_atomic; // @[L2TLB.scala 89:45]
  wire [1:0] PMPChecker_io_check_env_pma_5_cfg_a; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_5_cfg_x; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_5_cfg_w; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_5_cfg_r; // @[L2TLB.scala 89:45]
  wire [33:0] PMPChecker_io_check_env_pma_5_addr; // @[L2TLB.scala 89:45]
  wire [35:0] PMPChecker_io_check_env_pma_5_mask; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_6_cfg_c; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_6_cfg_atomic; // @[L2TLB.scala 89:45]
  wire [1:0] PMPChecker_io_check_env_pma_6_cfg_a; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_6_cfg_x; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_6_cfg_w; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_6_cfg_r; // @[L2TLB.scala 89:45]
  wire [33:0] PMPChecker_io_check_env_pma_6_addr; // @[L2TLB.scala 89:45]
  wire [35:0] PMPChecker_io_check_env_pma_6_mask; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_7_cfg_c; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_7_cfg_atomic; // @[L2TLB.scala 89:45]
  wire [1:0] PMPChecker_io_check_env_pma_7_cfg_a; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_7_cfg_x; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_7_cfg_w; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_7_cfg_r; // @[L2TLB.scala 89:45]
  wire [33:0] PMPChecker_io_check_env_pma_7_addr; // @[L2TLB.scala 89:45]
  wire [35:0] PMPChecker_io_check_env_pma_7_mask; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_8_cfg_c; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_8_cfg_atomic; // @[L2TLB.scala 89:45]
  wire [1:0] PMPChecker_io_check_env_pma_8_cfg_a; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_8_cfg_x; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_8_cfg_w; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_8_cfg_r; // @[L2TLB.scala 89:45]
  wire [33:0] PMPChecker_io_check_env_pma_8_addr; // @[L2TLB.scala 89:45]
  wire [35:0] PMPChecker_io_check_env_pma_8_mask; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_9_cfg_c; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_9_cfg_atomic; // @[L2TLB.scala 89:45]
  wire [1:0] PMPChecker_io_check_env_pma_9_cfg_a; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_9_cfg_x; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_9_cfg_w; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_9_cfg_r; // @[L2TLB.scala 89:45]
  wire [33:0] PMPChecker_io_check_env_pma_9_addr; // @[L2TLB.scala 89:45]
  wire [35:0] PMPChecker_io_check_env_pma_9_mask; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_10_cfg_c; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_10_cfg_atomic; // @[L2TLB.scala 89:45]
  wire [1:0] PMPChecker_io_check_env_pma_10_cfg_a; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_10_cfg_x; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_10_cfg_w; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_10_cfg_r; // @[L2TLB.scala 89:45]
  wire [33:0] PMPChecker_io_check_env_pma_10_addr; // @[L2TLB.scala 89:45]
  wire [35:0] PMPChecker_io_check_env_pma_10_mask; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_11_cfg_c; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_11_cfg_atomic; // @[L2TLB.scala 89:45]
  wire [1:0] PMPChecker_io_check_env_pma_11_cfg_a; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_11_cfg_x; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_11_cfg_w; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_11_cfg_r; // @[L2TLB.scala 89:45]
  wire [33:0] PMPChecker_io_check_env_pma_11_addr; // @[L2TLB.scala 89:45]
  wire [35:0] PMPChecker_io_check_env_pma_11_mask; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_12_cfg_c; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_12_cfg_atomic; // @[L2TLB.scala 89:45]
  wire [1:0] PMPChecker_io_check_env_pma_12_cfg_a; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_12_cfg_x; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_12_cfg_w; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_12_cfg_r; // @[L2TLB.scala 89:45]
  wire [33:0] PMPChecker_io_check_env_pma_12_addr; // @[L2TLB.scala 89:45]
  wire [35:0] PMPChecker_io_check_env_pma_12_mask; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_13_cfg_c; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_13_cfg_atomic; // @[L2TLB.scala 89:45]
  wire [1:0] PMPChecker_io_check_env_pma_13_cfg_a; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_13_cfg_x; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_13_cfg_w; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_13_cfg_r; // @[L2TLB.scala 89:45]
  wire [33:0] PMPChecker_io_check_env_pma_13_addr; // @[L2TLB.scala 89:45]
  wire [35:0] PMPChecker_io_check_env_pma_13_mask; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_14_cfg_c; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_14_cfg_atomic; // @[L2TLB.scala 89:45]
  wire [1:0] PMPChecker_io_check_env_pma_14_cfg_a; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_14_cfg_x; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_14_cfg_w; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_14_cfg_r; // @[L2TLB.scala 89:45]
  wire [33:0] PMPChecker_io_check_env_pma_14_addr; // @[L2TLB.scala 89:45]
  wire [35:0] PMPChecker_io_check_env_pma_14_mask; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_15_cfg_c; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_15_cfg_atomic; // @[L2TLB.scala 89:45]
  wire [1:0] PMPChecker_io_check_env_pma_15_cfg_a; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_15_cfg_x; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_15_cfg_w; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_check_env_pma_15_cfg_r; // @[L2TLB.scala 89:45]
  wire [33:0] PMPChecker_io_check_env_pma_15_addr; // @[L2TLB.scala 89:45]
  wire [35:0] PMPChecker_io_check_env_pma_15_mask; // @[L2TLB.scala 89:45]
  wire [35:0] PMPChecker_io_req_bits_addr; // @[L2TLB.scala 89:45]
  wire [2:0] PMPChecker_io_req_bits_cmd; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_resp_ld; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_resp_st; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_resp_instr; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_resp_mmio; // @[L2TLB.scala 89:45]
  wire  PMPChecker_io_resp_atomic; // @[L2TLB.scala 89:45]
  wire [1:0] PMPChecker_1_io_check_env_mode; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pmp_0_cfg_l; // @[L2TLB.scala 89:45]
  wire [1:0] PMPChecker_1_io_check_env_pmp_0_cfg_a; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pmp_0_cfg_x; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pmp_0_cfg_w; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pmp_0_cfg_r; // @[L2TLB.scala 89:45]
  wire [33:0] PMPChecker_1_io_check_env_pmp_0_addr; // @[L2TLB.scala 89:45]
  wire [35:0] PMPChecker_1_io_check_env_pmp_0_mask; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pmp_1_cfg_l; // @[L2TLB.scala 89:45]
  wire [1:0] PMPChecker_1_io_check_env_pmp_1_cfg_a; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pmp_1_cfg_x; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pmp_1_cfg_w; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pmp_1_cfg_r; // @[L2TLB.scala 89:45]
  wire [33:0] PMPChecker_1_io_check_env_pmp_1_addr; // @[L2TLB.scala 89:45]
  wire [35:0] PMPChecker_1_io_check_env_pmp_1_mask; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pmp_2_cfg_l; // @[L2TLB.scala 89:45]
  wire [1:0] PMPChecker_1_io_check_env_pmp_2_cfg_a; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pmp_2_cfg_x; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pmp_2_cfg_w; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pmp_2_cfg_r; // @[L2TLB.scala 89:45]
  wire [33:0] PMPChecker_1_io_check_env_pmp_2_addr; // @[L2TLB.scala 89:45]
  wire [35:0] PMPChecker_1_io_check_env_pmp_2_mask; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pmp_3_cfg_l; // @[L2TLB.scala 89:45]
  wire [1:0] PMPChecker_1_io_check_env_pmp_3_cfg_a; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pmp_3_cfg_x; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pmp_3_cfg_w; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pmp_3_cfg_r; // @[L2TLB.scala 89:45]
  wire [33:0] PMPChecker_1_io_check_env_pmp_3_addr; // @[L2TLB.scala 89:45]
  wire [35:0] PMPChecker_1_io_check_env_pmp_3_mask; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pmp_4_cfg_l; // @[L2TLB.scala 89:45]
  wire [1:0] PMPChecker_1_io_check_env_pmp_4_cfg_a; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pmp_4_cfg_x; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pmp_4_cfg_w; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pmp_4_cfg_r; // @[L2TLB.scala 89:45]
  wire [33:0] PMPChecker_1_io_check_env_pmp_4_addr; // @[L2TLB.scala 89:45]
  wire [35:0] PMPChecker_1_io_check_env_pmp_4_mask; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pmp_5_cfg_l; // @[L2TLB.scala 89:45]
  wire [1:0] PMPChecker_1_io_check_env_pmp_5_cfg_a; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pmp_5_cfg_x; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pmp_5_cfg_w; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pmp_5_cfg_r; // @[L2TLB.scala 89:45]
  wire [33:0] PMPChecker_1_io_check_env_pmp_5_addr; // @[L2TLB.scala 89:45]
  wire [35:0] PMPChecker_1_io_check_env_pmp_5_mask; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pmp_6_cfg_l; // @[L2TLB.scala 89:45]
  wire [1:0] PMPChecker_1_io_check_env_pmp_6_cfg_a; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pmp_6_cfg_x; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pmp_6_cfg_w; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pmp_6_cfg_r; // @[L2TLB.scala 89:45]
  wire [33:0] PMPChecker_1_io_check_env_pmp_6_addr; // @[L2TLB.scala 89:45]
  wire [35:0] PMPChecker_1_io_check_env_pmp_6_mask; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pmp_7_cfg_l; // @[L2TLB.scala 89:45]
  wire [1:0] PMPChecker_1_io_check_env_pmp_7_cfg_a; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pmp_7_cfg_x; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pmp_7_cfg_w; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pmp_7_cfg_r; // @[L2TLB.scala 89:45]
  wire [33:0] PMPChecker_1_io_check_env_pmp_7_addr; // @[L2TLB.scala 89:45]
  wire [35:0] PMPChecker_1_io_check_env_pmp_7_mask; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pmp_8_cfg_l; // @[L2TLB.scala 89:45]
  wire [1:0] PMPChecker_1_io_check_env_pmp_8_cfg_a; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pmp_8_cfg_x; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pmp_8_cfg_w; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pmp_8_cfg_r; // @[L2TLB.scala 89:45]
  wire [33:0] PMPChecker_1_io_check_env_pmp_8_addr; // @[L2TLB.scala 89:45]
  wire [35:0] PMPChecker_1_io_check_env_pmp_8_mask; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pmp_9_cfg_l; // @[L2TLB.scala 89:45]
  wire [1:0] PMPChecker_1_io_check_env_pmp_9_cfg_a; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pmp_9_cfg_x; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pmp_9_cfg_w; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pmp_9_cfg_r; // @[L2TLB.scala 89:45]
  wire [33:0] PMPChecker_1_io_check_env_pmp_9_addr; // @[L2TLB.scala 89:45]
  wire [35:0] PMPChecker_1_io_check_env_pmp_9_mask; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pmp_10_cfg_l; // @[L2TLB.scala 89:45]
  wire [1:0] PMPChecker_1_io_check_env_pmp_10_cfg_a; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pmp_10_cfg_x; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pmp_10_cfg_w; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pmp_10_cfg_r; // @[L2TLB.scala 89:45]
  wire [33:0] PMPChecker_1_io_check_env_pmp_10_addr; // @[L2TLB.scala 89:45]
  wire [35:0] PMPChecker_1_io_check_env_pmp_10_mask; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pmp_11_cfg_l; // @[L2TLB.scala 89:45]
  wire [1:0] PMPChecker_1_io_check_env_pmp_11_cfg_a; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pmp_11_cfg_x; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pmp_11_cfg_w; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pmp_11_cfg_r; // @[L2TLB.scala 89:45]
  wire [33:0] PMPChecker_1_io_check_env_pmp_11_addr; // @[L2TLB.scala 89:45]
  wire [35:0] PMPChecker_1_io_check_env_pmp_11_mask; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pmp_12_cfg_l; // @[L2TLB.scala 89:45]
  wire [1:0] PMPChecker_1_io_check_env_pmp_12_cfg_a; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pmp_12_cfg_x; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pmp_12_cfg_w; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pmp_12_cfg_r; // @[L2TLB.scala 89:45]
  wire [33:0] PMPChecker_1_io_check_env_pmp_12_addr; // @[L2TLB.scala 89:45]
  wire [35:0] PMPChecker_1_io_check_env_pmp_12_mask; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pmp_13_cfg_l; // @[L2TLB.scala 89:45]
  wire [1:0] PMPChecker_1_io_check_env_pmp_13_cfg_a; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pmp_13_cfg_x; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pmp_13_cfg_w; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pmp_13_cfg_r; // @[L2TLB.scala 89:45]
  wire [33:0] PMPChecker_1_io_check_env_pmp_13_addr; // @[L2TLB.scala 89:45]
  wire [35:0] PMPChecker_1_io_check_env_pmp_13_mask; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pmp_14_cfg_l; // @[L2TLB.scala 89:45]
  wire [1:0] PMPChecker_1_io_check_env_pmp_14_cfg_a; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pmp_14_cfg_x; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pmp_14_cfg_w; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pmp_14_cfg_r; // @[L2TLB.scala 89:45]
  wire [33:0] PMPChecker_1_io_check_env_pmp_14_addr; // @[L2TLB.scala 89:45]
  wire [35:0] PMPChecker_1_io_check_env_pmp_14_mask; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pmp_15_cfg_l; // @[L2TLB.scala 89:45]
  wire [1:0] PMPChecker_1_io_check_env_pmp_15_cfg_a; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pmp_15_cfg_x; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pmp_15_cfg_w; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pmp_15_cfg_r; // @[L2TLB.scala 89:45]
  wire [33:0] PMPChecker_1_io_check_env_pmp_15_addr; // @[L2TLB.scala 89:45]
  wire [35:0] PMPChecker_1_io_check_env_pmp_15_mask; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_0_cfg_c; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_0_cfg_atomic; // @[L2TLB.scala 89:45]
  wire [1:0] PMPChecker_1_io_check_env_pma_0_cfg_a; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_0_cfg_x; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_0_cfg_w; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_0_cfg_r; // @[L2TLB.scala 89:45]
  wire [33:0] PMPChecker_1_io_check_env_pma_0_addr; // @[L2TLB.scala 89:45]
  wire [35:0] PMPChecker_1_io_check_env_pma_0_mask; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_1_cfg_c; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_1_cfg_atomic; // @[L2TLB.scala 89:45]
  wire [1:0] PMPChecker_1_io_check_env_pma_1_cfg_a; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_1_cfg_x; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_1_cfg_w; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_1_cfg_r; // @[L2TLB.scala 89:45]
  wire [33:0] PMPChecker_1_io_check_env_pma_1_addr; // @[L2TLB.scala 89:45]
  wire [35:0] PMPChecker_1_io_check_env_pma_1_mask; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_2_cfg_c; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_2_cfg_atomic; // @[L2TLB.scala 89:45]
  wire [1:0] PMPChecker_1_io_check_env_pma_2_cfg_a; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_2_cfg_x; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_2_cfg_w; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_2_cfg_r; // @[L2TLB.scala 89:45]
  wire [33:0] PMPChecker_1_io_check_env_pma_2_addr; // @[L2TLB.scala 89:45]
  wire [35:0] PMPChecker_1_io_check_env_pma_2_mask; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_3_cfg_c; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_3_cfg_atomic; // @[L2TLB.scala 89:45]
  wire [1:0] PMPChecker_1_io_check_env_pma_3_cfg_a; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_3_cfg_x; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_3_cfg_w; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_3_cfg_r; // @[L2TLB.scala 89:45]
  wire [33:0] PMPChecker_1_io_check_env_pma_3_addr; // @[L2TLB.scala 89:45]
  wire [35:0] PMPChecker_1_io_check_env_pma_3_mask; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_4_cfg_c; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_4_cfg_atomic; // @[L2TLB.scala 89:45]
  wire [1:0] PMPChecker_1_io_check_env_pma_4_cfg_a; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_4_cfg_x; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_4_cfg_w; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_4_cfg_r; // @[L2TLB.scala 89:45]
  wire [33:0] PMPChecker_1_io_check_env_pma_4_addr; // @[L2TLB.scala 89:45]
  wire [35:0] PMPChecker_1_io_check_env_pma_4_mask; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_5_cfg_c; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_5_cfg_atomic; // @[L2TLB.scala 89:45]
  wire [1:0] PMPChecker_1_io_check_env_pma_5_cfg_a; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_5_cfg_x; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_5_cfg_w; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_5_cfg_r; // @[L2TLB.scala 89:45]
  wire [33:0] PMPChecker_1_io_check_env_pma_5_addr; // @[L2TLB.scala 89:45]
  wire [35:0] PMPChecker_1_io_check_env_pma_5_mask; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_6_cfg_c; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_6_cfg_atomic; // @[L2TLB.scala 89:45]
  wire [1:0] PMPChecker_1_io_check_env_pma_6_cfg_a; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_6_cfg_x; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_6_cfg_w; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_6_cfg_r; // @[L2TLB.scala 89:45]
  wire [33:0] PMPChecker_1_io_check_env_pma_6_addr; // @[L2TLB.scala 89:45]
  wire [35:0] PMPChecker_1_io_check_env_pma_6_mask; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_7_cfg_c; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_7_cfg_atomic; // @[L2TLB.scala 89:45]
  wire [1:0] PMPChecker_1_io_check_env_pma_7_cfg_a; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_7_cfg_x; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_7_cfg_w; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_7_cfg_r; // @[L2TLB.scala 89:45]
  wire [33:0] PMPChecker_1_io_check_env_pma_7_addr; // @[L2TLB.scala 89:45]
  wire [35:0] PMPChecker_1_io_check_env_pma_7_mask; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_8_cfg_c; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_8_cfg_atomic; // @[L2TLB.scala 89:45]
  wire [1:0] PMPChecker_1_io_check_env_pma_8_cfg_a; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_8_cfg_x; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_8_cfg_w; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_8_cfg_r; // @[L2TLB.scala 89:45]
  wire [33:0] PMPChecker_1_io_check_env_pma_8_addr; // @[L2TLB.scala 89:45]
  wire [35:0] PMPChecker_1_io_check_env_pma_8_mask; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_9_cfg_c; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_9_cfg_atomic; // @[L2TLB.scala 89:45]
  wire [1:0] PMPChecker_1_io_check_env_pma_9_cfg_a; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_9_cfg_x; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_9_cfg_w; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_9_cfg_r; // @[L2TLB.scala 89:45]
  wire [33:0] PMPChecker_1_io_check_env_pma_9_addr; // @[L2TLB.scala 89:45]
  wire [35:0] PMPChecker_1_io_check_env_pma_9_mask; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_10_cfg_c; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_10_cfg_atomic; // @[L2TLB.scala 89:45]
  wire [1:0] PMPChecker_1_io_check_env_pma_10_cfg_a; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_10_cfg_x; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_10_cfg_w; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_10_cfg_r; // @[L2TLB.scala 89:45]
  wire [33:0] PMPChecker_1_io_check_env_pma_10_addr; // @[L2TLB.scala 89:45]
  wire [35:0] PMPChecker_1_io_check_env_pma_10_mask; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_11_cfg_c; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_11_cfg_atomic; // @[L2TLB.scala 89:45]
  wire [1:0] PMPChecker_1_io_check_env_pma_11_cfg_a; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_11_cfg_x; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_11_cfg_w; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_11_cfg_r; // @[L2TLB.scala 89:45]
  wire [33:0] PMPChecker_1_io_check_env_pma_11_addr; // @[L2TLB.scala 89:45]
  wire [35:0] PMPChecker_1_io_check_env_pma_11_mask; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_12_cfg_c; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_12_cfg_atomic; // @[L2TLB.scala 89:45]
  wire [1:0] PMPChecker_1_io_check_env_pma_12_cfg_a; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_12_cfg_x; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_12_cfg_w; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_12_cfg_r; // @[L2TLB.scala 89:45]
  wire [33:0] PMPChecker_1_io_check_env_pma_12_addr; // @[L2TLB.scala 89:45]
  wire [35:0] PMPChecker_1_io_check_env_pma_12_mask; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_13_cfg_c; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_13_cfg_atomic; // @[L2TLB.scala 89:45]
  wire [1:0] PMPChecker_1_io_check_env_pma_13_cfg_a; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_13_cfg_x; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_13_cfg_w; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_13_cfg_r; // @[L2TLB.scala 89:45]
  wire [33:0] PMPChecker_1_io_check_env_pma_13_addr; // @[L2TLB.scala 89:45]
  wire [35:0] PMPChecker_1_io_check_env_pma_13_mask; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_14_cfg_c; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_14_cfg_atomic; // @[L2TLB.scala 89:45]
  wire [1:0] PMPChecker_1_io_check_env_pma_14_cfg_a; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_14_cfg_x; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_14_cfg_w; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_14_cfg_r; // @[L2TLB.scala 89:45]
  wire [33:0] PMPChecker_1_io_check_env_pma_14_addr; // @[L2TLB.scala 89:45]
  wire [35:0] PMPChecker_1_io_check_env_pma_14_mask; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_15_cfg_c; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_15_cfg_atomic; // @[L2TLB.scala 89:45]
  wire [1:0] PMPChecker_1_io_check_env_pma_15_cfg_a; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_15_cfg_x; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_15_cfg_w; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_check_env_pma_15_cfg_r; // @[L2TLB.scala 89:45]
  wire [33:0] PMPChecker_1_io_check_env_pma_15_addr; // @[L2TLB.scala 89:45]
  wire [35:0] PMPChecker_1_io_check_env_pma_15_mask; // @[L2TLB.scala 89:45]
  wire [35:0] PMPChecker_1_io_req_bits_addr; // @[L2TLB.scala 89:45]
  wire [2:0] PMPChecker_1_io_req_bits_cmd; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_resp_ld; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_resp_st; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_resp_instr; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_resp_mmio; // @[L2TLB.scala 89:45]
  wire  PMPChecker_1_io_resp_atomic; // @[L2TLB.scala 89:45]
  wire  missQueue_clock; // @[L2TLB.scala 93:25]
  wire  missQueue_reset; // @[L2TLB.scala 93:25]
  wire  missQueue_io_sfence_valid; // @[L2TLB.scala 93:25]
  wire  missQueue_io_csr_satp_changed; // @[L2TLB.scala 93:25]
  wire  missQueue_io_in_ready; // @[L2TLB.scala 93:25]
  wire  missQueue_io_in_valid; // @[L2TLB.scala 93:25]
  wire [26:0] missQueue_io_in_bits_vpn; // @[L2TLB.scala 93:25]
  wire [1:0] missQueue_io_in_bits_source; // @[L2TLB.scala 93:25]
  wire  missQueue_io_out_ready; // @[L2TLB.scala 93:25]
  wire  missQueue_io_out_valid; // @[L2TLB.scala 93:25]
  wire [26:0] missQueue_io_out_bits_vpn; // @[L2TLB.scala 93:25]
  wire [1:0] missQueue_io_out_bits_source; // @[L2TLB.scala 93:25]
  wire  cache_clock; // @[L2TLB.scala 94:21]
  wire  cache_reset; // @[L2TLB.scala 94:21]
  wire  cache_io_req_ready; // @[L2TLB.scala 94:21]
  wire  cache_io_req_valid; // @[L2TLB.scala 94:21]
  wire [26:0] cache_io_req_bits_req_info_vpn; // @[L2TLB.scala 94:21]
  wire [1:0] cache_io_req_bits_req_info_source; // @[L2TLB.scala 94:21]
  wire  cache_io_req_bits_isFirst; // @[L2TLB.scala 94:21]
  wire  cache_io_resp_ready; // @[L2TLB.scala 94:21]
  wire  cache_io_resp_valid; // @[L2TLB.scala 94:21]
  wire [26:0] cache_io_resp_bits_req_info_vpn; // @[L2TLB.scala 94:21]
  wire [1:0] cache_io_resp_bits_req_info_source; // @[L2TLB.scala 94:21]
  wire  cache_io_resp_bits_isFirst; // @[L2TLB.scala 94:21]
  wire  cache_io_resp_bits_hit; // @[L2TLB.scala 94:21]
  wire  cache_io_resp_bits_prefetch; // @[L2TLB.scala 94:21]
  wire  cache_io_resp_bits_bypassed; // @[L2TLB.scala 94:21]
  wire  cache_io_resp_bits_toFsm_l1Hit; // @[L2TLB.scala 94:21]
  wire  cache_io_resp_bits_toFsm_l2Hit; // @[L2TLB.scala 94:21]
  wire [23:0] cache_io_resp_bits_toFsm_ppn; // @[L2TLB.scala 94:21]
  wire [26:0] cache_io_resp_bits_toTlb_tag; // @[L2TLB.scala 94:21]
  wire [15:0] cache_io_resp_bits_toTlb_asid; // @[L2TLB.scala 94:21]
  wire [23:0] cache_io_resp_bits_toTlb_ppn; // @[L2TLB.scala 94:21]
  wire  cache_io_resp_bits_toTlb_perm_d; // @[L2TLB.scala 94:21]
  wire  cache_io_resp_bits_toTlb_perm_a; // @[L2TLB.scala 94:21]
  wire  cache_io_resp_bits_toTlb_perm_g; // @[L2TLB.scala 94:21]
  wire  cache_io_resp_bits_toTlb_perm_u; // @[L2TLB.scala 94:21]
  wire  cache_io_resp_bits_toTlb_perm_x; // @[L2TLB.scala 94:21]
  wire  cache_io_resp_bits_toTlb_perm_w; // @[L2TLB.scala 94:21]
  wire  cache_io_resp_bits_toTlb_perm_r; // @[L2TLB.scala 94:21]
  wire [1:0] cache_io_resp_bits_toTlb_level; // @[L2TLB.scala 94:21]
  wire  cache_io_resp_bits_toTlb_prefetch; // @[L2TLB.scala 94:21]
  wire  cache_io_resp_bits_toTlb_v; // @[L2TLB.scala 94:21]
  wire  cache_io_refill_valid; // @[L2TLB.scala 94:21]
  wire [511:0] cache_io_refill_bits_ptes; // @[L2TLB.scala 94:21]
  wire  cache_io_refill_bits_levelOH_sp; // @[L2TLB.scala 94:21]
  wire  cache_io_refill_bits_levelOH_l3; // @[L2TLB.scala 94:21]
  wire  cache_io_refill_bits_levelOH_l2; // @[L2TLB.scala 94:21]
  wire  cache_io_refill_bits_levelOH_l1; // @[L2TLB.scala 94:21]
  wire [26:0] cache_io_refill_bits_req_info_dup_0_vpn; // @[L2TLB.scala 94:21]
  wire [1:0] cache_io_refill_bits_req_info_dup_0_source; // @[L2TLB.scala 94:21]
  wire [26:0] cache_io_refill_bits_req_info_dup_1_vpn; // @[L2TLB.scala 94:21]
  wire [1:0] cache_io_refill_bits_req_info_dup_1_source; // @[L2TLB.scala 94:21]
  wire [26:0] cache_io_refill_bits_req_info_dup_2_vpn; // @[L2TLB.scala 94:21]
  wire [1:0] cache_io_refill_bits_req_info_dup_2_source; // @[L2TLB.scala 94:21]
  wire [1:0] cache_io_refill_bits_level_dup_0; // @[L2TLB.scala 94:21]
  wire [1:0] cache_io_refill_bits_level_dup_1; // @[L2TLB.scala 94:21]
  wire [1:0] cache_io_refill_bits_level_dup_2; // @[L2TLB.scala 94:21]
  wire [63:0] cache_io_refill_bits_sel_pte_dup_0; // @[L2TLB.scala 94:21]
  wire [63:0] cache_io_refill_bits_sel_pte_dup_1; // @[L2TLB.scala 94:21]
  wire [63:0] cache_io_refill_bits_sel_pte_dup_2; // @[L2TLB.scala 94:21]
  wire  cache_io_sfence_dup_0_valid; // @[L2TLB.scala 94:21]
  wire  cache_io_sfence_dup_0_bits_rs1; // @[L2TLB.scala 94:21]
  wire  cache_io_sfence_dup_0_bits_rs2; // @[L2TLB.scala 94:21]
  wire [38:0] cache_io_sfence_dup_0_bits_addr; // @[L2TLB.scala 94:21]
  wire [15:0] cache_io_sfence_dup_0_bits_asid; // @[L2TLB.scala 94:21]
  wire  cache_io_sfence_dup_1_valid; // @[L2TLB.scala 94:21]
  wire  cache_io_sfence_dup_2_valid; // @[L2TLB.scala 94:21]
  wire  cache_io_sfence_dup_3_valid; // @[L2TLB.scala 94:21]
  wire  cache_io_sfence_dup_3_bits_rs1; // @[L2TLB.scala 94:21]
  wire  cache_io_sfence_dup_3_bits_rs2; // @[L2TLB.scala 94:21]
  wire [38:0] cache_io_sfence_dup_3_bits_addr; // @[L2TLB.scala 94:21]
  wire [15:0] cache_io_csr_dup_0_satp_asid; // @[L2TLB.scala 94:21]
  wire  cache_io_csr_dup_0_satp_changed; // @[L2TLB.scala 94:21]
  wire [15:0] cache_io_csr_dup_1_satp_asid; // @[L2TLB.scala 94:21]
  wire  cache_io_csr_dup_1_satp_changed; // @[L2TLB.scala 94:21]
  wire [15:0] cache_io_csr_dup_2_satp_asid; // @[L2TLB.scala 94:21]
  wire  cache_io_csr_dup_2_satp_changed; // @[L2TLB.scala 94:21]
  wire [5:0] cache_io_perf_0_value; // @[L2TLB.scala 94:21]
  wire [5:0] cache_io_perf_1_value; // @[L2TLB.scala 94:21]
  wire [5:0] cache_io_perf_2_value; // @[L2TLB.scala 94:21]
  wire [5:0] cache_io_perf_3_value; // @[L2TLB.scala 94:21]
  wire [5:0] cache_io_perf_4_value; // @[L2TLB.scala 94:21]
  wire [5:0] cache_io_perf_5_value; // @[L2TLB.scala 94:21]
  wire [5:0] cache_io_perf_6_value; // @[L2TLB.scala 94:21]
  wire [5:0] cache_io_perf_7_value; // @[L2TLB.scala 94:21]
  wire  ptw_clock; // @[L2TLB.scala 95:19]
  wire  ptw_reset; // @[L2TLB.scala 95:19]
  wire  ptw_io_sfence_valid; // @[L2TLB.scala 95:19]
  wire [15:0] ptw_io_csr_satp_asid; // @[L2TLB.scala 95:19]
  wire [43:0] ptw_io_csr_satp_ppn; // @[L2TLB.scala 95:19]
  wire  ptw_io_req_ready; // @[L2TLB.scala 95:19]
  wire  ptw_io_req_valid; // @[L2TLB.scala 95:19]
  wire [26:0] ptw_io_req_bits_req_info_vpn; // @[L2TLB.scala 95:19]
  wire [1:0] ptw_io_req_bits_req_info_source; // @[L2TLB.scala 95:19]
  wire  ptw_io_req_bits_l1Hit; // @[L2TLB.scala 95:19]
  wire [23:0] ptw_io_req_bits_ppn; // @[L2TLB.scala 95:19]
  wire  ptw_io_resp_ready; // @[L2TLB.scala 95:19]
  wire  ptw_io_resp_valid; // @[L2TLB.scala 95:19]
  wire [1:0] ptw_io_resp_bits_source; // @[L2TLB.scala 95:19]
  wire [26:0] ptw_io_resp_bits_resp_entry_tag; // @[L2TLB.scala 95:19]
  wire [15:0] ptw_io_resp_bits_resp_entry_asid; // @[L2TLB.scala 95:19]
  wire [23:0] ptw_io_resp_bits_resp_entry_ppn; // @[L2TLB.scala 95:19]
  wire  ptw_io_resp_bits_resp_entry_perm_d; // @[L2TLB.scala 95:19]
  wire  ptw_io_resp_bits_resp_entry_perm_a; // @[L2TLB.scala 95:19]
  wire  ptw_io_resp_bits_resp_entry_perm_g; // @[L2TLB.scala 95:19]
  wire  ptw_io_resp_bits_resp_entry_perm_u; // @[L2TLB.scala 95:19]
  wire  ptw_io_resp_bits_resp_entry_perm_x; // @[L2TLB.scala 95:19]
  wire  ptw_io_resp_bits_resp_entry_perm_w; // @[L2TLB.scala 95:19]
  wire  ptw_io_resp_bits_resp_entry_perm_r; // @[L2TLB.scala 95:19]
  wire [1:0] ptw_io_resp_bits_resp_entry_level; // @[L2TLB.scala 95:19]
  wire  ptw_io_resp_bits_resp_pf; // @[L2TLB.scala 95:19]
  wire  ptw_io_resp_bits_resp_af; // @[L2TLB.scala 95:19]
  wire  ptw_io_llptw_ready; // @[L2TLB.scala 95:19]
  wire  ptw_io_llptw_valid; // @[L2TLB.scala 95:19]
  wire [26:0] ptw_io_llptw_bits_req_info_vpn; // @[L2TLB.scala 95:19]
  wire [1:0] ptw_io_llptw_bits_req_info_source; // @[L2TLB.scala 95:19]
  wire  ptw_io_mem_req_ready; // @[L2TLB.scala 95:19]
  wire  ptw_io_mem_req_valid; // @[L2TLB.scala 95:19]
  wire [35:0] ptw_io_mem_req_bits_addr; // @[L2TLB.scala 95:19]
  wire  ptw_io_mem_resp_valid; // @[L2TLB.scala 95:19]
  wire [63:0] ptw_io_mem_resp_bits; // @[L2TLB.scala 95:19]
  wire  ptw_io_mem_mask; // @[L2TLB.scala 95:19]
  wire [35:0] ptw_io_pmp_req_bits_addr; // @[L2TLB.scala 95:19]
  wire  ptw_io_pmp_resp_ld; // @[L2TLB.scala 95:19]
  wire  ptw_io_pmp_resp_mmio; // @[L2TLB.scala 95:19]
  wire [26:0] ptw_io_refill_req_info_vpn; // @[L2TLB.scala 95:19]
  wire [1:0] ptw_io_refill_req_info_source; // @[L2TLB.scala 95:19]
  wire [1:0] ptw_io_refill_level; // @[L2TLB.scala 95:19]
  wire [5:0] ptw_io_perf_0_value; // @[L2TLB.scala 95:19]
  wire [5:0] ptw_io_perf_1_value; // @[L2TLB.scala 95:19]
  wire [5:0] ptw_io_perf_2_value; // @[L2TLB.scala 95:19]
  wire [5:0] ptw_io_perf_3_value; // @[L2TLB.scala 95:19]
  wire [5:0] ptw_io_perf_4_value; // @[L2TLB.scala 95:19]
  wire [5:0] ptw_io_perf_5_value; // @[L2TLB.scala 95:19]
  wire [5:0] ptw_io_perf_6_value; // @[L2TLB.scala 95:19]
  wire  llptw_clock; // @[L2TLB.scala 96:21]
  wire  llptw_reset; // @[L2TLB.scala 96:21]
  wire  llptw_io_sfence_valid; // @[L2TLB.scala 96:21]
  wire  llptw_io_csr_satp_changed; // @[L2TLB.scala 96:21]
  wire  llptw_io_in_ready; // @[L2TLB.scala 96:21]
  wire  llptw_io_in_valid; // @[L2TLB.scala 96:21]
  wire [26:0] llptw_io_in_bits_req_info_vpn; // @[L2TLB.scala 96:21]
  wire [1:0] llptw_io_in_bits_req_info_source; // @[L2TLB.scala 96:21]
  wire [35:0] llptw_io_in_bits_ppn; // @[L2TLB.scala 96:21]
  wire  llptw_io_out_ready; // @[L2TLB.scala 96:21]
  wire  llptw_io_out_valid; // @[L2TLB.scala 96:21]
  wire [26:0] llptw_io_out_bits_req_info_vpn; // @[L2TLB.scala 96:21]
  wire [1:0] llptw_io_out_bits_req_info_source; // @[L2TLB.scala 96:21]
  wire [2:0] llptw_io_out_bits_id; // @[L2TLB.scala 96:21]
  wire  llptw_io_out_bits_af; // @[L2TLB.scala 96:21]
  wire  llptw_io_mem_req_ready; // @[L2TLB.scala 96:21]
  wire  llptw_io_mem_req_valid; // @[L2TLB.scala 96:21]
  wire [35:0] llptw_io_mem_req_bits_addr; // @[L2TLB.scala 96:21]
  wire [2:0] llptw_io_mem_req_bits_id; // @[L2TLB.scala 96:21]
  wire  llptw_io_mem_resp_valid; // @[L2TLB.scala 96:21]
  wire [2:0] llptw_io_mem_resp_bits_id; // @[L2TLB.scala 96:21]
  wire [2:0] llptw_io_mem_enq_ptr; // @[L2TLB.scala 96:21]
  wire  llptw_io_mem_buffer_it_0; // @[L2TLB.scala 96:21]
  wire  llptw_io_mem_buffer_it_1; // @[L2TLB.scala 96:21]
  wire  llptw_io_mem_buffer_it_2; // @[L2TLB.scala 96:21]
  wire  llptw_io_mem_buffer_it_3; // @[L2TLB.scala 96:21]
  wire  llptw_io_mem_buffer_it_4; // @[L2TLB.scala 96:21]
  wire  llptw_io_mem_buffer_it_5; // @[L2TLB.scala 96:21]
  wire [26:0] llptw_io_mem_refill_vpn; // @[L2TLB.scala 96:21]
  wire [1:0] llptw_io_mem_refill_source; // @[L2TLB.scala 96:21]
  wire  llptw_io_mem_req_mask_0; // @[L2TLB.scala 96:21]
  wire  llptw_io_mem_req_mask_1; // @[L2TLB.scala 96:21]
  wire  llptw_io_mem_req_mask_2; // @[L2TLB.scala 96:21]
  wire  llptw_io_mem_req_mask_3; // @[L2TLB.scala 96:21]
  wire  llptw_io_mem_req_mask_4; // @[L2TLB.scala 96:21]
  wire  llptw_io_mem_req_mask_5; // @[L2TLB.scala 96:21]
  wire  llptw_io_cache_ready; // @[L2TLB.scala 96:21]
  wire  llptw_io_cache_valid; // @[L2TLB.scala 96:21]
  wire [26:0] llptw_io_cache_bits_vpn; // @[L2TLB.scala 96:21]
  wire [1:0] llptw_io_cache_bits_source; // @[L2TLB.scala 96:21]
  wire  llptw_io_pmp_req_valid; // @[L2TLB.scala 96:21]
  wire [35:0] llptw_io_pmp_req_bits_addr; // @[L2TLB.scala 96:21]
  wire  llptw_io_pmp_resp_ld; // @[L2TLB.scala 96:21]
  wire  llptw_io_pmp_resp_mmio; // @[L2TLB.scala 96:21]
  wire [5:0] llptw_io_perf_0_value; // @[L2TLB.scala 96:21]
  wire [5:0] llptw_io_perf_1_value; // @[L2TLB.scala 96:21]
  wire [5:0] llptw_io_perf_2_value; // @[L2TLB.scala 96:21]
  wire [5:0] llptw_io_perf_3_value; // @[L2TLB.scala 96:21]
  wire  arb1_io_in_0_ready; // @[L2TLB.scala 98:20]
  wire  arb1_io_in_0_valid; // @[L2TLB.scala 98:20]
  wire [26:0] arb1_io_in_0_bits_vpn; // @[L2TLB.scala 98:20]
  wire  arb1_io_in_1_ready; // @[L2TLB.scala 98:20]
  wire  arb1_io_in_1_valid; // @[L2TLB.scala 98:20]
  wire [26:0] arb1_io_in_1_bits_vpn; // @[L2TLB.scala 98:20]
  wire  arb1_io_out_ready; // @[L2TLB.scala 98:20]
  wire  arb1_io_out_valid; // @[L2TLB.scala 98:20]
  wire [26:0] arb1_io_out_bits_vpn; // @[L2TLB.scala 98:20]
  wire  arb1_io_chosen; // @[L2TLB.scala 98:20]
  wire  arb2_io_in_0_ready; // @[L2TLB.scala 99:20]
  wire  arb2_io_in_0_valid; // @[L2TLB.scala 99:20]
  wire [26:0] arb2_io_in_0_bits_vpn; // @[L2TLB.scala 99:20]
  wire [1:0] arb2_io_in_0_bits_source; // @[L2TLB.scala 99:20]
  wire  arb2_io_in_1_ready; // @[L2TLB.scala 99:20]
  wire  arb2_io_in_1_valid; // @[L2TLB.scala 99:20]
  wire [26:0] arb2_io_in_1_bits_vpn; // @[L2TLB.scala 99:20]
  wire [1:0] arb2_io_in_1_bits_source; // @[L2TLB.scala 99:20]
  wire  arb2_io_in_2_ready; // @[L2TLB.scala 99:20]
  wire  arb2_io_in_2_valid; // @[L2TLB.scala 99:20]
  wire [26:0] arb2_io_in_2_bits_vpn; // @[L2TLB.scala 99:20]
  wire [1:0] arb2_io_in_2_bits_source; // @[L2TLB.scala 99:20]
  wire  arb2_io_in_3_ready; // @[L2TLB.scala 99:20]
  wire  arb2_io_in_3_valid; // @[L2TLB.scala 99:20]
  wire [26:0] arb2_io_in_3_bits_vpn; // @[L2TLB.scala 99:20]
  wire  arb2_io_out_ready; // @[L2TLB.scala 99:20]
  wire  arb2_io_out_valid; // @[L2TLB.scala 99:20]
  wire [26:0] arb2_io_out_bits_vpn; // @[L2TLB.scala 99:20]
  wire [1:0] arb2_io_out_bits_source; // @[L2TLB.scala 99:20]
  wire [1:0] arb2_io_chosen; // @[L2TLB.scala 99:20]
  wire  Arbiter_io_in_0_ready; // @[L2TLB.scala 103:50]
  wire  Arbiter_io_in_0_valid; // @[L2TLB.scala 103:50]
  wire [26:0] Arbiter_io_in_0_bits_entry_tag; // @[L2TLB.scala 103:50]
  wire [15:0] Arbiter_io_in_0_bits_entry_asid; // @[L2TLB.scala 103:50]
  wire [23:0] Arbiter_io_in_0_bits_entry_ppn; // @[L2TLB.scala 103:50]
  wire  Arbiter_io_in_0_bits_entry_perm_d; // @[L2TLB.scala 103:50]
  wire  Arbiter_io_in_0_bits_entry_perm_a; // @[L2TLB.scala 103:50]
  wire  Arbiter_io_in_0_bits_entry_perm_g; // @[L2TLB.scala 103:50]
  wire  Arbiter_io_in_0_bits_entry_perm_u; // @[L2TLB.scala 103:50]
  wire  Arbiter_io_in_0_bits_entry_perm_x; // @[L2TLB.scala 103:50]
  wire  Arbiter_io_in_0_bits_entry_perm_w; // @[L2TLB.scala 103:50]
  wire  Arbiter_io_in_0_bits_entry_perm_r; // @[L2TLB.scala 103:50]
  wire [1:0] Arbiter_io_in_0_bits_entry_level; // @[L2TLB.scala 103:50]
  wire  Arbiter_io_in_0_bits_pf; // @[L2TLB.scala 103:50]
  wire  Arbiter_io_in_1_ready; // @[L2TLB.scala 103:50]
  wire  Arbiter_io_in_1_valid; // @[L2TLB.scala 103:50]
  wire [26:0] Arbiter_io_in_1_bits_entry_tag; // @[L2TLB.scala 103:50]
  wire [15:0] Arbiter_io_in_1_bits_entry_asid; // @[L2TLB.scala 103:50]
  wire [23:0] Arbiter_io_in_1_bits_entry_ppn; // @[L2TLB.scala 103:50]
  wire  Arbiter_io_in_1_bits_entry_perm_d; // @[L2TLB.scala 103:50]
  wire  Arbiter_io_in_1_bits_entry_perm_a; // @[L2TLB.scala 103:50]
  wire  Arbiter_io_in_1_bits_entry_perm_g; // @[L2TLB.scala 103:50]
  wire  Arbiter_io_in_1_bits_entry_perm_u; // @[L2TLB.scala 103:50]
  wire  Arbiter_io_in_1_bits_entry_perm_x; // @[L2TLB.scala 103:50]
  wire  Arbiter_io_in_1_bits_entry_perm_w; // @[L2TLB.scala 103:50]
  wire  Arbiter_io_in_1_bits_entry_perm_r; // @[L2TLB.scala 103:50]
  wire [1:0] Arbiter_io_in_1_bits_entry_level; // @[L2TLB.scala 103:50]
  wire  Arbiter_io_in_1_bits_pf; // @[L2TLB.scala 103:50]
  wire  Arbiter_io_in_1_bits_af; // @[L2TLB.scala 103:50]
  wire  Arbiter_io_in_2_ready; // @[L2TLB.scala 103:50]
  wire  Arbiter_io_in_2_valid; // @[L2TLB.scala 103:50]
  wire [26:0] Arbiter_io_in_2_bits_entry_tag; // @[L2TLB.scala 103:50]
  wire [15:0] Arbiter_io_in_2_bits_entry_asid; // @[L2TLB.scala 103:50]
  wire [23:0] Arbiter_io_in_2_bits_entry_ppn; // @[L2TLB.scala 103:50]
  wire  Arbiter_io_in_2_bits_entry_perm_d; // @[L2TLB.scala 103:50]
  wire  Arbiter_io_in_2_bits_entry_perm_a; // @[L2TLB.scala 103:50]
  wire  Arbiter_io_in_2_bits_entry_perm_g; // @[L2TLB.scala 103:50]
  wire  Arbiter_io_in_2_bits_entry_perm_u; // @[L2TLB.scala 103:50]
  wire  Arbiter_io_in_2_bits_entry_perm_x; // @[L2TLB.scala 103:50]
  wire  Arbiter_io_in_2_bits_entry_perm_w; // @[L2TLB.scala 103:50]
  wire  Arbiter_io_in_2_bits_entry_perm_r; // @[L2TLB.scala 103:50]
  wire  Arbiter_io_in_2_bits_pf; // @[L2TLB.scala 103:50]
  wire  Arbiter_io_in_2_bits_af; // @[L2TLB.scala 103:50]
  wire  Arbiter_io_out_ready; // @[L2TLB.scala 103:50]
  wire  Arbiter_io_out_valid; // @[L2TLB.scala 103:50]
  wire [26:0] Arbiter_io_out_bits_entry_tag; // @[L2TLB.scala 103:50]
  wire [15:0] Arbiter_io_out_bits_entry_asid; // @[L2TLB.scala 103:50]
  wire [23:0] Arbiter_io_out_bits_entry_ppn; // @[L2TLB.scala 103:50]
  wire  Arbiter_io_out_bits_entry_perm_d; // @[L2TLB.scala 103:50]
  wire  Arbiter_io_out_bits_entry_perm_a; // @[L2TLB.scala 103:50]
  wire  Arbiter_io_out_bits_entry_perm_g; // @[L2TLB.scala 103:50]
  wire  Arbiter_io_out_bits_entry_perm_u; // @[L2TLB.scala 103:50]
  wire  Arbiter_io_out_bits_entry_perm_x; // @[L2TLB.scala 103:50]
  wire  Arbiter_io_out_bits_entry_perm_w; // @[L2TLB.scala 103:50]
  wire  Arbiter_io_out_bits_entry_perm_r; // @[L2TLB.scala 103:50]
  wire [1:0] Arbiter_io_out_bits_entry_level; // @[L2TLB.scala 103:50]
  wire  Arbiter_io_out_bits_pf; // @[L2TLB.scala 103:50]
  wire  Arbiter_io_out_bits_af; // @[L2TLB.scala 103:50]
  wire  Arbiter_1_io_in_0_ready; // @[L2TLB.scala 103:50]
  wire  Arbiter_1_io_in_0_valid; // @[L2TLB.scala 103:50]
  wire [26:0] Arbiter_1_io_in_0_bits_entry_tag; // @[L2TLB.scala 103:50]
  wire [15:0] Arbiter_1_io_in_0_bits_entry_asid; // @[L2TLB.scala 103:50]
  wire [23:0] Arbiter_1_io_in_0_bits_entry_ppn; // @[L2TLB.scala 103:50]
  wire  Arbiter_1_io_in_0_bits_entry_perm_d; // @[L2TLB.scala 103:50]
  wire  Arbiter_1_io_in_0_bits_entry_perm_a; // @[L2TLB.scala 103:50]
  wire  Arbiter_1_io_in_0_bits_entry_perm_g; // @[L2TLB.scala 103:50]
  wire  Arbiter_1_io_in_0_bits_entry_perm_u; // @[L2TLB.scala 103:50]
  wire  Arbiter_1_io_in_0_bits_entry_perm_x; // @[L2TLB.scala 103:50]
  wire  Arbiter_1_io_in_0_bits_entry_perm_w; // @[L2TLB.scala 103:50]
  wire  Arbiter_1_io_in_0_bits_entry_perm_r; // @[L2TLB.scala 103:50]
  wire [1:0] Arbiter_1_io_in_0_bits_entry_level; // @[L2TLB.scala 103:50]
  wire  Arbiter_1_io_in_0_bits_pf; // @[L2TLB.scala 103:50]
  wire  Arbiter_1_io_in_1_ready; // @[L2TLB.scala 103:50]
  wire  Arbiter_1_io_in_1_valid; // @[L2TLB.scala 103:50]
  wire [26:0] Arbiter_1_io_in_1_bits_entry_tag; // @[L2TLB.scala 103:50]
  wire [15:0] Arbiter_1_io_in_1_bits_entry_asid; // @[L2TLB.scala 103:50]
  wire [23:0] Arbiter_1_io_in_1_bits_entry_ppn; // @[L2TLB.scala 103:50]
  wire  Arbiter_1_io_in_1_bits_entry_perm_d; // @[L2TLB.scala 103:50]
  wire  Arbiter_1_io_in_1_bits_entry_perm_a; // @[L2TLB.scala 103:50]
  wire  Arbiter_1_io_in_1_bits_entry_perm_g; // @[L2TLB.scala 103:50]
  wire  Arbiter_1_io_in_1_bits_entry_perm_u; // @[L2TLB.scala 103:50]
  wire  Arbiter_1_io_in_1_bits_entry_perm_x; // @[L2TLB.scala 103:50]
  wire  Arbiter_1_io_in_1_bits_entry_perm_w; // @[L2TLB.scala 103:50]
  wire  Arbiter_1_io_in_1_bits_entry_perm_r; // @[L2TLB.scala 103:50]
  wire [1:0] Arbiter_1_io_in_1_bits_entry_level; // @[L2TLB.scala 103:50]
  wire  Arbiter_1_io_in_1_bits_pf; // @[L2TLB.scala 103:50]
  wire  Arbiter_1_io_in_1_bits_af; // @[L2TLB.scala 103:50]
  wire  Arbiter_1_io_in_2_ready; // @[L2TLB.scala 103:50]
  wire  Arbiter_1_io_in_2_valid; // @[L2TLB.scala 103:50]
  wire [26:0] Arbiter_1_io_in_2_bits_entry_tag; // @[L2TLB.scala 103:50]
  wire [15:0] Arbiter_1_io_in_2_bits_entry_asid; // @[L2TLB.scala 103:50]
  wire [23:0] Arbiter_1_io_in_2_bits_entry_ppn; // @[L2TLB.scala 103:50]
  wire  Arbiter_1_io_in_2_bits_entry_perm_d; // @[L2TLB.scala 103:50]
  wire  Arbiter_1_io_in_2_bits_entry_perm_a; // @[L2TLB.scala 103:50]
  wire  Arbiter_1_io_in_2_bits_entry_perm_g; // @[L2TLB.scala 103:50]
  wire  Arbiter_1_io_in_2_bits_entry_perm_u; // @[L2TLB.scala 103:50]
  wire  Arbiter_1_io_in_2_bits_entry_perm_x; // @[L2TLB.scala 103:50]
  wire  Arbiter_1_io_in_2_bits_entry_perm_w; // @[L2TLB.scala 103:50]
  wire  Arbiter_1_io_in_2_bits_entry_perm_r; // @[L2TLB.scala 103:50]
  wire  Arbiter_1_io_in_2_bits_pf; // @[L2TLB.scala 103:50]
  wire  Arbiter_1_io_in_2_bits_af; // @[L2TLB.scala 103:50]
  wire  Arbiter_1_io_out_ready; // @[L2TLB.scala 103:50]
  wire  Arbiter_1_io_out_valid; // @[L2TLB.scala 103:50]
  wire [26:0] Arbiter_1_io_out_bits_entry_tag; // @[L2TLB.scala 103:50]
  wire [15:0] Arbiter_1_io_out_bits_entry_asid; // @[L2TLB.scala 103:50]
  wire [23:0] Arbiter_1_io_out_bits_entry_ppn; // @[L2TLB.scala 103:50]
  wire  Arbiter_1_io_out_bits_entry_perm_d; // @[L2TLB.scala 103:50]
  wire  Arbiter_1_io_out_bits_entry_perm_a; // @[L2TLB.scala 103:50]
  wire  Arbiter_1_io_out_bits_entry_perm_g; // @[L2TLB.scala 103:50]
  wire  Arbiter_1_io_out_bits_entry_perm_u; // @[L2TLB.scala 103:50]
  wire  Arbiter_1_io_out_bits_entry_perm_x; // @[L2TLB.scala 103:50]
  wire  Arbiter_1_io_out_bits_entry_perm_w; // @[L2TLB.scala 103:50]
  wire  Arbiter_1_io_out_bits_entry_perm_r; // @[L2TLB.scala 103:50]
  wire [1:0] Arbiter_1_io_out_bits_entry_level; // @[L2TLB.scala 103:50]
  wire  Arbiter_1_io_out_bits_pf; // @[L2TLB.scala 103:50]
  wire  Arbiter_1_io_out_bits_af; // @[L2TLB.scala 103:50]
  wire  prefetch_clock; // @[L2TLB.scala 127:26]
  wire  prefetch_reset; // @[L2TLB.scala 127:26]
  wire  prefetch_io_sfence_valid; // @[L2TLB.scala 127:26]
  wire  prefetch_io_csr_satp_changed; // @[L2TLB.scala 127:26]
  wire  prefetch_io_in_valid; // @[L2TLB.scala 127:26]
  wire [26:0] prefetch_io_in_bits_vpn; // @[L2TLB.scala 127:26]
  wire  prefetch_io_out_ready; // @[L2TLB.scala 127:26]
  wire  prefetch_io_out_valid; // @[L2TLB.scala 127:26]
  wire [26:0] prefetch_io_out_bits_vpn; // @[L2TLB.scala 127:26]
  wire  writer_clock; // @[ChiselDB.scala 132:24]
  wire  writer_reset; // @[ChiselDB.scala 132:24]
  wire  writer_en; // @[ChiselDB.scala 132:24]
  wire [63:0] writer_stamp; // @[ChiselDB.scala 132:24]
  wire [26:0] writer_data_vpn; // @[ChiselDB.scala 132:24]
  wire  mq_arb_io_in_0_ready; // @[L2TLB.scala 146:22]
  wire  mq_arb_io_in_0_valid; // @[L2TLB.scala 146:22]
  wire [26:0] mq_arb_io_in_0_bits_vpn; // @[L2TLB.scala 146:22]
  wire [1:0] mq_arb_io_in_0_bits_source; // @[L2TLB.scala 146:22]
  wire  mq_arb_io_in_1_ready; // @[L2TLB.scala 146:22]
  wire  mq_arb_io_in_1_valid; // @[L2TLB.scala 146:22]
  wire [26:0] mq_arb_io_in_1_bits_vpn; // @[L2TLB.scala 146:22]
  wire [1:0] mq_arb_io_in_1_bits_source; // @[L2TLB.scala 146:22]
  wire  mq_arb_io_out_ready; // @[L2TLB.scala 146:22]
  wire  mq_arb_io_out_valid; // @[L2TLB.scala 146:22]
  wire [26:0] mq_arb_io_out_bits_vpn; // @[L2TLB.scala 146:22]
  wire [1:0] mq_arb_io_out_bits_source; // @[L2TLB.scala 146:22]
  wire  mem_arb_io_in_0_valid; // @[L2TLB.scala 215:23]
  wire [35:0] mem_arb_io_in_0_bits_addr; // @[L2TLB.scala 215:23]
  wire  mem_arb_io_in_1_ready; // @[L2TLB.scala 215:23]
  wire  mem_arb_io_in_1_valid; // @[L2TLB.scala 215:23]
  wire [35:0] mem_arb_io_in_1_bits_addr; // @[L2TLB.scala 215:23]
  wire [2:0] mem_arb_io_in_1_bits_id; // @[L2TLB.scala 215:23]
  wire  mem_arb_io_out_ready; // @[L2TLB.scala 215:23]
  wire  mem_arb_io_out_valid; // @[L2TLB.scala 215:23]
  wire [35:0] mem_arb_io_out_bits_addr; // @[L2TLB.scala 215:23]
  wire [2:0] mem_arb_io_out_bits_id; // @[L2TLB.scala 215:23]
  wire  writer_1_clock; // @[ChiselDB.scala 132:24]
  wire  writer_1_reset; // @[ChiselDB.scala 132:24]
  wire  writer_1_en; // @[ChiselDB.scala 132:24]
  wire [63:0] writer_1_stamp; // @[ChiselDB.scala 132:24]
  wire [26:0] writer_1_data_vpn; // @[ChiselDB.scala 132:24]
  wire  writer_2_clock; // @[ChiselDB.scala 132:24]
  wire  writer_2_reset; // @[ChiselDB.scala 132:24]
  wire  writer_2_en; // @[ChiselDB.scala 132:24]
  wire [63:0] writer_2_stamp; // @[ChiselDB.scala 132:24]
  wire [26:0] writer_2_data_vpn; // @[ChiselDB.scala 132:24]
  wire  writer_3_clock; // @[ChiselDB.scala 132:24]
  wire  writer_3_reset; // @[ChiselDB.scala 132:24]
  wire  writer_3_en; // @[ChiselDB.scala 132:24]
  wire [63:0] writer_3_stamp; // @[ChiselDB.scala 132:24]
  wire [26:0] writer_3_data_vpn; // @[ChiselDB.scala 132:24]
  wire  writer_4_clock; // @[ChiselDB.scala 132:24]
  wire  writer_4_reset; // @[ChiselDB.scala 132:24]
  wire  writer_4_en; // @[ChiselDB.scala 132:24]
  wire [63:0] writer_4_stamp; // @[ChiselDB.scala 132:24]
  wire [26:0] writer_4_data_vpn; // @[ChiselDB.scala 132:24]
  wire  writer_5_clock; // @[ChiselDB.scala 132:24]
  wire  writer_5_reset; // @[ChiselDB.scala 132:24]
  wire  writer_5_en; // @[ChiselDB.scala 132:24]
  wire [63:0] writer_5_stamp; // @[ChiselDB.scala 132:24]
  wire [26:0] writer_5_data_vpn; // @[ChiselDB.scala 132:24]
  wire [1:0] writer_5_data_source; // @[ChiselDB.scala 132:24]
  wire  writer_5_data_bypassed; // @[ChiselDB.scala 132:24]
  wire  writer_5_data_is_first; // @[ChiselDB.scala 132:24]
  wire  writer_5_data_prefetched; // @[ChiselDB.scala 132:24]
  wire  writer_5_data_prefetch; // @[ChiselDB.scala 132:24]
  wire  writer_5_data_l2Hit; // @[ChiselDB.scala 132:24]
  wire  writer_5_data_l1Hit; // @[ChiselDB.scala 132:24]
  wire  writer_5_data_hit; // @[ChiselDB.scala 132:24]
  wire  writer_6_clock; // @[ChiselDB.scala 132:24]
  wire  writer_6_reset; // @[ChiselDB.scala 132:24]
  wire  writer_6_en; // @[ChiselDB.scala 132:24]
  wire [63:0] writer_6_stamp; // @[ChiselDB.scala 132:24]
  wire [26:0] writer_6_data_vpn; // @[ChiselDB.scala 132:24]
  wire [1:0] writer_6_data_source; // @[ChiselDB.scala 132:24]
  wire  writer_7_clock; // @[ChiselDB.scala 132:24]
  wire  writer_7_reset; // @[ChiselDB.scala 132:24]
  wire  writer_7_en; // @[ChiselDB.scala 132:24]
  wire [63:0] writer_7_stamp; // @[ChiselDB.scala 132:24]
  wire [26:0] writer_7_data_vpn; // @[ChiselDB.scala 132:24]
  wire [1:0] writer_7_data_source; // @[ChiselDB.scala 132:24]
  wire  writer_8_clock; // @[ChiselDB.scala 132:24]
  wire  writer_8_reset; // @[ChiselDB.scala 132:24]
  wire  writer_8_en; // @[ChiselDB.scala 132:24]
  wire [63:0] writer_8_stamp; // @[ChiselDB.scala 132:24]
  wire [26:0] writer_8_data_vpn; // @[ChiselDB.scala 132:24]
  wire [1:0] writer_8_data_source; // @[ChiselDB.scala 132:24]
  wire  writer_9_clock; // @[ChiselDB.scala 132:24]
  wire  writer_9_reset; // @[ChiselDB.scala 132:24]
  wire  writer_9_en; // @[ChiselDB.scala 132:24]
  wire [63:0] writer_9_stamp; // @[ChiselDB.scala 132:24]
  wire [26:0] writer_9_data_vpn; // @[ChiselDB.scala 132:24]
  wire [1:0] writer_9_data_source; // @[ChiselDB.scala 132:24]
  wire  writer_10_clock; // @[ChiselDB.scala 132:24]
  wire  writer_10_reset; // @[ChiselDB.scala 132:24]
  wire  writer_10_en; // @[ChiselDB.scala 132:24]
  wire [63:0] writer_10_stamp; // @[ChiselDB.scala 132:24]
  wire [26:0] writer_10_data_vpn; // @[ChiselDB.scala 132:24]
  wire  writer_11_clock; // @[ChiselDB.scala 132:24]
  wire  writer_11_reset; // @[ChiselDB.scala 132:24]
  wire  writer_11_en; // @[ChiselDB.scala 132:24]
  wire [63:0] writer_11_stamp; // @[ChiselDB.scala 132:24]
  wire [26:0] writer_11_data_vpn; // @[ChiselDB.scala 132:24]
  reg  sfence_dup_0_valid; // @[L2TLB.scala 82:39]
  reg  sfence_dup_1_valid; // @[L2TLB.scala 82:39]
  reg  sfence_dup_2_valid; // @[L2TLB.scala 82:39]
  reg  sfence_dup_2_bits_rs1; // @[L2TLB.scala 82:39]
  reg  sfence_dup_2_bits_rs2; // @[L2TLB.scala 82:39]
  reg [38:0] sfence_dup_2_bits_addr; // @[L2TLB.scala 82:39]
  reg [15:0] sfence_dup_2_bits_asid; // @[L2TLB.scala 82:39]
  reg  sfence_dup_3_valid; // @[L2TLB.scala 82:39]
  reg  sfence_dup_4_valid; // @[L2TLB.scala 82:39]
  reg  sfence_dup_5_valid; // @[L2TLB.scala 82:39]
  reg  sfence_dup_5_bits_rs1; // @[L2TLB.scala 82:39]
  reg  sfence_dup_5_bits_rs2; // @[L2TLB.scala 82:39]
  reg [38:0] sfence_dup_5_bits_addr; // @[L2TLB.scala 82:39]
  reg  sfence_dup_6_valid; // @[L2TLB.scala 82:39]
  reg  sfence_dup_7_valid; // @[L2TLB.scala 82:39]
  reg [15:0] csr_dup_0_satp_asid; // @[L2TLB.scala 83:36]
  reg  csr_dup_0_satp_changed; // @[L2TLB.scala 83:36]
  reg  csr_dup_1_satp_changed; // @[L2TLB.scala 83:36]
  reg [15:0] csr_dup_2_satp_asid; // @[L2TLB.scala 83:36]
  reg  csr_dup_2_satp_changed; // @[L2TLB.scala 83:36]
  reg [15:0] csr_dup_3_satp_asid; // @[L2TLB.scala 83:36]
  reg  csr_dup_3_satp_changed; // @[L2TLB.scala 83:36]
  reg [15:0] csr_dup_4_satp_asid; // @[L2TLB.scala 83:36]
  reg  csr_dup_4_satp_changed; // @[L2TLB.scala 83:36]
  reg  csr_dup_5_satp_changed; // @[L2TLB.scala 83:36]
  reg [15:0] csr_dup_6_satp_asid; // @[L2TLB.scala 83:36]
  reg [43:0] csr_dup_6_satp_ppn; // @[L2TLB.scala 83:36]
  wire  flush = sfence_dup_0_valid | csr_dup_0_satp_changed; // @[L2TLB.scala 86:36]
  wire  _T = ~ptw_io_req_ready; // @[L2TLB.scala 121:69]
  wire  _arb2_io_in_1_valid_T = ~_T; // @[L2TLB.scala 365:37]
  wire  _prefetch_io_in_valid_T = cache_io_resp_ready & cache_io_resp_valid; // @[Decoupled.scala 50:35]
  wire  _prefetch_io_in_valid_T_1 = cache_io_resp_bits_req_info_source == 2'h2; // @[MMUConst.scala 254:13]
  wire  _prefetch_io_in_valid_T_2 = ~_prefetch_io_in_valid_T_1; // @[L2TLB.scala 131:44]
  wire  _prefetch_io_in_valid_T_4 = ~cache_io_resp_bits_hit; // @[L2TLB.scala 131:85]
  wire  _prefetch_io_in_valid_T_6 = _prefetch_io_in_valid_T & ~_prefetch_io_in_valid_T_1 & (~cache_io_resp_bits_hit |
    cache_io_resp_bits_prefetch); // @[L2TLB.scala 131:81]
  reg [63:0] cnt; // @[ChiselDB.scala 133:22]
  wire  _mq_arb_io_in_0_valid_T_1 = cache_io_resp_valid & _prefetch_io_in_valid_T_4; // @[L2TLB.scala 147:48]
  wire  _mq_arb_io_in_0_valid_T_2 = ~cache_io_resp_bits_toFsm_l2Hit; // @[L2TLB.scala 148:6]
  wire  _mq_arb_io_in_0_valid_T_3 = ~cache_io_resp_bits_toFsm_l2Hit | cache_io_resp_bits_bypassed; // @[L2TLB.scala 148:38]
  wire  _mq_arb_io_in_0_valid_T_4 = cache_io_resp_valid & _prefetch_io_in_valid_T_4 & _mq_arb_io_in_0_valid_T_3; // @[L2TLB.scala 147:75]
  wire  _mq_arb_io_in_0_valid_T_7 = _mq_arb_io_in_0_valid_T_4 & _prefetch_io_in_valid_T_2; // @[L2TLB.scala 148:70]
  wire  _mq_arb_io_in_0_valid_T_8 = cache_io_resp_bits_bypassed | cache_io_resp_bits_isFirst; // @[L2TLB.scala 150:34]
  wire  _mq_arb_io_in_0_valid_T_10 = cache_io_resp_bits_bypassed | cache_io_resp_bits_isFirst | _T; // @[L2TLB.scala 150:64]
  wire  _llptw_io_in_valid_T_3 = ~cache_io_resp_bits_bypassed; // @[L2TLB.scala 160:108]
  wire  _cache_io_resp_ready_T_1 = 2'h0 == cache_io_resp_bits_req_info_source ? Arbiter_io_in_0_ready : 1'h1; // @[Mux.scala 81:58]
  wire  _cache_io_resp_ready_T_3 = 2'h1 == cache_io_resp_bits_req_info_source ? Arbiter_1_io_in_0_ready :
    _cache_io_resp_ready_T_1; // @[Mux.scala 81:58]
  wire  _cache_io_resp_ready_T_8 = _mq_arb_io_in_0_valid_T_8 ? mq_arb_io_in_0_ready : mq_arb_io_in_0_ready |
    ptw_io_req_ready; // @[L2TLB.scala 178:8]
  wire  _cache_io_resp_ready_T_9 = cache_io_resp_bits_toFsm_l2Hit & _llptw_io_in_valid_T_3 ? llptw_io_in_ready :
    _cache_io_resp_ready_T_8; // @[L2TLB.scala 177:8]
  wire  _ptw_io_req_valid_T_5 = _mq_arb_io_in_0_valid_T_1 & _mq_arb_io_in_0_valid_T_2 & _llptw_io_in_valid_T_3; // @[L2TLB.scala 181:105]
  wire  _ptw_io_req_valid_T_6 = ~cache_io_resp_bits_isFirst; // @[L2TLB.scala 183:5]
  wire  _ptw_io_resp_ready_T_1 = 2'h0 == ptw_io_resp_bits_source ? Arbiter_io_in_1_ready : 1'h1; // @[Mux.scala 81:58]
  reg  waiting_resp_0; // @[L2TLB.scala 204:29]
  reg  waiting_resp_1; // @[L2TLB.scala 204:29]
  reg  waiting_resp_2; // @[L2TLB.scala 204:29]
  reg  waiting_resp_3; // @[L2TLB.scala 204:29]
  reg  waiting_resp_4; // @[L2TLB.scala 204:29]
  reg  waiting_resp_5; // @[L2TLB.scala 204:29]
  reg  waiting_resp_6; // @[L2TLB.scala 204:29]
  reg  flush_latch_0; // @[L2TLB.scala 205:28]
  reg  flush_latch_1; // @[L2TLB.scala 205:28]
  reg  flush_latch_2; // @[L2TLB.scala 205:28]
  reg  flush_latch_3; // @[L2TLB.scala 205:28]
  reg  flush_latch_4; // @[L2TLB.scala 205:28]
  reg  flush_latch_5; // @[L2TLB.scala 205:28]
  reg  flush_latch_6; // @[L2TLB.scala 205:28]
  wire  _mem_arb_io_out_ready_T = ~flush; // @[L2TLB.scala 218:42]
  reg [2:0] req_addr_low_0; // @[L2TLB.scala 235:25]
  reg [2:0] req_addr_low_1; // @[L2TLB.scala 235:25]
  reg [2:0] req_addr_low_2; // @[L2TLB.scala 235:25]
  reg [2:0] req_addr_low_3; // @[L2TLB.scala 235:25]
  reg [2:0] req_addr_low_4; // @[L2TLB.scala 235:25]
  reg [2:0] req_addr_low_5; // @[L2TLB.scala 235:25]
  reg [2:0] req_addr_low_6; // @[L2TLB.scala 235:25]
  wire  _T_42 = llptw_io_in_ready & llptw_io_in_valid; // @[Decoupled.scala 50:35]
  wire [2:0] _GEN_4 = 3'h0 == llptw_io_mem_enq_ptr ? llptw_io_in_bits_req_info_vpn[2:0] : req_addr_low_0; // @[L2TLB.scala 235:25 239:{37,37}]
  wire [2:0] _GEN_5 = 3'h1 == llptw_io_mem_enq_ptr ? llptw_io_in_bits_req_info_vpn[2:0] : req_addr_low_1; // @[L2TLB.scala 235:25 239:{37,37}]
  wire [2:0] _GEN_6 = 3'h2 == llptw_io_mem_enq_ptr ? llptw_io_in_bits_req_info_vpn[2:0] : req_addr_low_2; // @[L2TLB.scala 235:25 239:{37,37}]
  wire [2:0] _GEN_7 = 3'h3 == llptw_io_mem_enq_ptr ? llptw_io_in_bits_req_info_vpn[2:0] : req_addr_low_3; // @[L2TLB.scala 235:25 239:{37,37}]
  wire [2:0] _GEN_8 = 3'h4 == llptw_io_mem_enq_ptr ? llptw_io_in_bits_req_info_vpn[2:0] : req_addr_low_4; // @[L2TLB.scala 235:25 239:{37,37}]
  wire [2:0] _GEN_9 = 3'h5 == llptw_io_mem_enq_ptr ? llptw_io_in_bits_req_info_vpn[2:0] : req_addr_low_5; // @[L2TLB.scala 235:25 239:{37,37}]
  wire [2:0] _GEN_10 = 3'h6 == llptw_io_mem_enq_ptr ? llptw_io_in_bits_req_info_vpn[2:0] : req_addr_low_6; // @[L2TLB.scala 235:25 239:{37,37}]
  wire [2:0] _GEN_11 = _T_42 ? _GEN_4 : req_addr_low_0; // @[L2TLB.scala 235:25 237:29]
  wire [2:0] _GEN_12 = _T_42 ? _GEN_5 : req_addr_low_1; // @[L2TLB.scala 235:25 237:29]
  wire [2:0] _GEN_13 = _T_42 ? _GEN_6 : req_addr_low_2; // @[L2TLB.scala 235:25 237:29]
  wire [2:0] _GEN_14 = _T_42 ? _GEN_7 : req_addr_low_3; // @[L2TLB.scala 235:25 237:29]
  wire [2:0] _GEN_15 = _T_42 ? _GEN_8 : req_addr_low_4; // @[L2TLB.scala 235:25 237:29]
  wire [2:0] _GEN_16 = _T_42 ? _GEN_9 : req_addr_low_5; // @[L2TLB.scala 235:25 237:29]
  wire [2:0] _GEN_17 = _T_42 ? _GEN_10 : req_addr_low_6; // @[L2TLB.scala 235:25 237:29]
  wire  _T_43 = mem_arb_io_out_ready & mem_arb_io_out_valid; // @[Decoupled.scala 50:35]
  wire  _GEN_25 = 3'h0 == mem_arb_io_out_bits_id | waiting_resp_0; // @[L2TLB.scala 204:29 243:{42,42}]
  wire  _GEN_26 = 3'h1 == mem_arb_io_out_bits_id | waiting_resp_1; // @[L2TLB.scala 204:29 243:{42,42}]
  wire  _GEN_27 = 3'h2 == mem_arb_io_out_bits_id | waiting_resp_2; // @[L2TLB.scala 204:29 243:{42,42}]
  wire  _GEN_28 = 3'h3 == mem_arb_io_out_bits_id | waiting_resp_3; // @[L2TLB.scala 204:29 243:{42,42}]
  wire  _GEN_29 = 3'h4 == mem_arb_io_out_bits_id | waiting_resp_4; // @[L2TLB.scala 204:29 243:{42,42}]
  wire  _GEN_30 = 3'h5 == mem_arb_io_out_bits_id | waiting_resp_5; // @[L2TLB.scala 204:29 243:{42,42}]
  wire  _GEN_31 = 3'h6 == mem_arb_io_out_bits_id | waiting_resp_6; // @[L2TLB.scala 204:29 243:{42,42}]
  wire  _GEN_39 = _T_43 ? _GEN_25 : waiting_resp_0; // @[L2TLB.scala 204:29 241:32]
  wire  _GEN_40 = _T_43 ? _GEN_26 : waiting_resp_1; // @[L2TLB.scala 204:29 241:32]
  wire  _GEN_41 = _T_43 ? _GEN_27 : waiting_resp_2; // @[L2TLB.scala 204:29 241:32]
  wire  _GEN_42 = _T_43 ? _GEN_28 : waiting_resp_3; // @[L2TLB.scala 204:29 241:32]
  wire  _GEN_43 = _T_43 ? _GEN_29 : waiting_resp_4; // @[L2TLB.scala 204:29 241:32]
  wire  _GEN_44 = _T_43 ? _GEN_30 : waiting_resp_5; // @[L2TLB.scala 204:29 241:32]
  wire  _GEN_45 = _T_43 ? _GEN_31 : waiting_resp_6; // @[L2TLB.scala 204:29 241:32]
  reg [255:0] refill_data_0; // @[L2TLB.scala 256:24]
  reg [255:0] refill_data_1; // @[L2TLB.scala 256:24]
  wire [12:0] _beats1_decode_T_1 = 13'h3f << auto_out_d_bits_size; // @[package.scala 234:77]
  wire [5:0] _beats1_decode_T_3 = ~_beats1_decode_T_1[5:0]; // @[package.scala 234:46]
  wire  beats1_decode = _beats1_decode_T_3[5]; // @[Edges.scala 219:59]
  wire  beats1_opdata = auto_out_d_bits_opcode[0]; // @[Edges.scala 105:36]
  wire  beats1 = beats1_opdata & beats1_decode; // @[Edges.scala 220:14]
  reg  counter; // @[Edges.scala 228:27]
  wire  counter1 = counter - 1'h1; // @[Edges.scala 229:28]
  wire  first = ~counter; // @[Edges.scala 230:25]
  wire  last = counter | ~beats1; // @[Edges.scala 231:37]
  wire  mem_resp_done = last & auto_out_d_valid; // @[Edges.scala 232:22]
  wire  count = beats1 & ~counter1; // @[Edges.scala 233:25]
  wire  mem_resp_from_mq = auto_out_d_bits_source != 3'h6; // @[L2TLB.scala 202:9]
  wire [255:0] _GEN_47 = ~count ? auto_out_d_bits_data : refill_data_0; // @[L2TLB.scala 256:24 262:{35,35}]
  wire [255:0] _GEN_48 = count ? auto_out_d_bits_data : refill_data_1; // @[L2TLB.scala 256:24 262:{35,35}]
  wire [511:0] _resp_pte_inner_data_T = {refill_data_1,refill_data_0}; // @[L2TLB.scala 371:35]
  wire [63:0] inner_data__0 = _resp_pte_inner_data_T[63:0]; // @[L2TLB.scala 371:35]
  wire [63:0] inner_data__1 = _resp_pte_inner_data_T[127:64]; // @[L2TLB.scala 371:35]
  wire [63:0] inner_data__2 = _resp_pte_inner_data_T[191:128]; // @[L2TLB.scala 371:35]
  wire [63:0] inner_data__3 = _resp_pte_inner_data_T[255:192]; // @[L2TLB.scala 371:35]
  wire [63:0] inner_data__4 = _resp_pte_inner_data_T[319:256]; // @[L2TLB.scala 371:35]
  wire [63:0] inner_data__5 = _resp_pte_inner_data_T[383:320]; // @[L2TLB.scala 371:35]
  wire [63:0] inner_data__6 = _resp_pte_inner_data_T[447:384]; // @[L2TLB.scala 371:35]
  wire [63:0] inner_data__7 = _resp_pte_inner_data_T[511:448]; // @[L2TLB.scala 371:35]
  reg [63:0] resp_pte_r; // @[Reg.scala 16:16]
  wire [63:0] _GEN_54 = 3'h1 == req_addr_low_0 ? inner_data__1 : inner_data__0; // @[Reg.scala 17:{22,22}]
  wire [63:0] _GEN_55 = 3'h2 == req_addr_low_0 ? inner_data__2 : _GEN_54; // @[Reg.scala 17:{22,22}]
  wire [63:0] _GEN_56 = 3'h3 == req_addr_low_0 ? inner_data__3 : _GEN_55; // @[Reg.scala 17:{22,22}]
  wire [63:0] _GEN_57 = 3'h4 == req_addr_low_0 ? inner_data__4 : _GEN_56; // @[Reg.scala 17:{22,22}]
  wire [63:0] _GEN_58 = 3'h5 == req_addr_low_0 ? inner_data__5 : _GEN_57; // @[Reg.scala 17:{22,22}]
  wire [63:0] _GEN_59 = 3'h6 == req_addr_low_0 ? inner_data__6 : _GEN_58; // @[Reg.scala 17:{22,22}]
  wire [63:0] _GEN_60 = 3'h7 == req_addr_low_0 ? inner_data__7 : _GEN_59; // @[Reg.scala 17:{22,22}]
  wire [63:0] _GEN_61 = llptw_io_mem_buffer_it_0 ? _GEN_60 : resp_pte_r; // @[Reg.scala 16:16 17:{18,22}]
  reg [63:0] resp_pte_r1; // @[Reg.scala 16:16]
  wire [63:0] _GEN_63 = 3'h1 == req_addr_low_1 ? inner_data__1 : inner_data__0; // @[Reg.scala 17:{22,22}]
  wire [63:0] _GEN_64 = 3'h2 == req_addr_low_1 ? inner_data__2 : _GEN_63; // @[Reg.scala 17:{22,22}]
  wire [63:0] _GEN_65 = 3'h3 == req_addr_low_1 ? inner_data__3 : _GEN_64; // @[Reg.scala 17:{22,22}]
  wire [63:0] _GEN_66 = 3'h4 == req_addr_low_1 ? inner_data__4 : _GEN_65; // @[Reg.scala 17:{22,22}]
  wire [63:0] _GEN_67 = 3'h5 == req_addr_low_1 ? inner_data__5 : _GEN_66; // @[Reg.scala 17:{22,22}]
  wire [63:0] _GEN_68 = 3'h6 == req_addr_low_1 ? inner_data__6 : _GEN_67; // @[Reg.scala 17:{22,22}]
  wire [63:0] _GEN_69 = 3'h7 == req_addr_low_1 ? inner_data__7 : _GEN_68; // @[Reg.scala 17:{22,22}]
  wire [63:0] _GEN_70 = llptw_io_mem_buffer_it_1 ? _GEN_69 : resp_pte_r1; // @[Reg.scala 16:16 17:{18,22}]
  reg [63:0] resp_pte_r2; // @[Reg.scala 16:16]
  wire [63:0] _GEN_72 = 3'h1 == req_addr_low_2 ? inner_data__1 : inner_data__0; // @[Reg.scala 17:{22,22}]
  wire [63:0] _GEN_73 = 3'h2 == req_addr_low_2 ? inner_data__2 : _GEN_72; // @[Reg.scala 17:{22,22}]
  wire [63:0] _GEN_74 = 3'h3 == req_addr_low_2 ? inner_data__3 : _GEN_73; // @[Reg.scala 17:{22,22}]
  wire [63:0] _GEN_75 = 3'h4 == req_addr_low_2 ? inner_data__4 : _GEN_74; // @[Reg.scala 17:{22,22}]
  wire [63:0] _GEN_76 = 3'h5 == req_addr_low_2 ? inner_data__5 : _GEN_75; // @[Reg.scala 17:{22,22}]
  wire [63:0] _GEN_77 = 3'h6 == req_addr_low_2 ? inner_data__6 : _GEN_76; // @[Reg.scala 17:{22,22}]
  wire [63:0] _GEN_78 = 3'h7 == req_addr_low_2 ? inner_data__7 : _GEN_77; // @[Reg.scala 17:{22,22}]
  wire [63:0] _GEN_79 = llptw_io_mem_buffer_it_2 ? _GEN_78 : resp_pte_r2; // @[Reg.scala 16:16 17:{18,22}]
  reg [63:0] resp_pte_r3; // @[Reg.scala 16:16]
  wire [63:0] _GEN_81 = 3'h1 == req_addr_low_3 ? inner_data__1 : inner_data__0; // @[Reg.scala 17:{22,22}]
  wire [63:0] _GEN_82 = 3'h2 == req_addr_low_3 ? inner_data__2 : _GEN_81; // @[Reg.scala 17:{22,22}]
  wire [63:0] _GEN_83 = 3'h3 == req_addr_low_3 ? inner_data__3 : _GEN_82; // @[Reg.scala 17:{22,22}]
  wire [63:0] _GEN_84 = 3'h4 == req_addr_low_3 ? inner_data__4 : _GEN_83; // @[Reg.scala 17:{22,22}]
  wire [63:0] _GEN_85 = 3'h5 == req_addr_low_3 ? inner_data__5 : _GEN_84; // @[Reg.scala 17:{22,22}]
  wire [63:0] _GEN_86 = 3'h6 == req_addr_low_3 ? inner_data__6 : _GEN_85; // @[Reg.scala 17:{22,22}]
  wire [63:0] _GEN_87 = 3'h7 == req_addr_low_3 ? inner_data__7 : _GEN_86; // @[Reg.scala 17:{22,22}]
  wire [63:0] _GEN_88 = llptw_io_mem_buffer_it_3 ? _GEN_87 : resp_pte_r3; // @[Reg.scala 16:16 17:{18,22}]
  reg [63:0] resp_pte_r4; // @[Reg.scala 16:16]
  wire [63:0] _GEN_90 = 3'h1 == req_addr_low_4 ? inner_data__1 : inner_data__0; // @[Reg.scala 17:{22,22}]
  wire [63:0] _GEN_91 = 3'h2 == req_addr_low_4 ? inner_data__2 : _GEN_90; // @[Reg.scala 17:{22,22}]
  wire [63:0] _GEN_92 = 3'h3 == req_addr_low_4 ? inner_data__3 : _GEN_91; // @[Reg.scala 17:{22,22}]
  wire [63:0] _GEN_93 = 3'h4 == req_addr_low_4 ? inner_data__4 : _GEN_92; // @[Reg.scala 17:{22,22}]
  wire [63:0] _GEN_94 = 3'h5 == req_addr_low_4 ? inner_data__5 : _GEN_93; // @[Reg.scala 17:{22,22}]
  wire [63:0] _GEN_95 = 3'h6 == req_addr_low_4 ? inner_data__6 : _GEN_94; // @[Reg.scala 17:{22,22}]
  wire [63:0] _GEN_96 = 3'h7 == req_addr_low_4 ? inner_data__7 : _GEN_95; // @[Reg.scala 17:{22,22}]
  wire [63:0] _GEN_97 = llptw_io_mem_buffer_it_4 ? _GEN_96 : resp_pte_r4; // @[Reg.scala 16:16 17:{18,22}]
  reg [63:0] resp_pte_r5; // @[Reg.scala 16:16]
  wire [63:0] _GEN_99 = 3'h1 == req_addr_low_5 ? inner_data__1 : inner_data__0; // @[Reg.scala 17:{22,22}]
  wire [63:0] _GEN_100 = 3'h2 == req_addr_low_5 ? inner_data__2 : _GEN_99; // @[Reg.scala 17:{22,22}]
  wire [63:0] _GEN_101 = 3'h3 == req_addr_low_5 ? inner_data__3 : _GEN_100; // @[Reg.scala 17:{22,22}]
  wire [63:0] _GEN_102 = 3'h4 == req_addr_low_5 ? inner_data__4 : _GEN_101; // @[Reg.scala 17:{22,22}]
  wire [63:0] _GEN_103 = 3'h5 == req_addr_low_5 ? inner_data__5 : _GEN_102; // @[Reg.scala 17:{22,22}]
  wire [63:0] _GEN_104 = 3'h6 == req_addr_low_5 ? inner_data__6 : _GEN_103; // @[Reg.scala 17:{22,22}]
  wire [63:0] _GEN_105 = 3'h7 == req_addr_low_5 ? inner_data__7 : _GEN_104; // @[Reg.scala 17:{22,22}]
  wire [63:0] _GEN_106 = llptw_io_mem_buffer_it_5 ? _GEN_105 : resp_pte_r5; // @[Reg.scala 16:16 17:{18,22}]
  wire [511:0] _resp_pte_inner_data_T_54 = {_GEN_48,_GEN_47}; // @[L2TLB.scala 371:35]
  wire [63:0] inner_data_6_0 = _resp_pte_inner_data_T_54[63:0]; // @[L2TLB.scala 371:35]
  wire [63:0] inner_data_6_1 = _resp_pte_inner_data_T_54[127:64]; // @[L2TLB.scala 371:35]
  wire [63:0] inner_data_6_2 = _resp_pte_inner_data_T_54[191:128]; // @[L2TLB.scala 371:35]
  wire [63:0] inner_data_6_3 = _resp_pte_inner_data_T_54[255:192]; // @[L2TLB.scala 371:35]
  wire [63:0] inner_data_6_4 = _resp_pte_inner_data_T_54[319:256]; // @[L2TLB.scala 371:35]
  wire [63:0] inner_data_6_5 = _resp_pte_inner_data_T_54[383:320]; // @[L2TLB.scala 371:35]
  wire [63:0] inner_data_6_6 = _resp_pte_inner_data_T_54[447:384]; // @[L2TLB.scala 371:35]
  wire [63:0] inner_data_6_7 = _resp_pte_inner_data_T_54[511:448]; // @[L2TLB.scala 371:35]
  wire  _resp_pte_T_6 = ~mem_resp_from_mq; // @[L2TLB.scala 271:109]
  wire  _resp_pte_T_7 = mem_resp_done & ~mem_resp_from_mq; // @[L2TLB.scala 271:106]
  reg [63:0] resp_pte_r6; // @[Reg.scala 16:16]
  wire [63:0] _GEN_108 = 3'h1 == req_addr_low_6 ? inner_data_6_1 : inner_data_6_0; // @[Reg.scala 17:{22,22}]
  wire [63:0] _GEN_109 = 3'h2 == req_addr_low_6 ? inner_data_6_2 : _GEN_108; // @[Reg.scala 17:{22,22}]
  wire [63:0] _GEN_110 = 3'h3 == req_addr_low_6 ? inner_data_6_3 : _GEN_109; // @[Reg.scala 17:{22,22}]
  wire [63:0] _GEN_111 = 3'h4 == req_addr_low_6 ? inner_data_6_4 : _GEN_110; // @[Reg.scala 17:{22,22}]
  reg [2:0] llptw_io_mem_resp_bits_id_r; // @[Reg.scala 16:16]
  wire  _refill_level_T = ptw_io_mem_req_ready & ptw_io_mem_req_valid; // @[Decoupled.scala 50:35]
  reg [1:0] refill_level_r; // @[Reg.scala 28:20]
  wire [1:0] refill_level = mem_resp_from_mq ? 2'h2 : refill_level_r; // @[L2TLB.scala 285:25]
  wire  _GEN_119 = 3'h1 == auto_out_d_bits_source ? flush_latch_1 : flush_latch_0; // @[L2TLB.scala 286:{49,49}]
  wire  _GEN_120 = 3'h2 == auto_out_d_bits_source ? flush_latch_2 : _GEN_119; // @[L2TLB.scala 286:{49,49}]
  wire  _GEN_121 = 3'h3 == auto_out_d_bits_source ? flush_latch_3 : _GEN_120; // @[L2TLB.scala 286:{49,49}]
  wire  _GEN_122 = 3'h4 == auto_out_d_bits_source ? flush_latch_4 : _GEN_121; // @[L2TLB.scala 286:{49,49}]
  wire  _GEN_123 = 3'h5 == auto_out_d_bits_source ? flush_latch_5 : _GEN_122; // @[L2TLB.scala 286:{49,49}]
  wire  _GEN_124 = 3'h6 == auto_out_d_bits_source ? flush_latch_6 : _GEN_123; // @[L2TLB.scala 286:{49,49}]
  wire  refill_valid = mem_resp_done & _mem_arb_io_out_ready_T & ~_GEN_124; // @[L2TLB.scala 286:46]
  reg  cache_io_refill_valid_REG; // @[L2TLB.scala 288:35]
  reg [26:0] cache_io_refill_bits_req_info_dup_0_rvpn; // @[Reg.scala 16:16]
  reg [1:0] cache_io_refill_bits_req_info_dup_0_rsource; // @[Reg.scala 16:16]
  reg [26:0] cache_io_refill_bits_req_info_dup_1_rvpn; // @[Reg.scala 16:16]
  reg [1:0] cache_io_refill_bits_req_info_dup_1_rsource; // @[Reg.scala 16:16]
  reg [26:0] cache_io_refill_bits_req_info_dup_2_rvpn; // @[Reg.scala 16:16]
  reg [1:0] cache_io_refill_bits_req_info_dup_2_rsource; // @[Reg.scala 16:16]
  reg [1:0] cache_io_refill_bits_level_dup_0_r; // @[Reg.scala 16:16]
  reg [1:0] cache_io_refill_bits_level_dup_1_r; // @[Reg.scala 16:16]
  reg [1:0] cache_io_refill_bits_level_dup_2_r; // @[Reg.scala 16:16]
  wire  _cache_io_refill_bits_levelOH_sp_T = refill_level == 2'h0; // @[PageTableCache.scala 94:34]
  wire  _cache_io_refill_bits_levelOH_sp_T_1 = refill_level == 2'h1; // @[PageTableCache.scala 94:55]
  reg  cache_io_refill_bits_levelOH_sp_REG; // @[PageTableCache.scala 94:22]
  reg  cache_io_refill_bits_levelOH_l3_REG; // @[PageTableCache.scala 95:22]
  reg  cache_io_refill_bits_levelOH_l2_REG; // @[PageTableCache.scala 96:22]
  reg  cache_io_refill_bits_levelOH_l1_REG; // @[PageTableCache.scala 97:22]
  reg [63:0] cache_io_refill_bits_sel_pte_dup_0_REG; // @[L2TLB.scala 293:52]
  wire [2:0] _GEN_135 = 3'h1 == auto_out_d_bits_source ? req_addr_low_1 : req_addr_low_0; // @[L2TLB.scala 293:{52,52}]
  wire [2:0] _GEN_136 = 3'h2 == auto_out_d_bits_source ? req_addr_low_2 : _GEN_135; // @[L2TLB.scala 293:{52,52}]
  wire [2:0] _GEN_137 = 3'h3 == auto_out_d_bits_source ? req_addr_low_3 : _GEN_136; // @[L2TLB.scala 293:{52,52}]
  wire [2:0] _GEN_138 = 3'h4 == auto_out_d_bits_source ? req_addr_low_4 : _GEN_137; // @[L2TLB.scala 293:{52,52}]
  wire [2:0] _GEN_139 = 3'h5 == auto_out_d_bits_source ? req_addr_low_5 : _GEN_138; // @[L2TLB.scala 293:{52,52}]
  wire [2:0] _GEN_140 = 3'h6 == auto_out_d_bits_source ? req_addr_low_6 : _GEN_139; // @[L2TLB.scala 293:{52,52}]
  wire [63:0] _GEN_142 = 3'h1 == _GEN_140 ? inner_data_6_1 : inner_data_6_0; // @[L2TLB.scala 293:{52,52}]
  wire [63:0] _GEN_143 = 3'h2 == _GEN_140 ? inner_data_6_2 : _GEN_142; // @[L2TLB.scala 293:{52,52}]
  wire [63:0] _GEN_144 = 3'h3 == _GEN_140 ? inner_data_6_3 : _GEN_143; // @[L2TLB.scala 293:{52,52}]
  reg [63:0] cache_io_refill_bits_sel_pte_dup_1_REG; // @[L2TLB.scala 293:52]
  reg [63:0] cache_io_refill_bits_sel_pte_dup_2_REG; // @[L2TLB.scala 293:52]
  wire  _llptw_io_out_ready_T_1 = 2'h0 == llptw_io_out_bits_req_info_source ? Arbiter_io_in_2_ready : 1'h1; // @[Mux.scala 81:58]
  wire [63:0] _GEN_166 = 3'h1 == llptw_io_out_bits_id ? _GEN_70 : _GEN_61; // @[]
  wire [63:0] _GEN_167 = 3'h2 == llptw_io_out_bits_id ? _GEN_79 : _GEN_166; // @[]
  wire [63:0] _GEN_168 = 3'h3 == llptw_io_out_bits_id ? _GEN_88 : _GEN_167; // @[]
  wire [63:0] _GEN_169 = 3'h4 == llptw_io_out_bits_id ? _GEN_97 : _GEN_168; // @[]
  wire [63:0] _GEN_170 = 3'h5 == llptw_io_out_bits_id ? _GEN_106 : _GEN_169; // @[]
  wire [63:0] _GEN_171 = 3'h6 == llptw_io_out_bits_id ? resp_pte_r6 : _GEN_170; // @[]
  wire  pte_in_perm_v = _GEN_171[0]; // @[L2TLB.scala 376:30]
  wire  pte_in_perm_r = _GEN_171[1]; // @[L2TLB.scala 376:30]
  wire  pte_in_perm_w = _GEN_171[2]; // @[L2TLB.scala 376:30]
  wire [19:0] pte_in_ppn_high = _GEN_171[53:34]; // @[L2TLB.scala 376:30]
  wire  _ptw_resp_pf_T_4 = ~pte_in_perm_v | ~pte_in_perm_r & pte_in_perm_w; // @[MMUBundle.scala 522:13]
  wire  _ptw_resp_af_T_1 = ~(pte_in_ppn_high == 20'h0); // @[MMUBundle.scala 528:5]
  wire  _GEN_172 = waiting_resp_0 | flush_latch_0; // @[L2TLB.scala 352:30 353:24 205:28]
  wire  _GEN_173 = waiting_resp_1 | flush_latch_1; // @[L2TLB.scala 352:30 353:24 205:28]
  wire  _GEN_174 = waiting_resp_2 | flush_latch_2; // @[L2TLB.scala 352:30 353:24 205:28]
  wire  _GEN_175 = waiting_resp_3 | flush_latch_3; // @[L2TLB.scala 352:30 353:24 205:28]
  wire  _GEN_176 = waiting_resp_4 | flush_latch_4; // @[L2TLB.scala 352:30 353:24 205:28]
  wire  _GEN_177 = waiting_resp_5 | flush_latch_5; // @[L2TLB.scala 352:30 353:24 205:28]
  wire  _GEN_178 = waiting_resp_6 | flush_latch_6; // @[L2TLB.scala 352:30 353:24 205:28]
  wire  _GEN_179 = flush ? _GEN_172 : flush_latch_0; // @[L2TLB.scala 350:16 205:28]
  wire  _GEN_180 = flush ? _GEN_173 : flush_latch_1; // @[L2TLB.scala 350:16 205:28]
  wire  _GEN_181 = flush ? _GEN_174 : flush_latch_2; // @[L2TLB.scala 350:16 205:28]
  wire  _GEN_182 = flush ? _GEN_175 : flush_latch_3; // @[L2TLB.scala 350:16 205:28]
  wire  _GEN_183 = flush ? _GEN_176 : flush_latch_4; // @[L2TLB.scala 350:16 205:28]
  wire  _GEN_184 = flush ? _GEN_177 : flush_latch_5; // @[L2TLB.scala 350:16 205:28]
  wire  _GEN_185 = flush ? _GEN_178 : flush_latch_6; // @[L2TLB.scala 350:16 205:28]
  reg [5:0] io_perf_0_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg [5:0] io_perf_0_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg [5:0] io_perf_1_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg [5:0] io_perf_1_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg [5:0] io_perf_2_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg [5:0] io_perf_2_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg [5:0] io_perf_3_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg [5:0] io_perf_3_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg [5:0] io_perf_4_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg [5:0] io_perf_4_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg [5:0] io_perf_5_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg [5:0] io_perf_5_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg [5:0] io_perf_6_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg [5:0] io_perf_6_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg [5:0] io_perf_7_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg [5:0] io_perf_7_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg [5:0] io_perf_8_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg [5:0] io_perf_8_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg [5:0] io_perf_9_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg [5:0] io_perf_9_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg [5:0] io_perf_10_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg [5:0] io_perf_10_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg [5:0] io_perf_11_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg [5:0] io_perf_11_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg [5:0] io_perf_12_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg [5:0] io_perf_12_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg [5:0] io_perf_13_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg [5:0] io_perf_13_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg [5:0] io_perf_14_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg [5:0] io_perf_14_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg [5:0] io_perf_15_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg [5:0] io_perf_15_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg [5:0] io_perf_16_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg [5:0] io_perf_16_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg [5:0] io_perf_17_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg [5:0] io_perf_17_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg [5:0] io_perf_18_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg [5:0] io_perf_18_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg [63:0] cnt_1; // @[ChiselDB.scala 133:22]
  reg [63:0] cnt_2; // @[ChiselDB.scala 133:22]
  reg [63:0] cnt_3; // @[ChiselDB.scala 133:22]
  reg [63:0] cnt_4; // @[ChiselDB.scala 133:22]
  reg [63:0] cnt_5; // @[ChiselDB.scala 133:22]
  reg [63:0] cnt_6; // @[ChiselDB.scala 133:22]
  reg [63:0] cnt_7; // @[ChiselDB.scala 133:22]
  reg [63:0] cnt_8; // @[ChiselDB.scala 133:22]
  reg [63:0] cnt_9; // @[ChiselDB.scala 133:22]
  reg [63:0] cnt_10; // @[ChiselDB.scala 133:22]
  reg [63:0] cnt_11; // @[ChiselDB.scala 133:22]
  DelayN_23 sfence_tmp_delay ( // @[Hold.scala 97:23]
    .clock(sfence_tmp_delay_clock),
    .io_in_valid(sfence_tmp_delay_io_in_valid),
    .io_in_bits_rs1(sfence_tmp_delay_io_in_bits_rs1),
    .io_in_bits_rs2(sfence_tmp_delay_io_in_bits_rs2),
    .io_in_bits_addr(sfence_tmp_delay_io_in_bits_addr),
    .io_in_bits_asid(sfence_tmp_delay_io_in_bits_asid),
    .io_out_valid(sfence_tmp_delay_io_out_valid),
    .io_out_bits_rs1(sfence_tmp_delay_io_out_bits_rs1),
    .io_out_bits_rs2(sfence_tmp_delay_io_out_bits_rs2),
    .io_out_bits_addr(sfence_tmp_delay_io_out_bits_addr),
    .io_out_bits_asid(sfence_tmp_delay_io_out_bits_asid)
  );
  DelayN_24 csr_tmp_delay ( // @[Hold.scala 97:23]
    .clock(csr_tmp_delay_clock),
    .io_in_satp_asid(csr_tmp_delay_io_in_satp_asid),
    .io_in_satp_ppn(csr_tmp_delay_io_in_satp_ppn),
    .io_in_satp_changed(csr_tmp_delay_io_in_satp_changed),
    .io_out_satp_asid(csr_tmp_delay_io_out_satp_asid),
    .io_out_satp_ppn(csr_tmp_delay_io_out_satp_ppn),
    .io_out_satp_changed(csr_tmp_delay_io_out_satp_changed)
  );
  PMP pmp ( // @[L2TLB.scala 88:19]
    .clock(pmp_clock),
    .reset(pmp_reset),
    .io_distribute_csr_wvalid(pmp_io_distribute_csr_wvalid),
    .io_distribute_csr_waddr(pmp_io_distribute_csr_waddr),
    .io_distribute_csr_wdata(pmp_io_distribute_csr_wdata),
    .io_pmp_0_cfg_l(pmp_io_pmp_0_cfg_l),
    .io_pmp_0_cfg_a(pmp_io_pmp_0_cfg_a),
    .io_pmp_0_cfg_x(pmp_io_pmp_0_cfg_x),
    .io_pmp_0_cfg_w(pmp_io_pmp_0_cfg_w),
    .io_pmp_0_cfg_r(pmp_io_pmp_0_cfg_r),
    .io_pmp_0_addr(pmp_io_pmp_0_addr),
    .io_pmp_0_mask(pmp_io_pmp_0_mask),
    .io_pmp_1_cfg_l(pmp_io_pmp_1_cfg_l),
    .io_pmp_1_cfg_a(pmp_io_pmp_1_cfg_a),
    .io_pmp_1_cfg_x(pmp_io_pmp_1_cfg_x),
    .io_pmp_1_cfg_w(pmp_io_pmp_1_cfg_w),
    .io_pmp_1_cfg_r(pmp_io_pmp_1_cfg_r),
    .io_pmp_1_addr(pmp_io_pmp_1_addr),
    .io_pmp_1_mask(pmp_io_pmp_1_mask),
    .io_pmp_2_cfg_l(pmp_io_pmp_2_cfg_l),
    .io_pmp_2_cfg_a(pmp_io_pmp_2_cfg_a),
    .io_pmp_2_cfg_x(pmp_io_pmp_2_cfg_x),
    .io_pmp_2_cfg_w(pmp_io_pmp_2_cfg_w),
    .io_pmp_2_cfg_r(pmp_io_pmp_2_cfg_r),
    .io_pmp_2_addr(pmp_io_pmp_2_addr),
    .io_pmp_2_mask(pmp_io_pmp_2_mask),
    .io_pmp_3_cfg_l(pmp_io_pmp_3_cfg_l),
    .io_pmp_3_cfg_a(pmp_io_pmp_3_cfg_a),
    .io_pmp_3_cfg_x(pmp_io_pmp_3_cfg_x),
    .io_pmp_3_cfg_w(pmp_io_pmp_3_cfg_w),
    .io_pmp_3_cfg_r(pmp_io_pmp_3_cfg_r),
    .io_pmp_3_addr(pmp_io_pmp_3_addr),
    .io_pmp_3_mask(pmp_io_pmp_3_mask),
    .io_pmp_4_cfg_l(pmp_io_pmp_4_cfg_l),
    .io_pmp_4_cfg_a(pmp_io_pmp_4_cfg_a),
    .io_pmp_4_cfg_x(pmp_io_pmp_4_cfg_x),
    .io_pmp_4_cfg_w(pmp_io_pmp_4_cfg_w),
    .io_pmp_4_cfg_r(pmp_io_pmp_4_cfg_r),
    .io_pmp_4_addr(pmp_io_pmp_4_addr),
    .io_pmp_4_mask(pmp_io_pmp_4_mask),
    .io_pmp_5_cfg_l(pmp_io_pmp_5_cfg_l),
    .io_pmp_5_cfg_a(pmp_io_pmp_5_cfg_a),
    .io_pmp_5_cfg_x(pmp_io_pmp_5_cfg_x),
    .io_pmp_5_cfg_w(pmp_io_pmp_5_cfg_w),
    .io_pmp_5_cfg_r(pmp_io_pmp_5_cfg_r),
    .io_pmp_5_addr(pmp_io_pmp_5_addr),
    .io_pmp_5_mask(pmp_io_pmp_5_mask),
    .io_pmp_6_cfg_l(pmp_io_pmp_6_cfg_l),
    .io_pmp_6_cfg_a(pmp_io_pmp_6_cfg_a),
    .io_pmp_6_cfg_x(pmp_io_pmp_6_cfg_x),
    .io_pmp_6_cfg_w(pmp_io_pmp_6_cfg_w),
    .io_pmp_6_cfg_r(pmp_io_pmp_6_cfg_r),
    .io_pmp_6_addr(pmp_io_pmp_6_addr),
    .io_pmp_6_mask(pmp_io_pmp_6_mask),
    .io_pmp_7_cfg_l(pmp_io_pmp_7_cfg_l),
    .io_pmp_7_cfg_a(pmp_io_pmp_7_cfg_a),
    .io_pmp_7_cfg_x(pmp_io_pmp_7_cfg_x),
    .io_pmp_7_cfg_w(pmp_io_pmp_7_cfg_w),
    .io_pmp_7_cfg_r(pmp_io_pmp_7_cfg_r),
    .io_pmp_7_addr(pmp_io_pmp_7_addr),
    .io_pmp_7_mask(pmp_io_pmp_7_mask),
    .io_pmp_8_cfg_l(pmp_io_pmp_8_cfg_l),
    .io_pmp_8_cfg_a(pmp_io_pmp_8_cfg_a),
    .io_pmp_8_cfg_x(pmp_io_pmp_8_cfg_x),
    .io_pmp_8_cfg_w(pmp_io_pmp_8_cfg_w),
    .io_pmp_8_cfg_r(pmp_io_pmp_8_cfg_r),
    .io_pmp_8_addr(pmp_io_pmp_8_addr),
    .io_pmp_8_mask(pmp_io_pmp_8_mask),
    .io_pmp_9_cfg_l(pmp_io_pmp_9_cfg_l),
    .io_pmp_9_cfg_a(pmp_io_pmp_9_cfg_a),
    .io_pmp_9_cfg_x(pmp_io_pmp_9_cfg_x),
    .io_pmp_9_cfg_w(pmp_io_pmp_9_cfg_w),
    .io_pmp_9_cfg_r(pmp_io_pmp_9_cfg_r),
    .io_pmp_9_addr(pmp_io_pmp_9_addr),
    .io_pmp_9_mask(pmp_io_pmp_9_mask),
    .io_pmp_10_cfg_l(pmp_io_pmp_10_cfg_l),
    .io_pmp_10_cfg_a(pmp_io_pmp_10_cfg_a),
    .io_pmp_10_cfg_x(pmp_io_pmp_10_cfg_x),
    .io_pmp_10_cfg_w(pmp_io_pmp_10_cfg_w),
    .io_pmp_10_cfg_r(pmp_io_pmp_10_cfg_r),
    .io_pmp_10_addr(pmp_io_pmp_10_addr),
    .io_pmp_10_mask(pmp_io_pmp_10_mask),
    .io_pmp_11_cfg_l(pmp_io_pmp_11_cfg_l),
    .io_pmp_11_cfg_a(pmp_io_pmp_11_cfg_a),
    .io_pmp_11_cfg_x(pmp_io_pmp_11_cfg_x),
    .io_pmp_11_cfg_w(pmp_io_pmp_11_cfg_w),
    .io_pmp_11_cfg_r(pmp_io_pmp_11_cfg_r),
    .io_pmp_11_addr(pmp_io_pmp_11_addr),
    .io_pmp_11_mask(pmp_io_pmp_11_mask),
    .io_pmp_12_cfg_l(pmp_io_pmp_12_cfg_l),
    .io_pmp_12_cfg_a(pmp_io_pmp_12_cfg_a),
    .io_pmp_12_cfg_x(pmp_io_pmp_12_cfg_x),
    .io_pmp_12_cfg_w(pmp_io_pmp_12_cfg_w),
    .io_pmp_12_cfg_r(pmp_io_pmp_12_cfg_r),
    .io_pmp_12_addr(pmp_io_pmp_12_addr),
    .io_pmp_12_mask(pmp_io_pmp_12_mask),
    .io_pmp_13_cfg_l(pmp_io_pmp_13_cfg_l),
    .io_pmp_13_cfg_a(pmp_io_pmp_13_cfg_a),
    .io_pmp_13_cfg_x(pmp_io_pmp_13_cfg_x),
    .io_pmp_13_cfg_w(pmp_io_pmp_13_cfg_w),
    .io_pmp_13_cfg_r(pmp_io_pmp_13_cfg_r),
    .io_pmp_13_addr(pmp_io_pmp_13_addr),
    .io_pmp_13_mask(pmp_io_pmp_13_mask),
    .io_pmp_14_cfg_l(pmp_io_pmp_14_cfg_l),
    .io_pmp_14_cfg_a(pmp_io_pmp_14_cfg_a),
    .io_pmp_14_cfg_x(pmp_io_pmp_14_cfg_x),
    .io_pmp_14_cfg_w(pmp_io_pmp_14_cfg_w),
    .io_pmp_14_cfg_r(pmp_io_pmp_14_cfg_r),
    .io_pmp_14_addr(pmp_io_pmp_14_addr),
    .io_pmp_14_mask(pmp_io_pmp_14_mask),
    .io_pmp_15_cfg_l(pmp_io_pmp_15_cfg_l),
    .io_pmp_15_cfg_a(pmp_io_pmp_15_cfg_a),
    .io_pmp_15_cfg_x(pmp_io_pmp_15_cfg_x),
    .io_pmp_15_cfg_w(pmp_io_pmp_15_cfg_w),
    .io_pmp_15_cfg_r(pmp_io_pmp_15_cfg_r),
    .io_pmp_15_addr(pmp_io_pmp_15_addr),
    .io_pmp_15_mask(pmp_io_pmp_15_mask),
    .io_pma_0_cfg_c(pmp_io_pma_0_cfg_c),
    .io_pma_0_cfg_atomic(pmp_io_pma_0_cfg_atomic),
    .io_pma_0_cfg_a(pmp_io_pma_0_cfg_a),
    .io_pma_0_cfg_x(pmp_io_pma_0_cfg_x),
    .io_pma_0_cfg_w(pmp_io_pma_0_cfg_w),
    .io_pma_0_cfg_r(pmp_io_pma_0_cfg_r),
    .io_pma_0_addr(pmp_io_pma_0_addr),
    .io_pma_0_mask(pmp_io_pma_0_mask),
    .io_pma_1_cfg_c(pmp_io_pma_1_cfg_c),
    .io_pma_1_cfg_atomic(pmp_io_pma_1_cfg_atomic),
    .io_pma_1_cfg_a(pmp_io_pma_1_cfg_a),
    .io_pma_1_cfg_x(pmp_io_pma_1_cfg_x),
    .io_pma_1_cfg_w(pmp_io_pma_1_cfg_w),
    .io_pma_1_cfg_r(pmp_io_pma_1_cfg_r),
    .io_pma_1_addr(pmp_io_pma_1_addr),
    .io_pma_1_mask(pmp_io_pma_1_mask),
    .io_pma_2_cfg_c(pmp_io_pma_2_cfg_c),
    .io_pma_2_cfg_atomic(pmp_io_pma_2_cfg_atomic),
    .io_pma_2_cfg_a(pmp_io_pma_2_cfg_a),
    .io_pma_2_cfg_x(pmp_io_pma_2_cfg_x),
    .io_pma_2_cfg_w(pmp_io_pma_2_cfg_w),
    .io_pma_2_cfg_r(pmp_io_pma_2_cfg_r),
    .io_pma_2_addr(pmp_io_pma_2_addr),
    .io_pma_2_mask(pmp_io_pma_2_mask),
    .io_pma_3_cfg_c(pmp_io_pma_3_cfg_c),
    .io_pma_3_cfg_atomic(pmp_io_pma_3_cfg_atomic),
    .io_pma_3_cfg_a(pmp_io_pma_3_cfg_a),
    .io_pma_3_cfg_x(pmp_io_pma_3_cfg_x),
    .io_pma_3_cfg_w(pmp_io_pma_3_cfg_w),
    .io_pma_3_cfg_r(pmp_io_pma_3_cfg_r),
    .io_pma_3_addr(pmp_io_pma_3_addr),
    .io_pma_3_mask(pmp_io_pma_3_mask),
    .io_pma_4_cfg_c(pmp_io_pma_4_cfg_c),
    .io_pma_4_cfg_atomic(pmp_io_pma_4_cfg_atomic),
    .io_pma_4_cfg_a(pmp_io_pma_4_cfg_a),
    .io_pma_4_cfg_x(pmp_io_pma_4_cfg_x),
    .io_pma_4_cfg_w(pmp_io_pma_4_cfg_w),
    .io_pma_4_cfg_r(pmp_io_pma_4_cfg_r),
    .io_pma_4_addr(pmp_io_pma_4_addr),
    .io_pma_4_mask(pmp_io_pma_4_mask),
    .io_pma_5_cfg_c(pmp_io_pma_5_cfg_c),
    .io_pma_5_cfg_atomic(pmp_io_pma_5_cfg_atomic),
    .io_pma_5_cfg_a(pmp_io_pma_5_cfg_a),
    .io_pma_5_cfg_x(pmp_io_pma_5_cfg_x),
    .io_pma_5_cfg_w(pmp_io_pma_5_cfg_w),
    .io_pma_5_cfg_r(pmp_io_pma_5_cfg_r),
    .io_pma_5_addr(pmp_io_pma_5_addr),
    .io_pma_5_mask(pmp_io_pma_5_mask),
    .io_pma_6_cfg_c(pmp_io_pma_6_cfg_c),
    .io_pma_6_cfg_atomic(pmp_io_pma_6_cfg_atomic),
    .io_pma_6_cfg_a(pmp_io_pma_6_cfg_a),
    .io_pma_6_cfg_x(pmp_io_pma_6_cfg_x),
    .io_pma_6_cfg_w(pmp_io_pma_6_cfg_w),
    .io_pma_6_cfg_r(pmp_io_pma_6_cfg_r),
    .io_pma_6_addr(pmp_io_pma_6_addr),
    .io_pma_6_mask(pmp_io_pma_6_mask),
    .io_pma_7_cfg_c(pmp_io_pma_7_cfg_c),
    .io_pma_7_cfg_atomic(pmp_io_pma_7_cfg_atomic),
    .io_pma_7_cfg_a(pmp_io_pma_7_cfg_a),
    .io_pma_7_cfg_x(pmp_io_pma_7_cfg_x),
    .io_pma_7_cfg_w(pmp_io_pma_7_cfg_w),
    .io_pma_7_cfg_r(pmp_io_pma_7_cfg_r),
    .io_pma_7_addr(pmp_io_pma_7_addr),
    .io_pma_7_mask(pmp_io_pma_7_mask),
    .io_pma_8_cfg_c(pmp_io_pma_8_cfg_c),
    .io_pma_8_cfg_atomic(pmp_io_pma_8_cfg_atomic),
    .io_pma_8_cfg_a(pmp_io_pma_8_cfg_a),
    .io_pma_8_cfg_x(pmp_io_pma_8_cfg_x),
    .io_pma_8_cfg_w(pmp_io_pma_8_cfg_w),
    .io_pma_8_cfg_r(pmp_io_pma_8_cfg_r),
    .io_pma_8_addr(pmp_io_pma_8_addr),
    .io_pma_8_mask(pmp_io_pma_8_mask),
    .io_pma_9_cfg_c(pmp_io_pma_9_cfg_c),
    .io_pma_9_cfg_atomic(pmp_io_pma_9_cfg_atomic),
    .io_pma_9_cfg_a(pmp_io_pma_9_cfg_a),
    .io_pma_9_cfg_x(pmp_io_pma_9_cfg_x),
    .io_pma_9_cfg_w(pmp_io_pma_9_cfg_w),
    .io_pma_9_cfg_r(pmp_io_pma_9_cfg_r),
    .io_pma_9_addr(pmp_io_pma_9_addr),
    .io_pma_9_mask(pmp_io_pma_9_mask),
    .io_pma_10_cfg_c(pmp_io_pma_10_cfg_c),
    .io_pma_10_cfg_atomic(pmp_io_pma_10_cfg_atomic),
    .io_pma_10_cfg_a(pmp_io_pma_10_cfg_a),
    .io_pma_10_cfg_x(pmp_io_pma_10_cfg_x),
    .io_pma_10_cfg_w(pmp_io_pma_10_cfg_w),
    .io_pma_10_cfg_r(pmp_io_pma_10_cfg_r),
    .io_pma_10_addr(pmp_io_pma_10_addr),
    .io_pma_10_mask(pmp_io_pma_10_mask),
    .io_pma_11_cfg_c(pmp_io_pma_11_cfg_c),
    .io_pma_11_cfg_atomic(pmp_io_pma_11_cfg_atomic),
    .io_pma_11_cfg_a(pmp_io_pma_11_cfg_a),
    .io_pma_11_cfg_x(pmp_io_pma_11_cfg_x),
    .io_pma_11_cfg_w(pmp_io_pma_11_cfg_w),
    .io_pma_11_cfg_r(pmp_io_pma_11_cfg_r),
    .io_pma_11_addr(pmp_io_pma_11_addr),
    .io_pma_11_mask(pmp_io_pma_11_mask),
    .io_pma_12_cfg_c(pmp_io_pma_12_cfg_c),
    .io_pma_12_cfg_atomic(pmp_io_pma_12_cfg_atomic),
    .io_pma_12_cfg_a(pmp_io_pma_12_cfg_a),
    .io_pma_12_cfg_x(pmp_io_pma_12_cfg_x),
    .io_pma_12_cfg_w(pmp_io_pma_12_cfg_w),
    .io_pma_12_cfg_r(pmp_io_pma_12_cfg_r),
    .io_pma_12_addr(pmp_io_pma_12_addr),
    .io_pma_12_mask(pmp_io_pma_12_mask),
    .io_pma_13_cfg_c(pmp_io_pma_13_cfg_c),
    .io_pma_13_cfg_atomic(pmp_io_pma_13_cfg_atomic),
    .io_pma_13_cfg_a(pmp_io_pma_13_cfg_a),
    .io_pma_13_cfg_x(pmp_io_pma_13_cfg_x),
    .io_pma_13_cfg_w(pmp_io_pma_13_cfg_w),
    .io_pma_13_cfg_r(pmp_io_pma_13_cfg_r),
    .io_pma_13_addr(pmp_io_pma_13_addr),
    .io_pma_13_mask(pmp_io_pma_13_mask),
    .io_pma_14_cfg_c(pmp_io_pma_14_cfg_c),
    .io_pma_14_cfg_atomic(pmp_io_pma_14_cfg_atomic),
    .io_pma_14_cfg_a(pmp_io_pma_14_cfg_a),
    .io_pma_14_cfg_x(pmp_io_pma_14_cfg_x),
    .io_pma_14_cfg_w(pmp_io_pma_14_cfg_w),
    .io_pma_14_cfg_r(pmp_io_pma_14_cfg_r),
    .io_pma_14_addr(pmp_io_pma_14_addr),
    .io_pma_14_mask(pmp_io_pma_14_mask),
    .io_pma_15_cfg_c(pmp_io_pma_15_cfg_c),
    .io_pma_15_cfg_atomic(pmp_io_pma_15_cfg_atomic),
    .io_pma_15_cfg_a(pmp_io_pma_15_cfg_a),
    .io_pma_15_cfg_x(pmp_io_pma_15_cfg_x),
    .io_pma_15_cfg_w(pmp_io_pma_15_cfg_w),
    .io_pma_15_cfg_r(pmp_io_pma_15_cfg_r),
    .io_pma_15_addr(pmp_io_pma_15_addr),
    .io_pma_15_mask(pmp_io_pma_15_mask)
  );
  PMPChecker PMPChecker ( // @[L2TLB.scala 89:45]
    .io_check_env_mode(PMPChecker_io_check_env_mode),
    .io_check_env_pmp_0_cfg_l(PMPChecker_io_check_env_pmp_0_cfg_l),
    .io_check_env_pmp_0_cfg_a(PMPChecker_io_check_env_pmp_0_cfg_a),
    .io_check_env_pmp_0_cfg_x(PMPChecker_io_check_env_pmp_0_cfg_x),
    .io_check_env_pmp_0_cfg_w(PMPChecker_io_check_env_pmp_0_cfg_w),
    .io_check_env_pmp_0_cfg_r(PMPChecker_io_check_env_pmp_0_cfg_r),
    .io_check_env_pmp_0_addr(PMPChecker_io_check_env_pmp_0_addr),
    .io_check_env_pmp_0_mask(PMPChecker_io_check_env_pmp_0_mask),
    .io_check_env_pmp_1_cfg_l(PMPChecker_io_check_env_pmp_1_cfg_l),
    .io_check_env_pmp_1_cfg_a(PMPChecker_io_check_env_pmp_1_cfg_a),
    .io_check_env_pmp_1_cfg_x(PMPChecker_io_check_env_pmp_1_cfg_x),
    .io_check_env_pmp_1_cfg_w(PMPChecker_io_check_env_pmp_1_cfg_w),
    .io_check_env_pmp_1_cfg_r(PMPChecker_io_check_env_pmp_1_cfg_r),
    .io_check_env_pmp_1_addr(PMPChecker_io_check_env_pmp_1_addr),
    .io_check_env_pmp_1_mask(PMPChecker_io_check_env_pmp_1_mask),
    .io_check_env_pmp_2_cfg_l(PMPChecker_io_check_env_pmp_2_cfg_l),
    .io_check_env_pmp_2_cfg_a(PMPChecker_io_check_env_pmp_2_cfg_a),
    .io_check_env_pmp_2_cfg_x(PMPChecker_io_check_env_pmp_2_cfg_x),
    .io_check_env_pmp_2_cfg_w(PMPChecker_io_check_env_pmp_2_cfg_w),
    .io_check_env_pmp_2_cfg_r(PMPChecker_io_check_env_pmp_2_cfg_r),
    .io_check_env_pmp_2_addr(PMPChecker_io_check_env_pmp_2_addr),
    .io_check_env_pmp_2_mask(PMPChecker_io_check_env_pmp_2_mask),
    .io_check_env_pmp_3_cfg_l(PMPChecker_io_check_env_pmp_3_cfg_l),
    .io_check_env_pmp_3_cfg_a(PMPChecker_io_check_env_pmp_3_cfg_a),
    .io_check_env_pmp_3_cfg_x(PMPChecker_io_check_env_pmp_3_cfg_x),
    .io_check_env_pmp_3_cfg_w(PMPChecker_io_check_env_pmp_3_cfg_w),
    .io_check_env_pmp_3_cfg_r(PMPChecker_io_check_env_pmp_3_cfg_r),
    .io_check_env_pmp_3_addr(PMPChecker_io_check_env_pmp_3_addr),
    .io_check_env_pmp_3_mask(PMPChecker_io_check_env_pmp_3_mask),
    .io_check_env_pmp_4_cfg_l(PMPChecker_io_check_env_pmp_4_cfg_l),
    .io_check_env_pmp_4_cfg_a(PMPChecker_io_check_env_pmp_4_cfg_a),
    .io_check_env_pmp_4_cfg_x(PMPChecker_io_check_env_pmp_4_cfg_x),
    .io_check_env_pmp_4_cfg_w(PMPChecker_io_check_env_pmp_4_cfg_w),
    .io_check_env_pmp_4_cfg_r(PMPChecker_io_check_env_pmp_4_cfg_r),
    .io_check_env_pmp_4_addr(PMPChecker_io_check_env_pmp_4_addr),
    .io_check_env_pmp_4_mask(PMPChecker_io_check_env_pmp_4_mask),
    .io_check_env_pmp_5_cfg_l(PMPChecker_io_check_env_pmp_5_cfg_l),
    .io_check_env_pmp_5_cfg_a(PMPChecker_io_check_env_pmp_5_cfg_a),
    .io_check_env_pmp_5_cfg_x(PMPChecker_io_check_env_pmp_5_cfg_x),
    .io_check_env_pmp_5_cfg_w(PMPChecker_io_check_env_pmp_5_cfg_w),
    .io_check_env_pmp_5_cfg_r(PMPChecker_io_check_env_pmp_5_cfg_r),
    .io_check_env_pmp_5_addr(PMPChecker_io_check_env_pmp_5_addr),
    .io_check_env_pmp_5_mask(PMPChecker_io_check_env_pmp_5_mask),
    .io_check_env_pmp_6_cfg_l(PMPChecker_io_check_env_pmp_6_cfg_l),
    .io_check_env_pmp_6_cfg_a(PMPChecker_io_check_env_pmp_6_cfg_a),
    .io_check_env_pmp_6_cfg_x(PMPChecker_io_check_env_pmp_6_cfg_x),
    .io_check_env_pmp_6_cfg_w(PMPChecker_io_check_env_pmp_6_cfg_w),
    .io_check_env_pmp_6_cfg_r(PMPChecker_io_check_env_pmp_6_cfg_r),
    .io_check_env_pmp_6_addr(PMPChecker_io_check_env_pmp_6_addr),
    .io_check_env_pmp_6_mask(PMPChecker_io_check_env_pmp_6_mask),
    .io_check_env_pmp_7_cfg_l(PMPChecker_io_check_env_pmp_7_cfg_l),
    .io_check_env_pmp_7_cfg_a(PMPChecker_io_check_env_pmp_7_cfg_a),
    .io_check_env_pmp_7_cfg_x(PMPChecker_io_check_env_pmp_7_cfg_x),
    .io_check_env_pmp_7_cfg_w(PMPChecker_io_check_env_pmp_7_cfg_w),
    .io_check_env_pmp_7_cfg_r(PMPChecker_io_check_env_pmp_7_cfg_r),
    .io_check_env_pmp_7_addr(PMPChecker_io_check_env_pmp_7_addr),
    .io_check_env_pmp_7_mask(PMPChecker_io_check_env_pmp_7_mask),
    .io_check_env_pmp_8_cfg_l(PMPChecker_io_check_env_pmp_8_cfg_l),
    .io_check_env_pmp_8_cfg_a(PMPChecker_io_check_env_pmp_8_cfg_a),
    .io_check_env_pmp_8_cfg_x(PMPChecker_io_check_env_pmp_8_cfg_x),
    .io_check_env_pmp_8_cfg_w(PMPChecker_io_check_env_pmp_8_cfg_w),
    .io_check_env_pmp_8_cfg_r(PMPChecker_io_check_env_pmp_8_cfg_r),
    .io_check_env_pmp_8_addr(PMPChecker_io_check_env_pmp_8_addr),
    .io_check_env_pmp_8_mask(PMPChecker_io_check_env_pmp_8_mask),
    .io_check_env_pmp_9_cfg_l(PMPChecker_io_check_env_pmp_9_cfg_l),
    .io_check_env_pmp_9_cfg_a(PMPChecker_io_check_env_pmp_9_cfg_a),
    .io_check_env_pmp_9_cfg_x(PMPChecker_io_check_env_pmp_9_cfg_x),
    .io_check_env_pmp_9_cfg_w(PMPChecker_io_check_env_pmp_9_cfg_w),
    .io_check_env_pmp_9_cfg_r(PMPChecker_io_check_env_pmp_9_cfg_r),
    .io_check_env_pmp_9_addr(PMPChecker_io_check_env_pmp_9_addr),
    .io_check_env_pmp_9_mask(PMPChecker_io_check_env_pmp_9_mask),
    .io_check_env_pmp_10_cfg_l(PMPChecker_io_check_env_pmp_10_cfg_l),
    .io_check_env_pmp_10_cfg_a(PMPChecker_io_check_env_pmp_10_cfg_a),
    .io_check_env_pmp_10_cfg_x(PMPChecker_io_check_env_pmp_10_cfg_x),
    .io_check_env_pmp_10_cfg_w(PMPChecker_io_check_env_pmp_10_cfg_w),
    .io_check_env_pmp_10_cfg_r(PMPChecker_io_check_env_pmp_10_cfg_r),
    .io_check_env_pmp_10_addr(PMPChecker_io_check_env_pmp_10_addr),
    .io_check_env_pmp_10_mask(PMPChecker_io_check_env_pmp_10_mask),
    .io_check_env_pmp_11_cfg_l(PMPChecker_io_check_env_pmp_11_cfg_l),
    .io_check_env_pmp_11_cfg_a(PMPChecker_io_check_env_pmp_11_cfg_a),
    .io_check_env_pmp_11_cfg_x(PMPChecker_io_check_env_pmp_11_cfg_x),
    .io_check_env_pmp_11_cfg_w(PMPChecker_io_check_env_pmp_11_cfg_w),
    .io_check_env_pmp_11_cfg_r(PMPChecker_io_check_env_pmp_11_cfg_r),
    .io_check_env_pmp_11_addr(PMPChecker_io_check_env_pmp_11_addr),
    .io_check_env_pmp_11_mask(PMPChecker_io_check_env_pmp_11_mask),
    .io_check_env_pmp_12_cfg_l(PMPChecker_io_check_env_pmp_12_cfg_l),
    .io_check_env_pmp_12_cfg_a(PMPChecker_io_check_env_pmp_12_cfg_a),
    .io_check_env_pmp_12_cfg_x(PMPChecker_io_check_env_pmp_12_cfg_x),
    .io_check_env_pmp_12_cfg_w(PMPChecker_io_check_env_pmp_12_cfg_w),
    .io_check_env_pmp_12_cfg_r(PMPChecker_io_check_env_pmp_12_cfg_r),
    .io_check_env_pmp_12_addr(PMPChecker_io_check_env_pmp_12_addr),
    .io_check_env_pmp_12_mask(PMPChecker_io_check_env_pmp_12_mask),
    .io_check_env_pmp_13_cfg_l(PMPChecker_io_check_env_pmp_13_cfg_l),
    .io_check_env_pmp_13_cfg_a(PMPChecker_io_check_env_pmp_13_cfg_a),
    .io_check_env_pmp_13_cfg_x(PMPChecker_io_check_env_pmp_13_cfg_x),
    .io_check_env_pmp_13_cfg_w(PMPChecker_io_check_env_pmp_13_cfg_w),
    .io_check_env_pmp_13_cfg_r(PMPChecker_io_check_env_pmp_13_cfg_r),
    .io_check_env_pmp_13_addr(PMPChecker_io_check_env_pmp_13_addr),
    .io_check_env_pmp_13_mask(PMPChecker_io_check_env_pmp_13_mask),
    .io_check_env_pmp_14_cfg_l(PMPChecker_io_check_env_pmp_14_cfg_l),
    .io_check_env_pmp_14_cfg_a(PMPChecker_io_check_env_pmp_14_cfg_a),
    .io_check_env_pmp_14_cfg_x(PMPChecker_io_check_env_pmp_14_cfg_x),
    .io_check_env_pmp_14_cfg_w(PMPChecker_io_check_env_pmp_14_cfg_w),
    .io_check_env_pmp_14_cfg_r(PMPChecker_io_check_env_pmp_14_cfg_r),
    .io_check_env_pmp_14_addr(PMPChecker_io_check_env_pmp_14_addr),
    .io_check_env_pmp_14_mask(PMPChecker_io_check_env_pmp_14_mask),
    .io_check_env_pmp_15_cfg_l(PMPChecker_io_check_env_pmp_15_cfg_l),
    .io_check_env_pmp_15_cfg_a(PMPChecker_io_check_env_pmp_15_cfg_a),
    .io_check_env_pmp_15_cfg_x(PMPChecker_io_check_env_pmp_15_cfg_x),
    .io_check_env_pmp_15_cfg_w(PMPChecker_io_check_env_pmp_15_cfg_w),
    .io_check_env_pmp_15_cfg_r(PMPChecker_io_check_env_pmp_15_cfg_r),
    .io_check_env_pmp_15_addr(PMPChecker_io_check_env_pmp_15_addr),
    .io_check_env_pmp_15_mask(PMPChecker_io_check_env_pmp_15_mask),
    .io_check_env_pma_0_cfg_c(PMPChecker_io_check_env_pma_0_cfg_c),
    .io_check_env_pma_0_cfg_atomic(PMPChecker_io_check_env_pma_0_cfg_atomic),
    .io_check_env_pma_0_cfg_a(PMPChecker_io_check_env_pma_0_cfg_a),
    .io_check_env_pma_0_cfg_x(PMPChecker_io_check_env_pma_0_cfg_x),
    .io_check_env_pma_0_cfg_w(PMPChecker_io_check_env_pma_0_cfg_w),
    .io_check_env_pma_0_cfg_r(PMPChecker_io_check_env_pma_0_cfg_r),
    .io_check_env_pma_0_addr(PMPChecker_io_check_env_pma_0_addr),
    .io_check_env_pma_0_mask(PMPChecker_io_check_env_pma_0_mask),
    .io_check_env_pma_1_cfg_c(PMPChecker_io_check_env_pma_1_cfg_c),
    .io_check_env_pma_1_cfg_atomic(PMPChecker_io_check_env_pma_1_cfg_atomic),
    .io_check_env_pma_1_cfg_a(PMPChecker_io_check_env_pma_1_cfg_a),
    .io_check_env_pma_1_cfg_x(PMPChecker_io_check_env_pma_1_cfg_x),
    .io_check_env_pma_1_cfg_w(PMPChecker_io_check_env_pma_1_cfg_w),
    .io_check_env_pma_1_cfg_r(PMPChecker_io_check_env_pma_1_cfg_r),
    .io_check_env_pma_1_addr(PMPChecker_io_check_env_pma_1_addr),
    .io_check_env_pma_1_mask(PMPChecker_io_check_env_pma_1_mask),
    .io_check_env_pma_2_cfg_c(PMPChecker_io_check_env_pma_2_cfg_c),
    .io_check_env_pma_2_cfg_atomic(PMPChecker_io_check_env_pma_2_cfg_atomic),
    .io_check_env_pma_2_cfg_a(PMPChecker_io_check_env_pma_2_cfg_a),
    .io_check_env_pma_2_cfg_x(PMPChecker_io_check_env_pma_2_cfg_x),
    .io_check_env_pma_2_cfg_w(PMPChecker_io_check_env_pma_2_cfg_w),
    .io_check_env_pma_2_cfg_r(PMPChecker_io_check_env_pma_2_cfg_r),
    .io_check_env_pma_2_addr(PMPChecker_io_check_env_pma_2_addr),
    .io_check_env_pma_2_mask(PMPChecker_io_check_env_pma_2_mask),
    .io_check_env_pma_3_cfg_c(PMPChecker_io_check_env_pma_3_cfg_c),
    .io_check_env_pma_3_cfg_atomic(PMPChecker_io_check_env_pma_3_cfg_atomic),
    .io_check_env_pma_3_cfg_a(PMPChecker_io_check_env_pma_3_cfg_a),
    .io_check_env_pma_3_cfg_x(PMPChecker_io_check_env_pma_3_cfg_x),
    .io_check_env_pma_3_cfg_w(PMPChecker_io_check_env_pma_3_cfg_w),
    .io_check_env_pma_3_cfg_r(PMPChecker_io_check_env_pma_3_cfg_r),
    .io_check_env_pma_3_addr(PMPChecker_io_check_env_pma_3_addr),
    .io_check_env_pma_3_mask(PMPChecker_io_check_env_pma_3_mask),
    .io_check_env_pma_4_cfg_c(PMPChecker_io_check_env_pma_4_cfg_c),
    .io_check_env_pma_4_cfg_atomic(PMPChecker_io_check_env_pma_4_cfg_atomic),
    .io_check_env_pma_4_cfg_a(PMPChecker_io_check_env_pma_4_cfg_a),
    .io_check_env_pma_4_cfg_x(PMPChecker_io_check_env_pma_4_cfg_x),
    .io_check_env_pma_4_cfg_w(PMPChecker_io_check_env_pma_4_cfg_w),
    .io_check_env_pma_4_cfg_r(PMPChecker_io_check_env_pma_4_cfg_r),
    .io_check_env_pma_4_addr(PMPChecker_io_check_env_pma_4_addr),
    .io_check_env_pma_4_mask(PMPChecker_io_check_env_pma_4_mask),
    .io_check_env_pma_5_cfg_c(PMPChecker_io_check_env_pma_5_cfg_c),
    .io_check_env_pma_5_cfg_atomic(PMPChecker_io_check_env_pma_5_cfg_atomic),
    .io_check_env_pma_5_cfg_a(PMPChecker_io_check_env_pma_5_cfg_a),
    .io_check_env_pma_5_cfg_x(PMPChecker_io_check_env_pma_5_cfg_x),
    .io_check_env_pma_5_cfg_w(PMPChecker_io_check_env_pma_5_cfg_w),
    .io_check_env_pma_5_cfg_r(PMPChecker_io_check_env_pma_5_cfg_r),
    .io_check_env_pma_5_addr(PMPChecker_io_check_env_pma_5_addr),
    .io_check_env_pma_5_mask(PMPChecker_io_check_env_pma_5_mask),
    .io_check_env_pma_6_cfg_c(PMPChecker_io_check_env_pma_6_cfg_c),
    .io_check_env_pma_6_cfg_atomic(PMPChecker_io_check_env_pma_6_cfg_atomic),
    .io_check_env_pma_6_cfg_a(PMPChecker_io_check_env_pma_6_cfg_a),
    .io_check_env_pma_6_cfg_x(PMPChecker_io_check_env_pma_6_cfg_x),
    .io_check_env_pma_6_cfg_w(PMPChecker_io_check_env_pma_6_cfg_w),
    .io_check_env_pma_6_cfg_r(PMPChecker_io_check_env_pma_6_cfg_r),
    .io_check_env_pma_6_addr(PMPChecker_io_check_env_pma_6_addr),
    .io_check_env_pma_6_mask(PMPChecker_io_check_env_pma_6_mask),
    .io_check_env_pma_7_cfg_c(PMPChecker_io_check_env_pma_7_cfg_c),
    .io_check_env_pma_7_cfg_atomic(PMPChecker_io_check_env_pma_7_cfg_atomic),
    .io_check_env_pma_7_cfg_a(PMPChecker_io_check_env_pma_7_cfg_a),
    .io_check_env_pma_7_cfg_x(PMPChecker_io_check_env_pma_7_cfg_x),
    .io_check_env_pma_7_cfg_w(PMPChecker_io_check_env_pma_7_cfg_w),
    .io_check_env_pma_7_cfg_r(PMPChecker_io_check_env_pma_7_cfg_r),
    .io_check_env_pma_7_addr(PMPChecker_io_check_env_pma_7_addr),
    .io_check_env_pma_7_mask(PMPChecker_io_check_env_pma_7_mask),
    .io_check_env_pma_8_cfg_c(PMPChecker_io_check_env_pma_8_cfg_c),
    .io_check_env_pma_8_cfg_atomic(PMPChecker_io_check_env_pma_8_cfg_atomic),
    .io_check_env_pma_8_cfg_a(PMPChecker_io_check_env_pma_8_cfg_a),
    .io_check_env_pma_8_cfg_x(PMPChecker_io_check_env_pma_8_cfg_x),
    .io_check_env_pma_8_cfg_w(PMPChecker_io_check_env_pma_8_cfg_w),
    .io_check_env_pma_8_cfg_r(PMPChecker_io_check_env_pma_8_cfg_r),
    .io_check_env_pma_8_addr(PMPChecker_io_check_env_pma_8_addr),
    .io_check_env_pma_8_mask(PMPChecker_io_check_env_pma_8_mask),
    .io_check_env_pma_9_cfg_c(PMPChecker_io_check_env_pma_9_cfg_c),
    .io_check_env_pma_9_cfg_atomic(PMPChecker_io_check_env_pma_9_cfg_atomic),
    .io_check_env_pma_9_cfg_a(PMPChecker_io_check_env_pma_9_cfg_a),
    .io_check_env_pma_9_cfg_x(PMPChecker_io_check_env_pma_9_cfg_x),
    .io_check_env_pma_9_cfg_w(PMPChecker_io_check_env_pma_9_cfg_w),
    .io_check_env_pma_9_cfg_r(PMPChecker_io_check_env_pma_9_cfg_r),
    .io_check_env_pma_9_addr(PMPChecker_io_check_env_pma_9_addr),
    .io_check_env_pma_9_mask(PMPChecker_io_check_env_pma_9_mask),
    .io_check_env_pma_10_cfg_c(PMPChecker_io_check_env_pma_10_cfg_c),
    .io_check_env_pma_10_cfg_atomic(PMPChecker_io_check_env_pma_10_cfg_atomic),
    .io_check_env_pma_10_cfg_a(PMPChecker_io_check_env_pma_10_cfg_a),
    .io_check_env_pma_10_cfg_x(PMPChecker_io_check_env_pma_10_cfg_x),
    .io_check_env_pma_10_cfg_w(PMPChecker_io_check_env_pma_10_cfg_w),
    .io_check_env_pma_10_cfg_r(PMPChecker_io_check_env_pma_10_cfg_r),
    .io_check_env_pma_10_addr(PMPChecker_io_check_env_pma_10_addr),
    .io_check_env_pma_10_mask(PMPChecker_io_check_env_pma_10_mask),
    .io_check_env_pma_11_cfg_c(PMPChecker_io_check_env_pma_11_cfg_c),
    .io_check_env_pma_11_cfg_atomic(PMPChecker_io_check_env_pma_11_cfg_atomic),
    .io_check_env_pma_11_cfg_a(PMPChecker_io_check_env_pma_11_cfg_a),
    .io_check_env_pma_11_cfg_x(PMPChecker_io_check_env_pma_11_cfg_x),
    .io_check_env_pma_11_cfg_w(PMPChecker_io_check_env_pma_11_cfg_w),
    .io_check_env_pma_11_cfg_r(PMPChecker_io_check_env_pma_11_cfg_r),
    .io_check_env_pma_11_addr(PMPChecker_io_check_env_pma_11_addr),
    .io_check_env_pma_11_mask(PMPChecker_io_check_env_pma_11_mask),
    .io_check_env_pma_12_cfg_c(PMPChecker_io_check_env_pma_12_cfg_c),
    .io_check_env_pma_12_cfg_atomic(PMPChecker_io_check_env_pma_12_cfg_atomic),
    .io_check_env_pma_12_cfg_a(PMPChecker_io_check_env_pma_12_cfg_a),
    .io_check_env_pma_12_cfg_x(PMPChecker_io_check_env_pma_12_cfg_x),
    .io_check_env_pma_12_cfg_w(PMPChecker_io_check_env_pma_12_cfg_w),
    .io_check_env_pma_12_cfg_r(PMPChecker_io_check_env_pma_12_cfg_r),
    .io_check_env_pma_12_addr(PMPChecker_io_check_env_pma_12_addr),
    .io_check_env_pma_12_mask(PMPChecker_io_check_env_pma_12_mask),
    .io_check_env_pma_13_cfg_c(PMPChecker_io_check_env_pma_13_cfg_c),
    .io_check_env_pma_13_cfg_atomic(PMPChecker_io_check_env_pma_13_cfg_atomic),
    .io_check_env_pma_13_cfg_a(PMPChecker_io_check_env_pma_13_cfg_a),
    .io_check_env_pma_13_cfg_x(PMPChecker_io_check_env_pma_13_cfg_x),
    .io_check_env_pma_13_cfg_w(PMPChecker_io_check_env_pma_13_cfg_w),
    .io_check_env_pma_13_cfg_r(PMPChecker_io_check_env_pma_13_cfg_r),
    .io_check_env_pma_13_addr(PMPChecker_io_check_env_pma_13_addr),
    .io_check_env_pma_13_mask(PMPChecker_io_check_env_pma_13_mask),
    .io_check_env_pma_14_cfg_c(PMPChecker_io_check_env_pma_14_cfg_c),
    .io_check_env_pma_14_cfg_atomic(PMPChecker_io_check_env_pma_14_cfg_atomic),
    .io_check_env_pma_14_cfg_a(PMPChecker_io_check_env_pma_14_cfg_a),
    .io_check_env_pma_14_cfg_x(PMPChecker_io_check_env_pma_14_cfg_x),
    .io_check_env_pma_14_cfg_w(PMPChecker_io_check_env_pma_14_cfg_w),
    .io_check_env_pma_14_cfg_r(PMPChecker_io_check_env_pma_14_cfg_r),
    .io_check_env_pma_14_addr(PMPChecker_io_check_env_pma_14_addr),
    .io_check_env_pma_14_mask(PMPChecker_io_check_env_pma_14_mask),
    .io_check_env_pma_15_cfg_c(PMPChecker_io_check_env_pma_15_cfg_c),
    .io_check_env_pma_15_cfg_atomic(PMPChecker_io_check_env_pma_15_cfg_atomic),
    .io_check_env_pma_15_cfg_a(PMPChecker_io_check_env_pma_15_cfg_a),
    .io_check_env_pma_15_cfg_x(PMPChecker_io_check_env_pma_15_cfg_x),
    .io_check_env_pma_15_cfg_w(PMPChecker_io_check_env_pma_15_cfg_w),
    .io_check_env_pma_15_cfg_r(PMPChecker_io_check_env_pma_15_cfg_r),
    .io_check_env_pma_15_addr(PMPChecker_io_check_env_pma_15_addr),
    .io_check_env_pma_15_mask(PMPChecker_io_check_env_pma_15_mask),
    .io_req_bits_addr(PMPChecker_io_req_bits_addr),
    .io_req_bits_cmd(PMPChecker_io_req_bits_cmd),
    .io_resp_ld(PMPChecker_io_resp_ld),
    .io_resp_st(PMPChecker_io_resp_st),
    .io_resp_instr(PMPChecker_io_resp_instr),
    .io_resp_mmio(PMPChecker_io_resp_mmio),
    .io_resp_atomic(PMPChecker_io_resp_atomic)
  );
  PMPChecker PMPChecker_1 ( // @[L2TLB.scala 89:45]
    .io_check_env_mode(PMPChecker_1_io_check_env_mode),
    .io_check_env_pmp_0_cfg_l(PMPChecker_1_io_check_env_pmp_0_cfg_l),
    .io_check_env_pmp_0_cfg_a(PMPChecker_1_io_check_env_pmp_0_cfg_a),
    .io_check_env_pmp_0_cfg_x(PMPChecker_1_io_check_env_pmp_0_cfg_x),
    .io_check_env_pmp_0_cfg_w(PMPChecker_1_io_check_env_pmp_0_cfg_w),
    .io_check_env_pmp_0_cfg_r(PMPChecker_1_io_check_env_pmp_0_cfg_r),
    .io_check_env_pmp_0_addr(PMPChecker_1_io_check_env_pmp_0_addr),
    .io_check_env_pmp_0_mask(PMPChecker_1_io_check_env_pmp_0_mask),
    .io_check_env_pmp_1_cfg_l(PMPChecker_1_io_check_env_pmp_1_cfg_l),
    .io_check_env_pmp_1_cfg_a(PMPChecker_1_io_check_env_pmp_1_cfg_a),
    .io_check_env_pmp_1_cfg_x(PMPChecker_1_io_check_env_pmp_1_cfg_x),
    .io_check_env_pmp_1_cfg_w(PMPChecker_1_io_check_env_pmp_1_cfg_w),
    .io_check_env_pmp_1_cfg_r(PMPChecker_1_io_check_env_pmp_1_cfg_r),
    .io_check_env_pmp_1_addr(PMPChecker_1_io_check_env_pmp_1_addr),
    .io_check_env_pmp_1_mask(PMPChecker_1_io_check_env_pmp_1_mask),
    .io_check_env_pmp_2_cfg_l(PMPChecker_1_io_check_env_pmp_2_cfg_l),
    .io_check_env_pmp_2_cfg_a(PMPChecker_1_io_check_env_pmp_2_cfg_a),
    .io_check_env_pmp_2_cfg_x(PMPChecker_1_io_check_env_pmp_2_cfg_x),
    .io_check_env_pmp_2_cfg_w(PMPChecker_1_io_check_env_pmp_2_cfg_w),
    .io_check_env_pmp_2_cfg_r(PMPChecker_1_io_check_env_pmp_2_cfg_r),
    .io_check_env_pmp_2_addr(PMPChecker_1_io_check_env_pmp_2_addr),
    .io_check_env_pmp_2_mask(PMPChecker_1_io_check_env_pmp_2_mask),
    .io_check_env_pmp_3_cfg_l(PMPChecker_1_io_check_env_pmp_3_cfg_l),
    .io_check_env_pmp_3_cfg_a(PMPChecker_1_io_check_env_pmp_3_cfg_a),
    .io_check_env_pmp_3_cfg_x(PMPChecker_1_io_check_env_pmp_3_cfg_x),
    .io_check_env_pmp_3_cfg_w(PMPChecker_1_io_check_env_pmp_3_cfg_w),
    .io_check_env_pmp_3_cfg_r(PMPChecker_1_io_check_env_pmp_3_cfg_r),
    .io_check_env_pmp_3_addr(PMPChecker_1_io_check_env_pmp_3_addr),
    .io_check_env_pmp_3_mask(PMPChecker_1_io_check_env_pmp_3_mask),
    .io_check_env_pmp_4_cfg_l(PMPChecker_1_io_check_env_pmp_4_cfg_l),
    .io_check_env_pmp_4_cfg_a(PMPChecker_1_io_check_env_pmp_4_cfg_a),
    .io_check_env_pmp_4_cfg_x(PMPChecker_1_io_check_env_pmp_4_cfg_x),
    .io_check_env_pmp_4_cfg_w(PMPChecker_1_io_check_env_pmp_4_cfg_w),
    .io_check_env_pmp_4_cfg_r(PMPChecker_1_io_check_env_pmp_4_cfg_r),
    .io_check_env_pmp_4_addr(PMPChecker_1_io_check_env_pmp_4_addr),
    .io_check_env_pmp_4_mask(PMPChecker_1_io_check_env_pmp_4_mask),
    .io_check_env_pmp_5_cfg_l(PMPChecker_1_io_check_env_pmp_5_cfg_l),
    .io_check_env_pmp_5_cfg_a(PMPChecker_1_io_check_env_pmp_5_cfg_a),
    .io_check_env_pmp_5_cfg_x(PMPChecker_1_io_check_env_pmp_5_cfg_x),
    .io_check_env_pmp_5_cfg_w(PMPChecker_1_io_check_env_pmp_5_cfg_w),
    .io_check_env_pmp_5_cfg_r(PMPChecker_1_io_check_env_pmp_5_cfg_r),
    .io_check_env_pmp_5_addr(PMPChecker_1_io_check_env_pmp_5_addr),
    .io_check_env_pmp_5_mask(PMPChecker_1_io_check_env_pmp_5_mask),
    .io_check_env_pmp_6_cfg_l(PMPChecker_1_io_check_env_pmp_6_cfg_l),
    .io_check_env_pmp_6_cfg_a(PMPChecker_1_io_check_env_pmp_6_cfg_a),
    .io_check_env_pmp_6_cfg_x(PMPChecker_1_io_check_env_pmp_6_cfg_x),
    .io_check_env_pmp_6_cfg_w(PMPChecker_1_io_check_env_pmp_6_cfg_w),
    .io_check_env_pmp_6_cfg_r(PMPChecker_1_io_check_env_pmp_6_cfg_r),
    .io_check_env_pmp_6_addr(PMPChecker_1_io_check_env_pmp_6_addr),
    .io_check_env_pmp_6_mask(PMPChecker_1_io_check_env_pmp_6_mask),
    .io_check_env_pmp_7_cfg_l(PMPChecker_1_io_check_env_pmp_7_cfg_l),
    .io_check_env_pmp_7_cfg_a(PMPChecker_1_io_check_env_pmp_7_cfg_a),
    .io_check_env_pmp_7_cfg_x(PMPChecker_1_io_check_env_pmp_7_cfg_x),
    .io_check_env_pmp_7_cfg_w(PMPChecker_1_io_check_env_pmp_7_cfg_w),
    .io_check_env_pmp_7_cfg_r(PMPChecker_1_io_check_env_pmp_7_cfg_r),
    .io_check_env_pmp_7_addr(PMPChecker_1_io_check_env_pmp_7_addr),
    .io_check_env_pmp_7_mask(PMPChecker_1_io_check_env_pmp_7_mask),
    .io_check_env_pmp_8_cfg_l(PMPChecker_1_io_check_env_pmp_8_cfg_l),
    .io_check_env_pmp_8_cfg_a(PMPChecker_1_io_check_env_pmp_8_cfg_a),
    .io_check_env_pmp_8_cfg_x(PMPChecker_1_io_check_env_pmp_8_cfg_x),
    .io_check_env_pmp_8_cfg_w(PMPChecker_1_io_check_env_pmp_8_cfg_w),
    .io_check_env_pmp_8_cfg_r(PMPChecker_1_io_check_env_pmp_8_cfg_r),
    .io_check_env_pmp_8_addr(PMPChecker_1_io_check_env_pmp_8_addr),
    .io_check_env_pmp_8_mask(PMPChecker_1_io_check_env_pmp_8_mask),
    .io_check_env_pmp_9_cfg_l(PMPChecker_1_io_check_env_pmp_9_cfg_l),
    .io_check_env_pmp_9_cfg_a(PMPChecker_1_io_check_env_pmp_9_cfg_a),
    .io_check_env_pmp_9_cfg_x(PMPChecker_1_io_check_env_pmp_9_cfg_x),
    .io_check_env_pmp_9_cfg_w(PMPChecker_1_io_check_env_pmp_9_cfg_w),
    .io_check_env_pmp_9_cfg_r(PMPChecker_1_io_check_env_pmp_9_cfg_r),
    .io_check_env_pmp_9_addr(PMPChecker_1_io_check_env_pmp_9_addr),
    .io_check_env_pmp_9_mask(PMPChecker_1_io_check_env_pmp_9_mask),
    .io_check_env_pmp_10_cfg_l(PMPChecker_1_io_check_env_pmp_10_cfg_l),
    .io_check_env_pmp_10_cfg_a(PMPChecker_1_io_check_env_pmp_10_cfg_a),
    .io_check_env_pmp_10_cfg_x(PMPChecker_1_io_check_env_pmp_10_cfg_x),
    .io_check_env_pmp_10_cfg_w(PMPChecker_1_io_check_env_pmp_10_cfg_w),
    .io_check_env_pmp_10_cfg_r(PMPChecker_1_io_check_env_pmp_10_cfg_r),
    .io_check_env_pmp_10_addr(PMPChecker_1_io_check_env_pmp_10_addr),
    .io_check_env_pmp_10_mask(PMPChecker_1_io_check_env_pmp_10_mask),
    .io_check_env_pmp_11_cfg_l(PMPChecker_1_io_check_env_pmp_11_cfg_l),
    .io_check_env_pmp_11_cfg_a(PMPChecker_1_io_check_env_pmp_11_cfg_a),
    .io_check_env_pmp_11_cfg_x(PMPChecker_1_io_check_env_pmp_11_cfg_x),
    .io_check_env_pmp_11_cfg_w(PMPChecker_1_io_check_env_pmp_11_cfg_w),
    .io_check_env_pmp_11_cfg_r(PMPChecker_1_io_check_env_pmp_11_cfg_r),
    .io_check_env_pmp_11_addr(PMPChecker_1_io_check_env_pmp_11_addr),
    .io_check_env_pmp_11_mask(PMPChecker_1_io_check_env_pmp_11_mask),
    .io_check_env_pmp_12_cfg_l(PMPChecker_1_io_check_env_pmp_12_cfg_l),
    .io_check_env_pmp_12_cfg_a(PMPChecker_1_io_check_env_pmp_12_cfg_a),
    .io_check_env_pmp_12_cfg_x(PMPChecker_1_io_check_env_pmp_12_cfg_x),
    .io_check_env_pmp_12_cfg_w(PMPChecker_1_io_check_env_pmp_12_cfg_w),
    .io_check_env_pmp_12_cfg_r(PMPChecker_1_io_check_env_pmp_12_cfg_r),
    .io_check_env_pmp_12_addr(PMPChecker_1_io_check_env_pmp_12_addr),
    .io_check_env_pmp_12_mask(PMPChecker_1_io_check_env_pmp_12_mask),
    .io_check_env_pmp_13_cfg_l(PMPChecker_1_io_check_env_pmp_13_cfg_l),
    .io_check_env_pmp_13_cfg_a(PMPChecker_1_io_check_env_pmp_13_cfg_a),
    .io_check_env_pmp_13_cfg_x(PMPChecker_1_io_check_env_pmp_13_cfg_x),
    .io_check_env_pmp_13_cfg_w(PMPChecker_1_io_check_env_pmp_13_cfg_w),
    .io_check_env_pmp_13_cfg_r(PMPChecker_1_io_check_env_pmp_13_cfg_r),
    .io_check_env_pmp_13_addr(PMPChecker_1_io_check_env_pmp_13_addr),
    .io_check_env_pmp_13_mask(PMPChecker_1_io_check_env_pmp_13_mask),
    .io_check_env_pmp_14_cfg_l(PMPChecker_1_io_check_env_pmp_14_cfg_l),
    .io_check_env_pmp_14_cfg_a(PMPChecker_1_io_check_env_pmp_14_cfg_a),
    .io_check_env_pmp_14_cfg_x(PMPChecker_1_io_check_env_pmp_14_cfg_x),
    .io_check_env_pmp_14_cfg_w(PMPChecker_1_io_check_env_pmp_14_cfg_w),
    .io_check_env_pmp_14_cfg_r(PMPChecker_1_io_check_env_pmp_14_cfg_r),
    .io_check_env_pmp_14_addr(PMPChecker_1_io_check_env_pmp_14_addr),
    .io_check_env_pmp_14_mask(PMPChecker_1_io_check_env_pmp_14_mask),
    .io_check_env_pmp_15_cfg_l(PMPChecker_1_io_check_env_pmp_15_cfg_l),
    .io_check_env_pmp_15_cfg_a(PMPChecker_1_io_check_env_pmp_15_cfg_a),
    .io_check_env_pmp_15_cfg_x(PMPChecker_1_io_check_env_pmp_15_cfg_x),
    .io_check_env_pmp_15_cfg_w(PMPChecker_1_io_check_env_pmp_15_cfg_w),
    .io_check_env_pmp_15_cfg_r(PMPChecker_1_io_check_env_pmp_15_cfg_r),
    .io_check_env_pmp_15_addr(PMPChecker_1_io_check_env_pmp_15_addr),
    .io_check_env_pmp_15_mask(PMPChecker_1_io_check_env_pmp_15_mask),
    .io_check_env_pma_0_cfg_c(PMPChecker_1_io_check_env_pma_0_cfg_c),
    .io_check_env_pma_0_cfg_atomic(PMPChecker_1_io_check_env_pma_0_cfg_atomic),
    .io_check_env_pma_0_cfg_a(PMPChecker_1_io_check_env_pma_0_cfg_a),
    .io_check_env_pma_0_cfg_x(PMPChecker_1_io_check_env_pma_0_cfg_x),
    .io_check_env_pma_0_cfg_w(PMPChecker_1_io_check_env_pma_0_cfg_w),
    .io_check_env_pma_0_cfg_r(PMPChecker_1_io_check_env_pma_0_cfg_r),
    .io_check_env_pma_0_addr(PMPChecker_1_io_check_env_pma_0_addr),
    .io_check_env_pma_0_mask(PMPChecker_1_io_check_env_pma_0_mask),
    .io_check_env_pma_1_cfg_c(PMPChecker_1_io_check_env_pma_1_cfg_c),
    .io_check_env_pma_1_cfg_atomic(PMPChecker_1_io_check_env_pma_1_cfg_atomic),
    .io_check_env_pma_1_cfg_a(PMPChecker_1_io_check_env_pma_1_cfg_a),
    .io_check_env_pma_1_cfg_x(PMPChecker_1_io_check_env_pma_1_cfg_x),
    .io_check_env_pma_1_cfg_w(PMPChecker_1_io_check_env_pma_1_cfg_w),
    .io_check_env_pma_1_cfg_r(PMPChecker_1_io_check_env_pma_1_cfg_r),
    .io_check_env_pma_1_addr(PMPChecker_1_io_check_env_pma_1_addr),
    .io_check_env_pma_1_mask(PMPChecker_1_io_check_env_pma_1_mask),
    .io_check_env_pma_2_cfg_c(PMPChecker_1_io_check_env_pma_2_cfg_c),
    .io_check_env_pma_2_cfg_atomic(PMPChecker_1_io_check_env_pma_2_cfg_atomic),
    .io_check_env_pma_2_cfg_a(PMPChecker_1_io_check_env_pma_2_cfg_a),
    .io_check_env_pma_2_cfg_x(PMPChecker_1_io_check_env_pma_2_cfg_x),
    .io_check_env_pma_2_cfg_w(PMPChecker_1_io_check_env_pma_2_cfg_w),
    .io_check_env_pma_2_cfg_r(PMPChecker_1_io_check_env_pma_2_cfg_r),
    .io_check_env_pma_2_addr(PMPChecker_1_io_check_env_pma_2_addr),
    .io_check_env_pma_2_mask(PMPChecker_1_io_check_env_pma_2_mask),
    .io_check_env_pma_3_cfg_c(PMPChecker_1_io_check_env_pma_3_cfg_c),
    .io_check_env_pma_3_cfg_atomic(PMPChecker_1_io_check_env_pma_3_cfg_atomic),
    .io_check_env_pma_3_cfg_a(PMPChecker_1_io_check_env_pma_3_cfg_a),
    .io_check_env_pma_3_cfg_x(PMPChecker_1_io_check_env_pma_3_cfg_x),
    .io_check_env_pma_3_cfg_w(PMPChecker_1_io_check_env_pma_3_cfg_w),
    .io_check_env_pma_3_cfg_r(PMPChecker_1_io_check_env_pma_3_cfg_r),
    .io_check_env_pma_3_addr(PMPChecker_1_io_check_env_pma_3_addr),
    .io_check_env_pma_3_mask(PMPChecker_1_io_check_env_pma_3_mask),
    .io_check_env_pma_4_cfg_c(PMPChecker_1_io_check_env_pma_4_cfg_c),
    .io_check_env_pma_4_cfg_atomic(PMPChecker_1_io_check_env_pma_4_cfg_atomic),
    .io_check_env_pma_4_cfg_a(PMPChecker_1_io_check_env_pma_4_cfg_a),
    .io_check_env_pma_4_cfg_x(PMPChecker_1_io_check_env_pma_4_cfg_x),
    .io_check_env_pma_4_cfg_w(PMPChecker_1_io_check_env_pma_4_cfg_w),
    .io_check_env_pma_4_cfg_r(PMPChecker_1_io_check_env_pma_4_cfg_r),
    .io_check_env_pma_4_addr(PMPChecker_1_io_check_env_pma_4_addr),
    .io_check_env_pma_4_mask(PMPChecker_1_io_check_env_pma_4_mask),
    .io_check_env_pma_5_cfg_c(PMPChecker_1_io_check_env_pma_5_cfg_c),
    .io_check_env_pma_5_cfg_atomic(PMPChecker_1_io_check_env_pma_5_cfg_atomic),
    .io_check_env_pma_5_cfg_a(PMPChecker_1_io_check_env_pma_5_cfg_a),
    .io_check_env_pma_5_cfg_x(PMPChecker_1_io_check_env_pma_5_cfg_x),
    .io_check_env_pma_5_cfg_w(PMPChecker_1_io_check_env_pma_5_cfg_w),
    .io_check_env_pma_5_cfg_r(PMPChecker_1_io_check_env_pma_5_cfg_r),
    .io_check_env_pma_5_addr(PMPChecker_1_io_check_env_pma_5_addr),
    .io_check_env_pma_5_mask(PMPChecker_1_io_check_env_pma_5_mask),
    .io_check_env_pma_6_cfg_c(PMPChecker_1_io_check_env_pma_6_cfg_c),
    .io_check_env_pma_6_cfg_atomic(PMPChecker_1_io_check_env_pma_6_cfg_atomic),
    .io_check_env_pma_6_cfg_a(PMPChecker_1_io_check_env_pma_6_cfg_a),
    .io_check_env_pma_6_cfg_x(PMPChecker_1_io_check_env_pma_6_cfg_x),
    .io_check_env_pma_6_cfg_w(PMPChecker_1_io_check_env_pma_6_cfg_w),
    .io_check_env_pma_6_cfg_r(PMPChecker_1_io_check_env_pma_6_cfg_r),
    .io_check_env_pma_6_addr(PMPChecker_1_io_check_env_pma_6_addr),
    .io_check_env_pma_6_mask(PMPChecker_1_io_check_env_pma_6_mask),
    .io_check_env_pma_7_cfg_c(PMPChecker_1_io_check_env_pma_7_cfg_c),
    .io_check_env_pma_7_cfg_atomic(PMPChecker_1_io_check_env_pma_7_cfg_atomic),
    .io_check_env_pma_7_cfg_a(PMPChecker_1_io_check_env_pma_7_cfg_a),
    .io_check_env_pma_7_cfg_x(PMPChecker_1_io_check_env_pma_7_cfg_x),
    .io_check_env_pma_7_cfg_w(PMPChecker_1_io_check_env_pma_7_cfg_w),
    .io_check_env_pma_7_cfg_r(PMPChecker_1_io_check_env_pma_7_cfg_r),
    .io_check_env_pma_7_addr(PMPChecker_1_io_check_env_pma_7_addr),
    .io_check_env_pma_7_mask(PMPChecker_1_io_check_env_pma_7_mask),
    .io_check_env_pma_8_cfg_c(PMPChecker_1_io_check_env_pma_8_cfg_c),
    .io_check_env_pma_8_cfg_atomic(PMPChecker_1_io_check_env_pma_8_cfg_atomic),
    .io_check_env_pma_8_cfg_a(PMPChecker_1_io_check_env_pma_8_cfg_a),
    .io_check_env_pma_8_cfg_x(PMPChecker_1_io_check_env_pma_8_cfg_x),
    .io_check_env_pma_8_cfg_w(PMPChecker_1_io_check_env_pma_8_cfg_w),
    .io_check_env_pma_8_cfg_r(PMPChecker_1_io_check_env_pma_8_cfg_r),
    .io_check_env_pma_8_addr(PMPChecker_1_io_check_env_pma_8_addr),
    .io_check_env_pma_8_mask(PMPChecker_1_io_check_env_pma_8_mask),
    .io_check_env_pma_9_cfg_c(PMPChecker_1_io_check_env_pma_9_cfg_c),
    .io_check_env_pma_9_cfg_atomic(PMPChecker_1_io_check_env_pma_9_cfg_atomic),
    .io_check_env_pma_9_cfg_a(PMPChecker_1_io_check_env_pma_9_cfg_a),
    .io_check_env_pma_9_cfg_x(PMPChecker_1_io_check_env_pma_9_cfg_x),
    .io_check_env_pma_9_cfg_w(PMPChecker_1_io_check_env_pma_9_cfg_w),
    .io_check_env_pma_9_cfg_r(PMPChecker_1_io_check_env_pma_9_cfg_r),
    .io_check_env_pma_9_addr(PMPChecker_1_io_check_env_pma_9_addr),
    .io_check_env_pma_9_mask(PMPChecker_1_io_check_env_pma_9_mask),
    .io_check_env_pma_10_cfg_c(PMPChecker_1_io_check_env_pma_10_cfg_c),
    .io_check_env_pma_10_cfg_atomic(PMPChecker_1_io_check_env_pma_10_cfg_atomic),
    .io_check_env_pma_10_cfg_a(PMPChecker_1_io_check_env_pma_10_cfg_a),
    .io_check_env_pma_10_cfg_x(PMPChecker_1_io_check_env_pma_10_cfg_x),
    .io_check_env_pma_10_cfg_w(PMPChecker_1_io_check_env_pma_10_cfg_w),
    .io_check_env_pma_10_cfg_r(PMPChecker_1_io_check_env_pma_10_cfg_r),
    .io_check_env_pma_10_addr(PMPChecker_1_io_check_env_pma_10_addr),
    .io_check_env_pma_10_mask(PMPChecker_1_io_check_env_pma_10_mask),
    .io_check_env_pma_11_cfg_c(PMPChecker_1_io_check_env_pma_11_cfg_c),
    .io_check_env_pma_11_cfg_atomic(PMPChecker_1_io_check_env_pma_11_cfg_atomic),
    .io_check_env_pma_11_cfg_a(PMPChecker_1_io_check_env_pma_11_cfg_a),
    .io_check_env_pma_11_cfg_x(PMPChecker_1_io_check_env_pma_11_cfg_x),
    .io_check_env_pma_11_cfg_w(PMPChecker_1_io_check_env_pma_11_cfg_w),
    .io_check_env_pma_11_cfg_r(PMPChecker_1_io_check_env_pma_11_cfg_r),
    .io_check_env_pma_11_addr(PMPChecker_1_io_check_env_pma_11_addr),
    .io_check_env_pma_11_mask(PMPChecker_1_io_check_env_pma_11_mask),
    .io_check_env_pma_12_cfg_c(PMPChecker_1_io_check_env_pma_12_cfg_c),
    .io_check_env_pma_12_cfg_atomic(PMPChecker_1_io_check_env_pma_12_cfg_atomic),
    .io_check_env_pma_12_cfg_a(PMPChecker_1_io_check_env_pma_12_cfg_a),
    .io_check_env_pma_12_cfg_x(PMPChecker_1_io_check_env_pma_12_cfg_x),
    .io_check_env_pma_12_cfg_w(PMPChecker_1_io_check_env_pma_12_cfg_w),
    .io_check_env_pma_12_cfg_r(PMPChecker_1_io_check_env_pma_12_cfg_r),
    .io_check_env_pma_12_addr(PMPChecker_1_io_check_env_pma_12_addr),
    .io_check_env_pma_12_mask(PMPChecker_1_io_check_env_pma_12_mask),
    .io_check_env_pma_13_cfg_c(PMPChecker_1_io_check_env_pma_13_cfg_c),
    .io_check_env_pma_13_cfg_atomic(PMPChecker_1_io_check_env_pma_13_cfg_atomic),
    .io_check_env_pma_13_cfg_a(PMPChecker_1_io_check_env_pma_13_cfg_a),
    .io_check_env_pma_13_cfg_x(PMPChecker_1_io_check_env_pma_13_cfg_x),
    .io_check_env_pma_13_cfg_w(PMPChecker_1_io_check_env_pma_13_cfg_w),
    .io_check_env_pma_13_cfg_r(PMPChecker_1_io_check_env_pma_13_cfg_r),
    .io_check_env_pma_13_addr(PMPChecker_1_io_check_env_pma_13_addr),
    .io_check_env_pma_13_mask(PMPChecker_1_io_check_env_pma_13_mask),
    .io_check_env_pma_14_cfg_c(PMPChecker_1_io_check_env_pma_14_cfg_c),
    .io_check_env_pma_14_cfg_atomic(PMPChecker_1_io_check_env_pma_14_cfg_atomic),
    .io_check_env_pma_14_cfg_a(PMPChecker_1_io_check_env_pma_14_cfg_a),
    .io_check_env_pma_14_cfg_x(PMPChecker_1_io_check_env_pma_14_cfg_x),
    .io_check_env_pma_14_cfg_w(PMPChecker_1_io_check_env_pma_14_cfg_w),
    .io_check_env_pma_14_cfg_r(PMPChecker_1_io_check_env_pma_14_cfg_r),
    .io_check_env_pma_14_addr(PMPChecker_1_io_check_env_pma_14_addr),
    .io_check_env_pma_14_mask(PMPChecker_1_io_check_env_pma_14_mask),
    .io_check_env_pma_15_cfg_c(PMPChecker_1_io_check_env_pma_15_cfg_c),
    .io_check_env_pma_15_cfg_atomic(PMPChecker_1_io_check_env_pma_15_cfg_atomic),
    .io_check_env_pma_15_cfg_a(PMPChecker_1_io_check_env_pma_15_cfg_a),
    .io_check_env_pma_15_cfg_x(PMPChecker_1_io_check_env_pma_15_cfg_x),
    .io_check_env_pma_15_cfg_w(PMPChecker_1_io_check_env_pma_15_cfg_w),
    .io_check_env_pma_15_cfg_r(PMPChecker_1_io_check_env_pma_15_cfg_r),
    .io_check_env_pma_15_addr(PMPChecker_1_io_check_env_pma_15_addr),
    .io_check_env_pma_15_mask(PMPChecker_1_io_check_env_pma_15_mask),
    .io_req_bits_addr(PMPChecker_1_io_req_bits_addr),
    .io_req_bits_cmd(PMPChecker_1_io_req_bits_cmd),
    .io_resp_ld(PMPChecker_1_io_resp_ld),
    .io_resp_st(PMPChecker_1_io_resp_st),
    .io_resp_instr(PMPChecker_1_io_resp_instr),
    .io_resp_mmio(PMPChecker_1_io_resp_mmio),
    .io_resp_atomic(PMPChecker_1_io_resp_atomic)
  );
  L2TlbMissQueue missQueue ( // @[L2TLB.scala 93:25]
    .clock(missQueue_clock),
    .reset(missQueue_reset),
    .io_sfence_valid(missQueue_io_sfence_valid),
    .io_csr_satp_changed(missQueue_io_csr_satp_changed),
    .io_in_ready(missQueue_io_in_ready),
    .io_in_valid(missQueue_io_in_valid),
    .io_in_bits_vpn(missQueue_io_in_bits_vpn),
    .io_in_bits_source(missQueue_io_in_bits_source),
    .io_out_ready(missQueue_io_out_ready),
    .io_out_valid(missQueue_io_out_valid),
    .io_out_bits_vpn(missQueue_io_out_bits_vpn),
    .io_out_bits_source(missQueue_io_out_bits_source)
  );
  PtwCache cache ( // @[L2TLB.scala 94:21]
    .clock(cache_clock),
    .reset(cache_reset),
    .io_req_ready(cache_io_req_ready),
    .io_req_valid(cache_io_req_valid),
    .io_req_bits_req_info_vpn(cache_io_req_bits_req_info_vpn),
    .io_req_bits_req_info_source(cache_io_req_bits_req_info_source),
    .io_req_bits_isFirst(cache_io_req_bits_isFirst),
    .io_resp_ready(cache_io_resp_ready),
    .io_resp_valid(cache_io_resp_valid),
    .io_resp_bits_req_info_vpn(cache_io_resp_bits_req_info_vpn),
    .io_resp_bits_req_info_source(cache_io_resp_bits_req_info_source),
    .io_resp_bits_isFirst(cache_io_resp_bits_isFirst),
    .io_resp_bits_hit(cache_io_resp_bits_hit),
    .io_resp_bits_prefetch(cache_io_resp_bits_prefetch),
    .io_resp_bits_bypassed(cache_io_resp_bits_bypassed),
    .io_resp_bits_toFsm_l1Hit(cache_io_resp_bits_toFsm_l1Hit),
    .io_resp_bits_toFsm_l2Hit(cache_io_resp_bits_toFsm_l2Hit),
    .io_resp_bits_toFsm_ppn(cache_io_resp_bits_toFsm_ppn),
    .io_resp_bits_toTlb_tag(cache_io_resp_bits_toTlb_tag),
    .io_resp_bits_toTlb_asid(cache_io_resp_bits_toTlb_asid),
    .io_resp_bits_toTlb_ppn(cache_io_resp_bits_toTlb_ppn),
    .io_resp_bits_toTlb_perm_d(cache_io_resp_bits_toTlb_perm_d),
    .io_resp_bits_toTlb_perm_a(cache_io_resp_bits_toTlb_perm_a),
    .io_resp_bits_toTlb_perm_g(cache_io_resp_bits_toTlb_perm_g),
    .io_resp_bits_toTlb_perm_u(cache_io_resp_bits_toTlb_perm_u),
    .io_resp_bits_toTlb_perm_x(cache_io_resp_bits_toTlb_perm_x),
    .io_resp_bits_toTlb_perm_w(cache_io_resp_bits_toTlb_perm_w),
    .io_resp_bits_toTlb_perm_r(cache_io_resp_bits_toTlb_perm_r),
    .io_resp_bits_toTlb_level(cache_io_resp_bits_toTlb_level),
    .io_resp_bits_toTlb_prefetch(cache_io_resp_bits_toTlb_prefetch),
    .io_resp_bits_toTlb_v(cache_io_resp_bits_toTlb_v),
    .io_refill_valid(cache_io_refill_valid),
    .io_refill_bits_ptes(cache_io_refill_bits_ptes),
    .io_refill_bits_levelOH_sp(cache_io_refill_bits_levelOH_sp),
    .io_refill_bits_levelOH_l3(cache_io_refill_bits_levelOH_l3),
    .io_refill_bits_levelOH_l2(cache_io_refill_bits_levelOH_l2),
    .io_refill_bits_levelOH_l1(cache_io_refill_bits_levelOH_l1),
    .io_refill_bits_req_info_dup_0_vpn(cache_io_refill_bits_req_info_dup_0_vpn),
    .io_refill_bits_req_info_dup_0_source(cache_io_refill_bits_req_info_dup_0_source),
    .io_refill_bits_req_info_dup_1_vpn(cache_io_refill_bits_req_info_dup_1_vpn),
    .io_refill_bits_req_info_dup_1_source(cache_io_refill_bits_req_info_dup_1_source),
    .io_refill_bits_req_info_dup_2_vpn(cache_io_refill_bits_req_info_dup_2_vpn),
    .io_refill_bits_req_info_dup_2_source(cache_io_refill_bits_req_info_dup_2_source),
    .io_refill_bits_level_dup_0(cache_io_refill_bits_level_dup_0),
    .io_refill_bits_level_dup_1(cache_io_refill_bits_level_dup_1),
    .io_refill_bits_level_dup_2(cache_io_refill_bits_level_dup_2),
    .io_refill_bits_sel_pte_dup_0(cache_io_refill_bits_sel_pte_dup_0),
    .io_refill_bits_sel_pte_dup_1(cache_io_refill_bits_sel_pte_dup_1),
    .io_refill_bits_sel_pte_dup_2(cache_io_refill_bits_sel_pte_dup_2),
    .io_sfence_dup_0_valid(cache_io_sfence_dup_0_valid),
    .io_sfence_dup_0_bits_rs1(cache_io_sfence_dup_0_bits_rs1),
    .io_sfence_dup_0_bits_rs2(cache_io_sfence_dup_0_bits_rs2),
    .io_sfence_dup_0_bits_addr(cache_io_sfence_dup_0_bits_addr),
    .io_sfence_dup_0_bits_asid(cache_io_sfence_dup_0_bits_asid),
    .io_sfence_dup_1_valid(cache_io_sfence_dup_1_valid),
    .io_sfence_dup_2_valid(cache_io_sfence_dup_2_valid),
    .io_sfence_dup_3_valid(cache_io_sfence_dup_3_valid),
    .io_sfence_dup_3_bits_rs1(cache_io_sfence_dup_3_bits_rs1),
    .io_sfence_dup_3_bits_rs2(cache_io_sfence_dup_3_bits_rs2),
    .io_sfence_dup_3_bits_addr(cache_io_sfence_dup_3_bits_addr),
    .io_csr_dup_0_satp_asid(cache_io_csr_dup_0_satp_asid),
    .io_csr_dup_0_satp_changed(cache_io_csr_dup_0_satp_changed),
    .io_csr_dup_1_satp_asid(cache_io_csr_dup_1_satp_asid),
    .io_csr_dup_1_satp_changed(cache_io_csr_dup_1_satp_changed),
    .io_csr_dup_2_satp_asid(cache_io_csr_dup_2_satp_asid),
    .io_csr_dup_2_satp_changed(cache_io_csr_dup_2_satp_changed),
    .io_perf_0_value(cache_io_perf_0_value),
    .io_perf_1_value(cache_io_perf_1_value),
    .io_perf_2_value(cache_io_perf_2_value),
    .io_perf_3_value(cache_io_perf_3_value),
    .io_perf_4_value(cache_io_perf_4_value),
    .io_perf_5_value(cache_io_perf_5_value),
    .io_perf_6_value(cache_io_perf_6_value),
    .io_perf_7_value(cache_io_perf_7_value)
  );
  PTW ptw ( // @[L2TLB.scala 95:19]
    .clock(ptw_clock),
    .reset(ptw_reset),
    .io_sfence_valid(ptw_io_sfence_valid),
    .io_csr_satp_asid(ptw_io_csr_satp_asid),
    .io_csr_satp_ppn(ptw_io_csr_satp_ppn),
    .io_req_ready(ptw_io_req_ready),
    .io_req_valid(ptw_io_req_valid),
    .io_req_bits_req_info_vpn(ptw_io_req_bits_req_info_vpn),
    .io_req_bits_req_info_source(ptw_io_req_bits_req_info_source),
    .io_req_bits_l1Hit(ptw_io_req_bits_l1Hit),
    .io_req_bits_ppn(ptw_io_req_bits_ppn),
    .io_resp_ready(ptw_io_resp_ready),
    .io_resp_valid(ptw_io_resp_valid),
    .io_resp_bits_source(ptw_io_resp_bits_source),
    .io_resp_bits_resp_entry_tag(ptw_io_resp_bits_resp_entry_tag),
    .io_resp_bits_resp_entry_asid(ptw_io_resp_bits_resp_entry_asid),
    .io_resp_bits_resp_entry_ppn(ptw_io_resp_bits_resp_entry_ppn),
    .io_resp_bits_resp_entry_perm_d(ptw_io_resp_bits_resp_entry_perm_d),
    .io_resp_bits_resp_entry_perm_a(ptw_io_resp_bits_resp_entry_perm_a),
    .io_resp_bits_resp_entry_perm_g(ptw_io_resp_bits_resp_entry_perm_g),
    .io_resp_bits_resp_entry_perm_u(ptw_io_resp_bits_resp_entry_perm_u),
    .io_resp_bits_resp_entry_perm_x(ptw_io_resp_bits_resp_entry_perm_x),
    .io_resp_bits_resp_entry_perm_w(ptw_io_resp_bits_resp_entry_perm_w),
    .io_resp_bits_resp_entry_perm_r(ptw_io_resp_bits_resp_entry_perm_r),
    .io_resp_bits_resp_entry_level(ptw_io_resp_bits_resp_entry_level),
    .io_resp_bits_resp_pf(ptw_io_resp_bits_resp_pf),
    .io_resp_bits_resp_af(ptw_io_resp_bits_resp_af),
    .io_llptw_ready(ptw_io_llptw_ready),
    .io_llptw_valid(ptw_io_llptw_valid),
    .io_llptw_bits_req_info_vpn(ptw_io_llptw_bits_req_info_vpn),
    .io_llptw_bits_req_info_source(ptw_io_llptw_bits_req_info_source),
    .io_mem_req_ready(ptw_io_mem_req_ready),
    .io_mem_req_valid(ptw_io_mem_req_valid),
    .io_mem_req_bits_addr(ptw_io_mem_req_bits_addr),
    .io_mem_resp_valid(ptw_io_mem_resp_valid),
    .io_mem_resp_bits(ptw_io_mem_resp_bits),
    .io_mem_mask(ptw_io_mem_mask),
    .io_pmp_req_bits_addr(ptw_io_pmp_req_bits_addr),
    .io_pmp_resp_ld(ptw_io_pmp_resp_ld),
    .io_pmp_resp_mmio(ptw_io_pmp_resp_mmio),
    .io_refill_req_info_vpn(ptw_io_refill_req_info_vpn),
    .io_refill_req_info_source(ptw_io_refill_req_info_source),
    .io_refill_level(ptw_io_refill_level),
    .io_perf_0_value(ptw_io_perf_0_value),
    .io_perf_1_value(ptw_io_perf_1_value),
    .io_perf_2_value(ptw_io_perf_2_value),
    .io_perf_3_value(ptw_io_perf_3_value),
    .io_perf_4_value(ptw_io_perf_4_value),
    .io_perf_5_value(ptw_io_perf_5_value),
    .io_perf_6_value(ptw_io_perf_6_value)
  );
  LLPTW llptw ( // @[L2TLB.scala 96:21]
    .clock(llptw_clock),
    .reset(llptw_reset),
    .io_sfence_valid(llptw_io_sfence_valid),
    .io_csr_satp_changed(llptw_io_csr_satp_changed),
    .io_in_ready(llptw_io_in_ready),
    .io_in_valid(llptw_io_in_valid),
    .io_in_bits_req_info_vpn(llptw_io_in_bits_req_info_vpn),
    .io_in_bits_req_info_source(llptw_io_in_bits_req_info_source),
    .io_in_bits_ppn(llptw_io_in_bits_ppn),
    .io_out_ready(llptw_io_out_ready),
    .io_out_valid(llptw_io_out_valid),
    .io_out_bits_req_info_vpn(llptw_io_out_bits_req_info_vpn),
    .io_out_bits_req_info_source(llptw_io_out_bits_req_info_source),
    .io_out_bits_id(llptw_io_out_bits_id),
    .io_out_bits_af(llptw_io_out_bits_af),
    .io_mem_req_ready(llptw_io_mem_req_ready),
    .io_mem_req_valid(llptw_io_mem_req_valid),
    .io_mem_req_bits_addr(llptw_io_mem_req_bits_addr),
    .io_mem_req_bits_id(llptw_io_mem_req_bits_id),
    .io_mem_resp_valid(llptw_io_mem_resp_valid),
    .io_mem_resp_bits_id(llptw_io_mem_resp_bits_id),
    .io_mem_enq_ptr(llptw_io_mem_enq_ptr),
    .io_mem_buffer_it_0(llptw_io_mem_buffer_it_0),
    .io_mem_buffer_it_1(llptw_io_mem_buffer_it_1),
    .io_mem_buffer_it_2(llptw_io_mem_buffer_it_2),
    .io_mem_buffer_it_3(llptw_io_mem_buffer_it_3),
    .io_mem_buffer_it_4(llptw_io_mem_buffer_it_4),
    .io_mem_buffer_it_5(llptw_io_mem_buffer_it_5),
    .io_mem_refill_vpn(llptw_io_mem_refill_vpn),
    .io_mem_refill_source(llptw_io_mem_refill_source),
    .io_mem_req_mask_0(llptw_io_mem_req_mask_0),
    .io_mem_req_mask_1(llptw_io_mem_req_mask_1),
    .io_mem_req_mask_2(llptw_io_mem_req_mask_2),
    .io_mem_req_mask_3(llptw_io_mem_req_mask_3),
    .io_mem_req_mask_4(llptw_io_mem_req_mask_4),
    .io_mem_req_mask_5(llptw_io_mem_req_mask_5),
    .io_cache_ready(llptw_io_cache_ready),
    .io_cache_valid(llptw_io_cache_valid),
    .io_cache_bits_vpn(llptw_io_cache_bits_vpn),
    .io_cache_bits_source(llptw_io_cache_bits_source),
    .io_pmp_req_valid(llptw_io_pmp_req_valid),
    .io_pmp_req_bits_addr(llptw_io_pmp_req_bits_addr),
    .io_pmp_resp_ld(llptw_io_pmp_resp_ld),
    .io_pmp_resp_mmio(llptw_io_pmp_resp_mmio),
    .io_perf_0_value(llptw_io_perf_0_value),
    .io_perf_1_value(llptw_io_perf_1_value),
    .io_perf_2_value(llptw_io_perf_2_value),
    .io_perf_3_value(llptw_io_perf_3_value)
  );
  Arbiter_8 arb1 ( // @[L2TLB.scala 98:20]
    .io_in_0_ready(arb1_io_in_0_ready),
    .io_in_0_valid(arb1_io_in_0_valid),
    .io_in_0_bits_vpn(arb1_io_in_0_bits_vpn),
    .io_in_1_ready(arb1_io_in_1_ready),
    .io_in_1_valid(arb1_io_in_1_valid),
    .io_in_1_bits_vpn(arb1_io_in_1_bits_vpn),
    .io_out_ready(arb1_io_out_ready),
    .io_out_valid(arb1_io_out_valid),
    .io_out_bits_vpn(arb1_io_out_bits_vpn),
    .io_chosen(arb1_io_chosen)
  );
  Arbiter_9 arb2 ( // @[L2TLB.scala 99:20]
    .io_in_0_ready(arb2_io_in_0_ready),
    .io_in_0_valid(arb2_io_in_0_valid),
    .io_in_0_bits_vpn(arb2_io_in_0_bits_vpn),
    .io_in_0_bits_source(arb2_io_in_0_bits_source),
    .io_in_1_ready(arb2_io_in_1_ready),
    .io_in_1_valid(arb2_io_in_1_valid),
    .io_in_1_bits_vpn(arb2_io_in_1_bits_vpn),
    .io_in_1_bits_source(arb2_io_in_1_bits_source),
    .io_in_2_ready(arb2_io_in_2_ready),
    .io_in_2_valid(arb2_io_in_2_valid),
    .io_in_2_bits_vpn(arb2_io_in_2_bits_vpn),
    .io_in_2_bits_source(arb2_io_in_2_bits_source),
    .io_in_3_ready(arb2_io_in_3_ready),
    .io_in_3_valid(arb2_io_in_3_valid),
    .io_in_3_bits_vpn(arb2_io_in_3_bits_vpn),
    .io_out_ready(arb2_io_out_ready),
    .io_out_valid(arb2_io_out_valid),
    .io_out_bits_vpn(arb2_io_out_bits_vpn),
    .io_out_bits_source(arb2_io_out_bits_source),
    .io_chosen(arb2_io_chosen)
  );
  Arbiter_10 Arbiter ( // @[L2TLB.scala 103:50]
    .io_in_0_ready(Arbiter_io_in_0_ready),
    .io_in_0_valid(Arbiter_io_in_0_valid),
    .io_in_0_bits_entry_tag(Arbiter_io_in_0_bits_entry_tag),
    .io_in_0_bits_entry_asid(Arbiter_io_in_0_bits_entry_asid),
    .io_in_0_bits_entry_ppn(Arbiter_io_in_0_bits_entry_ppn),
    .io_in_0_bits_entry_perm_d(Arbiter_io_in_0_bits_entry_perm_d),
    .io_in_0_bits_entry_perm_a(Arbiter_io_in_0_bits_entry_perm_a),
    .io_in_0_bits_entry_perm_g(Arbiter_io_in_0_bits_entry_perm_g),
    .io_in_0_bits_entry_perm_u(Arbiter_io_in_0_bits_entry_perm_u),
    .io_in_0_bits_entry_perm_x(Arbiter_io_in_0_bits_entry_perm_x),
    .io_in_0_bits_entry_perm_w(Arbiter_io_in_0_bits_entry_perm_w),
    .io_in_0_bits_entry_perm_r(Arbiter_io_in_0_bits_entry_perm_r),
    .io_in_0_bits_entry_level(Arbiter_io_in_0_bits_entry_level),
    .io_in_0_bits_pf(Arbiter_io_in_0_bits_pf),
    .io_in_1_ready(Arbiter_io_in_1_ready),
    .io_in_1_valid(Arbiter_io_in_1_valid),
    .io_in_1_bits_entry_tag(Arbiter_io_in_1_bits_entry_tag),
    .io_in_1_bits_entry_asid(Arbiter_io_in_1_bits_entry_asid),
    .io_in_1_bits_entry_ppn(Arbiter_io_in_1_bits_entry_ppn),
    .io_in_1_bits_entry_perm_d(Arbiter_io_in_1_bits_entry_perm_d),
    .io_in_1_bits_entry_perm_a(Arbiter_io_in_1_bits_entry_perm_a),
    .io_in_1_bits_entry_perm_g(Arbiter_io_in_1_bits_entry_perm_g),
    .io_in_1_bits_entry_perm_u(Arbiter_io_in_1_bits_entry_perm_u),
    .io_in_1_bits_entry_perm_x(Arbiter_io_in_1_bits_entry_perm_x),
    .io_in_1_bits_entry_perm_w(Arbiter_io_in_1_bits_entry_perm_w),
    .io_in_1_bits_entry_perm_r(Arbiter_io_in_1_bits_entry_perm_r),
    .io_in_1_bits_entry_level(Arbiter_io_in_1_bits_entry_level),
    .io_in_1_bits_pf(Arbiter_io_in_1_bits_pf),
    .io_in_1_bits_af(Arbiter_io_in_1_bits_af),
    .io_in_2_ready(Arbiter_io_in_2_ready),
    .io_in_2_valid(Arbiter_io_in_2_valid),
    .io_in_2_bits_entry_tag(Arbiter_io_in_2_bits_entry_tag),
    .io_in_2_bits_entry_asid(Arbiter_io_in_2_bits_entry_asid),
    .io_in_2_bits_entry_ppn(Arbiter_io_in_2_bits_entry_ppn),
    .io_in_2_bits_entry_perm_d(Arbiter_io_in_2_bits_entry_perm_d),
    .io_in_2_bits_entry_perm_a(Arbiter_io_in_2_bits_entry_perm_a),
    .io_in_2_bits_entry_perm_g(Arbiter_io_in_2_bits_entry_perm_g),
    .io_in_2_bits_entry_perm_u(Arbiter_io_in_2_bits_entry_perm_u),
    .io_in_2_bits_entry_perm_x(Arbiter_io_in_2_bits_entry_perm_x),
    .io_in_2_bits_entry_perm_w(Arbiter_io_in_2_bits_entry_perm_w),
    .io_in_2_bits_entry_perm_r(Arbiter_io_in_2_bits_entry_perm_r),
    .io_in_2_bits_pf(Arbiter_io_in_2_bits_pf),
    .io_in_2_bits_af(Arbiter_io_in_2_bits_af),
    .io_out_ready(Arbiter_io_out_ready),
    .io_out_valid(Arbiter_io_out_valid),
    .io_out_bits_entry_tag(Arbiter_io_out_bits_entry_tag),
    .io_out_bits_entry_asid(Arbiter_io_out_bits_entry_asid),
    .io_out_bits_entry_ppn(Arbiter_io_out_bits_entry_ppn),
    .io_out_bits_entry_perm_d(Arbiter_io_out_bits_entry_perm_d),
    .io_out_bits_entry_perm_a(Arbiter_io_out_bits_entry_perm_a),
    .io_out_bits_entry_perm_g(Arbiter_io_out_bits_entry_perm_g),
    .io_out_bits_entry_perm_u(Arbiter_io_out_bits_entry_perm_u),
    .io_out_bits_entry_perm_x(Arbiter_io_out_bits_entry_perm_x),
    .io_out_bits_entry_perm_w(Arbiter_io_out_bits_entry_perm_w),
    .io_out_bits_entry_perm_r(Arbiter_io_out_bits_entry_perm_r),
    .io_out_bits_entry_level(Arbiter_io_out_bits_entry_level),
    .io_out_bits_pf(Arbiter_io_out_bits_pf),
    .io_out_bits_af(Arbiter_io_out_bits_af)
  );
  Arbiter_10 Arbiter_1 ( // @[L2TLB.scala 103:50]
    .io_in_0_ready(Arbiter_1_io_in_0_ready),
    .io_in_0_valid(Arbiter_1_io_in_0_valid),
    .io_in_0_bits_entry_tag(Arbiter_1_io_in_0_bits_entry_tag),
    .io_in_0_bits_entry_asid(Arbiter_1_io_in_0_bits_entry_asid),
    .io_in_0_bits_entry_ppn(Arbiter_1_io_in_0_bits_entry_ppn),
    .io_in_0_bits_entry_perm_d(Arbiter_1_io_in_0_bits_entry_perm_d),
    .io_in_0_bits_entry_perm_a(Arbiter_1_io_in_0_bits_entry_perm_a),
    .io_in_0_bits_entry_perm_g(Arbiter_1_io_in_0_bits_entry_perm_g),
    .io_in_0_bits_entry_perm_u(Arbiter_1_io_in_0_bits_entry_perm_u),
    .io_in_0_bits_entry_perm_x(Arbiter_1_io_in_0_bits_entry_perm_x),
    .io_in_0_bits_entry_perm_w(Arbiter_1_io_in_0_bits_entry_perm_w),
    .io_in_0_bits_entry_perm_r(Arbiter_1_io_in_0_bits_entry_perm_r),
    .io_in_0_bits_entry_level(Arbiter_1_io_in_0_bits_entry_level),
    .io_in_0_bits_pf(Arbiter_1_io_in_0_bits_pf),
    .io_in_1_ready(Arbiter_1_io_in_1_ready),
    .io_in_1_valid(Arbiter_1_io_in_1_valid),
    .io_in_1_bits_entry_tag(Arbiter_1_io_in_1_bits_entry_tag),
    .io_in_1_bits_entry_asid(Arbiter_1_io_in_1_bits_entry_asid),
    .io_in_1_bits_entry_ppn(Arbiter_1_io_in_1_bits_entry_ppn),
    .io_in_1_bits_entry_perm_d(Arbiter_1_io_in_1_bits_entry_perm_d),
    .io_in_1_bits_entry_perm_a(Arbiter_1_io_in_1_bits_entry_perm_a),
    .io_in_1_bits_entry_perm_g(Arbiter_1_io_in_1_bits_entry_perm_g),
    .io_in_1_bits_entry_perm_u(Arbiter_1_io_in_1_bits_entry_perm_u),
    .io_in_1_bits_entry_perm_x(Arbiter_1_io_in_1_bits_entry_perm_x),
    .io_in_1_bits_entry_perm_w(Arbiter_1_io_in_1_bits_entry_perm_w),
    .io_in_1_bits_entry_perm_r(Arbiter_1_io_in_1_bits_entry_perm_r),
    .io_in_1_bits_entry_level(Arbiter_1_io_in_1_bits_entry_level),
    .io_in_1_bits_pf(Arbiter_1_io_in_1_bits_pf),
    .io_in_1_bits_af(Arbiter_1_io_in_1_bits_af),
    .io_in_2_ready(Arbiter_1_io_in_2_ready),
    .io_in_2_valid(Arbiter_1_io_in_2_valid),
    .io_in_2_bits_entry_tag(Arbiter_1_io_in_2_bits_entry_tag),
    .io_in_2_bits_entry_asid(Arbiter_1_io_in_2_bits_entry_asid),
    .io_in_2_bits_entry_ppn(Arbiter_1_io_in_2_bits_entry_ppn),
    .io_in_2_bits_entry_perm_d(Arbiter_1_io_in_2_bits_entry_perm_d),
    .io_in_2_bits_entry_perm_a(Arbiter_1_io_in_2_bits_entry_perm_a),
    .io_in_2_bits_entry_perm_g(Arbiter_1_io_in_2_bits_entry_perm_g),
    .io_in_2_bits_entry_perm_u(Arbiter_1_io_in_2_bits_entry_perm_u),
    .io_in_2_bits_entry_perm_x(Arbiter_1_io_in_2_bits_entry_perm_x),
    .io_in_2_bits_entry_perm_w(Arbiter_1_io_in_2_bits_entry_perm_w),
    .io_in_2_bits_entry_perm_r(Arbiter_1_io_in_2_bits_entry_perm_r),
    .io_in_2_bits_pf(Arbiter_1_io_in_2_bits_pf),
    .io_in_2_bits_af(Arbiter_1_io_in_2_bits_af),
    .io_out_ready(Arbiter_1_io_out_ready),
    .io_out_valid(Arbiter_1_io_out_valid),
    .io_out_bits_entry_tag(Arbiter_1_io_out_bits_entry_tag),
    .io_out_bits_entry_asid(Arbiter_1_io_out_bits_entry_asid),
    .io_out_bits_entry_ppn(Arbiter_1_io_out_bits_entry_ppn),
    .io_out_bits_entry_perm_d(Arbiter_1_io_out_bits_entry_perm_d),
    .io_out_bits_entry_perm_a(Arbiter_1_io_out_bits_entry_perm_a),
    .io_out_bits_entry_perm_g(Arbiter_1_io_out_bits_entry_perm_g),
    .io_out_bits_entry_perm_u(Arbiter_1_io_out_bits_entry_perm_u),
    .io_out_bits_entry_perm_x(Arbiter_1_io_out_bits_entry_perm_x),
    .io_out_bits_entry_perm_w(Arbiter_1_io_out_bits_entry_perm_w),
    .io_out_bits_entry_perm_r(Arbiter_1_io_out_bits_entry_perm_r),
    .io_out_bits_entry_level(Arbiter_1_io_out_bits_entry_level),
    .io_out_bits_pf(Arbiter_1_io_out_bits_pf),
    .io_out_bits_af(Arbiter_1_io_out_bits_af)
  );
  L2TlbPrefetch prefetch ( // @[L2TLB.scala 127:26]
    .clock(prefetch_clock),
    .reset(prefetch_reset),
    .io_sfence_valid(prefetch_io_sfence_valid),
    .io_csr_satp_changed(prefetch_io_csr_satp_changed),
    .io_in_valid(prefetch_io_in_valid),
    .io_in_bits_vpn(prefetch_io_in_bits_vpn),
    .io_out_ready(prefetch_io_out_ready),
    .io_out_valid(prefetch_io_out_valid),
    .io_out_bits_vpn(prefetch_io_out_bits_vpn)
  );
  L2TlbPrefetch_hart0Writer #(.site("L2TlbPrefetch")) writer ( // @[ChiselDB.scala 132:24]
    .clock(writer_clock),
    .reset(writer_reset),
    .en(writer_en),
    .stamp(writer_stamp),
    .data_vpn(writer_data_vpn)
  );
  Arbiter_12 mq_arb ( // @[L2TLB.scala 146:22]
    .io_in_0_ready(mq_arb_io_in_0_ready),
    .io_in_0_valid(mq_arb_io_in_0_valid),
    .io_in_0_bits_vpn(mq_arb_io_in_0_bits_vpn),
    .io_in_0_bits_source(mq_arb_io_in_0_bits_source),
    .io_in_1_ready(mq_arb_io_in_1_ready),
    .io_in_1_valid(mq_arb_io_in_1_valid),
    .io_in_1_bits_vpn(mq_arb_io_in_1_bits_vpn),
    .io_in_1_bits_source(mq_arb_io_in_1_bits_source),
    .io_out_ready(mq_arb_io_out_ready),
    .io_out_valid(mq_arb_io_out_valid),
    .io_out_bits_vpn(mq_arb_io_out_bits_vpn),
    .io_out_bits_source(mq_arb_io_out_bits_source)
  );
  Arbiter_13 mem_arb ( // @[L2TLB.scala 215:23]
    .io_in_0_valid(mem_arb_io_in_0_valid),
    .io_in_0_bits_addr(mem_arb_io_in_0_bits_addr),
    .io_in_1_ready(mem_arb_io_in_1_ready),
    .io_in_1_valid(mem_arb_io_in_1_valid),
    .io_in_1_bits_addr(mem_arb_io_in_1_bits_addr),
    .io_in_1_bits_id(mem_arb_io_in_1_bits_id),
    .io_out_ready(mem_arb_io_out_ready),
    .io_out_valid(mem_arb_io_out_valid),
    .io_out_bits_addr(mem_arb_io_out_bits_addr),
    .io_out_bits_id(mem_arb_io_out_bits_id)
  );
  L1Tlb_hart0Writer #(.site("ITlbReq")) writer_1 ( // @[ChiselDB.scala 132:24]
    .clock(writer_1_clock),
    .reset(writer_1_reset),
    .en(writer_1_en),
    .stamp(writer_1_stamp),
    .data_vpn(writer_1_data_vpn)
  );
  L1Tlb_hart0Writer #(.site("DTlbReq")) writer_2 ( // @[ChiselDB.scala 132:24]
    .clock(writer_2_clock),
    .reset(writer_2_reset),
    .en(writer_2_en),
    .stamp(writer_2_stamp),
    .data_vpn(writer_2_data_vpn)
  );
  L1Tlb_hart0Writer #(.site("ITlbResp")) writer_3 ( // @[ChiselDB.scala 132:24]
    .clock(writer_3_clock),
    .reset(writer_3_reset),
    .en(writer_3_en),
    .stamp(writer_3_stamp),
    .data_vpn(writer_3_data_vpn)
  );
  L1Tlb_hart0Writer #(.site("DTlbResp")) writer_4 ( // @[ChiselDB.scala 132:24]
    .clock(writer_4_clock),
    .reset(writer_4_reset),
    .en(writer_4_en),
    .stamp(writer_4_stamp),
    .data_vpn(writer_4_data_vpn)
  );
  PageCache_hart0Writer #(.site("PageCache")) writer_5 ( // @[ChiselDB.scala 132:24]
    .clock(writer_5_clock),
    .reset(writer_5_reset),
    .en(writer_5_en),
    .stamp(writer_5_stamp),
    .data_vpn(writer_5_data_vpn),
    .data_source(writer_5_data_source),
    .data_bypassed(writer_5_data_bypassed),
    .data_is_first(writer_5_data_is_first),
    .data_prefetched(writer_5_data_prefetched),
    .data_prefetch(writer_5_data_prefetch),
    .data_l2Hit(writer_5_data_l2Hit),
    .data_l1Hit(writer_5_data_l1Hit),
    .data_hit(writer_5_data_hit)
  );
  PTW_hart0Writer #(.site("PTWReq")) writer_6 ( // @[ChiselDB.scala 132:24]
    .clock(writer_6_clock),
    .reset(writer_6_reset),
    .en(writer_6_en),
    .stamp(writer_6_stamp),
    .data_vpn(writer_6_data_vpn),
    .data_source(writer_6_data_source)
  );
  PTW_hart0Writer #(.site("PTWResp")) writer_7 ( // @[ChiselDB.scala 132:24]
    .clock(writer_7_clock),
    .reset(writer_7_reset),
    .en(writer_7_en),
    .stamp(writer_7_stamp),
    .data_vpn(writer_7_data_vpn),
    .data_source(writer_7_data_source)
  );
  PTW_hart0Writer #(.site("LLPTWReq")) writer_8 ( // @[ChiselDB.scala 132:24]
    .clock(writer_8_clock),
    .reset(writer_8_reset),
    .en(writer_8_en),
    .stamp(writer_8_stamp),
    .data_vpn(writer_8_data_vpn),
    .data_source(writer_8_data_source)
  );
  PTW_hart0Writer #(.site("LLPTWResp")) writer_9 ( // @[ChiselDB.scala 132:24]
    .clock(writer_9_clock),
    .reset(writer_9_reset),
    .en(writer_9_en),
    .stamp(writer_9_stamp),
    .data_vpn(writer_9_data_vpn),
    .data_source(writer_9_data_source)
  );
  L2TlbMissQueue_hart0Writer #(.site("L2TlbMissQueueIn")) writer_10 ( // @[ChiselDB.scala 132:24]
    .clock(writer_10_clock),
    .reset(writer_10_reset),
    .en(writer_10_en),
    .stamp(writer_10_stamp),
    .data_vpn(writer_10_data_vpn)
  );
  L2TlbMissQueue_hart0Writer #(.site("L2TlbMissQueueOut")) writer_11 ( // @[ChiselDB.scala 132:24]
    .clock(writer_11_clock),
    .reset(writer_11_reset),
    .en(writer_11_en),
    .stamp(writer_11_stamp),
    .data_vpn(writer_11_data_vpn)
  );
  assign auto_out_a_valid = mem_arb_io_out_valid & _mem_arb_io_out_ready_T; // @[L2TLB.scala 253:39]
  assign auto_out_a_bits_source = mem_arb_io_out_bits_id; // @[Edges.scala 447:17 451:15]
  assign auto_out_a_bits_address = {mem_arb_io_out_bits_addr[35:6],6'h0}; // @[Cat.scala 31:58]
  assign io_tlb_0_req_0_ready = arb1_io_in_0_ready; // @[L2TLB.scala 114:{14,24}]
  assign io_tlb_0_resp_valid = Arbiter_io_out_valid; // @[L2TLB.scala 346:30]
  assign io_tlb_0_resp_bits_entry_tag = Arbiter_io_out_bits_entry_tag; // @[L2TLB.scala 346:30]
  assign io_tlb_0_resp_bits_entry_asid = Arbiter_io_out_bits_entry_asid; // @[L2TLB.scala 346:30]
  assign io_tlb_0_resp_bits_entry_ppn = Arbiter_io_out_bits_entry_ppn; // @[L2TLB.scala 346:30]
  assign io_tlb_0_resp_bits_entry_perm_d = Arbiter_io_out_bits_entry_perm_d; // @[L2TLB.scala 346:30]
  assign io_tlb_0_resp_bits_entry_perm_a = Arbiter_io_out_bits_entry_perm_a; // @[L2TLB.scala 346:30]
  assign io_tlb_0_resp_bits_entry_perm_g = Arbiter_io_out_bits_entry_perm_g; // @[L2TLB.scala 346:30]
  assign io_tlb_0_resp_bits_entry_perm_u = Arbiter_io_out_bits_entry_perm_u; // @[L2TLB.scala 346:30]
  assign io_tlb_0_resp_bits_entry_perm_x = Arbiter_io_out_bits_entry_perm_x; // @[L2TLB.scala 346:30]
  assign io_tlb_0_resp_bits_entry_perm_w = Arbiter_io_out_bits_entry_perm_w; // @[L2TLB.scala 346:30]
  assign io_tlb_0_resp_bits_entry_perm_r = Arbiter_io_out_bits_entry_perm_r; // @[L2TLB.scala 346:30]
  assign io_tlb_0_resp_bits_entry_level = Arbiter_io_out_bits_entry_level; // @[L2TLB.scala 346:30]
  assign io_tlb_0_resp_bits_pf = Arbiter_io_out_bits_pf; // @[L2TLB.scala 346:30]
  assign io_tlb_0_resp_bits_af = Arbiter_io_out_bits_af; // @[L2TLB.scala 346:30]
  assign io_tlb_1_req_0_ready = arb1_io_in_1_ready; // @[L2TLB.scala 114:{14,24}]
  assign io_tlb_1_resp_valid = Arbiter_1_io_out_valid; // @[L2TLB.scala 346:30]
  assign io_tlb_1_resp_bits_entry_tag = Arbiter_1_io_out_bits_entry_tag; // @[L2TLB.scala 346:30]
  assign io_tlb_1_resp_bits_entry_asid = Arbiter_1_io_out_bits_entry_asid; // @[L2TLB.scala 346:30]
  assign io_tlb_1_resp_bits_entry_ppn = Arbiter_1_io_out_bits_entry_ppn; // @[L2TLB.scala 346:30]
  assign io_tlb_1_resp_bits_entry_perm_d = Arbiter_1_io_out_bits_entry_perm_d; // @[L2TLB.scala 346:30]
  assign io_tlb_1_resp_bits_entry_perm_a = Arbiter_1_io_out_bits_entry_perm_a; // @[L2TLB.scala 346:30]
  assign io_tlb_1_resp_bits_entry_perm_g = Arbiter_1_io_out_bits_entry_perm_g; // @[L2TLB.scala 346:30]
  assign io_tlb_1_resp_bits_entry_perm_u = Arbiter_1_io_out_bits_entry_perm_u; // @[L2TLB.scala 346:30]
  assign io_tlb_1_resp_bits_entry_perm_x = Arbiter_1_io_out_bits_entry_perm_x; // @[L2TLB.scala 346:30]
  assign io_tlb_1_resp_bits_entry_perm_w = Arbiter_1_io_out_bits_entry_perm_w; // @[L2TLB.scala 346:30]
  assign io_tlb_1_resp_bits_entry_perm_r = Arbiter_1_io_out_bits_entry_perm_r; // @[L2TLB.scala 346:30]
  assign io_tlb_1_resp_bits_entry_level = Arbiter_1_io_out_bits_entry_level; // @[L2TLB.scala 346:30]
  assign io_tlb_1_resp_bits_pf = Arbiter_1_io_out_bits_pf; // @[L2TLB.scala 346:30]
  assign io_tlb_1_resp_bits_af = Arbiter_1_io_out_bits_af; // @[L2TLB.scala 346:30]
  assign io_perf_0_value = io_perf_0_value_REG_1; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_1_value = io_perf_1_value_REG_1; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_2_value = io_perf_2_value_REG_1; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_3_value = io_perf_3_value_REG_1; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_4_value = io_perf_4_value_REG_1; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_5_value = io_perf_5_value_REG_1; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_6_value = io_perf_6_value_REG_1; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_7_value = io_perf_7_value_REG_1; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_8_value = io_perf_8_value_REG_1; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_9_value = io_perf_9_value_REG_1; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_10_value = io_perf_10_value_REG_1; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_11_value = io_perf_11_value_REG_1; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_12_value = io_perf_12_value_REG_1; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_13_value = io_perf_13_value_REG_1; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_14_value = io_perf_14_value_REG_1; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_15_value = io_perf_15_value_REG_1; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_16_value = io_perf_16_value_REG_1; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_17_value = io_perf_17_value_REG_1; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_18_value = io_perf_18_value_REG_1; // @[PerfCounterUtils.scala 188:17]
  assign sfence_tmp_delay_clock = clock;
  assign sfence_tmp_delay_io_in_valid = io_sfence_valid; // @[Hold.scala 98:17]
  assign sfence_tmp_delay_io_in_bits_rs1 = io_sfence_bits_rs1; // @[Hold.scala 98:17]
  assign sfence_tmp_delay_io_in_bits_rs2 = io_sfence_bits_rs2; // @[Hold.scala 98:17]
  assign sfence_tmp_delay_io_in_bits_addr = io_sfence_bits_addr; // @[Hold.scala 98:17]
  assign sfence_tmp_delay_io_in_bits_asid = io_sfence_bits_asid; // @[Hold.scala 98:17]
  assign csr_tmp_delay_clock = clock;
  assign csr_tmp_delay_io_in_satp_asid = io_csr_tlb_satp_asid; // @[Hold.scala 98:17]
  assign csr_tmp_delay_io_in_satp_ppn = io_csr_tlb_satp_ppn; // @[Hold.scala 98:17]
  assign csr_tmp_delay_io_in_satp_changed = io_csr_tlb_satp_changed; // @[Hold.scala 98:17]
  assign pmp_clock = clock;
  assign pmp_reset = reset;
  assign pmp_io_distribute_csr_wvalid = io_csr_distribute_csr_wvalid; // @[L2TLB.scala 90:25]
  assign pmp_io_distribute_csr_waddr = io_csr_distribute_csr_waddr; // @[L2TLB.scala 90:25]
  assign pmp_io_distribute_csr_wdata = io_csr_distribute_csr_wdata; // @[L2TLB.scala 90:25]
  assign PMPChecker_io_check_env_mode = 2'h1; // @[L2TLB.scala 89:26 PMP.scala 465:15]
  assign PMPChecker_io_check_env_pmp_0_cfg_l = pmp_io_pmp_0_cfg_l; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_0_cfg_a = pmp_io_pmp_0_cfg_a; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_0_cfg_x = pmp_io_pmp_0_cfg_x; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_0_cfg_w = pmp_io_pmp_0_cfg_w; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_0_cfg_r = pmp_io_pmp_0_cfg_r; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_0_addr = pmp_io_pmp_0_addr; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_0_mask = pmp_io_pmp_0_mask; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_1_cfg_l = pmp_io_pmp_1_cfg_l; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_1_cfg_a = pmp_io_pmp_1_cfg_a; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_1_cfg_x = pmp_io_pmp_1_cfg_x; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_1_cfg_w = pmp_io_pmp_1_cfg_w; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_1_cfg_r = pmp_io_pmp_1_cfg_r; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_1_addr = pmp_io_pmp_1_addr; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_1_mask = pmp_io_pmp_1_mask; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_2_cfg_l = pmp_io_pmp_2_cfg_l; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_2_cfg_a = pmp_io_pmp_2_cfg_a; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_2_cfg_x = pmp_io_pmp_2_cfg_x; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_2_cfg_w = pmp_io_pmp_2_cfg_w; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_2_cfg_r = pmp_io_pmp_2_cfg_r; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_2_addr = pmp_io_pmp_2_addr; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_2_mask = pmp_io_pmp_2_mask; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_3_cfg_l = pmp_io_pmp_3_cfg_l; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_3_cfg_a = pmp_io_pmp_3_cfg_a; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_3_cfg_x = pmp_io_pmp_3_cfg_x; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_3_cfg_w = pmp_io_pmp_3_cfg_w; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_3_cfg_r = pmp_io_pmp_3_cfg_r; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_3_addr = pmp_io_pmp_3_addr; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_3_mask = pmp_io_pmp_3_mask; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_4_cfg_l = pmp_io_pmp_4_cfg_l; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_4_cfg_a = pmp_io_pmp_4_cfg_a; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_4_cfg_x = pmp_io_pmp_4_cfg_x; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_4_cfg_w = pmp_io_pmp_4_cfg_w; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_4_cfg_r = pmp_io_pmp_4_cfg_r; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_4_addr = pmp_io_pmp_4_addr; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_4_mask = pmp_io_pmp_4_mask; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_5_cfg_l = pmp_io_pmp_5_cfg_l; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_5_cfg_a = pmp_io_pmp_5_cfg_a; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_5_cfg_x = pmp_io_pmp_5_cfg_x; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_5_cfg_w = pmp_io_pmp_5_cfg_w; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_5_cfg_r = pmp_io_pmp_5_cfg_r; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_5_addr = pmp_io_pmp_5_addr; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_5_mask = pmp_io_pmp_5_mask; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_6_cfg_l = pmp_io_pmp_6_cfg_l; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_6_cfg_a = pmp_io_pmp_6_cfg_a; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_6_cfg_x = pmp_io_pmp_6_cfg_x; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_6_cfg_w = pmp_io_pmp_6_cfg_w; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_6_cfg_r = pmp_io_pmp_6_cfg_r; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_6_addr = pmp_io_pmp_6_addr; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_6_mask = pmp_io_pmp_6_mask; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_7_cfg_l = pmp_io_pmp_7_cfg_l; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_7_cfg_a = pmp_io_pmp_7_cfg_a; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_7_cfg_x = pmp_io_pmp_7_cfg_x; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_7_cfg_w = pmp_io_pmp_7_cfg_w; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_7_cfg_r = pmp_io_pmp_7_cfg_r; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_7_addr = pmp_io_pmp_7_addr; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_7_mask = pmp_io_pmp_7_mask; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_8_cfg_l = pmp_io_pmp_8_cfg_l; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_8_cfg_a = pmp_io_pmp_8_cfg_a; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_8_cfg_x = pmp_io_pmp_8_cfg_x; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_8_cfg_w = pmp_io_pmp_8_cfg_w; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_8_cfg_r = pmp_io_pmp_8_cfg_r; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_8_addr = pmp_io_pmp_8_addr; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_8_mask = pmp_io_pmp_8_mask; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_9_cfg_l = pmp_io_pmp_9_cfg_l; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_9_cfg_a = pmp_io_pmp_9_cfg_a; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_9_cfg_x = pmp_io_pmp_9_cfg_x; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_9_cfg_w = pmp_io_pmp_9_cfg_w; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_9_cfg_r = pmp_io_pmp_9_cfg_r; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_9_addr = pmp_io_pmp_9_addr; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_9_mask = pmp_io_pmp_9_mask; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_10_cfg_l = pmp_io_pmp_10_cfg_l; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_10_cfg_a = pmp_io_pmp_10_cfg_a; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_10_cfg_x = pmp_io_pmp_10_cfg_x; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_10_cfg_w = pmp_io_pmp_10_cfg_w; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_10_cfg_r = pmp_io_pmp_10_cfg_r; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_10_addr = pmp_io_pmp_10_addr; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_10_mask = pmp_io_pmp_10_mask; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_11_cfg_l = pmp_io_pmp_11_cfg_l; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_11_cfg_a = pmp_io_pmp_11_cfg_a; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_11_cfg_x = pmp_io_pmp_11_cfg_x; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_11_cfg_w = pmp_io_pmp_11_cfg_w; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_11_cfg_r = pmp_io_pmp_11_cfg_r; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_11_addr = pmp_io_pmp_11_addr; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_11_mask = pmp_io_pmp_11_mask; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_12_cfg_l = pmp_io_pmp_12_cfg_l; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_12_cfg_a = pmp_io_pmp_12_cfg_a; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_12_cfg_x = pmp_io_pmp_12_cfg_x; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_12_cfg_w = pmp_io_pmp_12_cfg_w; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_12_cfg_r = pmp_io_pmp_12_cfg_r; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_12_addr = pmp_io_pmp_12_addr; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_12_mask = pmp_io_pmp_12_mask; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_13_cfg_l = pmp_io_pmp_13_cfg_l; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_13_cfg_a = pmp_io_pmp_13_cfg_a; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_13_cfg_x = pmp_io_pmp_13_cfg_x; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_13_cfg_w = pmp_io_pmp_13_cfg_w; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_13_cfg_r = pmp_io_pmp_13_cfg_r; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_13_addr = pmp_io_pmp_13_addr; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_13_mask = pmp_io_pmp_13_mask; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_14_cfg_l = pmp_io_pmp_14_cfg_l; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_14_cfg_a = pmp_io_pmp_14_cfg_a; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_14_cfg_x = pmp_io_pmp_14_cfg_x; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_14_cfg_w = pmp_io_pmp_14_cfg_w; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_14_cfg_r = pmp_io_pmp_14_cfg_r; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_14_addr = pmp_io_pmp_14_addr; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_14_mask = pmp_io_pmp_14_mask; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_15_cfg_l = pmp_io_pmp_15_cfg_l; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_15_cfg_a = pmp_io_pmp_15_cfg_a; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_15_cfg_x = pmp_io_pmp_15_cfg_x; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_15_cfg_w = pmp_io_pmp_15_cfg_w; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_15_cfg_r = pmp_io_pmp_15_cfg_r; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_15_addr = pmp_io_pmp_15_addr; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_15_mask = pmp_io_pmp_15_mask; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pma_0_cfg_c = pmp_io_pma_0_cfg_c; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_0_cfg_atomic = pmp_io_pma_0_cfg_atomic; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_0_cfg_a = pmp_io_pma_0_cfg_a; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_0_cfg_x = pmp_io_pma_0_cfg_x; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_0_cfg_w = pmp_io_pma_0_cfg_w; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_0_cfg_r = pmp_io_pma_0_cfg_r; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_0_addr = pmp_io_pma_0_addr; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_0_mask = pmp_io_pma_0_mask; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_1_cfg_c = pmp_io_pma_1_cfg_c; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_1_cfg_atomic = pmp_io_pma_1_cfg_atomic; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_1_cfg_a = pmp_io_pma_1_cfg_a; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_1_cfg_x = pmp_io_pma_1_cfg_x; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_1_cfg_w = pmp_io_pma_1_cfg_w; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_1_cfg_r = pmp_io_pma_1_cfg_r; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_1_addr = pmp_io_pma_1_addr; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_1_mask = pmp_io_pma_1_mask; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_2_cfg_c = pmp_io_pma_2_cfg_c; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_2_cfg_atomic = pmp_io_pma_2_cfg_atomic; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_2_cfg_a = pmp_io_pma_2_cfg_a; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_2_cfg_x = pmp_io_pma_2_cfg_x; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_2_cfg_w = pmp_io_pma_2_cfg_w; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_2_cfg_r = pmp_io_pma_2_cfg_r; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_2_addr = pmp_io_pma_2_addr; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_2_mask = pmp_io_pma_2_mask; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_3_cfg_c = pmp_io_pma_3_cfg_c; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_3_cfg_atomic = pmp_io_pma_3_cfg_atomic; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_3_cfg_a = pmp_io_pma_3_cfg_a; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_3_cfg_x = pmp_io_pma_3_cfg_x; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_3_cfg_w = pmp_io_pma_3_cfg_w; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_3_cfg_r = pmp_io_pma_3_cfg_r; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_3_addr = pmp_io_pma_3_addr; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_3_mask = pmp_io_pma_3_mask; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_4_cfg_c = pmp_io_pma_4_cfg_c; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_4_cfg_atomic = pmp_io_pma_4_cfg_atomic; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_4_cfg_a = pmp_io_pma_4_cfg_a; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_4_cfg_x = pmp_io_pma_4_cfg_x; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_4_cfg_w = pmp_io_pma_4_cfg_w; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_4_cfg_r = pmp_io_pma_4_cfg_r; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_4_addr = pmp_io_pma_4_addr; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_4_mask = pmp_io_pma_4_mask; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_5_cfg_c = pmp_io_pma_5_cfg_c; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_5_cfg_atomic = pmp_io_pma_5_cfg_atomic; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_5_cfg_a = pmp_io_pma_5_cfg_a; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_5_cfg_x = pmp_io_pma_5_cfg_x; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_5_cfg_w = pmp_io_pma_5_cfg_w; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_5_cfg_r = pmp_io_pma_5_cfg_r; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_5_addr = pmp_io_pma_5_addr; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_5_mask = pmp_io_pma_5_mask; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_6_cfg_c = pmp_io_pma_6_cfg_c; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_6_cfg_atomic = pmp_io_pma_6_cfg_atomic; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_6_cfg_a = pmp_io_pma_6_cfg_a; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_6_cfg_x = pmp_io_pma_6_cfg_x; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_6_cfg_w = pmp_io_pma_6_cfg_w; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_6_cfg_r = pmp_io_pma_6_cfg_r; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_6_addr = pmp_io_pma_6_addr; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_6_mask = pmp_io_pma_6_mask; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_7_cfg_c = pmp_io_pma_7_cfg_c; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_7_cfg_atomic = pmp_io_pma_7_cfg_atomic; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_7_cfg_a = pmp_io_pma_7_cfg_a; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_7_cfg_x = pmp_io_pma_7_cfg_x; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_7_cfg_w = pmp_io_pma_7_cfg_w; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_7_cfg_r = pmp_io_pma_7_cfg_r; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_7_addr = pmp_io_pma_7_addr; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_7_mask = pmp_io_pma_7_mask; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_8_cfg_c = pmp_io_pma_8_cfg_c; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_8_cfg_atomic = pmp_io_pma_8_cfg_atomic; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_8_cfg_a = pmp_io_pma_8_cfg_a; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_8_cfg_x = pmp_io_pma_8_cfg_x; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_8_cfg_w = pmp_io_pma_8_cfg_w; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_8_cfg_r = pmp_io_pma_8_cfg_r; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_8_addr = pmp_io_pma_8_addr; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_8_mask = pmp_io_pma_8_mask; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_9_cfg_c = pmp_io_pma_9_cfg_c; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_9_cfg_atomic = pmp_io_pma_9_cfg_atomic; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_9_cfg_a = pmp_io_pma_9_cfg_a; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_9_cfg_x = pmp_io_pma_9_cfg_x; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_9_cfg_w = pmp_io_pma_9_cfg_w; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_9_cfg_r = pmp_io_pma_9_cfg_r; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_9_addr = pmp_io_pma_9_addr; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_9_mask = pmp_io_pma_9_mask; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_10_cfg_c = pmp_io_pma_10_cfg_c; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_10_cfg_atomic = pmp_io_pma_10_cfg_atomic; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_10_cfg_a = pmp_io_pma_10_cfg_a; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_10_cfg_x = pmp_io_pma_10_cfg_x; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_10_cfg_w = pmp_io_pma_10_cfg_w; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_10_cfg_r = pmp_io_pma_10_cfg_r; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_10_addr = pmp_io_pma_10_addr; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_10_mask = pmp_io_pma_10_mask; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_11_cfg_c = pmp_io_pma_11_cfg_c; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_11_cfg_atomic = pmp_io_pma_11_cfg_atomic; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_11_cfg_a = pmp_io_pma_11_cfg_a; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_11_cfg_x = pmp_io_pma_11_cfg_x; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_11_cfg_w = pmp_io_pma_11_cfg_w; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_11_cfg_r = pmp_io_pma_11_cfg_r; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_11_addr = pmp_io_pma_11_addr; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_11_mask = pmp_io_pma_11_mask; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_12_cfg_c = pmp_io_pma_12_cfg_c; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_12_cfg_atomic = pmp_io_pma_12_cfg_atomic; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_12_cfg_a = pmp_io_pma_12_cfg_a; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_12_cfg_x = pmp_io_pma_12_cfg_x; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_12_cfg_w = pmp_io_pma_12_cfg_w; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_12_cfg_r = pmp_io_pma_12_cfg_r; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_12_addr = pmp_io_pma_12_addr; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_12_mask = pmp_io_pma_12_mask; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_13_cfg_c = pmp_io_pma_13_cfg_c; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_13_cfg_atomic = pmp_io_pma_13_cfg_atomic; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_13_cfg_a = pmp_io_pma_13_cfg_a; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_13_cfg_x = pmp_io_pma_13_cfg_x; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_13_cfg_w = pmp_io_pma_13_cfg_w; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_13_cfg_r = pmp_io_pma_13_cfg_r; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_13_addr = pmp_io_pma_13_addr; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_13_mask = pmp_io_pma_13_mask; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_14_cfg_c = pmp_io_pma_14_cfg_c; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_14_cfg_atomic = pmp_io_pma_14_cfg_atomic; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_14_cfg_a = pmp_io_pma_14_cfg_a; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_14_cfg_x = pmp_io_pma_14_cfg_x; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_14_cfg_w = pmp_io_pma_14_cfg_w; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_14_cfg_r = pmp_io_pma_14_cfg_r; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_14_addr = pmp_io_pma_14_addr; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_14_mask = pmp_io_pma_14_mask; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_15_cfg_c = pmp_io_pma_15_cfg_c; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_15_cfg_atomic = pmp_io_pma_15_cfg_atomic; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_15_cfg_a = pmp_io_pma_15_cfg_a; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_15_cfg_x = pmp_io_pma_15_cfg_x; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_15_cfg_w = pmp_io_pma_15_cfg_w; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_15_cfg_r = pmp_io_pma_15_cfg_r; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_15_addr = pmp_io_pma_15_addr; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_15_mask = pmp_io_pma_15_mask; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_io_req_bits_addr = ptw_io_pmp_req_bits_addr; // @[L2TLB.scala 327:20 89:26]
  assign PMPChecker_io_req_bits_cmd = 3'h0; // @[L2TLB.scala 327:20 89:26]
  assign PMPChecker_1_io_check_env_mode = 2'h1; // @[L2TLB.scala 89:26 PMP.scala 465:15]
  assign PMPChecker_1_io_check_env_pmp_0_cfg_l = pmp_io_pmp_0_cfg_l; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_0_cfg_a = pmp_io_pmp_0_cfg_a; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_0_cfg_x = pmp_io_pmp_0_cfg_x; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_0_cfg_w = pmp_io_pmp_0_cfg_w; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_0_cfg_r = pmp_io_pmp_0_cfg_r; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_0_addr = pmp_io_pmp_0_addr; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_0_mask = pmp_io_pmp_0_mask; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_1_cfg_l = pmp_io_pmp_1_cfg_l; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_1_cfg_a = pmp_io_pmp_1_cfg_a; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_1_cfg_x = pmp_io_pmp_1_cfg_x; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_1_cfg_w = pmp_io_pmp_1_cfg_w; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_1_cfg_r = pmp_io_pmp_1_cfg_r; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_1_addr = pmp_io_pmp_1_addr; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_1_mask = pmp_io_pmp_1_mask; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_2_cfg_l = pmp_io_pmp_2_cfg_l; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_2_cfg_a = pmp_io_pmp_2_cfg_a; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_2_cfg_x = pmp_io_pmp_2_cfg_x; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_2_cfg_w = pmp_io_pmp_2_cfg_w; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_2_cfg_r = pmp_io_pmp_2_cfg_r; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_2_addr = pmp_io_pmp_2_addr; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_2_mask = pmp_io_pmp_2_mask; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_3_cfg_l = pmp_io_pmp_3_cfg_l; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_3_cfg_a = pmp_io_pmp_3_cfg_a; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_3_cfg_x = pmp_io_pmp_3_cfg_x; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_3_cfg_w = pmp_io_pmp_3_cfg_w; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_3_cfg_r = pmp_io_pmp_3_cfg_r; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_3_addr = pmp_io_pmp_3_addr; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_3_mask = pmp_io_pmp_3_mask; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_4_cfg_l = pmp_io_pmp_4_cfg_l; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_4_cfg_a = pmp_io_pmp_4_cfg_a; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_4_cfg_x = pmp_io_pmp_4_cfg_x; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_4_cfg_w = pmp_io_pmp_4_cfg_w; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_4_cfg_r = pmp_io_pmp_4_cfg_r; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_4_addr = pmp_io_pmp_4_addr; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_4_mask = pmp_io_pmp_4_mask; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_5_cfg_l = pmp_io_pmp_5_cfg_l; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_5_cfg_a = pmp_io_pmp_5_cfg_a; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_5_cfg_x = pmp_io_pmp_5_cfg_x; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_5_cfg_w = pmp_io_pmp_5_cfg_w; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_5_cfg_r = pmp_io_pmp_5_cfg_r; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_5_addr = pmp_io_pmp_5_addr; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_5_mask = pmp_io_pmp_5_mask; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_6_cfg_l = pmp_io_pmp_6_cfg_l; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_6_cfg_a = pmp_io_pmp_6_cfg_a; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_6_cfg_x = pmp_io_pmp_6_cfg_x; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_6_cfg_w = pmp_io_pmp_6_cfg_w; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_6_cfg_r = pmp_io_pmp_6_cfg_r; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_6_addr = pmp_io_pmp_6_addr; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_6_mask = pmp_io_pmp_6_mask; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_7_cfg_l = pmp_io_pmp_7_cfg_l; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_7_cfg_a = pmp_io_pmp_7_cfg_a; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_7_cfg_x = pmp_io_pmp_7_cfg_x; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_7_cfg_w = pmp_io_pmp_7_cfg_w; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_7_cfg_r = pmp_io_pmp_7_cfg_r; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_7_addr = pmp_io_pmp_7_addr; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_7_mask = pmp_io_pmp_7_mask; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_8_cfg_l = pmp_io_pmp_8_cfg_l; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_8_cfg_a = pmp_io_pmp_8_cfg_a; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_8_cfg_x = pmp_io_pmp_8_cfg_x; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_8_cfg_w = pmp_io_pmp_8_cfg_w; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_8_cfg_r = pmp_io_pmp_8_cfg_r; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_8_addr = pmp_io_pmp_8_addr; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_8_mask = pmp_io_pmp_8_mask; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_9_cfg_l = pmp_io_pmp_9_cfg_l; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_9_cfg_a = pmp_io_pmp_9_cfg_a; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_9_cfg_x = pmp_io_pmp_9_cfg_x; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_9_cfg_w = pmp_io_pmp_9_cfg_w; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_9_cfg_r = pmp_io_pmp_9_cfg_r; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_9_addr = pmp_io_pmp_9_addr; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_9_mask = pmp_io_pmp_9_mask; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_10_cfg_l = pmp_io_pmp_10_cfg_l; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_10_cfg_a = pmp_io_pmp_10_cfg_a; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_10_cfg_x = pmp_io_pmp_10_cfg_x; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_10_cfg_w = pmp_io_pmp_10_cfg_w; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_10_cfg_r = pmp_io_pmp_10_cfg_r; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_10_addr = pmp_io_pmp_10_addr; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_10_mask = pmp_io_pmp_10_mask; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_11_cfg_l = pmp_io_pmp_11_cfg_l; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_11_cfg_a = pmp_io_pmp_11_cfg_a; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_11_cfg_x = pmp_io_pmp_11_cfg_x; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_11_cfg_w = pmp_io_pmp_11_cfg_w; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_11_cfg_r = pmp_io_pmp_11_cfg_r; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_11_addr = pmp_io_pmp_11_addr; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_11_mask = pmp_io_pmp_11_mask; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_12_cfg_l = pmp_io_pmp_12_cfg_l; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_12_cfg_a = pmp_io_pmp_12_cfg_a; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_12_cfg_x = pmp_io_pmp_12_cfg_x; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_12_cfg_w = pmp_io_pmp_12_cfg_w; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_12_cfg_r = pmp_io_pmp_12_cfg_r; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_12_addr = pmp_io_pmp_12_addr; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_12_mask = pmp_io_pmp_12_mask; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_13_cfg_l = pmp_io_pmp_13_cfg_l; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_13_cfg_a = pmp_io_pmp_13_cfg_a; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_13_cfg_x = pmp_io_pmp_13_cfg_x; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_13_cfg_w = pmp_io_pmp_13_cfg_w; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_13_cfg_r = pmp_io_pmp_13_cfg_r; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_13_addr = pmp_io_pmp_13_addr; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_13_mask = pmp_io_pmp_13_mask; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_14_cfg_l = pmp_io_pmp_14_cfg_l; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_14_cfg_a = pmp_io_pmp_14_cfg_a; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_14_cfg_x = pmp_io_pmp_14_cfg_x; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_14_cfg_w = pmp_io_pmp_14_cfg_w; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_14_cfg_r = pmp_io_pmp_14_cfg_r; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_14_addr = pmp_io_pmp_14_addr; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_14_mask = pmp_io_pmp_14_mask; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_15_cfg_l = pmp_io_pmp_15_cfg_l; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_15_cfg_a = pmp_io_pmp_15_cfg_a; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_15_cfg_x = pmp_io_pmp_15_cfg_x; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_15_cfg_w = pmp_io_pmp_15_cfg_w; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_15_cfg_r = pmp_io_pmp_15_cfg_r; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_15_addr = pmp_io_pmp_15_addr; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_15_mask = pmp_io_pmp_15_mask; // @[L2TLB.scala 89:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pma_0_cfg_c = pmp_io_pma_0_cfg_c; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_0_cfg_atomic = pmp_io_pma_0_cfg_atomic; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_0_cfg_a = pmp_io_pma_0_cfg_a; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_0_cfg_x = pmp_io_pma_0_cfg_x; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_0_cfg_w = pmp_io_pma_0_cfg_w; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_0_cfg_r = pmp_io_pma_0_cfg_r; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_0_addr = pmp_io_pma_0_addr; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_0_mask = pmp_io_pma_0_mask; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_1_cfg_c = pmp_io_pma_1_cfg_c; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_1_cfg_atomic = pmp_io_pma_1_cfg_atomic; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_1_cfg_a = pmp_io_pma_1_cfg_a; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_1_cfg_x = pmp_io_pma_1_cfg_x; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_1_cfg_w = pmp_io_pma_1_cfg_w; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_1_cfg_r = pmp_io_pma_1_cfg_r; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_1_addr = pmp_io_pma_1_addr; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_1_mask = pmp_io_pma_1_mask; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_2_cfg_c = pmp_io_pma_2_cfg_c; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_2_cfg_atomic = pmp_io_pma_2_cfg_atomic; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_2_cfg_a = pmp_io_pma_2_cfg_a; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_2_cfg_x = pmp_io_pma_2_cfg_x; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_2_cfg_w = pmp_io_pma_2_cfg_w; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_2_cfg_r = pmp_io_pma_2_cfg_r; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_2_addr = pmp_io_pma_2_addr; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_2_mask = pmp_io_pma_2_mask; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_3_cfg_c = pmp_io_pma_3_cfg_c; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_3_cfg_atomic = pmp_io_pma_3_cfg_atomic; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_3_cfg_a = pmp_io_pma_3_cfg_a; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_3_cfg_x = pmp_io_pma_3_cfg_x; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_3_cfg_w = pmp_io_pma_3_cfg_w; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_3_cfg_r = pmp_io_pma_3_cfg_r; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_3_addr = pmp_io_pma_3_addr; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_3_mask = pmp_io_pma_3_mask; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_4_cfg_c = pmp_io_pma_4_cfg_c; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_4_cfg_atomic = pmp_io_pma_4_cfg_atomic; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_4_cfg_a = pmp_io_pma_4_cfg_a; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_4_cfg_x = pmp_io_pma_4_cfg_x; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_4_cfg_w = pmp_io_pma_4_cfg_w; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_4_cfg_r = pmp_io_pma_4_cfg_r; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_4_addr = pmp_io_pma_4_addr; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_4_mask = pmp_io_pma_4_mask; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_5_cfg_c = pmp_io_pma_5_cfg_c; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_5_cfg_atomic = pmp_io_pma_5_cfg_atomic; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_5_cfg_a = pmp_io_pma_5_cfg_a; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_5_cfg_x = pmp_io_pma_5_cfg_x; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_5_cfg_w = pmp_io_pma_5_cfg_w; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_5_cfg_r = pmp_io_pma_5_cfg_r; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_5_addr = pmp_io_pma_5_addr; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_5_mask = pmp_io_pma_5_mask; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_6_cfg_c = pmp_io_pma_6_cfg_c; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_6_cfg_atomic = pmp_io_pma_6_cfg_atomic; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_6_cfg_a = pmp_io_pma_6_cfg_a; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_6_cfg_x = pmp_io_pma_6_cfg_x; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_6_cfg_w = pmp_io_pma_6_cfg_w; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_6_cfg_r = pmp_io_pma_6_cfg_r; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_6_addr = pmp_io_pma_6_addr; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_6_mask = pmp_io_pma_6_mask; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_7_cfg_c = pmp_io_pma_7_cfg_c; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_7_cfg_atomic = pmp_io_pma_7_cfg_atomic; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_7_cfg_a = pmp_io_pma_7_cfg_a; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_7_cfg_x = pmp_io_pma_7_cfg_x; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_7_cfg_w = pmp_io_pma_7_cfg_w; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_7_cfg_r = pmp_io_pma_7_cfg_r; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_7_addr = pmp_io_pma_7_addr; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_7_mask = pmp_io_pma_7_mask; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_8_cfg_c = pmp_io_pma_8_cfg_c; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_8_cfg_atomic = pmp_io_pma_8_cfg_atomic; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_8_cfg_a = pmp_io_pma_8_cfg_a; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_8_cfg_x = pmp_io_pma_8_cfg_x; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_8_cfg_w = pmp_io_pma_8_cfg_w; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_8_cfg_r = pmp_io_pma_8_cfg_r; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_8_addr = pmp_io_pma_8_addr; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_8_mask = pmp_io_pma_8_mask; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_9_cfg_c = pmp_io_pma_9_cfg_c; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_9_cfg_atomic = pmp_io_pma_9_cfg_atomic; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_9_cfg_a = pmp_io_pma_9_cfg_a; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_9_cfg_x = pmp_io_pma_9_cfg_x; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_9_cfg_w = pmp_io_pma_9_cfg_w; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_9_cfg_r = pmp_io_pma_9_cfg_r; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_9_addr = pmp_io_pma_9_addr; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_9_mask = pmp_io_pma_9_mask; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_10_cfg_c = pmp_io_pma_10_cfg_c; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_10_cfg_atomic = pmp_io_pma_10_cfg_atomic; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_10_cfg_a = pmp_io_pma_10_cfg_a; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_10_cfg_x = pmp_io_pma_10_cfg_x; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_10_cfg_w = pmp_io_pma_10_cfg_w; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_10_cfg_r = pmp_io_pma_10_cfg_r; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_10_addr = pmp_io_pma_10_addr; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_10_mask = pmp_io_pma_10_mask; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_11_cfg_c = pmp_io_pma_11_cfg_c; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_11_cfg_atomic = pmp_io_pma_11_cfg_atomic; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_11_cfg_a = pmp_io_pma_11_cfg_a; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_11_cfg_x = pmp_io_pma_11_cfg_x; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_11_cfg_w = pmp_io_pma_11_cfg_w; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_11_cfg_r = pmp_io_pma_11_cfg_r; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_11_addr = pmp_io_pma_11_addr; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_11_mask = pmp_io_pma_11_mask; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_12_cfg_c = pmp_io_pma_12_cfg_c; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_12_cfg_atomic = pmp_io_pma_12_cfg_atomic; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_12_cfg_a = pmp_io_pma_12_cfg_a; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_12_cfg_x = pmp_io_pma_12_cfg_x; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_12_cfg_w = pmp_io_pma_12_cfg_w; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_12_cfg_r = pmp_io_pma_12_cfg_r; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_12_addr = pmp_io_pma_12_addr; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_12_mask = pmp_io_pma_12_mask; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_13_cfg_c = pmp_io_pma_13_cfg_c; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_13_cfg_atomic = pmp_io_pma_13_cfg_atomic; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_13_cfg_a = pmp_io_pma_13_cfg_a; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_13_cfg_x = pmp_io_pma_13_cfg_x; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_13_cfg_w = pmp_io_pma_13_cfg_w; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_13_cfg_r = pmp_io_pma_13_cfg_r; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_13_addr = pmp_io_pma_13_addr; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_13_mask = pmp_io_pma_13_mask; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_14_cfg_c = pmp_io_pma_14_cfg_c; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_14_cfg_atomic = pmp_io_pma_14_cfg_atomic; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_14_cfg_a = pmp_io_pma_14_cfg_a; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_14_cfg_x = pmp_io_pma_14_cfg_x; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_14_cfg_w = pmp_io_pma_14_cfg_w; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_14_cfg_r = pmp_io_pma_14_cfg_r; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_14_addr = pmp_io_pma_14_addr; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_14_mask = pmp_io_pma_14_mask; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_15_cfg_c = pmp_io_pma_15_cfg_c; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_15_cfg_atomic = pmp_io_pma_15_cfg_atomic; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_15_cfg_a = pmp_io_pma_15_cfg_a; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_15_cfg_x = pmp_io_pma_15_cfg_x; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_15_cfg_w = pmp_io_pma_15_cfg_w; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_15_cfg_r = pmp_io_pma_15_cfg_r; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_15_addr = pmp_io_pma_15_addr; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_15_mask = pmp_io_pma_15_mask; // @[L2TLB.scala 89:26 PMP.scala 467:14]
  assign PMPChecker_1_io_req_bits_addr = llptw_io_pmp_req_bits_addr; // @[L2TLB.scala 329:20 89:26]
  assign PMPChecker_1_io_req_bits_cmd = 3'h0; // @[L2TLB.scala 329:20 89:26]
  assign missQueue_clock = clock;
  assign missQueue_reset = reset;
  assign missQueue_io_sfence_valid = sfence_dup_6_valid; // @[L2TLB.scala 154:24]
  assign missQueue_io_csr_satp_changed = csr_dup_5_satp_changed; // @[L2TLB.scala 155:20]
  assign missQueue_io_in_valid = mq_arb_io_out_valid; // @[L2TLB.scala 153:19]
  assign missQueue_io_in_bits_vpn = mq_arb_io_out_bits_vpn; // @[L2TLB.scala 153:19]
  assign missQueue_io_in_bits_source = mq_arb_io_out_bits_source; // @[L2TLB.scala 153:19]
  assign missQueue_io_out_ready = arb2_io_in_1_ready & _arb2_io_in_1_valid_T; // @[L2TLB.scala 366:34]
  assign cache_clock = clock;
  assign cache_reset = reset;
  assign cache_io_req_valid = arb2_io_out_valid; // @[L2TLB.scala 166:22]
  assign cache_io_req_bits_req_info_vpn = arb2_io_out_bits_vpn; // @[L2TLB.scala 167:34]
  assign cache_io_req_bits_req_info_source = arb2_io_out_bits_source; // @[L2TLB.scala 168:37]
  assign cache_io_req_bits_isFirst = arb2_io_chosen != 2'h1; // @[L2TLB.scala 169:47]
  assign cache_io_resp_ready = cache_io_resp_bits_hit ? _cache_io_resp_ready_T_3 : _cache_io_resp_ready_T_9; // @[L2TLB.scala 175:29]
  assign cache_io_refill_valid = cache_io_refill_valid_REG; // @[L2TLB.scala 288:25]
  assign cache_io_refill_bits_ptes = {refill_data_1,refill_data_0}; // @[L2TLB.scala 289:44]
  assign cache_io_refill_bits_levelOH_sp = cache_io_refill_bits_levelOH_sp_REG; // @[PageTableCache.scala 94:12]
  assign cache_io_refill_bits_levelOH_l3 = cache_io_refill_bits_levelOH_l3_REG; // @[PageTableCache.scala 95:12]
  assign cache_io_refill_bits_levelOH_l2 = cache_io_refill_bits_levelOH_l2_REG; // @[PageTableCache.scala 96:12]
  assign cache_io_refill_bits_levelOH_l1 = cache_io_refill_bits_levelOH_l1_REG; // @[PageTableCache.scala 97:12]
  assign cache_io_refill_bits_req_info_dup_0_vpn = cache_io_refill_bits_req_info_dup_0_rvpn; // @[L2TLB.scala 290:43]
  assign cache_io_refill_bits_req_info_dup_0_source = cache_io_refill_bits_req_info_dup_0_rsource; // @[L2TLB.scala 290:43]
  assign cache_io_refill_bits_req_info_dup_1_vpn = cache_io_refill_bits_req_info_dup_1_rvpn; // @[L2TLB.scala 290:43]
  assign cache_io_refill_bits_req_info_dup_1_source = cache_io_refill_bits_req_info_dup_1_rsource; // @[L2TLB.scala 290:43]
  assign cache_io_refill_bits_req_info_dup_2_vpn = cache_io_refill_bits_req_info_dup_2_rvpn; // @[L2TLB.scala 290:43]
  assign cache_io_refill_bits_req_info_dup_2_source = cache_io_refill_bits_req_info_dup_2_rsource; // @[L2TLB.scala 290:43]
  assign cache_io_refill_bits_level_dup_0 = cache_io_refill_bits_level_dup_0_r; // @[L2TLB.scala 291:40]
  assign cache_io_refill_bits_level_dup_1 = cache_io_refill_bits_level_dup_1_r; // @[L2TLB.scala 291:40]
  assign cache_io_refill_bits_level_dup_2 = cache_io_refill_bits_level_dup_2_r; // @[L2TLB.scala 291:40]
  assign cache_io_refill_bits_sel_pte_dup_0 = cache_io_refill_bits_sel_pte_dup_0_REG; // @[L2TLB.scala 293:42]
  assign cache_io_refill_bits_sel_pte_dup_1 = cache_io_refill_bits_sel_pte_dup_1_REG; // @[L2TLB.scala 293:42]
  assign cache_io_refill_bits_sel_pte_dup_2 = cache_io_refill_bits_sel_pte_dup_2_REG; // @[L2TLB.scala 293:42]
  assign cache_io_sfence_dup_0_valid = sfence_dup_2_valid; // @[L2TLB.scala 173:69]
  assign cache_io_sfence_dup_0_bits_rs1 = sfence_dup_2_bits_rs1; // @[L2TLB.scala 173:69]
  assign cache_io_sfence_dup_0_bits_rs2 = sfence_dup_2_bits_rs2; // @[L2TLB.scala 173:69]
  assign cache_io_sfence_dup_0_bits_addr = sfence_dup_2_bits_addr; // @[L2TLB.scala 173:69]
  assign cache_io_sfence_dup_0_bits_asid = sfence_dup_2_bits_asid; // @[L2TLB.scala 173:69]
  assign cache_io_sfence_dup_1_valid = sfence_dup_3_valid; // @[L2TLB.scala 173:69]
  assign cache_io_sfence_dup_2_valid = sfence_dup_4_valid; // @[L2TLB.scala 173:69]
  assign cache_io_sfence_dup_3_valid = sfence_dup_5_valid; // @[L2TLB.scala 173:69]
  assign cache_io_sfence_dup_3_bits_rs1 = sfence_dup_5_bits_rs1; // @[L2TLB.scala 173:69]
  assign cache_io_sfence_dup_3_bits_rs2 = sfence_dup_5_bits_rs2; // @[L2TLB.scala 173:69]
  assign cache_io_sfence_dup_3_bits_addr = sfence_dup_5_bits_addr; // @[L2TLB.scala 173:69]
  assign cache_io_csr_dup_0_satp_asid = csr_dup_2_satp_asid; // @[L2TLB.scala 174:63]
  assign cache_io_csr_dup_0_satp_changed = csr_dup_2_satp_changed; // @[L2TLB.scala 174:63]
  assign cache_io_csr_dup_1_satp_asid = csr_dup_3_satp_asid; // @[L2TLB.scala 174:63]
  assign cache_io_csr_dup_1_satp_changed = csr_dup_3_satp_changed; // @[L2TLB.scala 174:63]
  assign cache_io_csr_dup_2_satp_asid = csr_dup_4_satp_asid; // @[L2TLB.scala 174:63]
  assign cache_io_csr_dup_2_satp_changed = csr_dup_4_satp_changed; // @[L2TLB.scala 174:63]
  assign ptw_clock = clock;
  assign ptw_reset = reset;
  assign ptw_io_sfence_valid = sfence_dup_7_valid; // @[L2TLB.scala 187:17]
  assign ptw_io_csr_satp_asid = csr_dup_6_satp_asid; // @[L2TLB.scala 188:14]
  assign ptw_io_csr_satp_ppn = csr_dup_6_satp_ppn; // @[L2TLB.scala 188:14]
  assign ptw_io_req_valid = _ptw_io_req_valid_T_5 & _ptw_io_req_valid_T_6; // @[L2TLB.scala 182:34]
  assign ptw_io_req_bits_req_info_vpn = cache_io_resp_bits_req_info_vpn; // @[L2TLB.scala 184:28]
  assign ptw_io_req_bits_req_info_source = cache_io_resp_bits_req_info_source; // @[L2TLB.scala 184:28]
  assign ptw_io_req_bits_l1Hit = cache_io_resp_bits_toFsm_l1Hit; // @[L2TLB.scala 185:25]
  assign ptw_io_req_bits_ppn = cache_io_resp_bits_toFsm_ppn; // @[L2TLB.scala 186:23]
  assign ptw_io_resp_ready = 2'h1 == ptw_io_resp_bits_source ? Arbiter_1_io_in_1_ready : _ptw_io_resp_ready_T_1; // @[Mux.scala 81:58]
  assign ptw_io_llptw_ready = arb2_io_in_0_ready; // @[L2TLB.scala 120:22]
  assign ptw_io_mem_req_ready = auto_out_a_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign ptw_io_mem_resp_valid = mem_resp_done & _resp_pte_T_6; // @[L2TLB.scala 281:42]
  assign ptw_io_mem_resp_bits = resp_pte_r6; // @[L2TLB.scala 270:{25,25}]
  assign ptw_io_mem_mask = waiting_resp_6; // @[L2TLB.scala 213:19]
  assign ptw_io_pmp_resp_ld = PMPChecker_io_resp_ld; // @[L2TLB.scala 89:{26,26}]
  assign ptw_io_pmp_resp_mmio = PMPChecker_io_resp_mmio; // @[L2TLB.scala 89:{26,26}]
  assign llptw_clock = clock;
  assign llptw_reset = reset;
  assign llptw_io_sfence_valid = sfence_dup_1_valid; // @[L2TLB.scala 163:19]
  assign llptw_io_csr_satp_changed = csr_dup_1_satp_changed; // @[L2TLB.scala 164:16]
  assign llptw_io_in_valid = _mq_arb_io_in_0_valid_T_1 & cache_io_resp_bits_toFsm_l2Hit & ~cache_io_resp_bits_bypassed; // @[L2TLB.scala 160:105]
  assign llptw_io_in_bits_req_info_vpn = cache_io_resp_bits_req_info_vpn; // @[L2TLB.scala 161:29]
  assign llptw_io_in_bits_req_info_source = cache_io_resp_bits_req_info_source; // @[L2TLB.scala 161:29]
  assign llptw_io_in_bits_ppn = {{12'd0}, cache_io_resp_bits_toFsm_ppn}; // @[L2TLB.scala 162:24]
  assign llptw_io_out_ready = 2'h1 == llptw_io_out_bits_req_info_source ? Arbiter_1_io_in_2_ready :
    _llptw_io_out_ready_T_1; // @[Mux.scala 81:58]
  assign llptw_io_mem_req_ready = mem_arb_io_in_1_ready; // @[L2TLB.scala 217:20]
  assign llptw_io_mem_resp_valid = mem_resp_done & mem_resp_from_mq; // @[L2TLB.scala 277:41]
  assign llptw_io_mem_resp_bits_id = auto_out_d_valid ? auto_out_d_bits_source : llptw_io_mem_resp_bits_id_r; // @[Hold.scala 67:8]
  assign llptw_io_mem_req_mask_0 = waiting_resp_0; // @[L2TLB.scala 212:22]
  assign llptw_io_mem_req_mask_1 = waiting_resp_1; // @[L2TLB.scala 212:22]
  assign llptw_io_mem_req_mask_2 = waiting_resp_2; // @[L2TLB.scala 212:22]
  assign llptw_io_mem_req_mask_3 = waiting_resp_3; // @[L2TLB.scala 212:22]
  assign llptw_io_mem_req_mask_4 = waiting_resp_4; // @[L2TLB.scala 212:22]
  assign llptw_io_mem_req_mask_5 = waiting_resp_5; // @[L2TLB.scala 212:22]
  assign llptw_io_cache_ready = mq_arb_io_in_1_ready; // @[L2TLB.scala 152:19]
  assign llptw_io_pmp_resp_ld = PMPChecker_1_io_resp_ld; // @[L2TLB.scala 89:{26,26}]
  assign llptw_io_pmp_resp_mmio = PMPChecker_1_io_resp_mmio; // @[L2TLB.scala 89:{26,26}]
  assign arb1_io_in_0_valid = io_tlb_0_req_0_valid; // @[L2TLB.scala 114:{24,24}]
  assign arb1_io_in_0_bits_vpn = io_tlb_0_req_0_bits_vpn; // @[L2TLB.scala 114:{24,24}]
  assign arb1_io_in_1_valid = io_tlb_1_req_0_valid; // @[L2TLB.scala 114:{24,24}]
  assign arb1_io_in_1_bits_vpn = io_tlb_1_req_0_bits_vpn; // @[L2TLB.scala 114:{24,24}]
  assign arb1_io_out_ready = arb2_io_in_2_ready; // @[L2TLB.scala 115:21]
  assign arb2_io_in_0_valid = ptw_io_llptw_valid; // @[L2TLB.scala 117:34]
  assign arb2_io_in_0_bits_vpn = ptw_io_llptw_bits_req_info_vpn; // @[L2TLB.scala 118:37]
  assign arb2_io_in_0_bits_source = ptw_io_llptw_bits_req_info_source; // @[L2TLB.scala 119:40]
  assign arb2_io_in_1_valid = missQueue_io_out_valid & ~_T; // @[L2TLB.scala 365:34]
  assign arb2_io_in_1_bits_vpn = missQueue_io_out_bits_vpn; // @[L2TLB.scala 367:18]
  assign arb2_io_in_1_bits_source = missQueue_io_out_bits_source; // @[L2TLB.scala 367:18]
  assign arb2_io_in_2_valid = arb1_io_out_valid; // @[L2TLB.scala 123:34]
  assign arb2_io_in_2_bits_vpn = arb1_io_out_bits_vpn; // @[L2TLB.scala 124:37]
  assign arb2_io_in_2_bits_source = {{1'd0}, arb1_io_chosen}; // @[L2TLB.scala 125:40]
  assign arb2_io_in_3_valid = prefetch_io_out_valid; // @[L2TLB.scala 136:35]
  assign arb2_io_in_3_bits_vpn = prefetch_io_out_bits_vpn; // @[L2TLB.scala 136:35]
  assign arb2_io_out_ready = cache_io_req_ready; // @[L2TLB.scala 143:21]
  assign Arbiter_io_in_0_valid = cache_io_resp_valid & cache_io_resp_bits_hit & cache_io_resp_bits_req_info_source == 2'h0
    ; // @[L2TLB.scala 334:90]
  assign Arbiter_io_in_0_bits_entry_tag = cache_io_resp_bits_toTlb_tag; // @[L2TLB.scala 335:46]
  assign Arbiter_io_in_0_bits_entry_asid = cache_io_resp_bits_toTlb_asid; // @[L2TLB.scala 335:46]
  assign Arbiter_io_in_0_bits_entry_ppn = cache_io_resp_bits_toTlb_ppn; // @[L2TLB.scala 335:46]
  assign Arbiter_io_in_0_bits_entry_perm_d = cache_io_resp_bits_toTlb_perm_d; // @[L2TLB.scala 335:46]
  assign Arbiter_io_in_0_bits_entry_perm_a = cache_io_resp_bits_toTlb_perm_a; // @[L2TLB.scala 335:46]
  assign Arbiter_io_in_0_bits_entry_perm_g = cache_io_resp_bits_toTlb_perm_g; // @[L2TLB.scala 335:46]
  assign Arbiter_io_in_0_bits_entry_perm_u = cache_io_resp_bits_toTlb_perm_u; // @[L2TLB.scala 335:46]
  assign Arbiter_io_in_0_bits_entry_perm_x = cache_io_resp_bits_toTlb_perm_x; // @[L2TLB.scala 335:46]
  assign Arbiter_io_in_0_bits_entry_perm_w = cache_io_resp_bits_toTlb_perm_w; // @[L2TLB.scala 335:46]
  assign Arbiter_io_in_0_bits_entry_perm_r = cache_io_resp_bits_toTlb_perm_r; // @[L2TLB.scala 335:46]
  assign Arbiter_io_in_0_bits_entry_level = cache_io_resp_bits_toTlb_level; // @[L2TLB.scala 335:46]
  assign Arbiter_io_in_0_bits_pf = ~cache_io_resp_bits_toTlb_v; // @[L2TLB.scala 336:46]
  assign Arbiter_io_in_1_valid = ptw_io_resp_valid & ptw_io_resp_bits_source == 2'h0; // @[L2TLB.scala 338:60]
  assign Arbiter_io_in_1_bits_entry_tag = ptw_io_resp_bits_resp_entry_tag; // @[L2TLB.scala 339:38]
  assign Arbiter_io_in_1_bits_entry_asid = ptw_io_resp_bits_resp_entry_asid; // @[L2TLB.scala 339:38]
  assign Arbiter_io_in_1_bits_entry_ppn = ptw_io_resp_bits_resp_entry_ppn; // @[L2TLB.scala 339:38]
  assign Arbiter_io_in_1_bits_entry_perm_d = ptw_io_resp_bits_resp_entry_perm_d; // @[L2TLB.scala 339:38]
  assign Arbiter_io_in_1_bits_entry_perm_a = ptw_io_resp_bits_resp_entry_perm_a; // @[L2TLB.scala 339:38]
  assign Arbiter_io_in_1_bits_entry_perm_g = ptw_io_resp_bits_resp_entry_perm_g; // @[L2TLB.scala 339:38]
  assign Arbiter_io_in_1_bits_entry_perm_u = ptw_io_resp_bits_resp_entry_perm_u; // @[L2TLB.scala 339:38]
  assign Arbiter_io_in_1_bits_entry_perm_x = ptw_io_resp_bits_resp_entry_perm_x; // @[L2TLB.scala 339:38]
  assign Arbiter_io_in_1_bits_entry_perm_w = ptw_io_resp_bits_resp_entry_perm_w; // @[L2TLB.scala 339:38]
  assign Arbiter_io_in_1_bits_entry_perm_r = ptw_io_resp_bits_resp_entry_perm_r; // @[L2TLB.scala 339:38]
  assign Arbiter_io_in_1_bits_entry_level = ptw_io_resp_bits_resp_entry_level; // @[L2TLB.scala 339:38]
  assign Arbiter_io_in_1_bits_pf = ptw_io_resp_bits_resp_pf; // @[L2TLB.scala 339:38]
  assign Arbiter_io_in_1_bits_af = ptw_io_resp_bits_resp_af; // @[L2TLB.scala 339:38]
  assign Arbiter_io_in_2_valid = llptw_io_out_valid & llptw_io_out_bits_req_info_source == 2'h0; // @[L2TLB.scala 340:57]
  assign Arbiter_io_in_2_bits_entry_tag = llptw_io_out_bits_req_info_vpn; // @[L2TLB.scala 377:24 381:24]
  assign Arbiter_io_in_2_bits_entry_asid = csr_dup_0_satp_asid; // @[L2TLB.scala 377:24 386:25]
  assign Arbiter_io_in_2_bits_entry_ppn = _GEN_171[33:10]; // @[L2TLB.scala 376:30]
  assign Arbiter_io_in_2_bits_entry_perm_d = _GEN_171[7]; // @[L2TLB.scala 376:30]
  assign Arbiter_io_in_2_bits_entry_perm_a = _GEN_171[6]; // @[L2TLB.scala 376:30]
  assign Arbiter_io_in_2_bits_entry_perm_g = _GEN_171[5]; // @[L2TLB.scala 376:30]
  assign Arbiter_io_in_2_bits_entry_perm_u = _GEN_171[4]; // @[L2TLB.scala 376:30]
  assign Arbiter_io_in_2_bits_entry_perm_x = _GEN_171[3]; // @[L2TLB.scala 376:30]
  assign Arbiter_io_in_2_bits_entry_perm_w = _GEN_171[2]; // @[L2TLB.scala 376:30]
  assign Arbiter_io_in_2_bits_entry_perm_r = _GEN_171[1]; // @[L2TLB.scala 376:30]
  assign Arbiter_io_in_2_bits_pf = ~llptw_io_out_bits_af & _ptw_resp_pf_T_4; // @[L2TLB.scala 382:52]
  assign Arbiter_io_in_2_bits_af = llptw_io_out_bits_af | _ptw_resp_af_T_1; // @[L2TLB.scala 383:73]
  assign Arbiter_io_out_ready = io_tlb_0_resp_ready; // @[L2TLB.scala 346:30]
  assign Arbiter_1_io_in_0_valid = cache_io_resp_valid & cache_io_resp_bits_hit & cache_io_resp_bits_req_info_source == 2'h1
    ; // @[L2TLB.scala 334:90]
  assign Arbiter_1_io_in_0_bits_entry_tag = cache_io_resp_bits_toTlb_tag; // @[L2TLB.scala 335:46]
  assign Arbiter_1_io_in_0_bits_entry_asid = cache_io_resp_bits_toTlb_asid; // @[L2TLB.scala 335:46]
  assign Arbiter_1_io_in_0_bits_entry_ppn = cache_io_resp_bits_toTlb_ppn; // @[L2TLB.scala 335:46]
  assign Arbiter_1_io_in_0_bits_entry_perm_d = cache_io_resp_bits_toTlb_perm_d; // @[L2TLB.scala 335:46]
  assign Arbiter_1_io_in_0_bits_entry_perm_a = cache_io_resp_bits_toTlb_perm_a; // @[L2TLB.scala 335:46]
  assign Arbiter_1_io_in_0_bits_entry_perm_g = cache_io_resp_bits_toTlb_perm_g; // @[L2TLB.scala 335:46]
  assign Arbiter_1_io_in_0_bits_entry_perm_u = cache_io_resp_bits_toTlb_perm_u; // @[L2TLB.scala 335:46]
  assign Arbiter_1_io_in_0_bits_entry_perm_x = cache_io_resp_bits_toTlb_perm_x; // @[L2TLB.scala 335:46]
  assign Arbiter_1_io_in_0_bits_entry_perm_w = cache_io_resp_bits_toTlb_perm_w; // @[L2TLB.scala 335:46]
  assign Arbiter_1_io_in_0_bits_entry_perm_r = cache_io_resp_bits_toTlb_perm_r; // @[L2TLB.scala 335:46]
  assign Arbiter_1_io_in_0_bits_entry_level = cache_io_resp_bits_toTlb_level; // @[L2TLB.scala 335:46]
  assign Arbiter_1_io_in_0_bits_pf = ~cache_io_resp_bits_toTlb_v; // @[L2TLB.scala 336:46]
  assign Arbiter_1_io_in_1_valid = ptw_io_resp_valid & ptw_io_resp_bits_source == 2'h1; // @[L2TLB.scala 338:60]
  assign Arbiter_1_io_in_1_bits_entry_tag = ptw_io_resp_bits_resp_entry_tag; // @[L2TLB.scala 339:38]
  assign Arbiter_1_io_in_1_bits_entry_asid = ptw_io_resp_bits_resp_entry_asid; // @[L2TLB.scala 339:38]
  assign Arbiter_1_io_in_1_bits_entry_ppn = ptw_io_resp_bits_resp_entry_ppn; // @[L2TLB.scala 339:38]
  assign Arbiter_1_io_in_1_bits_entry_perm_d = ptw_io_resp_bits_resp_entry_perm_d; // @[L2TLB.scala 339:38]
  assign Arbiter_1_io_in_1_bits_entry_perm_a = ptw_io_resp_bits_resp_entry_perm_a; // @[L2TLB.scala 339:38]
  assign Arbiter_1_io_in_1_bits_entry_perm_g = ptw_io_resp_bits_resp_entry_perm_g; // @[L2TLB.scala 339:38]
  assign Arbiter_1_io_in_1_bits_entry_perm_u = ptw_io_resp_bits_resp_entry_perm_u; // @[L2TLB.scala 339:38]
  assign Arbiter_1_io_in_1_bits_entry_perm_x = ptw_io_resp_bits_resp_entry_perm_x; // @[L2TLB.scala 339:38]
  assign Arbiter_1_io_in_1_bits_entry_perm_w = ptw_io_resp_bits_resp_entry_perm_w; // @[L2TLB.scala 339:38]
  assign Arbiter_1_io_in_1_bits_entry_perm_r = ptw_io_resp_bits_resp_entry_perm_r; // @[L2TLB.scala 339:38]
  assign Arbiter_1_io_in_1_bits_entry_level = ptw_io_resp_bits_resp_entry_level; // @[L2TLB.scala 339:38]
  assign Arbiter_1_io_in_1_bits_pf = ptw_io_resp_bits_resp_pf; // @[L2TLB.scala 339:38]
  assign Arbiter_1_io_in_1_bits_af = ptw_io_resp_bits_resp_af; // @[L2TLB.scala 339:38]
  assign Arbiter_1_io_in_2_valid = llptw_io_out_valid & llptw_io_out_bits_req_info_source == 2'h1; // @[L2TLB.scala 340:57]
  assign Arbiter_1_io_in_2_bits_entry_tag = llptw_io_out_bits_req_info_vpn; // @[L2TLB.scala 377:24 381:24]
  assign Arbiter_1_io_in_2_bits_entry_asid = csr_dup_0_satp_asid; // @[L2TLB.scala 377:24 386:25]
  assign Arbiter_1_io_in_2_bits_entry_ppn = _GEN_171[33:10]; // @[L2TLB.scala 376:30]
  assign Arbiter_1_io_in_2_bits_entry_perm_d = _GEN_171[7]; // @[L2TLB.scala 376:30]
  assign Arbiter_1_io_in_2_bits_entry_perm_a = _GEN_171[6]; // @[L2TLB.scala 376:30]
  assign Arbiter_1_io_in_2_bits_entry_perm_g = _GEN_171[5]; // @[L2TLB.scala 376:30]
  assign Arbiter_1_io_in_2_bits_entry_perm_u = _GEN_171[4]; // @[L2TLB.scala 376:30]
  assign Arbiter_1_io_in_2_bits_entry_perm_x = _GEN_171[3]; // @[L2TLB.scala 376:30]
  assign Arbiter_1_io_in_2_bits_entry_perm_w = _GEN_171[2]; // @[L2TLB.scala 376:30]
  assign Arbiter_1_io_in_2_bits_entry_perm_r = _GEN_171[1]; // @[L2TLB.scala 376:30]
  assign Arbiter_1_io_in_2_bits_pf = ~llptw_io_out_bits_af & _ptw_resp_pf_T_4; // @[L2TLB.scala 382:52]
  assign Arbiter_1_io_in_2_bits_af = llptw_io_out_bits_af | _ptw_resp_af_T_1; // @[L2TLB.scala 383:73]
  assign Arbiter_1_io_out_ready = io_tlb_1_resp_ready; // @[L2TLB.scala 346:30]
  assign prefetch_clock = clock;
  assign prefetch_reset = reset;
  assign prefetch_io_sfence_valid = sfence_dup_0_valid; // @[L2TLB.scala 134:24]
  assign prefetch_io_csr_satp_changed = csr_dup_0_satp_changed; // @[L2TLB.scala 135:21]
  assign prefetch_io_in_valid = _prefetch_io_in_valid_T_6 & cache_io_resp_bits_isFirst; // @[L2TLB.scala 132:27]
  assign prefetch_io_in_bits_vpn = cache_io_resp_bits_req_info_vpn; // @[L2TLB.scala 133:29]
  assign prefetch_io_out_ready = arb2_io_in_3_ready; // @[L2TLB.scala 136:35]
  assign writer_clock = clock; // @[ChiselDB.scala 135:21]
  assign writer_reset = reset; // @[ChiselDB.scala 136:21]
  assign writer_en = prefetch_io_out_ready & prefetch_io_out_valid; // @[Decoupled.scala 50:35]
  assign writer_stamp = cnt; // @[ChiselDB.scala 138:21]
  assign writer_data_vpn = prefetch_io_out_bits_vpn; // @[L2TLB.scala 139:31 140:25]
  assign mq_arb_io_in_0_valid = _mq_arb_io_in_0_valid_T_7 & _mq_arb_io_in_0_valid_T_10; // @[L2TLB.scala 149:51]
  assign mq_arb_io_in_0_bits_vpn = cache_io_resp_bits_req_info_vpn; // @[L2TLB.scala 151:24]
  assign mq_arb_io_in_0_bits_source = cache_io_resp_bits_req_info_source; // @[L2TLB.scala 151:24]
  assign mq_arb_io_in_1_valid = llptw_io_cache_valid; // @[L2TLB.scala 152:19]
  assign mq_arb_io_in_1_bits_vpn = llptw_io_cache_bits_vpn; // @[L2TLB.scala 152:19]
  assign mq_arb_io_in_1_bits_source = llptw_io_cache_bits_source; // @[L2TLB.scala 152:19]
  assign mq_arb_io_out_ready = missQueue_io_in_ready; // @[L2TLB.scala 153:19]
  assign mem_arb_io_in_0_valid = ptw_io_mem_req_valid; // @[L2TLB.scala 216:20]
  assign mem_arb_io_in_0_bits_addr = ptw_io_mem_req_bits_addr; // @[L2TLB.scala 216:20]
  assign mem_arb_io_in_1_valid = llptw_io_mem_req_valid; // @[L2TLB.scala 217:20]
  assign mem_arb_io_in_1_bits_addr = llptw_io_mem_req_bits_addr; // @[L2TLB.scala 217:20]
  assign mem_arb_io_in_1_bits_id = llptw_io_mem_req_bits_id; // @[L2TLB.scala 217:20]
  assign mem_arb_io_out_ready = auto_out_a_ready & ~flush; // @[L2TLB.scala 218:39]
  assign writer_1_clock = clock; // @[ChiselDB.scala 135:21]
  assign writer_1_reset = reset; // @[ChiselDB.scala 136:21]
  assign writer_1_en = io_tlb_0_req_0_ready & io_tlb_0_req_0_valid; // @[Decoupled.scala 50:35]
  assign writer_1_stamp = cnt_1; // @[ChiselDB.scala 138:21]
  assign writer_1_data_vpn = io_tlb_0_req_0_bits_vpn; // @[L2TLB.scala 431:58 432:17]
  assign writer_2_clock = clock; // @[ChiselDB.scala 135:21]
  assign writer_2_reset = reset; // @[ChiselDB.scala 136:21]
  assign writer_2_en = io_tlb_1_req_0_ready & io_tlb_1_req_0_valid; // @[Decoupled.scala 50:35]
  assign writer_2_stamp = cnt_2; // @[ChiselDB.scala 138:21]
  assign writer_2_data_vpn = io_tlb_1_req_0_bits_vpn; // @[L2TLB.scala 431:58 433:17]
  assign writer_3_clock = clock; // @[ChiselDB.scala 135:21]
  assign writer_3_reset = reset; // @[ChiselDB.scala 136:21]
  assign writer_3_en = io_tlb_0_resp_ready & io_tlb_0_resp_valid; // @[Decoupled.scala 50:35]
  assign writer_3_stamp = cnt_3; // @[ChiselDB.scala 138:21]
  assign writer_3_data_vpn = io_tlb_0_resp_bits_entry_tag; // @[L2TLB.scala 431:58 434:18]
  assign writer_4_clock = clock; // @[ChiselDB.scala 135:21]
  assign writer_4_reset = reset; // @[ChiselDB.scala 136:21]
  assign writer_4_en = io_tlb_1_resp_ready & io_tlb_1_resp_valid; // @[Decoupled.scala 50:35]
  assign writer_4_stamp = cnt_4; // @[ChiselDB.scala 138:21]
  assign writer_4_data_vpn = io_tlb_1_resp_bits_entry_tag; // @[L2TLB.scala 431:58 435:18]
  assign writer_5_clock = clock; // @[ChiselDB.scala 135:21]
  assign writer_5_reset = reset; // @[ChiselDB.scala 136:21]
  assign writer_5_en = cache_io_resp_ready & cache_io_resp_valid; // @[Decoupled.scala 50:35]
  assign writer_5_stamp = cnt_5; // @[ChiselDB.scala 138:21]
  assign writer_5_data_vpn = cache_io_resp_bits_toTlb_tag; // @[L2TLB.scala 442:25 443:19]
  assign writer_5_data_source = cache_io_resp_bits_req_info_source; // @[L2TLB.scala 442:25 444:22]
  assign writer_5_data_bypassed = cache_io_resp_bits_bypassed; // @[L2TLB.scala 442:25 445:24]
  assign writer_5_data_is_first = cache_io_resp_bits_isFirst; // @[L2TLB.scala 442:25 446:24]
  assign writer_5_data_prefetched = cache_io_resp_bits_toTlb_prefetch; // @[L2TLB.scala 442:25 447:26]
  assign writer_5_data_prefetch = cache_io_resp_bits_prefetch; // @[L2TLB.scala 442:25 448:24]
  assign writer_5_data_l2Hit = cache_io_resp_bits_toFsm_l2Hit; // @[L2TLB.scala 442:25 449:21]
  assign writer_5_data_l1Hit = cache_io_resp_bits_toFsm_l1Hit; // @[L2TLB.scala 442:25 450:21]
  assign writer_5_data_hit = cache_io_resp_bits_hit; // @[L2TLB.scala 442:25 451:19]
  assign writer_6_clock = clock; // @[ChiselDB.scala 135:21]
  assign writer_6_reset = reset; // @[ChiselDB.scala 136:21]
  assign writer_6_en = ptw_io_req_ready & ptw_io_req_valid; // @[Decoupled.scala 50:35]
  assign writer_6_stamp = cnt_6; // @[ChiselDB.scala 138:21]
  assign writer_6_data_vpn = ptw_io_req_bits_req_info_vpn; // @[L2TLB.scala 455:58 456:16]
  assign writer_6_data_source = ptw_io_req_bits_req_info_source; // @[L2TLB.scala 455:58 457:19]
  assign writer_7_clock = clock; // @[ChiselDB.scala 135:21]
  assign writer_7_reset = reset; // @[ChiselDB.scala 136:21]
  assign writer_7_en = ptw_io_mem_resp_valid; // @[ChiselDB.scala 137:18]
  assign writer_7_stamp = cnt_7; // @[ChiselDB.scala 138:21]
  assign writer_7_data_vpn = ptw_io_refill_req_info_vpn; // @[L2TLB.scala 455:58 458:17]
  assign writer_7_data_source = ptw_io_refill_req_info_source; // @[L2TLB.scala 455:58 459:20]
  assign writer_8_clock = clock; // @[ChiselDB.scala 135:21]
  assign writer_8_reset = reset; // @[ChiselDB.scala 136:21]
  assign writer_8_en = llptw_io_in_ready & llptw_io_in_valid; // @[Decoupled.scala 50:35]
  assign writer_8_stamp = cnt_8; // @[ChiselDB.scala 138:21]
  assign writer_8_data_vpn = llptw_io_in_bits_req_info_vpn; // @[L2TLB.scala 455:58 460:18]
  assign writer_8_data_source = llptw_io_in_bits_req_info_source; // @[L2TLB.scala 455:58 461:21]
  assign writer_9_clock = clock; // @[ChiselDB.scala 135:21]
  assign writer_9_reset = reset; // @[ChiselDB.scala 136:21]
  assign writer_9_en = llptw_io_mem_resp_valid; // @[ChiselDB.scala 137:18]
  assign writer_9_stamp = cnt_9; // @[ChiselDB.scala 138:21]
  assign writer_9_data_vpn = llptw_io_mem_refill_vpn; // @[L2TLB.scala 455:58 462:19]
  assign writer_9_data_source = llptw_io_mem_refill_source; // @[L2TLB.scala 455:58 463:22]
  assign writer_10_clock = clock; // @[ChiselDB.scala 135:21]
  assign writer_10_reset = reset; // @[ChiselDB.scala 136:21]
  assign writer_10_en = missQueue_io_in_ready & missQueue_io_in_valid; // @[Decoupled.scala 50:35]
  assign writer_10_stamp = cnt_10; // @[ChiselDB.scala 138:21]
  assign writer_10_data_vpn = missQueue_io_in_bits_vpn; // @[L2TLB.scala 470:53 471:26]
  assign writer_11_clock = clock; // @[ChiselDB.scala 135:21]
  assign writer_11_reset = reset; // @[ChiselDB.scala 136:21]
  assign writer_11_en = missQueue_io_out_ready & missQueue_io_out_valid; // @[Decoupled.scala 50:35]
  assign writer_11_stamp = cnt_11; // @[ChiselDB.scala 138:21]
  assign writer_11_data_vpn = missQueue_io_out_bits_vpn; // @[L2TLB.scala 470:53 472:27]
  always @(posedge clock) begin
    sfence_dup_0_valid <= sfence_tmp_delay_io_out_valid; // @[L2TLB.scala 82:39]
    sfence_dup_1_valid <= sfence_tmp_delay_io_out_valid; // @[L2TLB.scala 82:39]
    sfence_dup_2_valid <= sfence_tmp_delay_io_out_valid; // @[L2TLB.scala 82:39]
    sfence_dup_2_bits_rs1 <= sfence_tmp_delay_io_out_bits_rs1; // @[L2TLB.scala 82:39]
    sfence_dup_2_bits_rs2 <= sfence_tmp_delay_io_out_bits_rs2; // @[L2TLB.scala 82:39]
    sfence_dup_2_bits_addr <= sfence_tmp_delay_io_out_bits_addr; // @[L2TLB.scala 82:39]
    sfence_dup_2_bits_asid <= sfence_tmp_delay_io_out_bits_asid; // @[L2TLB.scala 82:39]
    sfence_dup_3_valid <= sfence_tmp_delay_io_out_valid; // @[L2TLB.scala 82:39]
    sfence_dup_4_valid <= sfence_tmp_delay_io_out_valid; // @[L2TLB.scala 82:39]
    sfence_dup_5_valid <= sfence_tmp_delay_io_out_valid; // @[L2TLB.scala 82:39]
    sfence_dup_5_bits_rs1 <= sfence_tmp_delay_io_out_bits_rs1; // @[L2TLB.scala 82:39]
    sfence_dup_5_bits_rs2 <= sfence_tmp_delay_io_out_bits_rs2; // @[L2TLB.scala 82:39]
    sfence_dup_5_bits_addr <= sfence_tmp_delay_io_out_bits_addr; // @[L2TLB.scala 82:39]
    sfence_dup_6_valid <= sfence_tmp_delay_io_out_valid; // @[L2TLB.scala 82:39]
    sfence_dup_7_valid <= sfence_tmp_delay_io_out_valid; // @[L2TLB.scala 82:39]
    csr_dup_0_satp_asid <= csr_tmp_delay_io_out_satp_asid; // @[L2TLB.scala 83:36]
    csr_dup_0_satp_changed <= csr_tmp_delay_io_out_satp_changed; // @[L2TLB.scala 83:36]
    csr_dup_1_satp_changed <= csr_tmp_delay_io_out_satp_changed; // @[L2TLB.scala 83:36]
    csr_dup_2_satp_asid <= csr_tmp_delay_io_out_satp_asid; // @[L2TLB.scala 83:36]
    csr_dup_2_satp_changed <= csr_tmp_delay_io_out_satp_changed; // @[L2TLB.scala 83:36]
    csr_dup_3_satp_asid <= csr_tmp_delay_io_out_satp_asid; // @[L2TLB.scala 83:36]
    csr_dup_3_satp_changed <= csr_tmp_delay_io_out_satp_changed; // @[L2TLB.scala 83:36]
    csr_dup_4_satp_asid <= csr_tmp_delay_io_out_satp_asid; // @[L2TLB.scala 83:36]
    csr_dup_4_satp_changed <= csr_tmp_delay_io_out_satp_changed; // @[L2TLB.scala 83:36]
    csr_dup_5_satp_changed <= csr_tmp_delay_io_out_satp_changed; // @[L2TLB.scala 83:36]
    csr_dup_6_satp_asid <= csr_tmp_delay_io_out_satp_asid; // @[L2TLB.scala 83:36]
    csr_dup_6_satp_ppn <= csr_tmp_delay_io_out_satp_ppn; // @[L2TLB.scala 83:36]
    if (_T_43) begin // @[L2TLB.scala 241:32]
      if (3'h0 == mem_arb_io_out_bits_id) begin // @[L2TLB.scala 242:42]
        req_addr_low_0 <= mem_arb_io_out_bits_addr[5:3]; // @[L2TLB.scala 242:42]
      end else begin
        req_addr_low_0 <= _GEN_11;
      end
    end else begin
      req_addr_low_0 <= _GEN_11;
    end
    if (_T_43) begin // @[L2TLB.scala 241:32]
      if (3'h1 == mem_arb_io_out_bits_id) begin // @[L2TLB.scala 242:42]
        req_addr_low_1 <= mem_arb_io_out_bits_addr[5:3]; // @[L2TLB.scala 242:42]
      end else begin
        req_addr_low_1 <= _GEN_12;
      end
    end else begin
      req_addr_low_1 <= _GEN_12;
    end
    if (_T_43) begin // @[L2TLB.scala 241:32]
      if (3'h2 == mem_arb_io_out_bits_id) begin // @[L2TLB.scala 242:42]
        req_addr_low_2 <= mem_arb_io_out_bits_addr[5:3]; // @[L2TLB.scala 242:42]
      end else begin
        req_addr_low_2 <= _GEN_13;
      end
    end else begin
      req_addr_low_2 <= _GEN_13;
    end
    if (_T_43) begin // @[L2TLB.scala 241:32]
      if (3'h3 == mem_arb_io_out_bits_id) begin // @[L2TLB.scala 242:42]
        req_addr_low_3 <= mem_arb_io_out_bits_addr[5:3]; // @[L2TLB.scala 242:42]
      end else begin
        req_addr_low_3 <= _GEN_14;
      end
    end else begin
      req_addr_low_3 <= _GEN_14;
    end
    if (_T_43) begin // @[L2TLB.scala 241:32]
      if (3'h4 == mem_arb_io_out_bits_id) begin // @[L2TLB.scala 242:42]
        req_addr_low_4 <= mem_arb_io_out_bits_addr[5:3]; // @[L2TLB.scala 242:42]
      end else begin
        req_addr_low_4 <= _GEN_15;
      end
    end else begin
      req_addr_low_4 <= _GEN_15;
    end
    if (_T_43) begin // @[L2TLB.scala 241:32]
      if (3'h5 == mem_arb_io_out_bits_id) begin // @[L2TLB.scala 242:42]
        req_addr_low_5 <= mem_arb_io_out_bits_addr[5:3]; // @[L2TLB.scala 242:42]
      end else begin
        req_addr_low_5 <= _GEN_16;
      end
    end else begin
      req_addr_low_5 <= _GEN_16;
    end
    if (_T_43) begin // @[L2TLB.scala 241:32]
      if (3'h6 == mem_arb_io_out_bits_id) begin // @[L2TLB.scala 242:42]
        req_addr_low_6 <= mem_arb_io_out_bits_addr[5:3]; // @[L2TLB.scala 242:42]
      end else begin
        req_addr_low_6 <= _GEN_17;
      end
    end else begin
      req_addr_low_6 <= _GEN_17;
    end
    if (auto_out_d_valid) begin // @[L2TLB.scala 260:22]
      if (~count) begin // @[L2TLB.scala 262:35]
        refill_data_0 <= auto_out_d_bits_data; // @[L2TLB.scala 262:35]
      end
    end
    if (auto_out_d_valid) begin // @[L2TLB.scala 260:22]
      if (count) begin // @[L2TLB.scala 262:35]
        refill_data_1 <= auto_out_d_bits_data; // @[L2TLB.scala 262:35]
      end
    end
    if (llptw_io_mem_buffer_it_0) begin // @[Reg.scala 17:18]
      if (3'h7 == req_addr_low_0) begin // @[Reg.scala 17:22]
        resp_pte_r <= inner_data__7; // @[Reg.scala 17:22]
      end else if (3'h6 == req_addr_low_0) begin // @[Reg.scala 17:22]
        resp_pte_r <= inner_data__6; // @[Reg.scala 17:22]
      end else if (3'h5 == req_addr_low_0) begin // @[Reg.scala 17:22]
        resp_pte_r <= inner_data__5; // @[Reg.scala 17:22]
      end else begin
        resp_pte_r <= _GEN_57;
      end
    end
    if (llptw_io_mem_buffer_it_1) begin // @[Reg.scala 17:18]
      if (3'h7 == req_addr_low_1) begin // @[Reg.scala 17:22]
        resp_pte_r1 <= inner_data__7; // @[Reg.scala 17:22]
      end else if (3'h6 == req_addr_low_1) begin // @[Reg.scala 17:22]
        resp_pte_r1 <= inner_data__6; // @[Reg.scala 17:22]
      end else if (3'h5 == req_addr_low_1) begin // @[Reg.scala 17:22]
        resp_pte_r1 <= inner_data__5; // @[Reg.scala 17:22]
      end else begin
        resp_pte_r1 <= _GEN_66;
      end
    end
    if (llptw_io_mem_buffer_it_2) begin // @[Reg.scala 17:18]
      if (3'h7 == req_addr_low_2) begin // @[Reg.scala 17:22]
        resp_pte_r2 <= inner_data__7; // @[Reg.scala 17:22]
      end else if (3'h6 == req_addr_low_2) begin // @[Reg.scala 17:22]
        resp_pte_r2 <= inner_data__6; // @[Reg.scala 17:22]
      end else if (3'h5 == req_addr_low_2) begin // @[Reg.scala 17:22]
        resp_pte_r2 <= inner_data__5; // @[Reg.scala 17:22]
      end else begin
        resp_pte_r2 <= _GEN_75;
      end
    end
    if (llptw_io_mem_buffer_it_3) begin // @[Reg.scala 17:18]
      if (3'h7 == req_addr_low_3) begin // @[Reg.scala 17:22]
        resp_pte_r3 <= inner_data__7; // @[Reg.scala 17:22]
      end else if (3'h6 == req_addr_low_3) begin // @[Reg.scala 17:22]
        resp_pte_r3 <= inner_data__6; // @[Reg.scala 17:22]
      end else if (3'h5 == req_addr_low_3) begin // @[Reg.scala 17:22]
        resp_pte_r3 <= inner_data__5; // @[Reg.scala 17:22]
      end else begin
        resp_pte_r3 <= _GEN_84;
      end
    end
    if (llptw_io_mem_buffer_it_4) begin // @[Reg.scala 17:18]
      if (3'h7 == req_addr_low_4) begin // @[Reg.scala 17:22]
        resp_pte_r4 <= inner_data__7; // @[Reg.scala 17:22]
      end else if (3'h6 == req_addr_low_4) begin // @[Reg.scala 17:22]
        resp_pte_r4 <= inner_data__6; // @[Reg.scala 17:22]
      end else if (3'h5 == req_addr_low_4) begin // @[Reg.scala 17:22]
        resp_pte_r4 <= inner_data__5; // @[Reg.scala 17:22]
      end else begin
        resp_pte_r4 <= _GEN_93;
      end
    end
    if (llptw_io_mem_buffer_it_5) begin // @[Reg.scala 17:18]
      if (3'h7 == req_addr_low_5) begin // @[Reg.scala 17:22]
        resp_pte_r5 <= inner_data__7; // @[Reg.scala 17:22]
      end else if (3'h6 == req_addr_low_5) begin // @[Reg.scala 17:22]
        resp_pte_r5 <= inner_data__6; // @[Reg.scala 17:22]
      end else if (3'h5 == req_addr_low_5) begin // @[Reg.scala 17:22]
        resp_pte_r5 <= inner_data__5; // @[Reg.scala 17:22]
      end else begin
        resp_pte_r5 <= _GEN_102;
      end
    end
    if (_resp_pte_T_7) begin // @[Reg.scala 17:18]
      if (3'h7 == req_addr_low_6) begin // @[Reg.scala 17:22]
        resp_pte_r6 <= inner_data_6_7; // @[Reg.scala 17:22]
      end else if (3'h6 == req_addr_low_6) begin // @[Reg.scala 17:22]
        resp_pte_r6 <= inner_data_6_6; // @[Reg.scala 17:22]
      end else if (3'h5 == req_addr_low_6) begin // @[Reg.scala 17:22]
        resp_pte_r6 <= inner_data_6_5; // @[Reg.scala 17:22]
      end else begin
        resp_pte_r6 <= _GEN_111;
      end
    end
    if (auto_out_d_valid) begin // @[Reg.scala 17:18]
      llptw_io_mem_resp_bits_id_r <= auto_out_d_bits_source; // @[Reg.scala 17:22]
    end
    if (refill_valid) begin // @[Reg.scala 17:18]
      if (mem_resp_from_mq) begin // @[L2TLB.scala 290:59]
        cache_io_refill_bits_req_info_dup_0_rvpn <= llptw_io_mem_refill_vpn;
      end else begin
        cache_io_refill_bits_req_info_dup_0_rvpn <= ptw_io_refill_req_info_vpn;
      end
    end
    if (refill_valid) begin // @[Reg.scala 17:18]
      if (mem_resp_from_mq) begin // @[L2TLB.scala 290:59]
        cache_io_refill_bits_req_info_dup_0_rsource <= llptw_io_mem_refill_source;
      end else begin
        cache_io_refill_bits_req_info_dup_0_rsource <= ptw_io_refill_req_info_source;
      end
    end
    if (refill_valid) begin // @[Reg.scala 17:18]
      if (mem_resp_from_mq) begin // @[L2TLB.scala 290:59]
        cache_io_refill_bits_req_info_dup_1_rvpn <= llptw_io_mem_refill_vpn;
      end else begin
        cache_io_refill_bits_req_info_dup_1_rvpn <= ptw_io_refill_req_info_vpn;
      end
    end
    if (refill_valid) begin // @[Reg.scala 17:18]
      if (mem_resp_from_mq) begin // @[L2TLB.scala 290:59]
        cache_io_refill_bits_req_info_dup_1_rsource <= llptw_io_mem_refill_source;
      end else begin
        cache_io_refill_bits_req_info_dup_1_rsource <= ptw_io_refill_req_info_source;
      end
    end
    if (refill_valid) begin // @[Reg.scala 17:18]
      if (mem_resp_from_mq) begin // @[L2TLB.scala 290:59]
        cache_io_refill_bits_req_info_dup_2_rvpn <= llptw_io_mem_refill_vpn;
      end else begin
        cache_io_refill_bits_req_info_dup_2_rvpn <= ptw_io_refill_req_info_vpn;
      end
    end
    if (refill_valid) begin // @[Reg.scala 17:18]
      if (mem_resp_from_mq) begin // @[L2TLB.scala 290:59]
        cache_io_refill_bits_req_info_dup_2_rsource <= llptw_io_mem_refill_source;
      end else begin
        cache_io_refill_bits_req_info_dup_2_rsource <= ptw_io_refill_req_info_source;
      end
    end
    if (refill_valid) begin // @[Reg.scala 17:18]
      if (mem_resp_from_mq) begin // @[L2TLB.scala 285:25]
        cache_io_refill_bits_level_dup_0_r <= 2'h2;
      end else begin
        cache_io_refill_bits_level_dup_0_r <= refill_level_r;
      end
    end
    if (refill_valid) begin // @[Reg.scala 17:18]
      if (mem_resp_from_mq) begin // @[L2TLB.scala 285:25]
        cache_io_refill_bits_level_dup_1_r <= 2'h2;
      end else begin
        cache_io_refill_bits_level_dup_1_r <= refill_level_r;
      end
    end
    if (refill_valid) begin // @[Reg.scala 17:18]
      if (mem_resp_from_mq) begin // @[L2TLB.scala 285:25]
        cache_io_refill_bits_level_dup_2_r <= 2'h2;
      end else begin
        cache_io_refill_bits_level_dup_2_r <= refill_level_r;
      end
    end
    if (3'h7 == _GEN_140) begin // @[L2TLB.scala 293:52]
      cache_io_refill_bits_sel_pte_dup_0_REG <= inner_data_6_7; // @[L2TLB.scala 293:52]
    end else if (3'h6 == _GEN_140) begin // @[L2TLB.scala 293:52]
      cache_io_refill_bits_sel_pte_dup_0_REG <= inner_data_6_6; // @[L2TLB.scala 293:52]
    end else if (3'h5 == _GEN_140) begin // @[L2TLB.scala 293:52]
      cache_io_refill_bits_sel_pte_dup_0_REG <= inner_data_6_5; // @[L2TLB.scala 293:52]
    end else if (3'h4 == _GEN_140) begin // @[L2TLB.scala 293:52]
      cache_io_refill_bits_sel_pte_dup_0_REG <= inner_data_6_4; // @[L2TLB.scala 293:52]
    end else begin
      cache_io_refill_bits_sel_pte_dup_0_REG <= _GEN_144;
    end
    if (3'h7 == _GEN_140) begin // @[L2TLB.scala 293:52]
      cache_io_refill_bits_sel_pte_dup_1_REG <= inner_data_6_7; // @[L2TLB.scala 293:52]
    end else if (3'h6 == _GEN_140) begin // @[L2TLB.scala 293:52]
      cache_io_refill_bits_sel_pte_dup_1_REG <= inner_data_6_6; // @[L2TLB.scala 293:52]
    end else if (3'h5 == _GEN_140) begin // @[L2TLB.scala 293:52]
      cache_io_refill_bits_sel_pte_dup_1_REG <= inner_data_6_5; // @[L2TLB.scala 293:52]
    end else if (3'h4 == _GEN_140) begin // @[L2TLB.scala 293:52]
      cache_io_refill_bits_sel_pte_dup_1_REG <= inner_data_6_4; // @[L2TLB.scala 293:52]
    end else begin
      cache_io_refill_bits_sel_pte_dup_1_REG <= _GEN_144;
    end
    if (3'h7 == _GEN_140) begin // @[L2TLB.scala 293:52]
      cache_io_refill_bits_sel_pte_dup_2_REG <= inner_data_6_7; // @[L2TLB.scala 293:52]
    end else if (3'h6 == _GEN_140) begin // @[L2TLB.scala 293:52]
      cache_io_refill_bits_sel_pte_dup_2_REG <= inner_data_6_6; // @[L2TLB.scala 293:52]
    end else if (3'h5 == _GEN_140) begin // @[L2TLB.scala 293:52]
      cache_io_refill_bits_sel_pte_dup_2_REG <= inner_data_6_5; // @[L2TLB.scala 293:52]
    end else if (3'h4 == _GEN_140) begin // @[L2TLB.scala 293:52]
      cache_io_refill_bits_sel_pte_dup_2_REG <= inner_data_6_4; // @[L2TLB.scala 293:52]
    end else begin
      cache_io_refill_bits_sel_pte_dup_2_REG <= _GEN_144;
    end
    io_perf_0_value_REG <= llptw_io_perf_0_value; // @[PerfCounterUtils.scala 188:35]
    io_perf_0_value_REG_1 <= io_perf_0_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_1_value_REG <= llptw_io_perf_1_value; // @[PerfCounterUtils.scala 188:35]
    io_perf_1_value_REG_1 <= io_perf_1_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_2_value_REG <= llptw_io_perf_2_value; // @[PerfCounterUtils.scala 188:35]
    io_perf_2_value_REG_1 <= io_perf_2_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_3_value_REG <= llptw_io_perf_3_value; // @[PerfCounterUtils.scala 188:35]
    io_perf_3_value_REG_1 <= io_perf_3_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_4_value_REG <= cache_io_perf_0_value; // @[PerfCounterUtils.scala 188:35]
    io_perf_4_value_REG_1 <= io_perf_4_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_5_value_REG <= cache_io_perf_1_value; // @[PerfCounterUtils.scala 188:35]
    io_perf_5_value_REG_1 <= io_perf_5_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_6_value_REG <= cache_io_perf_2_value; // @[PerfCounterUtils.scala 188:35]
    io_perf_6_value_REG_1 <= io_perf_6_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_7_value_REG <= cache_io_perf_3_value; // @[PerfCounterUtils.scala 188:35]
    io_perf_7_value_REG_1 <= io_perf_7_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_8_value_REG <= cache_io_perf_4_value; // @[PerfCounterUtils.scala 188:35]
    io_perf_8_value_REG_1 <= io_perf_8_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_9_value_REG <= cache_io_perf_5_value; // @[PerfCounterUtils.scala 188:35]
    io_perf_9_value_REG_1 <= io_perf_9_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_10_value_REG <= cache_io_perf_6_value; // @[PerfCounterUtils.scala 188:35]
    io_perf_10_value_REG_1 <= io_perf_10_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_11_value_REG <= cache_io_perf_7_value; // @[PerfCounterUtils.scala 188:35]
    io_perf_11_value_REG_1 <= io_perf_11_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_12_value_REG <= ptw_io_perf_0_value; // @[PerfCounterUtils.scala 188:35]
    io_perf_12_value_REG_1 <= io_perf_12_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_13_value_REG <= ptw_io_perf_1_value; // @[PerfCounterUtils.scala 188:35]
    io_perf_13_value_REG_1 <= io_perf_13_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_14_value_REG <= ptw_io_perf_2_value; // @[PerfCounterUtils.scala 188:35]
    io_perf_14_value_REG_1 <= io_perf_14_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_15_value_REG <= ptw_io_perf_3_value; // @[PerfCounterUtils.scala 188:35]
    io_perf_15_value_REG_1 <= io_perf_15_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_16_value_REG <= ptw_io_perf_4_value; // @[PerfCounterUtils.scala 188:35]
    io_perf_16_value_REG_1 <= io_perf_16_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_17_value_REG <= ptw_io_perf_5_value; // @[PerfCounterUtils.scala 188:35]
    io_perf_17_value_REG_1 <= io_perf_17_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_18_value_REG <= ptw_io_perf_6_value; // @[PerfCounterUtils.scala 188:35]
    io_perf_18_value_REG_1 <= io_perf_18_value_REG; // @[PerfCounterUtils.scala 188:27]
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ChiselDB.scala 134:16]
      cnt <= 64'h0;
    end else begin
      cnt <= cnt + 64'h1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[L2TLB.scala 359:24]
      waiting_resp_0 <= 1'h0; // @[L2TLB.scala 360:{37,37}]
    end else if (mem_resp_done) begin
      if (3'h0 == auto_out_d_bits_source) begin
        waiting_resp_0 <= 1'h0;
      end else begin
        waiting_resp_0 <= _GEN_39;
      end
    end else begin
      waiting_resp_0 <= _GEN_39;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[L2TLB.scala 359:24]
      waiting_resp_1 <= 1'h0; // @[L2TLB.scala 360:{37,37}]
    end else if (mem_resp_done) begin
      if (3'h1 == auto_out_d_bits_source) begin
        waiting_resp_1 <= 1'h0;
      end else begin
        waiting_resp_1 <= _GEN_40;
      end
    end else begin
      waiting_resp_1 <= _GEN_40;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[L2TLB.scala 359:24]
      waiting_resp_2 <= 1'h0; // @[L2TLB.scala 360:{37,37}]
    end else if (mem_resp_done) begin
      if (3'h2 == auto_out_d_bits_source) begin
        waiting_resp_2 <= 1'h0;
      end else begin
        waiting_resp_2 <= _GEN_41;
      end
    end else begin
      waiting_resp_2 <= _GEN_41;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[L2TLB.scala 359:24]
      waiting_resp_3 <= 1'h0; // @[L2TLB.scala 360:{37,37}]
    end else if (mem_resp_done) begin
      if (3'h3 == auto_out_d_bits_source) begin
        waiting_resp_3 <= 1'h0;
      end else begin
        waiting_resp_3 <= _GEN_42;
      end
    end else begin
      waiting_resp_3 <= _GEN_42;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[L2TLB.scala 359:24]
      waiting_resp_4 <= 1'h0; // @[L2TLB.scala 360:{37,37}]
    end else if (mem_resp_done) begin
      if (3'h4 == auto_out_d_bits_source) begin
        waiting_resp_4 <= 1'h0;
      end else begin
        waiting_resp_4 <= _GEN_43;
      end
    end else begin
      waiting_resp_4 <= _GEN_43;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[L2TLB.scala 359:24]
      waiting_resp_5 <= 1'h0; // @[L2TLB.scala 360:{37,37}]
    end else if (mem_resp_done) begin
      if (3'h5 == auto_out_d_bits_source) begin
        waiting_resp_5 <= 1'h0;
      end else begin
        waiting_resp_5 <= _GEN_44;
      end
    end else begin
      waiting_resp_5 <= _GEN_44;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[L2TLB.scala 359:24]
      waiting_resp_6 <= 1'h0; // @[L2TLB.scala 360:{37,37}]
    end else if (mem_resp_done) begin
      if (3'h6 == auto_out_d_bits_source) begin
        waiting_resp_6 <= 1'h0;
      end else begin
        waiting_resp_6 <= _GEN_45;
      end
    end else begin
      waiting_resp_6 <= _GEN_45;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[L2TLB.scala 359:24]
      flush_latch_0 <= 1'h0; // @[L2TLB.scala 361:{36,36}]
    end else if (mem_resp_done) begin
      if (3'h0 == auto_out_d_bits_source) begin
        flush_latch_0 <= 1'h0;
      end else begin
        flush_latch_0 <= _GEN_179;
      end
    end else begin
      flush_latch_0 <= _GEN_179;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[L2TLB.scala 359:24]
      flush_latch_1 <= 1'h0; // @[L2TLB.scala 361:{36,36}]
    end else if (mem_resp_done) begin
      if (3'h1 == auto_out_d_bits_source) begin
        flush_latch_1 <= 1'h0;
      end else begin
        flush_latch_1 <= _GEN_180;
      end
    end else begin
      flush_latch_1 <= _GEN_180;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[L2TLB.scala 359:24]
      flush_latch_2 <= 1'h0; // @[L2TLB.scala 361:{36,36}]
    end else if (mem_resp_done) begin
      if (3'h2 == auto_out_d_bits_source) begin
        flush_latch_2 <= 1'h0;
      end else begin
        flush_latch_2 <= _GEN_181;
      end
    end else begin
      flush_latch_2 <= _GEN_181;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[L2TLB.scala 359:24]
      flush_latch_3 <= 1'h0; // @[L2TLB.scala 361:{36,36}]
    end else if (mem_resp_done) begin
      if (3'h3 == auto_out_d_bits_source) begin
        flush_latch_3 <= 1'h0;
      end else begin
        flush_latch_3 <= _GEN_182;
      end
    end else begin
      flush_latch_3 <= _GEN_182;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[L2TLB.scala 359:24]
      flush_latch_4 <= 1'h0; // @[L2TLB.scala 361:{36,36}]
    end else if (mem_resp_done) begin
      if (3'h4 == auto_out_d_bits_source) begin
        flush_latch_4 <= 1'h0;
      end else begin
        flush_latch_4 <= _GEN_183;
      end
    end else begin
      flush_latch_4 <= _GEN_183;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[L2TLB.scala 359:24]
      flush_latch_5 <= 1'h0; // @[L2TLB.scala 361:{36,36}]
    end else if (mem_resp_done) begin
      if (3'h5 == auto_out_d_bits_source) begin
        flush_latch_5 <= 1'h0;
      end else begin
        flush_latch_5 <= _GEN_184;
      end
    end else begin
      flush_latch_5 <= _GEN_184;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[L2TLB.scala 359:24]
      flush_latch_6 <= 1'h0; // @[L2TLB.scala 361:{36,36}]
    end else if (mem_resp_done) begin
      if (3'h6 == auto_out_d_bits_source) begin
        flush_latch_6 <= 1'h0;
      end else begin
        flush_latch_6 <= _GEN_185;
      end
    end else begin
      flush_latch_6 <= _GEN_185;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Edges.scala 234:17]
      counter <= 1'h0; // @[Edges.scala 235:21]
    end else if (auto_out_d_valid) begin // @[Edges.scala 228:27]
      if (first) begin
        counter <= beats1;
      end else begin
        counter <= counter1;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      refill_level_r <= 2'h0; // @[Reg.scala 29:22]
    end else if (_refill_level_T) begin // @[Reg.scala 28:20]
      refill_level_r <= ptw_io_refill_level;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[L2TLB.scala 286:46]
      cache_io_refill_valid_REG <= 1'h0;
    end else begin
      cache_io_refill_valid_REG <= mem_resp_done & _mem_arb_io_out_ready_T & ~_GEN_124;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PageTableCache.scala 94:64]
      cache_io_refill_bits_levelOH_sp_REG <= 1'h0;
    end else begin
      cache_io_refill_bits_levelOH_sp_REG <= (refill_level == 2'h0 | refill_level == 2'h1) & refill_valid;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PageTableCache.scala 95:43]
      cache_io_refill_bits_levelOH_l3_REG <= 1'h0;
    end else begin
      cache_io_refill_bits_levelOH_l3_REG <= refill_level == 2'h2 & refill_valid;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PageTableCache.scala 96:43]
      cache_io_refill_bits_levelOH_l2_REG <= 1'h0;
    end else begin
      cache_io_refill_bits_levelOH_l2_REG <= _cache_io_refill_bits_levelOH_sp_T_1 & refill_valid;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PageTableCache.scala 97:43]
      cache_io_refill_bits_levelOH_l1_REG <= 1'h0;
    end else begin
      cache_io_refill_bits_levelOH_l1_REG <= _cache_io_refill_bits_levelOH_sp_T & refill_valid;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ChiselDB.scala 134:16]
      cnt_1 <= 64'h0;
    end else begin
      cnt_1 <= cnt_1 + 64'h1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ChiselDB.scala 134:16]
      cnt_2 <= 64'h0;
    end else begin
      cnt_2 <= cnt_2 + 64'h1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ChiselDB.scala 134:16]
      cnt_3 <= 64'h0;
    end else begin
      cnt_3 <= cnt_3 + 64'h1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ChiselDB.scala 134:16]
      cnt_4 <= 64'h0;
    end else begin
      cnt_4 <= cnt_4 + 64'h1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ChiselDB.scala 134:16]
      cnt_5 <= 64'h0;
    end else begin
      cnt_5 <= cnt_5 + 64'h1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ChiselDB.scala 134:16]
      cnt_6 <= 64'h0;
    end else begin
      cnt_6 <= cnt_6 + 64'h1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ChiselDB.scala 134:16]
      cnt_7 <= 64'h0;
    end else begin
      cnt_7 <= cnt_7 + 64'h1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ChiselDB.scala 134:16]
      cnt_8 <= 64'h0;
    end else begin
      cnt_8 <= cnt_8 + 64'h1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ChiselDB.scala 134:16]
      cnt_9 <= 64'h0;
    end else begin
      cnt_9 <= cnt_9 + 64'h1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ChiselDB.scala 134:16]
      cnt_10 <= 64'h0;
    end else begin
      cnt_10 <= cnt_10 + 64'h1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ChiselDB.scala 134:16]
      cnt_11 <= 64'h0;
    end else begin
      cnt_11 <= cnt_11 + 64'h1;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  sfence_dup_0_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  sfence_dup_1_valid = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  sfence_dup_2_valid = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  sfence_dup_2_bits_rs1 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  sfence_dup_2_bits_rs2 = _RAND_4[0:0];
  _RAND_5 = {2{`RANDOM}};
  sfence_dup_2_bits_addr = _RAND_5[38:0];
  _RAND_6 = {1{`RANDOM}};
  sfence_dup_2_bits_asid = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  sfence_dup_3_valid = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  sfence_dup_4_valid = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  sfence_dup_5_valid = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  sfence_dup_5_bits_rs1 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  sfence_dup_5_bits_rs2 = _RAND_11[0:0];
  _RAND_12 = {2{`RANDOM}};
  sfence_dup_5_bits_addr = _RAND_12[38:0];
  _RAND_13 = {1{`RANDOM}};
  sfence_dup_6_valid = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  sfence_dup_7_valid = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  csr_dup_0_satp_asid = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  csr_dup_0_satp_changed = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  csr_dup_1_satp_changed = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  csr_dup_2_satp_asid = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  csr_dup_2_satp_changed = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  csr_dup_3_satp_asid = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  csr_dup_3_satp_changed = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  csr_dup_4_satp_asid = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  csr_dup_4_satp_changed = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  csr_dup_5_satp_changed = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  csr_dup_6_satp_asid = _RAND_25[15:0];
  _RAND_26 = {2{`RANDOM}};
  csr_dup_6_satp_ppn = _RAND_26[43:0];
  _RAND_27 = {2{`RANDOM}};
  cnt = _RAND_27[63:0];
  _RAND_28 = {1{`RANDOM}};
  waiting_resp_0 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  waiting_resp_1 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  waiting_resp_2 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  waiting_resp_3 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  waiting_resp_4 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  waiting_resp_5 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  waiting_resp_6 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  flush_latch_0 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  flush_latch_1 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  flush_latch_2 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  flush_latch_3 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  flush_latch_4 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  flush_latch_5 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  flush_latch_6 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  req_addr_low_0 = _RAND_42[2:0];
  _RAND_43 = {1{`RANDOM}};
  req_addr_low_1 = _RAND_43[2:0];
  _RAND_44 = {1{`RANDOM}};
  req_addr_low_2 = _RAND_44[2:0];
  _RAND_45 = {1{`RANDOM}};
  req_addr_low_3 = _RAND_45[2:0];
  _RAND_46 = {1{`RANDOM}};
  req_addr_low_4 = _RAND_46[2:0];
  _RAND_47 = {1{`RANDOM}};
  req_addr_low_5 = _RAND_47[2:0];
  _RAND_48 = {1{`RANDOM}};
  req_addr_low_6 = _RAND_48[2:0];
  _RAND_49 = {8{`RANDOM}};
  refill_data_0 = _RAND_49[255:0];
  _RAND_50 = {8{`RANDOM}};
  refill_data_1 = _RAND_50[255:0];
  _RAND_51 = {1{`RANDOM}};
  counter = _RAND_51[0:0];
  _RAND_52 = {2{`RANDOM}};
  resp_pte_r = _RAND_52[63:0];
  _RAND_53 = {2{`RANDOM}};
  resp_pte_r1 = _RAND_53[63:0];
  _RAND_54 = {2{`RANDOM}};
  resp_pte_r2 = _RAND_54[63:0];
  _RAND_55 = {2{`RANDOM}};
  resp_pte_r3 = _RAND_55[63:0];
  _RAND_56 = {2{`RANDOM}};
  resp_pte_r4 = _RAND_56[63:0];
  _RAND_57 = {2{`RANDOM}};
  resp_pte_r5 = _RAND_57[63:0];
  _RAND_58 = {2{`RANDOM}};
  resp_pte_r6 = _RAND_58[63:0];
  _RAND_59 = {1{`RANDOM}};
  llptw_io_mem_resp_bits_id_r = _RAND_59[2:0];
  _RAND_60 = {1{`RANDOM}};
  refill_level_r = _RAND_60[1:0];
  _RAND_61 = {1{`RANDOM}};
  cache_io_refill_valid_REG = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  cache_io_refill_bits_req_info_dup_0_rvpn = _RAND_62[26:0];
  _RAND_63 = {1{`RANDOM}};
  cache_io_refill_bits_req_info_dup_0_rsource = _RAND_63[1:0];
  _RAND_64 = {1{`RANDOM}};
  cache_io_refill_bits_req_info_dup_1_rvpn = _RAND_64[26:0];
  _RAND_65 = {1{`RANDOM}};
  cache_io_refill_bits_req_info_dup_1_rsource = _RAND_65[1:0];
  _RAND_66 = {1{`RANDOM}};
  cache_io_refill_bits_req_info_dup_2_rvpn = _RAND_66[26:0];
  _RAND_67 = {1{`RANDOM}};
  cache_io_refill_bits_req_info_dup_2_rsource = _RAND_67[1:0];
  _RAND_68 = {1{`RANDOM}};
  cache_io_refill_bits_level_dup_0_r = _RAND_68[1:0];
  _RAND_69 = {1{`RANDOM}};
  cache_io_refill_bits_level_dup_1_r = _RAND_69[1:0];
  _RAND_70 = {1{`RANDOM}};
  cache_io_refill_bits_level_dup_2_r = _RAND_70[1:0];
  _RAND_71 = {1{`RANDOM}};
  cache_io_refill_bits_levelOH_sp_REG = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  cache_io_refill_bits_levelOH_l3_REG = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  cache_io_refill_bits_levelOH_l2_REG = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  cache_io_refill_bits_levelOH_l1_REG = _RAND_74[0:0];
  _RAND_75 = {2{`RANDOM}};
  cache_io_refill_bits_sel_pte_dup_0_REG = _RAND_75[63:0];
  _RAND_76 = {2{`RANDOM}};
  cache_io_refill_bits_sel_pte_dup_1_REG = _RAND_76[63:0];
  _RAND_77 = {2{`RANDOM}};
  cache_io_refill_bits_sel_pte_dup_2_REG = _RAND_77[63:0];
  _RAND_78 = {1{`RANDOM}};
  io_perf_0_value_REG = _RAND_78[5:0];
  _RAND_79 = {1{`RANDOM}};
  io_perf_0_value_REG_1 = _RAND_79[5:0];
  _RAND_80 = {1{`RANDOM}};
  io_perf_1_value_REG = _RAND_80[5:0];
  _RAND_81 = {1{`RANDOM}};
  io_perf_1_value_REG_1 = _RAND_81[5:0];
  _RAND_82 = {1{`RANDOM}};
  io_perf_2_value_REG = _RAND_82[5:0];
  _RAND_83 = {1{`RANDOM}};
  io_perf_2_value_REG_1 = _RAND_83[5:0];
  _RAND_84 = {1{`RANDOM}};
  io_perf_3_value_REG = _RAND_84[5:0];
  _RAND_85 = {1{`RANDOM}};
  io_perf_3_value_REG_1 = _RAND_85[5:0];
  _RAND_86 = {1{`RANDOM}};
  io_perf_4_value_REG = _RAND_86[5:0];
  _RAND_87 = {1{`RANDOM}};
  io_perf_4_value_REG_1 = _RAND_87[5:0];
  _RAND_88 = {1{`RANDOM}};
  io_perf_5_value_REG = _RAND_88[5:0];
  _RAND_89 = {1{`RANDOM}};
  io_perf_5_value_REG_1 = _RAND_89[5:0];
  _RAND_90 = {1{`RANDOM}};
  io_perf_6_value_REG = _RAND_90[5:0];
  _RAND_91 = {1{`RANDOM}};
  io_perf_6_value_REG_1 = _RAND_91[5:0];
  _RAND_92 = {1{`RANDOM}};
  io_perf_7_value_REG = _RAND_92[5:0];
  _RAND_93 = {1{`RANDOM}};
  io_perf_7_value_REG_1 = _RAND_93[5:0];
  _RAND_94 = {1{`RANDOM}};
  io_perf_8_value_REG = _RAND_94[5:0];
  _RAND_95 = {1{`RANDOM}};
  io_perf_8_value_REG_1 = _RAND_95[5:0];
  _RAND_96 = {1{`RANDOM}};
  io_perf_9_value_REG = _RAND_96[5:0];
  _RAND_97 = {1{`RANDOM}};
  io_perf_9_value_REG_1 = _RAND_97[5:0];
  _RAND_98 = {1{`RANDOM}};
  io_perf_10_value_REG = _RAND_98[5:0];
  _RAND_99 = {1{`RANDOM}};
  io_perf_10_value_REG_1 = _RAND_99[5:0];
  _RAND_100 = {1{`RANDOM}};
  io_perf_11_value_REG = _RAND_100[5:0];
  _RAND_101 = {1{`RANDOM}};
  io_perf_11_value_REG_1 = _RAND_101[5:0];
  _RAND_102 = {1{`RANDOM}};
  io_perf_12_value_REG = _RAND_102[5:0];
  _RAND_103 = {1{`RANDOM}};
  io_perf_12_value_REG_1 = _RAND_103[5:0];
  _RAND_104 = {1{`RANDOM}};
  io_perf_13_value_REG = _RAND_104[5:0];
  _RAND_105 = {1{`RANDOM}};
  io_perf_13_value_REG_1 = _RAND_105[5:0];
  _RAND_106 = {1{`RANDOM}};
  io_perf_14_value_REG = _RAND_106[5:0];
  _RAND_107 = {1{`RANDOM}};
  io_perf_14_value_REG_1 = _RAND_107[5:0];
  _RAND_108 = {1{`RANDOM}};
  io_perf_15_value_REG = _RAND_108[5:0];
  _RAND_109 = {1{`RANDOM}};
  io_perf_15_value_REG_1 = _RAND_109[5:0];
  _RAND_110 = {1{`RANDOM}};
  io_perf_16_value_REG = _RAND_110[5:0];
  _RAND_111 = {1{`RANDOM}};
  io_perf_16_value_REG_1 = _RAND_111[5:0];
  _RAND_112 = {1{`RANDOM}};
  io_perf_17_value_REG = _RAND_112[5:0];
  _RAND_113 = {1{`RANDOM}};
  io_perf_17_value_REG_1 = _RAND_113[5:0];
  _RAND_114 = {1{`RANDOM}};
  io_perf_18_value_REG = _RAND_114[5:0];
  _RAND_115 = {1{`RANDOM}};
  io_perf_18_value_REG_1 = _RAND_115[5:0];
  _RAND_116 = {2{`RANDOM}};
  cnt_1 = _RAND_116[63:0];
  _RAND_117 = {2{`RANDOM}};
  cnt_2 = _RAND_117[63:0];
  _RAND_118 = {2{`RANDOM}};
  cnt_3 = _RAND_118[63:0];
  _RAND_119 = {2{`RANDOM}};
  cnt_4 = _RAND_119[63:0];
  _RAND_120 = {2{`RANDOM}};
  cnt_5 = _RAND_120[63:0];
  _RAND_121 = {2{`RANDOM}};
  cnt_6 = _RAND_121[63:0];
  _RAND_122 = {2{`RANDOM}};
  cnt_7 = _RAND_122[63:0];
  _RAND_123 = {2{`RANDOM}};
  cnt_8 = _RAND_123[63:0];
  _RAND_124 = {2{`RANDOM}};
  cnt_9 = _RAND_124[63:0];
  _RAND_125 = {2{`RANDOM}};
  cnt_10 = _RAND_125[63:0];
  _RAND_126 = {2{`RANDOM}};
  cnt_11 = _RAND_126[63:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    cnt = 64'h0;
  end
  if (reset) begin
    waiting_resp_0 = 1'h0;
  end
  if (reset) begin
    waiting_resp_1 = 1'h0;
  end
  if (reset) begin
    waiting_resp_2 = 1'h0;
  end
  if (reset) begin
    waiting_resp_3 = 1'h0;
  end
  if (reset) begin
    waiting_resp_4 = 1'h0;
  end
  if (reset) begin
    waiting_resp_5 = 1'h0;
  end
  if (reset) begin
    waiting_resp_6 = 1'h0;
  end
  if (reset) begin
    flush_latch_0 = 1'h0;
  end
  if (reset) begin
    flush_latch_1 = 1'h0;
  end
  if (reset) begin
    flush_latch_2 = 1'h0;
  end
  if (reset) begin
    flush_latch_3 = 1'h0;
  end
  if (reset) begin
    flush_latch_4 = 1'h0;
  end
  if (reset) begin
    flush_latch_5 = 1'h0;
  end
  if (reset) begin
    flush_latch_6 = 1'h0;
  end
  if (reset) begin
    counter = 1'h0;
  end
  if (reset) begin
    refill_level_r = 2'h0;
  end
  if (reset) begin
    cache_io_refill_valid_REG = 1'h0;
  end
  if (reset) begin
    cache_io_refill_bits_levelOH_sp_REG = 1'h0;
  end
  if (reset) begin
    cache_io_refill_bits_levelOH_l3_REG = 1'h0;
  end
  if (reset) begin
    cache_io_refill_bits_levelOH_l2_REG = 1'h0;
  end
  if (reset) begin
    cache_io_refill_bits_levelOH_l1_REG = 1'h0;
  end
  if (reset) begin
    cnt_1 = 64'h0;
  end
  if (reset) begin
    cnt_2 = 64'h0;
  end
  if (reset) begin
    cnt_3 = 64'h0;
  end
  if (reset) begin
    cnt_4 = 64'h0;
  end
  if (reset) begin
    cnt_5 = 64'h0;
  end
  if (reset) begin
    cnt_6 = 64'h0;
  end
  if (reset) begin
    cnt_7 = 64'h0;
  end
  if (reset) begin
    cnt_8 = 64'h0;
  end
  if (reset) begin
    cnt_9 = 64'h0;
  end
  if (reset) begin
    cnt_10 = 64'h0;
  end
  if (reset) begin
    cnt_11 = 64'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule

