module ArrayMulDataModule(
  input          clock,
  input  [64:0]  io_a,
  input  [64:0]  io_b,
  input          io_regEnables_0,
  input          io_regEnables_1,
  output [129:0] io_result
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_786;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_789;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_793;
  reg [31:0] _RAND_794;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [31:0] _RAND_798;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_801;
  reg [31:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_804;
  reg [31:0] _RAND_805;
  reg [31:0] _RAND_806;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [31:0] _RAND_810;
  reg [31:0] _RAND_811;
  reg [31:0] _RAND_812;
  reg [31:0] _RAND_813;
  reg [31:0] _RAND_814;
  reg [31:0] _RAND_815;
  reg [31:0] _RAND_816;
  reg [31:0] _RAND_817;
  reg [31:0] _RAND_818;
  reg [31:0] _RAND_819;
  reg [31:0] _RAND_820;
  reg [31:0] _RAND_821;
  reg [31:0] _RAND_822;
  reg [31:0] _RAND_823;
  reg [31:0] _RAND_824;
  reg [31:0] _RAND_825;
  reg [31:0] _RAND_826;
  reg [31:0] _RAND_827;
  reg [31:0] _RAND_828;
  reg [31:0] _RAND_829;
  reg [31:0] _RAND_830;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
  reg [31:0] _RAND_834;
  reg [31:0] _RAND_835;
  reg [31:0] _RAND_836;
  reg [31:0] _RAND_837;
  reg [31:0] _RAND_838;
  reg [31:0] _RAND_839;
  reg [31:0] _RAND_840;
  reg [31:0] _RAND_841;
  reg [31:0] _RAND_842;
  reg [31:0] _RAND_843;
  reg [31:0] _RAND_844;
  reg [31:0] _RAND_845;
  reg [31:0] _RAND_846;
  reg [31:0] _RAND_847;
  reg [31:0] _RAND_848;
  reg [31:0] _RAND_849;
  reg [31:0] _RAND_850;
  reg [31:0] _RAND_851;
  reg [31:0] _RAND_852;
  reg [31:0] _RAND_853;
  reg [31:0] _RAND_854;
  reg [31:0] _RAND_855;
  reg [31:0] _RAND_856;
  reg [31:0] _RAND_857;
  reg [31:0] _RAND_858;
  reg [31:0] _RAND_859;
  reg [31:0] _RAND_860;
  reg [31:0] _RAND_861;
  reg [31:0] _RAND_862;
  reg [31:0] _RAND_863;
  reg [31:0] _RAND_864;
  reg [31:0] _RAND_865;
  reg [31:0] _RAND_866;
  reg [31:0] _RAND_867;
  reg [31:0] _RAND_868;
  reg [31:0] _RAND_869;
  reg [31:0] _RAND_870;
  reg [31:0] _RAND_871;
  reg [31:0] _RAND_872;
  reg [31:0] _RAND_873;
  reg [31:0] _RAND_874;
  reg [31:0] _RAND_875;
  reg [31:0] _RAND_876;
  reg [31:0] _RAND_877;
  reg [31:0] _RAND_878;
  reg [31:0] _RAND_879;
  reg [31:0] _RAND_880;
  reg [31:0] _RAND_881;
  reg [31:0] _RAND_882;
  reg [31:0] _RAND_883;
  reg [31:0] _RAND_884;
  reg [31:0] _RAND_885;
  reg [31:0] _RAND_886;
  reg [31:0] _RAND_887;
  reg [31:0] _RAND_888;
  reg [31:0] _RAND_889;
  reg [31:0] _RAND_890;
  reg [31:0] _RAND_891;
  reg [31:0] _RAND_892;
  reg [31:0] _RAND_893;
  reg [31:0] _RAND_894;
  reg [31:0] _RAND_895;
  reg [31:0] _RAND_896;
  reg [31:0] _RAND_897;
  reg [31:0] _RAND_898;
  reg [31:0] _RAND_899;
  reg [31:0] _RAND_900;
  reg [31:0] _RAND_901;
  reg [31:0] _RAND_902;
  reg [31:0] _RAND_903;
  reg [31:0] _RAND_904;
  reg [31:0] _RAND_905;
  reg [31:0] _RAND_906;
  reg [31:0] _RAND_907;
  reg [31:0] _RAND_908;
  reg [31:0] _RAND_909;
  reg [31:0] _RAND_910;
  reg [31:0] _RAND_911;
  reg [31:0] _RAND_912;
  reg [31:0] _RAND_913;
  reg [31:0] _RAND_914;
  reg [31:0] _RAND_915;
  reg [31:0] _RAND_916;
  reg [31:0] _RAND_917;
  reg [31:0] _RAND_918;
  reg [31:0] _RAND_919;
  reg [31:0] _RAND_920;
  reg [31:0] _RAND_921;
  reg [31:0] _RAND_922;
  reg [31:0] _RAND_923;
  reg [31:0] _RAND_924;
  reg [31:0] _RAND_925;
  reg [31:0] _RAND_926;
  reg [31:0] _RAND_927;
  reg [31:0] _RAND_928;
  reg [31:0] _RAND_929;
  reg [31:0] _RAND_930;
  reg [31:0] _RAND_931;
  reg [31:0] _RAND_932;
  reg [31:0] _RAND_933;
  reg [31:0] _RAND_934;
  reg [31:0] _RAND_935;
  reg [31:0] _RAND_936;
  reg [31:0] _RAND_937;
  reg [31:0] _RAND_938;
  reg [31:0] _RAND_939;
  reg [31:0] _RAND_940;
  reg [31:0] _RAND_941;
  reg [31:0] _RAND_942;
  reg [31:0] _RAND_943;
  reg [31:0] _RAND_944;
  reg [31:0] _RAND_945;
  reg [31:0] _RAND_946;
  reg [31:0] _RAND_947;
  reg [31:0] _RAND_948;
  reg [31:0] _RAND_949;
  reg [31:0] _RAND_950;
  reg [31:0] _RAND_951;
  reg [31:0] _RAND_952;
  reg [31:0] _RAND_953;
  reg [31:0] _RAND_954;
  reg [31:0] _RAND_955;
  reg [31:0] _RAND_956;
  reg [31:0] _RAND_957;
  reg [31:0] _RAND_958;
  reg [31:0] _RAND_959;
  reg [31:0] _RAND_960;
  reg [31:0] _RAND_961;
  reg [31:0] _RAND_962;
  reg [31:0] _RAND_963;
  reg [31:0] _RAND_964;
  reg [31:0] _RAND_965;
  reg [31:0] _RAND_966;
  reg [31:0] _RAND_967;
  reg [31:0] _RAND_968;
  reg [31:0] _RAND_969;
  reg [31:0] _RAND_970;
  reg [31:0] _RAND_971;
  reg [31:0] _RAND_972;
  reg [31:0] _RAND_973;
  reg [31:0] _RAND_974;
  reg [31:0] _RAND_975;
  reg [31:0] _RAND_976;
  reg [31:0] _RAND_977;
  reg [31:0] _RAND_978;
  reg [31:0] _RAND_979;
  reg [31:0] _RAND_980;
  reg [31:0] _RAND_981;
  reg [31:0] _RAND_982;
  reg [31:0] _RAND_983;
  reg [31:0] _RAND_984;
  reg [31:0] _RAND_985;
  reg [31:0] _RAND_986;
  reg [31:0] _RAND_987;
  reg [31:0] _RAND_988;
  reg [31:0] _RAND_989;
  reg [31:0] _RAND_990;
  reg [31:0] _RAND_991;
  reg [31:0] _RAND_992;
  reg [31:0] _RAND_993;
  reg [31:0] _RAND_994;
  reg [31:0] _RAND_995;
  reg [31:0] _RAND_996;
  reg [31:0] _RAND_997;
  reg [31:0] _RAND_998;
  reg [31:0] _RAND_999;
  reg [31:0] _RAND_1000;
  reg [31:0] _RAND_1001;
  reg [31:0] _RAND_1002;
  reg [31:0] _RAND_1003;
  reg [31:0] _RAND_1004;
  reg [31:0] _RAND_1005;
  reg [31:0] _RAND_1006;
  reg [31:0] _RAND_1007;
  reg [31:0] _RAND_1008;
  reg [31:0] _RAND_1009;
  reg [31:0] _RAND_1010;
  reg [31:0] _RAND_1011;
  reg [31:0] _RAND_1012;
  reg [31:0] _RAND_1013;
  reg [31:0] _RAND_1014;
  reg [31:0] _RAND_1015;
  reg [31:0] _RAND_1016;
  reg [31:0] _RAND_1017;
  reg [31:0] _RAND_1018;
  reg [31:0] _RAND_1019;
  reg [31:0] _RAND_1020;
  reg [31:0] _RAND_1021;
  reg [31:0] _RAND_1022;
  reg [31:0] _RAND_1023;
  reg [31:0] _RAND_1024;
  reg [31:0] _RAND_1025;
  reg [31:0] _RAND_1026;
  reg [31:0] _RAND_1027;
  reg [31:0] _RAND_1028;
  reg [31:0] _RAND_1029;
  reg [31:0] _RAND_1030;
  reg [31:0] _RAND_1031;
  reg [31:0] _RAND_1032;
  reg [31:0] _RAND_1033;
  reg [31:0] _RAND_1034;
  reg [31:0] _RAND_1035;
  reg [31:0] _RAND_1036;
  reg [31:0] _RAND_1037;
  reg [31:0] _RAND_1038;
  reg [31:0] _RAND_1039;
  reg [31:0] _RAND_1040;
  reg [31:0] _RAND_1041;
  reg [31:0] _RAND_1042;
  reg [31:0] _RAND_1043;
  reg [31:0] _RAND_1044;
  reg [31:0] _RAND_1045;
  reg [31:0] _RAND_1046;
  reg [31:0] _RAND_1047;
  reg [31:0] _RAND_1048;
  reg [31:0] _RAND_1049;
  reg [31:0] _RAND_1050;
  reg [31:0] _RAND_1051;
  reg [31:0] _RAND_1052;
  reg [31:0] _RAND_1053;
  reg [31:0] _RAND_1054;
  reg [31:0] _RAND_1055;
  reg [31:0] _RAND_1056;
  reg [31:0] _RAND_1057;
  reg [31:0] _RAND_1058;
  reg [31:0] _RAND_1059;
  reg [31:0] _RAND_1060;
  reg [31:0] _RAND_1061;
  reg [31:0] _RAND_1062;
  reg [31:0] _RAND_1063;
  reg [31:0] _RAND_1064;
  reg [31:0] _RAND_1065;
  reg [31:0] _RAND_1066;
  reg [31:0] _RAND_1067;
  reg [31:0] _RAND_1068;
  reg [31:0] _RAND_1069;
  reg [31:0] _RAND_1070;
  reg [31:0] _RAND_1071;
  reg [31:0] _RAND_1072;
  reg [31:0] _RAND_1073;
  reg [31:0] _RAND_1074;
  reg [31:0] _RAND_1075;
  reg [31:0] _RAND_1076;
  reg [31:0] _RAND_1077;
  reg [31:0] _RAND_1078;
  reg [31:0] _RAND_1079;
  reg [31:0] _RAND_1080;
  reg [31:0] _RAND_1081;
  reg [31:0] _RAND_1082;
  reg [31:0] _RAND_1083;
  reg [31:0] _RAND_1084;
  reg [31:0] _RAND_1085;
  reg [31:0] _RAND_1086;
  reg [31:0] _RAND_1087;
  reg [31:0] _RAND_1088;
  reg [31:0] _RAND_1089;
  reg [31:0] _RAND_1090;
  reg [31:0] _RAND_1091;
  reg [31:0] _RAND_1092;
  reg [31:0] _RAND_1093;
  reg [31:0] _RAND_1094;
  reg [31:0] _RAND_1095;
  reg [31:0] _RAND_1096;
  reg [31:0] _RAND_1097;
  reg [31:0] _RAND_1098;
  reg [31:0] _RAND_1099;
  reg [31:0] _RAND_1100;
  reg [31:0] _RAND_1101;
  reg [31:0] _RAND_1102;
  reg [31:0] _RAND_1103;
  reg [31:0] _RAND_1104;
  reg [31:0] _RAND_1105;
  reg [31:0] _RAND_1106;
  reg [31:0] _RAND_1107;
  reg [31:0] _RAND_1108;
  reg [31:0] _RAND_1109;
  reg [31:0] _RAND_1110;
  reg [31:0] _RAND_1111;
  reg [31:0] _RAND_1112;
  reg [31:0] _RAND_1113;
  reg [31:0] _RAND_1114;
  reg [31:0] _RAND_1115;
  reg [31:0] _RAND_1116;
  reg [31:0] _RAND_1117;
  reg [31:0] _RAND_1118;
  reg [31:0] _RAND_1119;
  reg [31:0] _RAND_1120;
  reg [31:0] _RAND_1121;
  reg [31:0] _RAND_1122;
  reg [31:0] _RAND_1123;
  reg [31:0] _RAND_1124;
  reg [31:0] _RAND_1125;
  reg [31:0] _RAND_1126;
  reg [31:0] _RAND_1127;
  reg [31:0] _RAND_1128;
  reg [31:0] _RAND_1129;
  reg [31:0] _RAND_1130;
  reg [31:0] _RAND_1131;
  reg [31:0] _RAND_1132;
  reg [31:0] _RAND_1133;
  reg [31:0] _RAND_1134;
  reg [31:0] _RAND_1135;
  reg [31:0] _RAND_1136;
  reg [31:0] _RAND_1137;
  reg [31:0] _RAND_1138;
  reg [31:0] _RAND_1139;
  reg [31:0] _RAND_1140;
  reg [31:0] _RAND_1141;
  reg [31:0] _RAND_1142;
  reg [31:0] _RAND_1143;
  reg [31:0] _RAND_1144;
  reg [31:0] _RAND_1145;
  reg [31:0] _RAND_1146;
  reg [31:0] _RAND_1147;
  reg [31:0] _RAND_1148;
  reg [31:0] _RAND_1149;
  reg [31:0] _RAND_1150;
  reg [31:0] _RAND_1151;
  reg [31:0] _RAND_1152;
  reg [31:0] _RAND_1153;
  reg [31:0] _RAND_1154;
  reg [31:0] _RAND_1155;
  reg [31:0] _RAND_1156;
  reg [31:0] _RAND_1157;
  reg [31:0] _RAND_1158;
  reg [31:0] _RAND_1159;
  reg [31:0] _RAND_1160;
  reg [31:0] _RAND_1161;
  reg [31:0] _RAND_1162;
  reg [31:0] _RAND_1163;
  reg [31:0] _RAND_1164;
  reg [31:0] _RAND_1165;
  reg [31:0] _RAND_1166;
  reg [31:0] _RAND_1167;
  reg [31:0] _RAND_1168;
  reg [31:0] _RAND_1169;
  reg [31:0] _RAND_1170;
  reg [31:0] _RAND_1171;
  reg [31:0] _RAND_1172;
  reg [31:0] _RAND_1173;
  reg [31:0] _RAND_1174;
  reg [31:0] _RAND_1175;
  reg [31:0] _RAND_1176;
  reg [31:0] _RAND_1177;
  reg [31:0] _RAND_1178;
  reg [31:0] _RAND_1179;
  reg [31:0] _RAND_1180;
  reg [31:0] _RAND_1181;
  reg [31:0] _RAND_1182;
  reg [31:0] _RAND_1183;
  reg [31:0] _RAND_1184;
  reg [31:0] _RAND_1185;
  reg [31:0] _RAND_1186;
  reg [31:0] _RAND_1187;
  reg [31:0] _RAND_1188;
  reg [31:0] _RAND_1189;
  reg [31:0] _RAND_1190;
  reg [31:0] _RAND_1191;
  reg [31:0] _RAND_1192;
  reg [31:0] _RAND_1193;
  reg [31:0] _RAND_1194;
  reg [31:0] _RAND_1195;
  reg [31:0] _RAND_1196;
  reg [31:0] _RAND_1197;
  reg [31:0] _RAND_1198;
  reg [31:0] _RAND_1199;
  reg [31:0] _RAND_1200;
  reg [31:0] _RAND_1201;
  reg [31:0] _RAND_1202;
  reg [31:0] _RAND_1203;
  reg [31:0] _RAND_1204;
  reg [31:0] _RAND_1205;
  reg [31:0] _RAND_1206;
  reg [31:0] _RAND_1207;
  reg [31:0] _RAND_1208;
  reg [31:0] _RAND_1209;
  reg [31:0] _RAND_1210;
  reg [31:0] _RAND_1211;
  reg [31:0] _RAND_1212;
  reg [31:0] _RAND_1213;
  reg [31:0] _RAND_1214;
  reg [31:0] _RAND_1215;
  reg [31:0] _RAND_1216;
  reg [31:0] _RAND_1217;
  reg [31:0] _RAND_1218;
  reg [31:0] _RAND_1219;
  reg [31:0] _RAND_1220;
  reg [31:0] _RAND_1221;
  reg [31:0] _RAND_1222;
  reg [31:0] _RAND_1223;
  reg [31:0] _RAND_1224;
  reg [31:0] _RAND_1225;
  reg [31:0] _RAND_1226;
  reg [31:0] _RAND_1227;
  reg [31:0] _RAND_1228;
  reg [31:0] _RAND_1229;
  reg [31:0] _RAND_1230;
  reg [31:0] _RAND_1231;
  reg [31:0] _RAND_1232;
  reg [31:0] _RAND_1233;
  reg [31:0] _RAND_1234;
  reg [31:0] _RAND_1235;
  reg [31:0] _RAND_1236;
  reg [31:0] _RAND_1237;
  reg [31:0] _RAND_1238;
  reg [31:0] _RAND_1239;
  reg [31:0] _RAND_1240;
  reg [31:0] _RAND_1241;
  reg [31:0] _RAND_1242;
  reg [31:0] _RAND_1243;
  reg [31:0] _RAND_1244;
  reg [31:0] _RAND_1245;
  reg [31:0] _RAND_1246;
  reg [31:0] _RAND_1247;
  reg [31:0] _RAND_1248;
  reg [31:0] _RAND_1249;
  reg [31:0] _RAND_1250;
  reg [31:0] _RAND_1251;
  reg [31:0] _RAND_1252;
  reg [31:0] _RAND_1253;
  reg [31:0] _RAND_1254;
  reg [31:0] _RAND_1255;
  reg [31:0] _RAND_1256;
  reg [31:0] _RAND_1257;
  reg [31:0] _RAND_1258;
  reg [31:0] _RAND_1259;
  reg [31:0] _RAND_1260;
  reg [31:0] _RAND_1261;
  reg [31:0] _RAND_1262;
  reg [31:0] _RAND_1263;
  reg [31:0] _RAND_1264;
  reg [31:0] _RAND_1265;
  reg [31:0] _RAND_1266;
  reg [31:0] _RAND_1267;
  reg [31:0] _RAND_1268;
  reg [31:0] _RAND_1269;
  reg [31:0] _RAND_1270;
  reg [31:0] _RAND_1271;
  reg [31:0] _RAND_1272;
  reg [31:0] _RAND_1273;
  reg [31:0] _RAND_1274;
  reg [31:0] _RAND_1275;
  reg [31:0] _RAND_1276;
  reg [31:0] _RAND_1277;
  reg [31:0] _RAND_1278;
  reg [31:0] _RAND_1279;
  reg [31:0] _RAND_1280;
  reg [31:0] _RAND_1281;
  reg [31:0] _RAND_1282;
  reg [31:0] _RAND_1283;
  reg [31:0] _RAND_1284;
  reg [31:0] _RAND_1285;
  reg [31:0] _RAND_1286;
  reg [31:0] _RAND_1287;
  reg [31:0] _RAND_1288;
  reg [31:0] _RAND_1289;
  reg [31:0] _RAND_1290;
  reg [31:0] _RAND_1291;
  reg [31:0] _RAND_1292;
  reg [31:0] _RAND_1293;
  reg [31:0] _RAND_1294;
  reg [31:0] _RAND_1295;
  reg [31:0] _RAND_1296;
  reg [31:0] _RAND_1297;
  reg [31:0] _RAND_1298;
  reg [31:0] _RAND_1299;
  reg [31:0] _RAND_1300;
  reg [31:0] _RAND_1301;
  reg [31:0] _RAND_1302;
  reg [31:0] _RAND_1303;
  reg [31:0] _RAND_1304;
  reg [31:0] _RAND_1305;
  reg [31:0] _RAND_1306;
  reg [31:0] _RAND_1307;
  reg [31:0] _RAND_1308;
  reg [31:0] _RAND_1309;
  reg [31:0] _RAND_1310;
  reg [31:0] _RAND_1311;
  reg [31:0] _RAND_1312;
  reg [31:0] _RAND_1313;
  reg [31:0] _RAND_1314;
  reg [31:0] _RAND_1315;
  reg [31:0] _RAND_1316;
  reg [31:0] _RAND_1317;
  reg [31:0] _RAND_1318;
  reg [31:0] _RAND_1319;
  reg [31:0] _RAND_1320;
  reg [31:0] _RAND_1321;
  reg [31:0] _RAND_1322;
  reg [31:0] _RAND_1323;
  reg [31:0] _RAND_1324;
  reg [31:0] _RAND_1325;
  reg [31:0] _RAND_1326;
  reg [31:0] _RAND_1327;
  reg [31:0] _RAND_1328;
  reg [31:0] _RAND_1329;
  reg [31:0] _RAND_1330;
  reg [31:0] _RAND_1331;
  reg [31:0] _RAND_1332;
  reg [31:0] _RAND_1333;
  reg [31:0] _RAND_1334;
  reg [31:0] _RAND_1335;
  reg [31:0] _RAND_1336;
  reg [31:0] _RAND_1337;
  reg [31:0] _RAND_1338;
  reg [31:0] _RAND_1339;
  reg [31:0] _RAND_1340;
  reg [31:0] _RAND_1341;
  reg [31:0] _RAND_1342;
  reg [31:0] _RAND_1343;
  reg [31:0] _RAND_1344;
  reg [31:0] _RAND_1345;
  reg [31:0] _RAND_1346;
  reg [31:0] _RAND_1347;
  reg [31:0] _RAND_1348;
  reg [31:0] _RAND_1349;
  reg [31:0] _RAND_1350;
  reg [31:0] _RAND_1351;
  reg [31:0] _RAND_1352;
  reg [31:0] _RAND_1353;
  reg [31:0] _RAND_1354;
  reg [31:0] _RAND_1355;
  reg [31:0] _RAND_1356;
  reg [31:0] _RAND_1357;
  reg [31:0] _RAND_1358;
  reg [31:0] _RAND_1359;
  reg [31:0] _RAND_1360;
  reg [31:0] _RAND_1361;
  reg [31:0] _RAND_1362;
  reg [31:0] _RAND_1363;
  reg [31:0] _RAND_1364;
  reg [31:0] _RAND_1365;
  reg [31:0] _RAND_1366;
  reg [31:0] _RAND_1367;
  reg [31:0] _RAND_1368;
  reg [31:0] _RAND_1369;
  reg [31:0] _RAND_1370;
  reg [31:0] _RAND_1371;
  reg [31:0] _RAND_1372;
  reg [31:0] _RAND_1373;
  reg [31:0] _RAND_1374;
  reg [31:0] _RAND_1375;
  reg [31:0] _RAND_1376;
  reg [31:0] _RAND_1377;
  reg [31:0] _RAND_1378;
  reg [31:0] _RAND_1379;
  reg [31:0] _RAND_1380;
  reg [31:0] _RAND_1381;
  reg [31:0] _RAND_1382;
  reg [31:0] _RAND_1383;
  reg [31:0] _RAND_1384;
  reg [31:0] _RAND_1385;
  reg [31:0] _RAND_1386;
  reg [31:0] _RAND_1387;
  reg [31:0] _RAND_1388;
  reg [31:0] _RAND_1389;
  reg [31:0] _RAND_1390;
  reg [31:0] _RAND_1391;
  reg [31:0] _RAND_1392;
  reg [31:0] _RAND_1393;
  reg [31:0] _RAND_1394;
  reg [31:0] _RAND_1395;
  reg [31:0] _RAND_1396;
  reg [31:0] _RAND_1397;
  reg [31:0] _RAND_1398;
  reg [31:0] _RAND_1399;
  reg [31:0] _RAND_1400;
  reg [31:0] _RAND_1401;
  reg [31:0] _RAND_1402;
  reg [31:0] _RAND_1403;
  reg [31:0] _RAND_1404;
  reg [31:0] _RAND_1405;
  reg [31:0] _RAND_1406;
  reg [31:0] _RAND_1407;
  reg [31:0] _RAND_1408;
  reg [31:0] _RAND_1409;
  reg [31:0] _RAND_1410;
  reg [31:0] _RAND_1411;
  reg [31:0] _RAND_1412;
  reg [31:0] _RAND_1413;
  reg [31:0] _RAND_1414;
  reg [31:0] _RAND_1415;
  reg [31:0] _RAND_1416;
  reg [31:0] _RAND_1417;
  reg [31:0] _RAND_1418;
  reg [31:0] _RAND_1419;
  reg [31:0] _RAND_1420;
  reg [31:0] _RAND_1421;
  reg [31:0] _RAND_1422;
  reg [31:0] _RAND_1423;
  reg [31:0] _RAND_1424;
  reg [31:0] _RAND_1425;
  reg [31:0] _RAND_1426;
  reg [31:0] _RAND_1427;
  reg [31:0] _RAND_1428;
  reg [31:0] _RAND_1429;
  reg [31:0] _RAND_1430;
  reg [31:0] _RAND_1431;
  reg [31:0] _RAND_1432;
  reg [31:0] _RAND_1433;
  reg [31:0] _RAND_1434;
  reg [31:0] _RAND_1435;
  reg [31:0] _RAND_1436;
  reg [31:0] _RAND_1437;
  reg [31:0] _RAND_1438;
  reg [31:0] _RAND_1439;
  reg [31:0] _RAND_1440;
  reg [31:0] _RAND_1441;
  reg [31:0] _RAND_1442;
  reg [31:0] _RAND_1443;
  reg [31:0] _RAND_1444;
  reg [31:0] _RAND_1445;
  reg [31:0] _RAND_1446;
  reg [31:0] _RAND_1447;
  reg [31:0] _RAND_1448;
  reg [31:0] _RAND_1449;
  reg [31:0] _RAND_1450;
  reg [31:0] _RAND_1451;
  reg [31:0] _RAND_1452;
  reg [31:0] _RAND_1453;
  reg [31:0] _RAND_1454;
  reg [31:0] _RAND_1455;
  reg [31:0] _RAND_1456;
  reg [31:0] _RAND_1457;
  reg [31:0] _RAND_1458;
  reg [31:0] _RAND_1459;
  reg [31:0] _RAND_1460;
  reg [31:0] _RAND_1461;
  reg [31:0] _RAND_1462;
  reg [31:0] _RAND_1463;
  reg [31:0] _RAND_1464;
  reg [31:0] _RAND_1465;
  reg [31:0] _RAND_1466;
  reg [31:0] _RAND_1467;
  reg [31:0] _RAND_1468;
  reg [31:0] _RAND_1469;
  reg [31:0] _RAND_1470;
  reg [31:0] _RAND_1471;
  reg [31:0] _RAND_1472;
  reg [31:0] _RAND_1473;
  reg [31:0] _RAND_1474;
  reg [31:0] _RAND_1475;
  reg [31:0] _RAND_1476;
  reg [31:0] _RAND_1477;
  reg [31:0] _RAND_1478;
  reg [31:0] _RAND_1479;
  reg [31:0] _RAND_1480;
  reg [31:0] _RAND_1481;
  reg [31:0] _RAND_1482;
  reg [31:0] _RAND_1483;
  reg [31:0] _RAND_1484;
  reg [31:0] _RAND_1485;
  reg [31:0] _RAND_1486;
  reg [31:0] _RAND_1487;
  reg [31:0] _RAND_1488;
  reg [31:0] _RAND_1489;
  reg [31:0] _RAND_1490;
  reg [31:0] _RAND_1491;
  reg [31:0] _RAND_1492;
  reg [31:0] _RAND_1493;
  reg [31:0] _RAND_1494;
  reg [31:0] _RAND_1495;
  reg [31:0] _RAND_1496;
  reg [31:0] _RAND_1497;
  reg [31:0] _RAND_1498;
  reg [31:0] _RAND_1499;
  reg [31:0] _RAND_1500;
  reg [31:0] _RAND_1501;
  reg [31:0] _RAND_1502;
  reg [31:0] _RAND_1503;
  reg [31:0] _RAND_1504;
  reg [31:0] _RAND_1505;
  reg [31:0] _RAND_1506;
  reg [31:0] _RAND_1507;
  reg [31:0] _RAND_1508;
  reg [31:0] _RAND_1509;
  reg [31:0] _RAND_1510;
  reg [31:0] _RAND_1511;
  reg [31:0] _RAND_1512;
  reg [31:0] _RAND_1513;
  reg [31:0] _RAND_1514;
  reg [31:0] _RAND_1515;
  reg [31:0] _RAND_1516;
  reg [31:0] _RAND_1517;
  reg [31:0] _RAND_1518;
  reg [31:0] _RAND_1519;
  reg [31:0] _RAND_1520;
  reg [31:0] _RAND_1521;
  reg [31:0] _RAND_1522;
  reg [31:0] _RAND_1523;
  reg [31:0] _RAND_1524;
  reg [31:0] _RAND_1525;
  reg [31:0] _RAND_1526;
  reg [31:0] _RAND_1527;
  reg [31:0] _RAND_1528;
  reg [31:0] _RAND_1529;
  reg [31:0] _RAND_1530;
  reg [31:0] _RAND_1531;
  reg [31:0] _RAND_1532;
  reg [31:0] _RAND_1533;
  reg [31:0] _RAND_1534;
  reg [31:0] _RAND_1535;
  reg [31:0] _RAND_1536;
  reg [31:0] _RAND_1537;
  reg [31:0] _RAND_1538;
  reg [31:0] _RAND_1539;
  reg [31:0] _RAND_1540;
  reg [31:0] _RAND_1541;
  reg [31:0] _RAND_1542;
  reg [31:0] _RAND_1543;
  reg [31:0] _RAND_1544;
  reg [31:0] _RAND_1545;
  reg [31:0] _RAND_1546;
  reg [31:0] _RAND_1547;
  reg [31:0] _RAND_1548;
  reg [31:0] _RAND_1549;
  reg [31:0] _RAND_1550;
  reg [31:0] _RAND_1551;
  reg [31:0] _RAND_1552;
  reg [31:0] _RAND_1553;
  reg [31:0] _RAND_1554;
  reg [31:0] _RAND_1555;
  reg [31:0] _RAND_1556;
  reg [31:0] _RAND_1557;
  reg [31:0] _RAND_1558;
  reg [31:0] _RAND_1559;
  reg [31:0] _RAND_1560;
  reg [31:0] _RAND_1561;
  reg [31:0] _RAND_1562;
  reg [31:0] _RAND_1563;
  reg [31:0] _RAND_1564;
  reg [31:0] _RAND_1565;
  reg [31:0] _RAND_1566;
  reg [31:0] _RAND_1567;
  reg [31:0] _RAND_1568;
  reg [31:0] _RAND_1569;
  reg [31:0] _RAND_1570;
  reg [31:0] _RAND_1571;
  reg [31:0] _RAND_1572;
  reg [31:0] _RAND_1573;
  reg [31:0] _RAND_1574;
  reg [31:0] _RAND_1575;
  reg [31:0] _RAND_1576;
  reg [31:0] _RAND_1577;
  reg [31:0] _RAND_1578;
  reg [31:0] _RAND_1579;
  reg [31:0] _RAND_1580;
  reg [31:0] _RAND_1581;
  reg [31:0] _RAND_1582;
  reg [31:0] _RAND_1583;
  reg [31:0] _RAND_1584;
  reg [31:0] _RAND_1585;
  reg [31:0] _RAND_1586;
  reg [31:0] _RAND_1587;
  reg [31:0] _RAND_1588;
  reg [31:0] _RAND_1589;
  reg [31:0] _RAND_1590;
  reg [31:0] _RAND_1591;
  reg [31:0] _RAND_1592;
  reg [31:0] _RAND_1593;
  reg [31:0] _RAND_1594;
  reg [31:0] _RAND_1595;
  reg [31:0] _RAND_1596;
  reg [31:0] _RAND_1597;
  reg [31:0] _RAND_1598;
  reg [31:0] _RAND_1599;
  reg [31:0] _RAND_1600;
  reg [31:0] _RAND_1601;
  reg [31:0] _RAND_1602;
  reg [31:0] _RAND_1603;
  reg [31:0] _RAND_1604;
  reg [31:0] _RAND_1605;
  reg [31:0] _RAND_1606;
  reg [31:0] _RAND_1607;
  reg [31:0] _RAND_1608;
  reg [31:0] _RAND_1609;
  reg [31:0] _RAND_1610;
  reg [31:0] _RAND_1611;
  reg [31:0] _RAND_1612;
  reg [31:0] _RAND_1613;
  reg [31:0] _RAND_1614;
  reg [31:0] _RAND_1615;
  reg [31:0] _RAND_1616;
  reg [31:0] _RAND_1617;
  reg [31:0] _RAND_1618;
  reg [31:0] _RAND_1619;
  reg [31:0] _RAND_1620;
  reg [31:0] _RAND_1621;
  reg [31:0] _RAND_1622;
  reg [31:0] _RAND_1623;
  reg [31:0] _RAND_1624;
  reg [31:0] _RAND_1625;
  reg [31:0] _RAND_1626;
  reg [31:0] _RAND_1627;
  reg [31:0] _RAND_1628;
  reg [31:0] _RAND_1629;
  reg [31:0] _RAND_1630;
  reg [31:0] _RAND_1631;
  reg [31:0] _RAND_1632;
  reg [31:0] _RAND_1633;
  reg [31:0] _RAND_1634;
  reg [31:0] _RAND_1635;
  reg [31:0] _RAND_1636;
  reg [31:0] _RAND_1637;
  reg [31:0] _RAND_1638;
  reg [31:0] _RAND_1639;
  reg [31:0] _RAND_1640;
  reg [31:0] _RAND_1641;
  reg [31:0] _RAND_1642;
  reg [31:0] _RAND_1643;
  reg [31:0] _RAND_1644;
  reg [31:0] _RAND_1645;
  reg [31:0] _RAND_1646;
  reg [31:0] _RAND_1647;
  reg [31:0] _RAND_1648;
  reg [31:0] _RAND_1649;
  reg [31:0] _RAND_1650;
  reg [31:0] _RAND_1651;
  reg [31:0] _RAND_1652;
  reg [31:0] _RAND_1653;
  reg [31:0] _RAND_1654;
  reg [31:0] _RAND_1655;
  reg [31:0] _RAND_1656;
  reg [31:0] _RAND_1657;
  reg [31:0] _RAND_1658;
  reg [31:0] _RAND_1659;
  reg [31:0] _RAND_1660;
  reg [31:0] _RAND_1661;
  reg [31:0] _RAND_1662;
  reg [31:0] _RAND_1663;
  reg [31:0] _RAND_1664;
  reg [31:0] _RAND_1665;
  reg [31:0] _RAND_1666;
  reg [31:0] _RAND_1667;
  reg [31:0] _RAND_1668;
  reg [31:0] _RAND_1669;
  reg [31:0] _RAND_1670;
  reg [31:0] _RAND_1671;
  reg [31:0] _RAND_1672;
  reg [31:0] _RAND_1673;
  reg [31:0] _RAND_1674;
  reg [31:0] _RAND_1675;
  reg [31:0] _RAND_1676;
  reg [31:0] _RAND_1677;
  reg [31:0] _RAND_1678;
  reg [31:0] _RAND_1679;
  reg [31:0] _RAND_1680;
  reg [31:0] _RAND_1681;
  reg [31:0] _RAND_1682;
  reg [31:0] _RAND_1683;
  reg [31:0] _RAND_1684;
  reg [31:0] _RAND_1685;
  reg [31:0] _RAND_1686;
  reg [31:0] _RAND_1687;
  reg [31:0] _RAND_1688;
  reg [31:0] _RAND_1689;
  reg [31:0] _RAND_1690;
  reg [31:0] _RAND_1691;
  reg [31:0] _RAND_1692;
  reg [31:0] _RAND_1693;
  reg [31:0] _RAND_1694;
  reg [31:0] _RAND_1695;
  reg [31:0] _RAND_1696;
  reg [31:0] _RAND_1697;
  reg [31:0] _RAND_1698;
  reg [31:0] _RAND_1699;
  reg [31:0] _RAND_1700;
  reg [31:0] _RAND_1701;
  reg [31:0] _RAND_1702;
  reg [31:0] _RAND_1703;
  reg [31:0] _RAND_1704;
  reg [31:0] _RAND_1705;
  reg [31:0] _RAND_1706;
  reg [31:0] _RAND_1707;
  reg [31:0] _RAND_1708;
  reg [31:0] _RAND_1709;
  reg [31:0] _RAND_1710;
  reg [31:0] _RAND_1711;
  reg [31:0] _RAND_1712;
  reg [31:0] _RAND_1713;
  reg [31:0] _RAND_1714;
  reg [31:0] _RAND_1715;
  reg [31:0] _RAND_1716;
  reg [31:0] _RAND_1717;
  reg [31:0] _RAND_1718;
  reg [31:0] _RAND_1719;
  reg [31:0] _RAND_1720;
  reg [31:0] _RAND_1721;
  reg [31:0] _RAND_1722;
  reg [31:0] _RAND_1723;
  reg [31:0] _RAND_1724;
  reg [31:0] _RAND_1725;
  reg [31:0] _RAND_1726;
  reg [31:0] _RAND_1727;
  reg [31:0] _RAND_1728;
  reg [31:0] _RAND_1729;
  reg [31:0] _RAND_1730;
  reg [31:0] _RAND_1731;
  reg [31:0] _RAND_1732;
  reg [31:0] _RAND_1733;
  reg [31:0] _RAND_1734;
  reg [31:0] _RAND_1735;
  reg [31:0] _RAND_1736;
  reg [31:0] _RAND_1737;
  reg [31:0] _RAND_1738;
  reg [31:0] _RAND_1739;
  reg [31:0] _RAND_1740;
  reg [31:0] _RAND_1741;
  reg [31:0] _RAND_1742;
  reg [31:0] _RAND_1743;
  reg [31:0] _RAND_1744;
  reg [31:0] _RAND_1745;
  reg [31:0] _RAND_1746;
  reg [31:0] _RAND_1747;
  reg [31:0] _RAND_1748;
  reg [31:0] _RAND_1749;
  reg [31:0] _RAND_1750;
  reg [31:0] _RAND_1751;
  reg [31:0] _RAND_1752;
  reg [31:0] _RAND_1753;
  reg [31:0] _RAND_1754;
  reg [31:0] _RAND_1755;
  reg [31:0] _RAND_1756;
  reg [31:0] _RAND_1757;
  reg [31:0] _RAND_1758;
  reg [31:0] _RAND_1759;
  reg [31:0] _RAND_1760;
  reg [31:0] _RAND_1761;
  reg [31:0] _RAND_1762;
  reg [31:0] _RAND_1763;
  reg [31:0] _RAND_1764;
  reg [31:0] _RAND_1765;
  reg [31:0] _RAND_1766;
  reg [31:0] _RAND_1767;
  reg [31:0] _RAND_1768;
  reg [31:0] _RAND_1769;
  reg [31:0] _RAND_1770;
  reg [31:0] _RAND_1771;
  reg [31:0] _RAND_1772;
  reg [31:0] _RAND_1773;
  reg [31:0] _RAND_1774;
  reg [31:0] _RAND_1775;
  reg [31:0] _RAND_1776;
  reg [31:0] _RAND_1777;
  reg [31:0] _RAND_1778;
  reg [31:0] _RAND_1779;
  reg [31:0] _RAND_1780;
  reg [31:0] _RAND_1781;
  reg [31:0] _RAND_1782;
  reg [31:0] _RAND_1783;
  reg [31:0] _RAND_1784;
  reg [31:0] _RAND_1785;
  reg [31:0] _RAND_1786;
  reg [31:0] _RAND_1787;
  reg [31:0] _RAND_1788;
  reg [31:0] _RAND_1789;
  reg [31:0] _RAND_1790;
  reg [31:0] _RAND_1791;
  reg [31:0] _RAND_1792;
  reg [31:0] _RAND_1793;
  reg [31:0] _RAND_1794;
  reg [31:0] _RAND_1795;
  reg [31:0] _RAND_1796;
  reg [31:0] _RAND_1797;
  reg [31:0] _RAND_1798;
  reg [31:0] _RAND_1799;
  reg [31:0] _RAND_1800;
  reg [31:0] _RAND_1801;
  reg [31:0] _RAND_1802;
  reg [31:0] _RAND_1803;
  reg [31:0] _RAND_1804;
  reg [31:0] _RAND_1805;
  reg [31:0] _RAND_1806;
  reg [31:0] _RAND_1807;
  reg [31:0] _RAND_1808;
  reg [31:0] _RAND_1809;
  reg [31:0] _RAND_1810;
  reg [31:0] _RAND_1811;
  reg [31:0] _RAND_1812;
  reg [31:0] _RAND_1813;
  reg [31:0] _RAND_1814;
  reg [31:0] _RAND_1815;
  reg [31:0] _RAND_1816;
  reg [31:0] _RAND_1817;
  reg [31:0] _RAND_1818;
  reg [31:0] _RAND_1819;
  reg [31:0] _RAND_1820;
  reg [31:0] _RAND_1821;
  reg [31:0] _RAND_1822;
  reg [31:0] _RAND_1823;
  reg [31:0] _RAND_1824;
  reg [31:0] _RAND_1825;
  reg [31:0] _RAND_1826;
  reg [31:0] _RAND_1827;
  reg [31:0] _RAND_1828;
  reg [31:0] _RAND_1829;
  reg [31:0] _RAND_1830;
  reg [31:0] _RAND_1831;
  reg [31:0] _RAND_1832;
  reg [31:0] _RAND_1833;
  reg [31:0] _RAND_1834;
  reg [31:0] _RAND_1835;
  reg [31:0] _RAND_1836;
  reg [31:0] _RAND_1837;
  reg [31:0] _RAND_1838;
  reg [31:0] _RAND_1839;
  reg [31:0] _RAND_1840;
  reg [31:0] _RAND_1841;
  reg [31:0] _RAND_1842;
  reg [31:0] _RAND_1843;
  reg [31:0] _RAND_1844;
  reg [31:0] _RAND_1845;
  reg [31:0] _RAND_1846;
  reg [31:0] _RAND_1847;
  reg [31:0] _RAND_1848;
  reg [31:0] _RAND_1849;
  reg [31:0] _RAND_1850;
  reg [31:0] _RAND_1851;
  reg [31:0] _RAND_1852;
  reg [31:0] _RAND_1853;
  reg [31:0] _RAND_1854;
  reg [31:0] _RAND_1855;
  reg [31:0] _RAND_1856;
  reg [31:0] _RAND_1857;
  reg [31:0] _RAND_1858;
  reg [31:0] _RAND_1859;
  reg [31:0] _RAND_1860;
  reg [31:0] _RAND_1861;
  reg [31:0] _RAND_1862;
  reg [31:0] _RAND_1863;
  reg [31:0] _RAND_1864;
  reg [31:0] _RAND_1865;
  reg [31:0] _RAND_1866;
  reg [31:0] _RAND_1867;
  reg [31:0] _RAND_1868;
  reg [31:0] _RAND_1869;
  reg [31:0] _RAND_1870;
  reg [31:0] _RAND_1871;
  reg [31:0] _RAND_1872;
  reg [31:0] _RAND_1873;
  reg [31:0] _RAND_1874;
  reg [31:0] _RAND_1875;
  reg [31:0] _RAND_1876;
  reg [31:0] _RAND_1877;
  reg [31:0] _RAND_1878;
  reg [31:0] _RAND_1879;
  reg [31:0] _RAND_1880;
  reg [31:0] _RAND_1881;
  reg [31:0] _RAND_1882;
  reg [31:0] _RAND_1883;
  reg [31:0] _RAND_1884;
  reg [31:0] _RAND_1885;
  reg [31:0] _RAND_1886;
  reg [31:0] _RAND_1887;
  reg [31:0] _RAND_1888;
  reg [31:0] _RAND_1889;
  reg [31:0] _RAND_1890;
  reg [31:0] _RAND_1891;
  reg [31:0] _RAND_1892;
  reg [31:0] _RAND_1893;
  reg [31:0] _RAND_1894;
  reg [31:0] _RAND_1895;
  reg [31:0] _RAND_1896;
  reg [31:0] _RAND_1897;
  reg [31:0] _RAND_1898;
  reg [31:0] _RAND_1899;
  reg [31:0] _RAND_1900;
  reg [31:0] _RAND_1901;
  reg [31:0] _RAND_1902;
  reg [31:0] _RAND_1903;
  reg [31:0] _RAND_1904;
  reg [31:0] _RAND_1905;
  reg [31:0] _RAND_1906;
  reg [31:0] _RAND_1907;
  reg [31:0] _RAND_1908;
  reg [31:0] _RAND_1909;
  reg [31:0] _RAND_1910;
  reg [31:0] _RAND_1911;
  reg [31:0] _RAND_1912;
  reg [31:0] _RAND_1913;
  reg [31:0] _RAND_1914;
  reg [31:0] _RAND_1915;
  reg [31:0] _RAND_1916;
  reg [31:0] _RAND_1917;
  reg [31:0] _RAND_1918;
  reg [31:0] _RAND_1919;
  reg [31:0] _RAND_1920;
  reg [31:0] _RAND_1921;
  reg [31:0] _RAND_1922;
  reg [31:0] _RAND_1923;
  reg [31:0] _RAND_1924;
  reg [31:0] _RAND_1925;
  reg [31:0] _RAND_1926;
  reg [31:0] _RAND_1927;
  reg [31:0] _RAND_1928;
  reg [31:0] _RAND_1929;
  reg [31:0] _RAND_1930;
  reg [31:0] _RAND_1931;
  reg [31:0] _RAND_1932;
  reg [31:0] _RAND_1933;
  reg [31:0] _RAND_1934;
  reg [31:0] _RAND_1935;
  reg [31:0] _RAND_1936;
  reg [31:0] _RAND_1937;
  reg [31:0] _RAND_1938;
  reg [31:0] _RAND_1939;
  reg [31:0] _RAND_1940;
  reg [31:0] _RAND_1941;
  reg [31:0] _RAND_1942;
  reg [31:0] _RAND_1943;
  reg [31:0] _RAND_1944;
  reg [31:0] _RAND_1945;
  reg [31:0] _RAND_1946;
  reg [31:0] _RAND_1947;
  reg [31:0] _RAND_1948;
  reg [31:0] _RAND_1949;
  reg [31:0] _RAND_1950;
  reg [31:0] _RAND_1951;
  reg [31:0] _RAND_1952;
  reg [31:0] _RAND_1953;
  reg [31:0] _RAND_1954;
  reg [31:0] _RAND_1955;
  reg [31:0] _RAND_1956;
  reg [31:0] _RAND_1957;
  reg [31:0] _RAND_1958;
  reg [31:0] _RAND_1959;
  reg [31:0] _RAND_1960;
  reg [31:0] _RAND_1961;
  reg [31:0] _RAND_1962;
  reg [31:0] _RAND_1963;
  reg [31:0] _RAND_1964;
  reg [31:0] _RAND_1965;
  reg [31:0] _RAND_1966;
  reg [31:0] _RAND_1967;
  reg [31:0] _RAND_1968;
  reg [31:0] _RAND_1969;
  reg [31:0] _RAND_1970;
  reg [31:0] _RAND_1971;
  reg [31:0] _RAND_1972;
  reg [31:0] _RAND_1973;
  reg [31:0] _RAND_1974;
  reg [31:0] _RAND_1975;
  reg [31:0] _RAND_1976;
  reg [31:0] _RAND_1977;
  reg [31:0] _RAND_1978;
  reg [31:0] _RAND_1979;
  reg [31:0] _RAND_1980;
  reg [31:0] _RAND_1981;
  reg [31:0] _RAND_1982;
  reg [31:0] _RAND_1983;
  reg [31:0] _RAND_1984;
  reg [31:0] _RAND_1985;
  reg [31:0] _RAND_1986;
  reg [31:0] _RAND_1987;
  reg [31:0] _RAND_1988;
  reg [31:0] _RAND_1989;
  reg [31:0] _RAND_1990;
  reg [31:0] _RAND_1991;
  reg [31:0] _RAND_1992;
  reg [31:0] _RAND_1993;
  reg [31:0] _RAND_1994;
  reg [31:0] _RAND_1995;
  reg [31:0] _RAND_1996;
  reg [31:0] _RAND_1997;
  reg [31:0] _RAND_1998;
  reg [31:0] _RAND_1999;
  reg [31:0] _RAND_2000;
  reg [31:0] _RAND_2001;
  reg [31:0] _RAND_2002;
  reg [31:0] _RAND_2003;
  reg [31:0] _RAND_2004;
  reg [31:0] _RAND_2005;
  reg [31:0] _RAND_2006;
  reg [31:0] _RAND_2007;
  reg [31:0] _RAND_2008;
  reg [31:0] _RAND_2009;
  reg [31:0] _RAND_2010;
  reg [31:0] _RAND_2011;
  reg [31:0] _RAND_2012;
  reg [31:0] _RAND_2013;
  reg [31:0] _RAND_2014;
  reg [31:0] _RAND_2015;
  reg [31:0] _RAND_2016;
  reg [31:0] _RAND_2017;
  reg [31:0] _RAND_2018;
  reg [31:0] _RAND_2019;
  reg [31:0] _RAND_2020;
  reg [31:0] _RAND_2021;
  reg [31:0] _RAND_2022;
  reg [31:0] _RAND_2023;
  reg [31:0] _RAND_2024;
  reg [31:0] _RAND_2025;
  reg [31:0] _RAND_2026;
  reg [31:0] _RAND_2027;
  reg [31:0] _RAND_2028;
  reg [31:0] _RAND_2029;
  reg [31:0] _RAND_2030;
  reg [31:0] _RAND_2031;
  reg [31:0] _RAND_2032;
  reg [31:0] _RAND_2033;
  reg [31:0] _RAND_2034;
  reg [31:0] _RAND_2035;
  reg [31:0] _RAND_2036;
  reg [31:0] _RAND_2037;
  reg [31:0] _RAND_2038;
  reg [31:0] _RAND_2039;
  reg [31:0] _RAND_2040;
  reg [31:0] _RAND_2041;
  reg [31:0] _RAND_2042;
  reg [31:0] _RAND_2043;
  reg [31:0] _RAND_2044;
  reg [31:0] _RAND_2045;
  reg [31:0] _RAND_2046;
  reg [31:0] _RAND_2047;
  reg [31:0] _RAND_2048;
  reg [31:0] _RAND_2049;
  reg [31:0] _RAND_2050;
  reg [31:0] _RAND_2051;
  reg [31:0] _RAND_2052;
  reg [31:0] _RAND_2053;
  reg [31:0] _RAND_2054;
  reg [31:0] _RAND_2055;
  reg [31:0] _RAND_2056;
  reg [31:0] _RAND_2057;
  reg [31:0] _RAND_2058;
  reg [31:0] _RAND_2059;
  reg [31:0] _RAND_2060;
  reg [31:0] _RAND_2061;
  reg [31:0] _RAND_2062;
  reg [31:0] _RAND_2063;
  reg [31:0] _RAND_2064;
  reg [31:0] _RAND_2065;
  reg [31:0] _RAND_2066;
  reg [31:0] _RAND_2067;
  reg [31:0] _RAND_2068;
  reg [31:0] _RAND_2069;
  reg [31:0] _RAND_2070;
  reg [31:0] _RAND_2071;
  reg [31:0] _RAND_2072;
  reg [31:0] _RAND_2073;
  reg [31:0] _RAND_2074;
  reg [31:0] _RAND_2075;
  reg [31:0] _RAND_2076;
  reg [31:0] _RAND_2077;
  reg [31:0] _RAND_2078;
  reg [31:0] _RAND_2079;
  reg [31:0] _RAND_2080;
  reg [31:0] _RAND_2081;
  reg [31:0] _RAND_2082;
  reg [31:0] _RAND_2083;
  reg [31:0] _RAND_2084;
  reg [31:0] _RAND_2085;
  reg [31:0] _RAND_2086;
  reg [31:0] _RAND_2087;
  reg [31:0] _RAND_2088;
  reg [31:0] _RAND_2089;
  reg [31:0] _RAND_2090;
  reg [31:0] _RAND_2091;
  reg [31:0] _RAND_2092;
  reg [31:0] _RAND_2093;
  reg [31:0] _RAND_2094;
  reg [31:0] _RAND_2095;
  reg [31:0] _RAND_2096;
  reg [31:0] _RAND_2097;
  reg [31:0] _RAND_2098;
  reg [31:0] _RAND_2099;
  reg [31:0] _RAND_2100;
  reg [31:0] _RAND_2101;
  reg [31:0] _RAND_2102;
  reg [31:0] _RAND_2103;
  reg [31:0] _RAND_2104;
  reg [31:0] _RAND_2105;
  reg [31:0] _RAND_2106;
  reg [31:0] _RAND_2107;
  reg [31:0] _RAND_2108;
  reg [31:0] _RAND_2109;
  reg [31:0] _RAND_2110;
  reg [31:0] _RAND_2111;
  reg [31:0] _RAND_2112;
  reg [31:0] _RAND_2113;
  reg [31:0] _RAND_2114;
  reg [31:0] _RAND_2115;
  reg [31:0] _RAND_2116;
  reg [31:0] _RAND_2117;
  reg [31:0] _RAND_2118;
  reg [31:0] _RAND_2119;
  reg [31:0] _RAND_2120;
  reg [31:0] _RAND_2121;
  reg [31:0] _RAND_2122;
  reg [31:0] _RAND_2123;
  reg [31:0] _RAND_2124;
  reg [31:0] _RAND_2125;
  reg [31:0] _RAND_2126;
  reg [31:0] _RAND_2127;
  reg [31:0] _RAND_2128;
  reg [31:0] _RAND_2129;
  reg [31:0] _RAND_2130;
  reg [31:0] _RAND_2131;
  reg [31:0] _RAND_2132;
  reg [31:0] _RAND_2133;
  reg [31:0] _RAND_2134;
  reg [31:0] _RAND_2135;
  reg [31:0] _RAND_2136;
  reg [31:0] _RAND_2137;
  reg [31:0] _RAND_2138;
  reg [31:0] _RAND_2139;
  reg [31:0] _RAND_2140;
  reg [31:0] _RAND_2141;
  reg [31:0] _RAND_2142;
  reg [31:0] _RAND_2143;
  reg [31:0] _RAND_2144;
  reg [31:0] _RAND_2145;
  reg [31:0] _RAND_2146;
  reg [31:0] _RAND_2147;
  reg [31:0] _RAND_2148;
  reg [31:0] _RAND_2149;
  reg [31:0] _RAND_2150;
  reg [31:0] _RAND_2151;
  reg [31:0] _RAND_2152;
  reg [31:0] _RAND_2153;
  reg [31:0] _RAND_2154;
  reg [31:0] _RAND_2155;
  reg [31:0] _RAND_2156;
  reg [31:0] _RAND_2157;
  reg [31:0] _RAND_2158;
  reg [31:0] _RAND_2159;
  reg [31:0] _RAND_2160;
  reg [31:0] _RAND_2161;
  reg [31:0] _RAND_2162;
  reg [31:0] _RAND_2163;
  reg [31:0] _RAND_2164;
  reg [31:0] _RAND_2165;
  reg [31:0] _RAND_2166;
  reg [31:0] _RAND_2167;
  reg [31:0] _RAND_2168;
  reg [31:0] _RAND_2169;
  reg [31:0] _RAND_2170;
  reg [31:0] _RAND_2171;
  reg [31:0] _RAND_2172;
  reg [31:0] _RAND_2173;
  reg [31:0] _RAND_2174;
  reg [31:0] _RAND_2175;
  reg [31:0] _RAND_2176;
  reg [31:0] _RAND_2177;
  reg [31:0] _RAND_2178;
  reg [31:0] _RAND_2179;
  reg [31:0] _RAND_2180;
  reg [31:0] _RAND_2181;
  reg [31:0] _RAND_2182;
  reg [31:0] _RAND_2183;
  reg [31:0] _RAND_2184;
  reg [31:0] _RAND_2185;
  reg [31:0] _RAND_2186;
  reg [31:0] _RAND_2187;
  reg [31:0] _RAND_2188;
  reg [31:0] _RAND_2189;
  reg [31:0] _RAND_2190;
  reg [31:0] _RAND_2191;
  reg [31:0] _RAND_2192;
  reg [31:0] _RAND_2193;
  reg [31:0] _RAND_2194;
  reg [31:0] _RAND_2195;
  reg [31:0] _RAND_2196;
  reg [31:0] _RAND_2197;
  reg [31:0] _RAND_2198;
  reg [31:0] _RAND_2199;
  reg [31:0] _RAND_2200;
  reg [31:0] _RAND_2201;
  reg [31:0] _RAND_2202;
  reg [31:0] _RAND_2203;
  reg [31:0] _RAND_2204;
  reg [31:0] _RAND_2205;
  reg [31:0] _RAND_2206;
  reg [31:0] _RAND_2207;
  reg [31:0] _RAND_2208;
  reg [31:0] _RAND_2209;
  reg [31:0] _RAND_2210;
  reg [31:0] _RAND_2211;
  reg [31:0] _RAND_2212;
  reg [31:0] _RAND_2213;
  reg [31:0] _RAND_2214;
  reg [31:0] _RAND_2215;
  reg [31:0] _RAND_2216;
  reg [31:0] _RAND_2217;
  reg [31:0] _RAND_2218;
  reg [31:0] _RAND_2219;
  reg [31:0] _RAND_2220;
  reg [31:0] _RAND_2221;
  reg [31:0] _RAND_2222;
  reg [31:0] _RAND_2223;
  reg [31:0] _RAND_2224;
  reg [31:0] _RAND_2225;
  reg [31:0] _RAND_2226;
  reg [31:0] _RAND_2227;
  reg [31:0] _RAND_2228;
  reg [31:0] _RAND_2229;
  reg [31:0] _RAND_2230;
  reg [31:0] _RAND_2231;
  reg [31:0] _RAND_2232;
  reg [31:0] _RAND_2233;
  reg [31:0] _RAND_2234;
  reg [31:0] _RAND_2235;
  reg [31:0] _RAND_2236;
  reg [31:0] _RAND_2237;
  reg [31:0] _RAND_2238;
  reg [31:0] _RAND_2239;
  reg [31:0] _RAND_2240;
  reg [31:0] _RAND_2241;
  reg [31:0] _RAND_2242;
  reg [31:0] _RAND_2243;
  reg [31:0] _RAND_2244;
  reg [31:0] _RAND_2245;
  reg [31:0] _RAND_2246;
  reg [31:0] _RAND_2247;
  reg [31:0] _RAND_2248;
  reg [31:0] _RAND_2249;
  reg [31:0] _RAND_2250;
  reg [31:0] _RAND_2251;
  reg [31:0] _RAND_2252;
  reg [31:0] _RAND_2253;
  reg [31:0] _RAND_2254;
  reg [31:0] _RAND_2255;
  reg [31:0] _RAND_2256;
  reg [31:0] _RAND_2257;
  reg [31:0] _RAND_2258;
  reg [31:0] _RAND_2259;
  reg [31:0] _RAND_2260;
  reg [31:0] _RAND_2261;
  reg [31:0] _RAND_2262;
  reg [31:0] _RAND_2263;
  reg [31:0] _RAND_2264;
  reg [31:0] _RAND_2265;
  reg [31:0] _RAND_2266;
  reg [31:0] _RAND_2267;
  reg [31:0] _RAND_2268;
  reg [31:0] _RAND_2269;
  reg [31:0] _RAND_2270;
  reg [31:0] _RAND_2271;
  reg [31:0] _RAND_2272;
  reg [31:0] _RAND_2273;
  reg [31:0] _RAND_2274;
  reg [31:0] _RAND_2275;
  reg [31:0] _RAND_2276;
  reg [31:0] _RAND_2277;
  reg [31:0] _RAND_2278;
  reg [31:0] _RAND_2279;
  reg [31:0] _RAND_2280;
  reg [31:0] _RAND_2281;
  reg [31:0] _RAND_2282;
  reg [31:0] _RAND_2283;
  reg [31:0] _RAND_2284;
  reg [31:0] _RAND_2285;
  reg [31:0] _RAND_2286;
  reg [31:0] _RAND_2287;
  reg [31:0] _RAND_2288;
  reg [31:0] _RAND_2289;
  reg [31:0] _RAND_2290;
  reg [31:0] _RAND_2291;
  reg [31:0] _RAND_2292;
  reg [31:0] _RAND_2293;
  reg [31:0] _RAND_2294;
  reg [31:0] _RAND_2295;
  reg [31:0] _RAND_2296;
  reg [31:0] _RAND_2297;
  reg [31:0] _RAND_2298;
  reg [31:0] _RAND_2299;
  reg [31:0] _RAND_2300;
  reg [31:0] _RAND_2301;
  reg [31:0] _RAND_2302;
  reg [31:0] _RAND_2303;
  reg [31:0] _RAND_2304;
  reg [31:0] _RAND_2305;
  reg [31:0] _RAND_2306;
  reg [31:0] _RAND_2307;
  reg [31:0] _RAND_2308;
  reg [31:0] _RAND_2309;
  reg [31:0] _RAND_2310;
  reg [31:0] _RAND_2311;
  reg [31:0] _RAND_2312;
  reg [31:0] _RAND_2313;
  reg [31:0] _RAND_2314;
  reg [31:0] _RAND_2315;
  reg [31:0] _RAND_2316;
  reg [31:0] _RAND_2317;
  reg [31:0] _RAND_2318;
  reg [31:0] _RAND_2319;
  reg [31:0] _RAND_2320;
  reg [31:0] _RAND_2321;
  reg [31:0] _RAND_2322;
  reg [31:0] _RAND_2323;
  reg [31:0] _RAND_2324;
  reg [31:0] _RAND_2325;
  reg [31:0] _RAND_2326;
  reg [31:0] _RAND_2327;
  reg [31:0] _RAND_2328;
  reg [31:0] _RAND_2329;
  reg [31:0] _RAND_2330;
  reg [31:0] _RAND_2331;
  reg [31:0] _RAND_2332;
  reg [31:0] _RAND_2333;
  reg [31:0] _RAND_2334;
  reg [31:0] _RAND_2335;
  reg [31:0] _RAND_2336;
  reg [31:0] _RAND_2337;
  reg [31:0] _RAND_2338;
  reg [31:0] _RAND_2339;
  reg [31:0] _RAND_2340;
  reg [31:0] _RAND_2341;
  reg [31:0] _RAND_2342;
  reg [31:0] _RAND_2343;
  reg [31:0] _RAND_2344;
  reg [31:0] _RAND_2345;
  reg [31:0] _RAND_2346;
  reg [31:0] _RAND_2347;
  reg [31:0] _RAND_2348;
  reg [31:0] _RAND_2349;
  reg [31:0] _RAND_2350;
  reg [31:0] _RAND_2351;
  reg [31:0] _RAND_2352;
  reg [31:0] _RAND_2353;
  reg [31:0] _RAND_2354;
  reg [31:0] _RAND_2355;
  reg [31:0] _RAND_2356;
  reg [31:0] _RAND_2357;
  reg [31:0] _RAND_2358;
  reg [31:0] _RAND_2359;
  reg [31:0] _RAND_2360;
  reg [31:0] _RAND_2361;
  reg [31:0] _RAND_2362;
  reg [31:0] _RAND_2363;
  reg [31:0] _RAND_2364;
  reg [31:0] _RAND_2365;
  reg [31:0] _RAND_2366;
  reg [31:0] _RAND_2367;
  reg [31:0] _RAND_2368;
  reg [31:0] _RAND_2369;
  reg [31:0] _RAND_2370;
  reg [31:0] _RAND_2371;
  reg [31:0] _RAND_2372;
  reg [31:0] _RAND_2373;
  reg [31:0] _RAND_2374;
  reg [31:0] _RAND_2375;
  reg [31:0] _RAND_2376;
  reg [31:0] _RAND_2377;
  reg [31:0] _RAND_2378;
  reg [31:0] _RAND_2379;
  reg [31:0] _RAND_2380;
  reg [31:0] _RAND_2381;
  reg [31:0] _RAND_2382;
  reg [31:0] _RAND_2383;
  reg [31:0] _RAND_2384;
  reg [31:0] _RAND_2385;
  reg [31:0] _RAND_2386;
  reg [31:0] _RAND_2387;
  reg [31:0] _RAND_2388;
  reg [31:0] _RAND_2389;
  reg [31:0] _RAND_2390;
  reg [31:0] _RAND_2391;
  reg [31:0] _RAND_2392;
  reg [31:0] _RAND_2393;
  reg [31:0] _RAND_2394;
  reg [31:0] _RAND_2395;
  reg [31:0] _RAND_2396;
  reg [31:0] _RAND_2397;
  reg [31:0] _RAND_2398;
  reg [31:0] _RAND_2399;
  reg [31:0] _RAND_2400;
  reg [31:0] _RAND_2401;
  reg [31:0] _RAND_2402;
  reg [31:0] _RAND_2403;
  reg [31:0] _RAND_2404;
  reg [31:0] _RAND_2405;
  reg [31:0] _RAND_2406;
  reg [31:0] _RAND_2407;
  reg [31:0] _RAND_2408;
  reg [31:0] _RAND_2409;
  reg [31:0] _RAND_2410;
  reg [31:0] _RAND_2411;
  reg [31:0] _RAND_2412;
  reg [31:0] _RAND_2413;
  reg [31:0] _RAND_2414;
  reg [31:0] _RAND_2415;
  reg [31:0] _RAND_2416;
  reg [31:0] _RAND_2417;
  reg [31:0] _RAND_2418;
  reg [31:0] _RAND_2419;
  reg [31:0] _RAND_2420;
  reg [31:0] _RAND_2421;
  reg [31:0] _RAND_2422;
  reg [31:0] _RAND_2423;
  reg [31:0] _RAND_2424;
  reg [31:0] _RAND_2425;
  reg [31:0] _RAND_2426;
  reg [31:0] _RAND_2427;
  reg [31:0] _RAND_2428;
  reg [31:0] _RAND_2429;
  reg [31:0] _RAND_2430;
  reg [31:0] _RAND_2431;
  reg [31:0] _RAND_2432;
  reg [31:0] _RAND_2433;
  reg [31:0] _RAND_2434;
  reg [31:0] _RAND_2435;
  reg [31:0] _RAND_2436;
  reg [31:0] _RAND_2437;
  reg [31:0] _RAND_2438;
  reg [31:0] _RAND_2439;
  reg [31:0] _RAND_2440;
  reg [31:0] _RAND_2441;
  reg [31:0] _RAND_2442;
  reg [31:0] _RAND_2443;
  reg [31:0] _RAND_2444;
  reg [31:0] _RAND_2445;
  reg [31:0] _RAND_2446;
  reg [31:0] _RAND_2447;
  reg [31:0] _RAND_2448;
  reg [31:0] _RAND_2449;
  reg [31:0] _RAND_2450;
  reg [31:0] _RAND_2451;
  reg [31:0] _RAND_2452;
  reg [31:0] _RAND_2453;
  reg [31:0] _RAND_2454;
  reg [31:0] _RAND_2455;
  reg [31:0] _RAND_2456;
  reg [31:0] _RAND_2457;
  reg [31:0] _RAND_2458;
  reg [31:0] _RAND_2459;
  reg [31:0] _RAND_2460;
  reg [31:0] _RAND_2461;
  reg [31:0] _RAND_2462;
  reg [31:0] _RAND_2463;
  reg [31:0] _RAND_2464;
  reg [31:0] _RAND_2465;
  reg [31:0] _RAND_2466;
  reg [31:0] _RAND_2467;
  reg [31:0] _RAND_2468;
  reg [31:0] _RAND_2469;
  reg [31:0] _RAND_2470;
  reg [31:0] _RAND_2471;
  reg [31:0] _RAND_2472;
  reg [31:0] _RAND_2473;
  reg [31:0] _RAND_2474;
  reg [31:0] _RAND_2475;
  reg [31:0] _RAND_2476;
  reg [31:0] _RAND_2477;
  reg [31:0] _RAND_2478;
  reg [31:0] _RAND_2479;
  reg [31:0] _RAND_2480;
  reg [31:0] _RAND_2481;
  reg [31:0] _RAND_2482;
  reg [31:0] _RAND_2483;
  reg [31:0] _RAND_2484;
  reg [31:0] _RAND_2485;
  reg [31:0] _RAND_2486;
  reg [31:0] _RAND_2487;
  reg [31:0] _RAND_2488;
  reg [31:0] _RAND_2489;
  reg [31:0] _RAND_2490;
  reg [31:0] _RAND_2491;
  reg [31:0] _RAND_2492;
  reg [31:0] _RAND_2493;
  reg [31:0] _RAND_2494;
  reg [31:0] _RAND_2495;
  reg [31:0] _RAND_2496;
  reg [31:0] _RAND_2497;
  reg [31:0] _RAND_2498;
  reg [31:0] _RAND_2499;
  reg [31:0] _RAND_2500;
  reg [31:0] _RAND_2501;
  reg [31:0] _RAND_2502;
  reg [31:0] _RAND_2503;
  reg [31:0] _RAND_2504;
  reg [31:0] _RAND_2505;
  reg [31:0] _RAND_2506;
  reg [31:0] _RAND_2507;
  reg [31:0] _RAND_2508;
  reg [31:0] _RAND_2509;
  reg [31:0] _RAND_2510;
  reg [31:0] _RAND_2511;
  reg [31:0] _RAND_2512;
  reg [31:0] _RAND_2513;
  reg [31:0] _RAND_2514;
  reg [31:0] _RAND_2515;
  reg [31:0] _RAND_2516;
  reg [31:0] _RAND_2517;
  reg [31:0] _RAND_2518;
  reg [31:0] _RAND_2519;
  reg [31:0] _RAND_2520;
  reg [31:0] _RAND_2521;
  reg [31:0] _RAND_2522;
  reg [31:0] _RAND_2523;
  reg [31:0] _RAND_2524;
  reg [31:0] _RAND_2525;
  reg [31:0] _RAND_2526;
  reg [31:0] _RAND_2527;
  reg [31:0] _RAND_2528;
  reg [31:0] _RAND_2529;
  reg [31:0] _RAND_2530;
  reg [31:0] _RAND_2531;
  reg [31:0] _RAND_2532;
  reg [31:0] _RAND_2533;
  reg [31:0] _RAND_2534;
  reg [31:0] _RAND_2535;
  reg [31:0] _RAND_2536;
  reg [31:0] _RAND_2537;
  reg [31:0] _RAND_2538;
  reg [31:0] _RAND_2539;
  reg [31:0] _RAND_2540;
  reg [31:0] _RAND_2541;
  reg [31:0] _RAND_2542;
  reg [31:0] _RAND_2543;
  reg [31:0] _RAND_2544;
  reg [31:0] _RAND_2545;
  reg [31:0] _RAND_2546;
  reg [31:0] _RAND_2547;
  reg [31:0] _RAND_2548;
  reg [31:0] _RAND_2549;
  reg [31:0] _RAND_2550;
  reg [31:0] _RAND_2551;
  reg [31:0] _RAND_2552;
  reg [31:0] _RAND_2553;
  reg [31:0] _RAND_2554;
  reg [31:0] _RAND_2555;
  reg [31:0] _RAND_2556;
  reg [31:0] _RAND_2557;
  reg [31:0] _RAND_2558;
  reg [31:0] _RAND_2559;
  reg [31:0] _RAND_2560;
  reg [31:0] _RAND_2561;
`endif // RANDOMIZE_REG_INIT
  wire  c22_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_1_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_1_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_1_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_1_io_out_1; // @[Multiplier.scala 120:25]
  wire  c32_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_io_out_1; // @[Multiplier.scala 125:25]
  wire  c32_1_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_1_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_1_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_1_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_1_io_out_1; // @[Multiplier.scala 125:25]
  wire  c53_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_1_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_1_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_1_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_1_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_1_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_1_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_1_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_1_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_2_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_2_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_2_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_2_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_2_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_2_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_2_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_2_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_3_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_3_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_3_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_3_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_3_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_3_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_3_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_3_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_4_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_4_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_4_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_4_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_4_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_4_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_4_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_4_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_2_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_2_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_2_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_2_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_5_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_5_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_5_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_5_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_5_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_5_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_5_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_5_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_3_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_3_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_3_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_3_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_6_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_6_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_6_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_6_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_6_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_6_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_6_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_6_io_out_2; // @[Multiplier.scala 130:25]
  wire  c32_2_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_2_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_2_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_2_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_2_io_out_1; // @[Multiplier.scala 125:25]
  wire  c53_7_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_7_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_7_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_7_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_7_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_7_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_7_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_7_io_out_2; // @[Multiplier.scala 130:25]
  wire  c32_3_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_3_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_3_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_3_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_3_io_out_1; // @[Multiplier.scala 125:25]
  wire  c53_8_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_8_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_8_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_8_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_8_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_8_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_8_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_8_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_9_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_9_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_9_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_9_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_9_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_9_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_9_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_9_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_10_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_10_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_10_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_10_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_10_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_10_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_10_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_10_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_11_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_11_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_11_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_11_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_11_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_11_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_11_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_11_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_12_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_12_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_12_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_12_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_12_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_12_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_12_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_12_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_13_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_13_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_13_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_13_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_13_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_13_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_13_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_13_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_14_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_14_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_14_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_14_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_14_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_14_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_14_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_14_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_15_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_15_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_15_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_15_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_15_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_15_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_15_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_15_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_16_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_16_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_16_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_16_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_16_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_16_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_16_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_16_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_17_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_17_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_17_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_17_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_17_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_17_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_17_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_17_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_4_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_4_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_4_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_4_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_18_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_18_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_18_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_18_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_18_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_18_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_18_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_18_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_19_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_19_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_19_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_19_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_19_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_19_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_19_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_19_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_5_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_5_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_5_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_5_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_20_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_20_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_20_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_20_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_20_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_20_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_20_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_20_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_21_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_21_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_21_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_21_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_21_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_21_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_21_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_21_io_out_2; // @[Multiplier.scala 130:25]
  wire  c32_4_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_4_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_4_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_4_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_4_io_out_1; // @[Multiplier.scala 125:25]
  wire  c53_22_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_22_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_22_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_22_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_22_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_22_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_22_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_22_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_23_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_23_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_23_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_23_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_23_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_23_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_23_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_23_io_out_2; // @[Multiplier.scala 130:25]
  wire  c32_5_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_5_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_5_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_5_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_5_io_out_1; // @[Multiplier.scala 125:25]
  wire  c53_24_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_24_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_24_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_24_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_24_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_24_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_24_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_24_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_25_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_25_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_25_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_25_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_25_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_25_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_25_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_25_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_26_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_26_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_26_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_26_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_26_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_26_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_26_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_26_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_27_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_27_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_27_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_27_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_27_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_27_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_27_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_27_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_28_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_28_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_28_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_28_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_28_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_28_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_28_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_28_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_29_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_29_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_29_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_29_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_29_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_29_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_29_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_29_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_30_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_30_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_30_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_30_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_30_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_30_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_30_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_30_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_31_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_31_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_31_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_31_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_31_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_31_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_31_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_31_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_32_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_32_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_32_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_32_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_32_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_32_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_32_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_32_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_33_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_33_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_33_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_33_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_33_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_33_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_33_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_33_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_34_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_34_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_34_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_34_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_34_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_34_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_34_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_34_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_35_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_35_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_35_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_35_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_35_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_35_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_35_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_35_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_36_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_36_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_36_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_36_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_36_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_36_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_36_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_36_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_37_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_37_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_37_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_37_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_37_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_37_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_37_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_37_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_38_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_38_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_38_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_38_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_38_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_38_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_38_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_38_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_6_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_6_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_6_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_6_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_39_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_39_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_39_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_39_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_39_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_39_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_39_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_39_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_40_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_40_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_40_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_40_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_40_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_40_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_40_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_40_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_41_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_41_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_41_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_41_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_41_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_41_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_41_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_41_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_7_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_7_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_7_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_7_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_42_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_42_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_42_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_42_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_42_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_42_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_42_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_42_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_43_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_43_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_43_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_43_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_43_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_43_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_43_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_43_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_44_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_44_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_44_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_44_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_44_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_44_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_44_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_44_io_out_2; // @[Multiplier.scala 130:25]
  wire  c32_6_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_6_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_6_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_6_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_6_io_out_1; // @[Multiplier.scala 125:25]
  wire  c53_45_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_45_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_45_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_45_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_45_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_45_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_45_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_45_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_46_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_46_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_46_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_46_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_46_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_46_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_46_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_46_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_47_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_47_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_47_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_47_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_47_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_47_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_47_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_47_io_out_2; // @[Multiplier.scala 130:25]
  wire  c32_7_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_7_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_7_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_7_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_7_io_out_1; // @[Multiplier.scala 125:25]
  wire  c53_48_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_48_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_48_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_48_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_48_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_48_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_48_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_48_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_49_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_49_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_49_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_49_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_49_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_49_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_49_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_49_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_50_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_50_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_50_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_50_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_50_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_50_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_50_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_50_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_51_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_51_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_51_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_51_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_51_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_51_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_51_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_51_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_52_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_52_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_52_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_52_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_52_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_52_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_52_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_52_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_53_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_53_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_53_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_53_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_53_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_53_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_53_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_53_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_54_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_54_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_54_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_54_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_54_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_54_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_54_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_54_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_55_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_55_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_55_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_55_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_55_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_55_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_55_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_55_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_56_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_56_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_56_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_56_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_56_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_56_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_56_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_56_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_57_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_57_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_57_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_57_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_57_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_57_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_57_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_57_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_58_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_58_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_58_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_58_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_58_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_58_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_58_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_58_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_59_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_59_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_59_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_59_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_59_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_59_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_59_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_59_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_60_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_60_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_60_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_60_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_60_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_60_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_60_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_60_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_61_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_61_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_61_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_61_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_61_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_61_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_61_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_61_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_62_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_62_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_62_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_62_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_62_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_62_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_62_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_62_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_63_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_63_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_63_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_63_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_63_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_63_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_63_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_63_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_64_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_64_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_64_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_64_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_64_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_64_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_64_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_64_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_65_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_65_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_65_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_65_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_65_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_65_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_65_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_65_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_66_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_66_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_66_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_66_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_66_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_66_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_66_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_66_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_67_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_67_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_67_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_67_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_67_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_67_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_67_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_67_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_8_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_8_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_8_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_8_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_68_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_68_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_68_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_68_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_68_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_68_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_68_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_68_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_69_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_69_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_69_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_69_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_69_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_69_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_69_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_69_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_70_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_70_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_70_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_70_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_70_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_70_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_70_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_70_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_71_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_71_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_71_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_71_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_71_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_71_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_71_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_71_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_9_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_9_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_9_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_9_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_72_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_72_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_72_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_72_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_72_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_72_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_72_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_72_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_73_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_73_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_73_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_73_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_73_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_73_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_73_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_73_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_74_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_74_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_74_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_74_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_74_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_74_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_74_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_74_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_75_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_75_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_75_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_75_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_75_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_75_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_75_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_75_io_out_2; // @[Multiplier.scala 130:25]
  wire  c32_8_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_8_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_8_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_8_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_8_io_out_1; // @[Multiplier.scala 125:25]
  wire  c53_76_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_76_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_76_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_76_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_76_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_76_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_76_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_76_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_77_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_77_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_77_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_77_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_77_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_77_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_77_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_77_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_78_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_78_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_78_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_78_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_78_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_78_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_78_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_78_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_79_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_79_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_79_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_79_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_79_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_79_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_79_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_79_io_out_2; // @[Multiplier.scala 130:25]
  wire  c32_9_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_9_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_9_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_9_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_9_io_out_1; // @[Multiplier.scala 125:25]
  wire  c53_80_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_80_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_80_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_80_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_80_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_80_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_80_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_80_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_81_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_81_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_81_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_81_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_81_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_81_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_81_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_81_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_82_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_82_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_82_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_82_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_82_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_82_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_82_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_82_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_83_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_83_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_83_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_83_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_83_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_83_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_83_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_83_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_84_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_84_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_84_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_84_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_84_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_84_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_84_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_84_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_85_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_85_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_85_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_85_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_85_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_85_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_85_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_85_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_86_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_86_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_86_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_86_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_86_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_86_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_86_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_86_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_87_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_87_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_87_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_87_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_87_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_87_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_87_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_87_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_88_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_88_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_88_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_88_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_88_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_88_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_88_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_88_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_89_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_89_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_89_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_89_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_89_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_89_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_89_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_89_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_90_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_90_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_90_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_90_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_90_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_90_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_90_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_90_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_91_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_91_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_91_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_91_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_91_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_91_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_91_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_91_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_92_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_92_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_92_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_92_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_92_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_92_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_92_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_92_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_93_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_93_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_93_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_93_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_93_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_93_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_93_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_93_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_94_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_94_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_94_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_94_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_94_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_94_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_94_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_94_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_95_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_95_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_95_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_95_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_95_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_95_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_95_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_95_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_96_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_96_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_96_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_96_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_96_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_96_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_96_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_96_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_97_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_97_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_97_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_97_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_97_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_97_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_97_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_97_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_98_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_98_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_98_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_98_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_98_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_98_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_98_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_98_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_99_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_99_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_99_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_99_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_99_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_99_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_99_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_99_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_100_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_100_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_100_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_100_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_100_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_100_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_100_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_100_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_101_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_101_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_101_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_101_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_101_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_101_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_101_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_101_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_102_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_102_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_102_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_102_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_102_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_102_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_102_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_102_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_103_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_103_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_103_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_103_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_103_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_103_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_103_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_103_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_104_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_104_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_104_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_104_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_104_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_104_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_104_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_104_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_10_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_10_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_10_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_10_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_105_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_105_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_105_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_105_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_105_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_105_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_105_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_105_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_106_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_106_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_106_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_106_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_106_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_106_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_106_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_106_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_107_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_107_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_107_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_107_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_107_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_107_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_107_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_107_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_108_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_108_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_108_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_108_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_108_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_108_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_108_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_108_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_109_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_109_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_109_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_109_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_109_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_109_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_109_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_109_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_11_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_11_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_11_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_11_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_110_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_110_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_110_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_110_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_110_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_110_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_110_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_110_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_111_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_111_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_111_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_111_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_111_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_111_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_111_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_111_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_112_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_112_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_112_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_112_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_112_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_112_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_112_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_112_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_113_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_113_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_113_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_113_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_113_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_113_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_113_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_113_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_114_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_114_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_114_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_114_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_114_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_114_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_114_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_114_io_out_2; // @[Multiplier.scala 130:25]
  wire  c32_10_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_10_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_10_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_10_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_10_io_out_1; // @[Multiplier.scala 125:25]
  wire  c53_115_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_115_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_115_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_115_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_115_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_115_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_115_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_115_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_116_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_116_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_116_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_116_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_116_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_116_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_116_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_116_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_117_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_117_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_117_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_117_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_117_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_117_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_117_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_117_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_118_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_118_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_118_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_118_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_118_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_118_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_118_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_118_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_119_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_119_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_119_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_119_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_119_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_119_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_119_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_119_io_out_2; // @[Multiplier.scala 130:25]
  wire  c32_11_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_11_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_11_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_11_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_11_io_out_1; // @[Multiplier.scala 125:25]
  wire  c53_120_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_120_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_120_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_120_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_120_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_120_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_120_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_120_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_121_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_121_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_121_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_121_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_121_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_121_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_121_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_121_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_122_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_122_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_122_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_122_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_122_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_122_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_122_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_122_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_123_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_123_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_123_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_123_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_123_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_123_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_123_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_123_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_124_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_124_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_124_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_124_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_124_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_124_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_124_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_124_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_125_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_125_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_125_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_125_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_125_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_125_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_125_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_125_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_126_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_126_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_126_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_126_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_126_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_126_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_126_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_126_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_127_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_127_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_127_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_127_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_127_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_127_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_127_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_127_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_128_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_128_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_128_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_128_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_128_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_128_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_128_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_128_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_129_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_129_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_129_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_129_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_129_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_129_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_129_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_129_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_130_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_130_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_130_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_130_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_130_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_130_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_130_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_130_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_131_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_131_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_131_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_131_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_131_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_131_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_131_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_131_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_132_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_132_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_132_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_132_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_132_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_132_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_132_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_132_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_133_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_133_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_133_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_133_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_133_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_133_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_133_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_133_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_134_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_134_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_134_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_134_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_134_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_134_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_134_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_134_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_135_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_135_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_135_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_135_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_135_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_135_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_135_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_135_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_136_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_136_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_136_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_136_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_136_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_136_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_136_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_136_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_137_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_137_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_137_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_137_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_137_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_137_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_137_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_137_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_138_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_138_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_138_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_138_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_138_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_138_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_138_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_138_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_139_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_139_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_139_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_139_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_139_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_139_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_139_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_139_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_140_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_140_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_140_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_140_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_140_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_140_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_140_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_140_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_141_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_141_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_141_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_141_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_141_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_141_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_141_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_141_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_142_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_142_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_142_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_142_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_142_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_142_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_142_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_142_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_143_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_143_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_143_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_143_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_143_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_143_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_143_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_143_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_144_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_144_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_144_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_144_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_144_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_144_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_144_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_144_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_145_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_145_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_145_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_145_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_145_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_145_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_145_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_145_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_146_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_146_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_146_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_146_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_146_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_146_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_146_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_146_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_147_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_147_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_147_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_147_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_147_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_147_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_147_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_147_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_148_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_148_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_148_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_148_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_148_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_148_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_148_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_148_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_149_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_149_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_149_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_149_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_149_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_149_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_149_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_149_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_12_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_12_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_12_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_12_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_150_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_150_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_150_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_150_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_150_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_150_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_150_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_150_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_151_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_151_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_151_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_151_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_151_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_151_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_151_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_151_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_152_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_152_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_152_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_152_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_152_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_152_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_152_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_152_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_153_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_153_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_153_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_153_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_153_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_153_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_153_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_153_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_154_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_154_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_154_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_154_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_154_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_154_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_154_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_154_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_155_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_155_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_155_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_155_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_155_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_155_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_155_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_155_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_13_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_13_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_13_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_13_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_156_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_156_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_156_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_156_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_156_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_156_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_156_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_156_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_157_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_157_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_157_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_157_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_157_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_157_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_157_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_157_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_158_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_158_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_158_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_158_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_158_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_158_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_158_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_158_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_159_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_159_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_159_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_159_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_159_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_159_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_159_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_159_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_160_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_160_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_160_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_160_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_160_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_160_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_160_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_160_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_161_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_161_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_161_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_161_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_161_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_161_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_161_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_161_io_out_2; // @[Multiplier.scala 130:25]
  wire  c32_12_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_12_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_12_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_12_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_12_io_out_1; // @[Multiplier.scala 125:25]
  wire  c53_162_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_162_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_162_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_162_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_162_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_162_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_162_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_162_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_163_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_163_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_163_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_163_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_163_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_163_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_163_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_163_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_164_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_164_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_164_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_164_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_164_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_164_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_164_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_164_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_165_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_165_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_165_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_165_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_165_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_165_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_165_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_165_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_166_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_166_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_166_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_166_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_166_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_166_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_166_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_166_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_167_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_167_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_167_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_167_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_167_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_167_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_167_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_167_io_out_2; // @[Multiplier.scala 130:25]
  wire  c32_13_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_13_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_13_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_13_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_13_io_out_1; // @[Multiplier.scala 125:25]
  wire  c53_168_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_168_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_168_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_168_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_168_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_168_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_168_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_168_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_169_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_169_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_169_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_169_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_169_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_169_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_169_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_169_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_170_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_170_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_170_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_170_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_170_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_170_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_170_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_170_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_171_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_171_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_171_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_171_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_171_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_171_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_171_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_171_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_172_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_172_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_172_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_172_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_172_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_172_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_172_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_172_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_173_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_173_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_173_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_173_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_173_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_173_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_173_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_173_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_174_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_174_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_174_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_174_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_174_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_174_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_174_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_174_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_175_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_175_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_175_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_175_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_175_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_175_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_175_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_175_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_176_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_176_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_176_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_176_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_176_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_176_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_176_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_176_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_177_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_177_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_177_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_177_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_177_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_177_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_177_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_177_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_178_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_178_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_178_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_178_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_178_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_178_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_178_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_178_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_179_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_179_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_179_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_179_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_179_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_179_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_179_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_179_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_180_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_180_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_180_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_180_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_180_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_180_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_180_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_180_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_181_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_181_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_181_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_181_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_181_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_181_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_181_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_181_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_182_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_182_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_182_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_182_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_182_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_182_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_182_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_182_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_183_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_183_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_183_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_183_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_183_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_183_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_183_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_183_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_184_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_184_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_184_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_184_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_184_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_184_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_184_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_184_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_185_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_185_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_185_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_185_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_185_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_185_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_185_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_185_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_186_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_186_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_186_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_186_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_186_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_186_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_186_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_186_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_187_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_187_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_187_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_187_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_187_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_187_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_187_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_187_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_188_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_188_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_188_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_188_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_188_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_188_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_188_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_188_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_189_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_189_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_189_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_189_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_189_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_189_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_189_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_189_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_190_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_190_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_190_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_190_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_190_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_190_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_190_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_190_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_191_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_191_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_191_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_191_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_191_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_191_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_191_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_191_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_192_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_192_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_192_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_192_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_192_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_192_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_192_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_192_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_193_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_193_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_193_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_193_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_193_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_193_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_193_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_193_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_194_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_194_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_194_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_194_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_194_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_194_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_194_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_194_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_195_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_195_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_195_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_195_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_195_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_195_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_195_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_195_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_196_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_196_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_196_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_196_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_196_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_196_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_196_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_196_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_197_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_197_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_197_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_197_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_197_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_197_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_197_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_197_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_198_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_198_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_198_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_198_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_198_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_198_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_198_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_198_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_199_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_199_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_199_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_199_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_199_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_199_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_199_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_199_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_200_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_200_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_200_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_200_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_200_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_200_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_200_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_200_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_201_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_201_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_201_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_201_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_201_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_201_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_201_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_201_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_202_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_202_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_202_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_202_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_202_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_202_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_202_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_202_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_14_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_14_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_14_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_14_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_203_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_203_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_203_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_203_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_203_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_203_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_203_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_203_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_204_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_204_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_204_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_204_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_204_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_204_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_204_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_204_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_205_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_205_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_205_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_205_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_205_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_205_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_205_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_205_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_206_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_206_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_206_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_206_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_206_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_206_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_206_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_206_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_207_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_207_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_207_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_207_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_207_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_207_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_207_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_207_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_208_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_208_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_208_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_208_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_208_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_208_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_208_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_208_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_209_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_209_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_209_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_209_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_209_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_209_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_209_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_209_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_15_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_15_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_15_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_15_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_210_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_210_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_210_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_210_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_210_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_210_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_210_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_210_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_211_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_211_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_211_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_211_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_211_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_211_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_211_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_211_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_212_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_212_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_212_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_212_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_212_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_212_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_212_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_212_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_213_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_213_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_213_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_213_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_213_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_213_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_213_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_213_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_214_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_214_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_214_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_214_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_214_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_214_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_214_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_214_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_215_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_215_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_215_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_215_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_215_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_215_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_215_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_215_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_216_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_216_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_216_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_216_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_216_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_216_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_216_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_216_io_out_2; // @[Multiplier.scala 130:25]
  wire  c32_14_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_14_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_14_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_14_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_14_io_out_1; // @[Multiplier.scala 125:25]
  wire  c53_217_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_217_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_217_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_217_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_217_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_217_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_217_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_217_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_218_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_218_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_218_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_218_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_218_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_218_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_218_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_218_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_219_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_219_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_219_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_219_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_219_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_219_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_219_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_219_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_220_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_220_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_220_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_220_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_220_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_220_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_220_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_220_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_221_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_221_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_221_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_221_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_221_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_221_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_221_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_221_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_222_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_222_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_222_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_222_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_222_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_222_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_222_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_222_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_223_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_223_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_223_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_223_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_223_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_223_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_223_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_223_io_out_2; // @[Multiplier.scala 130:25]
  wire  c32_15_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_15_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_15_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_15_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_15_io_out_1; // @[Multiplier.scala 125:25]
  wire  c53_224_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_224_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_224_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_224_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_224_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_224_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_224_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_224_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_225_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_225_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_225_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_225_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_225_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_225_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_225_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_225_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_226_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_226_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_226_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_226_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_226_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_226_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_226_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_226_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_227_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_227_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_227_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_227_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_227_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_227_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_227_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_227_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_228_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_228_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_228_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_228_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_228_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_228_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_228_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_228_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_229_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_229_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_229_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_229_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_229_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_229_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_229_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_229_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_230_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_230_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_230_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_230_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_230_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_230_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_230_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_230_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_231_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_231_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_231_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_231_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_231_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_231_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_231_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_231_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_232_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_232_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_232_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_232_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_232_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_232_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_232_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_232_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_233_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_233_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_233_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_233_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_233_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_233_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_233_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_233_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_234_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_234_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_234_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_234_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_234_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_234_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_234_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_234_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_235_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_235_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_235_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_235_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_235_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_235_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_235_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_235_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_236_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_236_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_236_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_236_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_236_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_236_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_236_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_236_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_237_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_237_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_237_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_237_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_237_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_237_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_237_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_237_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_238_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_238_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_238_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_238_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_238_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_238_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_238_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_238_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_239_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_239_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_239_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_239_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_239_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_239_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_239_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_239_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_240_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_240_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_240_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_240_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_240_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_240_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_240_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_240_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_241_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_241_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_241_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_241_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_241_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_241_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_241_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_241_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_242_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_242_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_242_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_242_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_242_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_242_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_242_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_242_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_243_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_243_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_243_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_243_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_243_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_243_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_243_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_243_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_244_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_244_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_244_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_244_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_244_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_244_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_244_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_244_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_245_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_245_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_245_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_245_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_245_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_245_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_245_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_245_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_246_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_246_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_246_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_246_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_246_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_246_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_246_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_246_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_247_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_247_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_247_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_247_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_247_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_247_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_247_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_247_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_248_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_248_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_248_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_248_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_248_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_248_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_248_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_248_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_249_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_249_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_249_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_249_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_249_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_249_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_249_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_249_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_250_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_250_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_250_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_250_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_250_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_250_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_250_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_250_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_251_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_251_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_251_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_251_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_251_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_251_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_251_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_251_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_252_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_252_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_252_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_252_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_252_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_252_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_252_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_252_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_253_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_253_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_253_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_253_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_253_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_253_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_253_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_253_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_254_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_254_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_254_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_254_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_254_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_254_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_254_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_254_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_255_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_255_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_255_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_255_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_255_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_255_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_255_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_255_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_256_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_256_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_256_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_256_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_256_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_256_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_256_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_256_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_257_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_257_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_257_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_257_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_257_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_257_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_257_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_257_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_258_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_258_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_258_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_258_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_258_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_258_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_258_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_258_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_259_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_259_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_259_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_259_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_259_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_259_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_259_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_259_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_260_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_260_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_260_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_260_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_260_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_260_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_260_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_260_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_261_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_261_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_261_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_261_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_261_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_261_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_261_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_261_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_262_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_262_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_262_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_262_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_262_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_262_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_262_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_262_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_263_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_263_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_263_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_263_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_263_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_263_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_263_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_263_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_264_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_264_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_264_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_264_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_264_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_264_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_264_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_264_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_265_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_265_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_265_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_265_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_265_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_265_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_265_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_265_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_266_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_266_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_266_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_266_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_266_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_266_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_266_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_266_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_267_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_267_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_267_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_267_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_267_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_267_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_267_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_267_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_268_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_268_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_268_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_268_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_268_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_268_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_268_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_268_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_269_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_269_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_269_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_269_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_269_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_269_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_269_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_269_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_270_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_270_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_270_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_270_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_270_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_270_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_270_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_270_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_271_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_271_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_271_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_271_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_271_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_271_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_271_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_271_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_272_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_272_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_272_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_272_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_272_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_272_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_272_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_272_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_273_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_273_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_273_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_273_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_273_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_273_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_273_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_273_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_274_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_274_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_274_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_274_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_274_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_274_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_274_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_274_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_275_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_275_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_275_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_275_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_275_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_275_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_275_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_275_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_276_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_276_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_276_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_276_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_276_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_276_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_276_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_276_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_277_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_277_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_277_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_277_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_277_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_277_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_277_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_277_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_278_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_278_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_278_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_278_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_278_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_278_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_278_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_278_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_279_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_279_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_279_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_279_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_279_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_279_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_279_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_279_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_280_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_280_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_280_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_280_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_280_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_280_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_280_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_280_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_281_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_281_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_281_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_281_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_281_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_281_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_281_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_281_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_282_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_282_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_282_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_282_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_282_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_282_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_282_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_282_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_283_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_283_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_283_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_283_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_283_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_283_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_283_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_283_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_284_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_284_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_284_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_284_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_284_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_284_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_284_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_284_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_285_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_285_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_285_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_285_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_285_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_285_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_285_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_285_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_286_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_286_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_286_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_286_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_286_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_286_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_286_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_286_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_287_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_287_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_287_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_287_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_287_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_287_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_287_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_287_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_288_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_288_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_288_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_288_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_288_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_288_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_288_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_288_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_289_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_289_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_289_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_289_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_289_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_289_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_289_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_289_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_290_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_290_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_290_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_290_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_290_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_290_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_290_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_290_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_291_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_291_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_291_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_291_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_291_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_291_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_291_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_291_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_292_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_292_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_292_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_292_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_292_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_292_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_292_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_292_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_293_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_293_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_293_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_293_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_293_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_293_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_293_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_293_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_294_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_294_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_294_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_294_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_294_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_294_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_294_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_294_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_295_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_295_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_295_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_295_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_295_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_295_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_295_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_295_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_296_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_296_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_296_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_296_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_296_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_296_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_296_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_296_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_297_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_297_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_297_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_297_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_297_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_297_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_297_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_297_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_298_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_298_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_298_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_298_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_298_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_298_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_298_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_298_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_299_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_299_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_299_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_299_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_299_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_299_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_299_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_299_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_300_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_300_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_300_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_300_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_300_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_300_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_300_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_300_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_301_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_301_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_301_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_301_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_301_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_301_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_301_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_301_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_302_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_302_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_302_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_302_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_302_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_302_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_302_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_302_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_303_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_303_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_303_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_303_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_303_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_303_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_303_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_303_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_304_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_304_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_304_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_304_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_304_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_304_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_304_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_304_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_305_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_305_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_305_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_305_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_305_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_305_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_305_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_305_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_306_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_306_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_306_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_306_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_306_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_306_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_306_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_306_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_307_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_307_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_307_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_307_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_307_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_307_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_307_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_307_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_308_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_308_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_308_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_308_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_308_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_308_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_308_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_308_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_309_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_309_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_309_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_309_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_309_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_309_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_309_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_309_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_310_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_310_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_310_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_310_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_310_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_310_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_310_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_310_io_out_2; // @[Multiplier.scala 130:25]
  wire  c32_16_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_16_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_16_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_16_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_16_io_out_1; // @[Multiplier.scala 125:25]
  wire  c53_311_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_311_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_311_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_311_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_311_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_311_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_311_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_311_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_312_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_312_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_312_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_312_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_312_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_312_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_312_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_312_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_313_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_313_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_313_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_313_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_313_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_313_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_313_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_313_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_314_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_314_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_314_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_314_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_314_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_314_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_314_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_314_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_315_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_315_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_315_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_315_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_315_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_315_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_315_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_315_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_316_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_316_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_316_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_316_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_316_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_316_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_316_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_316_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_317_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_317_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_317_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_317_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_317_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_317_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_317_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_317_io_out_2; // @[Multiplier.scala 130:25]
  wire  c32_17_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_17_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_17_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_17_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_17_io_out_1; // @[Multiplier.scala 125:25]
  wire  c53_318_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_318_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_318_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_318_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_318_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_318_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_318_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_318_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_319_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_319_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_319_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_319_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_319_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_319_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_319_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_319_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_320_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_320_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_320_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_320_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_320_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_320_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_320_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_320_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_321_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_321_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_321_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_321_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_321_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_321_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_321_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_321_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_322_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_322_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_322_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_322_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_322_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_322_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_322_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_322_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_323_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_323_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_323_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_323_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_323_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_323_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_323_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_323_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_324_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_324_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_324_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_324_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_324_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_324_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_324_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_324_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_16_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_16_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_16_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_16_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_325_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_325_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_325_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_325_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_325_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_325_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_325_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_325_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_326_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_326_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_326_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_326_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_326_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_326_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_326_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_326_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_327_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_327_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_327_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_327_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_327_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_327_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_327_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_327_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_328_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_328_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_328_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_328_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_328_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_328_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_328_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_328_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_329_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_329_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_329_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_329_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_329_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_329_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_329_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_329_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_330_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_330_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_330_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_330_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_330_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_330_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_330_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_330_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_331_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_331_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_331_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_331_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_331_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_331_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_331_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_331_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_17_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_17_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_17_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_17_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_332_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_332_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_332_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_332_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_332_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_332_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_332_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_332_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_333_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_333_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_333_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_333_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_333_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_333_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_333_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_333_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_334_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_334_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_334_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_334_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_334_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_334_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_334_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_334_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_335_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_335_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_335_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_335_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_335_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_335_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_335_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_335_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_336_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_336_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_336_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_336_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_336_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_336_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_336_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_336_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_337_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_337_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_337_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_337_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_337_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_337_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_337_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_337_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_338_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_338_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_338_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_338_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_338_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_338_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_338_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_338_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_339_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_339_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_339_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_339_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_339_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_339_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_339_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_339_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_340_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_340_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_340_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_340_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_340_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_340_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_340_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_340_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_341_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_341_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_341_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_341_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_341_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_341_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_341_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_341_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_342_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_342_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_342_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_342_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_342_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_342_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_342_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_342_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_343_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_343_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_343_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_343_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_343_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_343_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_343_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_343_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_344_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_344_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_344_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_344_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_344_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_344_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_344_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_344_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_345_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_345_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_345_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_345_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_345_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_345_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_345_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_345_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_346_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_346_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_346_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_346_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_346_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_346_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_346_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_346_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_347_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_347_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_347_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_347_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_347_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_347_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_347_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_347_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_348_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_348_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_348_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_348_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_348_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_348_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_348_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_348_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_349_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_349_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_349_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_349_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_349_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_349_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_349_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_349_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_350_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_350_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_350_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_350_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_350_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_350_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_350_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_350_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_351_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_351_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_351_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_351_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_351_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_351_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_351_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_351_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_352_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_352_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_352_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_352_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_352_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_352_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_352_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_352_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_353_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_353_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_353_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_353_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_353_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_353_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_353_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_353_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_354_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_354_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_354_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_354_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_354_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_354_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_354_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_354_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_355_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_355_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_355_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_355_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_355_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_355_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_355_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_355_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_356_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_356_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_356_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_356_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_356_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_356_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_356_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_356_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_357_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_357_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_357_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_357_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_357_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_357_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_357_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_357_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_358_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_358_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_358_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_358_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_358_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_358_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_358_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_358_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_359_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_359_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_359_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_359_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_359_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_359_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_359_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_359_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_360_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_360_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_360_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_360_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_360_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_360_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_360_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_360_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_361_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_361_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_361_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_361_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_361_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_361_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_361_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_361_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_362_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_362_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_362_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_362_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_362_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_362_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_362_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_362_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_363_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_363_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_363_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_363_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_363_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_363_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_363_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_363_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_364_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_364_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_364_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_364_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_364_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_364_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_364_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_364_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_365_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_365_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_365_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_365_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_365_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_365_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_365_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_365_io_out_2; // @[Multiplier.scala 130:25]
  wire  c32_18_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_18_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_18_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_18_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_18_io_out_1; // @[Multiplier.scala 125:25]
  wire  c53_366_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_366_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_366_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_366_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_366_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_366_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_366_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_366_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_367_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_367_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_367_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_367_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_367_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_367_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_367_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_367_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_368_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_368_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_368_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_368_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_368_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_368_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_368_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_368_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_369_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_369_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_369_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_369_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_369_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_369_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_369_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_369_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_370_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_370_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_370_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_370_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_370_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_370_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_370_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_370_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_371_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_371_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_371_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_371_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_371_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_371_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_371_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_371_io_out_2; // @[Multiplier.scala 130:25]
  wire  c32_19_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_19_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_19_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_19_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_19_io_out_1; // @[Multiplier.scala 125:25]
  wire  c53_372_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_372_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_372_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_372_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_372_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_372_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_372_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_372_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_373_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_373_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_373_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_373_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_373_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_373_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_373_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_373_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_374_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_374_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_374_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_374_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_374_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_374_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_374_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_374_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_375_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_375_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_375_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_375_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_375_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_375_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_375_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_375_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_376_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_376_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_376_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_376_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_376_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_376_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_376_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_376_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_377_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_377_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_377_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_377_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_377_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_377_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_377_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_377_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_18_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_18_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_18_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_18_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_378_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_378_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_378_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_378_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_378_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_378_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_378_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_378_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_379_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_379_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_379_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_379_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_379_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_379_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_379_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_379_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_380_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_380_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_380_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_380_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_380_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_380_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_380_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_380_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_381_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_381_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_381_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_381_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_381_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_381_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_381_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_381_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_382_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_382_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_382_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_382_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_382_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_382_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_382_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_382_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_383_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_383_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_383_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_383_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_383_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_383_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_383_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_383_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_19_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_19_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_19_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_19_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_384_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_384_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_384_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_384_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_384_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_384_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_384_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_384_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_385_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_385_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_385_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_385_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_385_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_385_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_385_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_385_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_386_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_386_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_386_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_386_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_386_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_386_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_386_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_386_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_387_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_387_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_387_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_387_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_387_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_387_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_387_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_387_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_388_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_388_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_388_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_388_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_388_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_388_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_388_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_388_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_389_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_389_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_389_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_389_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_389_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_389_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_389_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_389_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_390_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_390_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_390_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_390_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_390_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_390_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_390_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_390_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_391_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_391_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_391_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_391_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_391_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_391_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_391_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_391_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_392_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_392_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_392_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_392_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_392_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_392_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_392_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_392_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_393_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_393_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_393_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_393_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_393_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_393_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_393_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_393_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_394_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_394_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_394_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_394_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_394_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_394_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_394_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_394_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_395_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_395_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_395_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_395_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_395_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_395_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_395_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_395_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_396_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_396_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_396_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_396_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_396_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_396_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_396_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_396_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_397_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_397_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_397_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_397_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_397_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_397_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_397_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_397_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_398_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_398_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_398_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_398_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_398_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_398_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_398_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_398_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_399_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_399_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_399_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_399_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_399_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_399_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_399_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_399_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_400_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_400_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_400_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_400_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_400_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_400_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_400_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_400_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_401_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_401_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_401_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_401_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_401_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_401_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_401_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_401_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_402_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_402_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_402_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_402_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_402_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_402_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_402_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_402_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_403_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_403_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_403_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_403_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_403_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_403_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_403_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_403_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_404_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_404_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_404_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_404_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_404_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_404_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_404_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_404_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_405_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_405_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_405_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_405_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_405_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_405_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_405_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_405_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_406_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_406_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_406_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_406_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_406_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_406_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_406_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_406_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_407_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_407_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_407_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_407_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_407_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_407_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_407_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_407_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_408_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_408_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_408_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_408_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_408_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_408_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_408_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_408_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_409_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_409_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_409_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_409_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_409_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_409_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_409_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_409_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_410_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_410_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_410_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_410_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_410_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_410_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_410_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_410_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_411_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_411_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_411_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_411_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_411_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_411_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_411_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_411_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_412_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_412_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_412_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_412_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_412_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_412_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_412_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_412_io_out_2; // @[Multiplier.scala 130:25]
  wire  c32_20_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_20_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_20_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_20_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_20_io_out_1; // @[Multiplier.scala 125:25]
  wire  c53_413_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_413_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_413_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_413_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_413_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_413_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_413_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_413_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_414_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_414_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_414_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_414_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_414_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_414_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_414_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_414_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_415_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_415_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_415_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_415_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_415_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_415_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_415_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_415_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_416_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_416_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_416_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_416_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_416_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_416_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_416_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_416_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_417_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_417_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_417_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_417_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_417_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_417_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_417_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_417_io_out_2; // @[Multiplier.scala 130:25]
  wire  c32_21_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_21_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_21_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_21_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_21_io_out_1; // @[Multiplier.scala 125:25]
  wire  c53_418_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_418_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_418_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_418_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_418_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_418_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_418_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_418_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_419_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_419_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_419_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_419_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_419_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_419_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_419_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_419_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_420_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_420_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_420_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_420_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_420_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_420_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_420_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_420_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_421_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_421_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_421_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_421_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_421_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_421_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_421_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_421_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_422_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_422_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_422_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_422_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_422_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_422_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_422_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_422_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_20_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_20_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_20_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_20_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_423_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_423_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_423_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_423_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_423_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_423_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_423_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_423_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_424_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_424_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_424_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_424_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_424_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_424_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_424_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_424_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_425_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_425_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_425_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_425_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_425_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_425_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_425_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_425_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_426_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_426_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_426_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_426_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_426_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_426_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_426_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_426_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_427_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_427_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_427_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_427_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_427_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_427_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_427_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_427_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_21_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_21_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_21_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_21_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_428_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_428_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_428_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_428_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_428_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_428_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_428_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_428_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_429_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_429_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_429_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_429_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_429_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_429_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_429_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_429_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_430_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_430_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_430_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_430_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_430_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_430_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_430_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_430_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_431_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_431_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_431_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_431_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_431_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_431_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_431_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_431_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_432_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_432_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_432_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_432_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_432_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_432_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_432_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_432_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_433_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_433_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_433_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_433_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_433_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_433_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_433_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_433_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_434_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_434_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_434_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_434_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_434_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_434_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_434_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_434_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_435_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_435_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_435_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_435_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_435_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_435_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_435_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_435_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_436_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_436_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_436_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_436_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_436_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_436_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_436_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_436_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_437_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_437_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_437_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_437_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_437_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_437_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_437_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_437_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_438_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_438_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_438_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_438_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_438_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_438_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_438_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_438_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_439_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_439_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_439_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_439_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_439_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_439_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_439_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_439_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_440_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_440_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_440_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_440_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_440_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_440_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_440_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_440_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_441_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_441_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_441_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_441_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_441_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_441_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_441_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_441_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_442_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_442_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_442_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_442_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_442_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_442_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_442_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_442_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_443_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_443_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_443_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_443_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_443_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_443_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_443_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_443_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_444_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_444_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_444_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_444_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_444_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_444_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_444_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_444_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_445_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_445_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_445_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_445_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_445_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_445_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_445_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_445_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_446_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_446_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_446_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_446_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_446_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_446_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_446_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_446_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_447_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_447_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_447_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_447_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_447_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_447_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_447_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_447_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_448_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_448_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_448_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_448_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_448_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_448_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_448_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_448_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_449_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_449_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_449_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_449_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_449_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_449_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_449_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_449_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_450_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_450_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_450_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_450_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_450_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_450_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_450_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_450_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_451_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_451_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_451_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_451_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_451_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_451_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_451_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_451_io_out_2; // @[Multiplier.scala 130:25]
  wire  c32_22_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_22_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_22_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_22_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_22_io_out_1; // @[Multiplier.scala 125:25]
  wire  c53_452_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_452_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_452_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_452_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_452_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_452_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_452_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_452_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_453_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_453_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_453_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_453_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_453_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_453_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_453_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_453_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_454_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_454_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_454_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_454_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_454_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_454_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_454_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_454_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_455_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_455_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_455_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_455_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_455_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_455_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_455_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_455_io_out_2; // @[Multiplier.scala 130:25]
  wire  c32_23_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_23_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_23_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_23_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_23_io_out_1; // @[Multiplier.scala 125:25]
  wire  c53_456_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_456_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_456_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_456_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_456_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_456_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_456_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_456_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_457_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_457_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_457_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_457_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_457_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_457_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_457_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_457_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_458_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_458_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_458_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_458_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_458_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_458_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_458_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_458_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_459_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_459_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_459_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_459_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_459_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_459_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_459_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_459_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_22_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_22_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_22_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_22_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_460_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_460_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_460_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_460_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_460_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_460_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_460_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_460_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_461_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_461_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_461_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_461_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_461_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_461_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_461_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_461_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_462_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_462_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_462_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_462_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_462_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_462_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_462_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_462_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_463_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_463_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_463_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_463_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_463_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_463_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_463_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_463_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_23_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_23_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_23_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_23_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_464_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_464_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_464_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_464_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_464_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_464_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_464_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_464_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_465_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_465_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_465_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_465_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_465_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_465_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_465_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_465_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_466_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_466_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_466_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_466_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_466_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_466_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_466_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_466_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_467_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_467_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_467_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_467_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_467_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_467_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_467_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_467_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_468_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_468_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_468_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_468_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_468_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_468_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_468_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_468_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_469_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_469_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_469_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_469_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_469_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_469_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_469_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_469_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_470_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_470_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_470_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_470_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_470_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_470_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_470_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_470_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_471_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_471_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_471_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_471_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_471_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_471_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_471_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_471_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_472_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_472_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_472_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_472_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_472_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_472_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_472_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_472_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_473_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_473_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_473_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_473_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_473_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_473_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_473_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_473_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_474_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_474_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_474_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_474_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_474_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_474_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_474_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_474_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_475_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_475_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_475_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_475_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_475_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_475_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_475_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_475_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_476_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_476_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_476_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_476_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_476_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_476_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_476_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_476_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_477_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_477_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_477_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_477_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_477_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_477_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_477_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_477_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_478_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_478_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_478_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_478_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_478_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_478_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_478_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_478_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_479_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_479_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_479_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_479_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_479_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_479_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_479_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_479_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_480_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_480_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_480_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_480_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_480_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_480_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_480_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_480_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_481_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_481_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_481_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_481_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_481_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_481_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_481_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_481_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_482_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_482_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_482_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_482_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_482_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_482_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_482_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_482_io_out_2; // @[Multiplier.scala 130:25]
  wire  c32_24_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_24_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_24_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_24_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_24_io_out_1; // @[Multiplier.scala 125:25]
  wire  c53_483_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_483_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_483_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_483_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_483_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_483_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_483_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_483_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_484_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_484_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_484_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_484_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_484_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_484_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_484_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_484_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_485_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_485_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_485_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_485_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_485_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_485_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_485_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_485_io_out_2; // @[Multiplier.scala 130:25]
  wire  c32_25_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_25_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_25_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_25_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_25_io_out_1; // @[Multiplier.scala 125:25]
  wire  c53_486_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_486_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_486_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_486_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_486_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_486_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_486_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_486_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_487_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_487_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_487_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_487_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_487_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_487_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_487_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_487_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_488_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_488_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_488_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_488_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_488_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_488_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_488_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_488_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_24_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_24_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_24_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_24_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_489_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_489_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_489_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_489_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_489_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_489_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_489_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_489_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_490_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_490_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_490_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_490_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_490_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_490_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_490_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_490_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_491_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_491_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_491_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_491_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_491_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_491_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_491_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_491_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_25_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_25_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_25_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_25_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_492_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_492_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_492_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_492_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_492_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_492_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_492_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_492_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_493_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_493_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_493_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_493_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_493_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_493_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_493_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_493_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_494_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_494_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_494_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_494_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_494_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_494_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_494_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_494_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_495_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_495_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_495_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_495_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_495_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_495_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_495_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_495_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_496_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_496_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_496_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_496_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_496_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_496_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_496_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_496_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_497_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_497_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_497_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_497_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_497_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_497_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_497_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_497_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_498_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_498_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_498_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_498_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_498_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_498_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_498_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_498_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_499_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_499_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_499_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_499_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_499_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_499_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_499_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_499_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_500_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_500_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_500_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_500_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_500_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_500_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_500_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_500_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_501_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_501_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_501_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_501_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_501_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_501_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_501_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_501_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_502_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_502_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_502_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_502_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_502_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_502_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_502_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_502_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_503_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_503_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_503_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_503_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_503_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_503_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_503_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_503_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_504_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_504_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_504_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_504_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_504_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_504_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_504_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_504_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_505_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_505_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_505_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_505_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_505_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_505_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_505_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_505_io_out_2; // @[Multiplier.scala 130:25]
  wire  c32_26_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_26_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_26_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_26_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_26_io_out_1; // @[Multiplier.scala 125:25]
  wire  c53_506_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_506_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_506_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_506_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_506_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_506_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_506_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_506_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_507_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_507_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_507_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_507_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_507_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_507_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_507_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_507_io_out_2; // @[Multiplier.scala 130:25]
  wire  c32_27_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_27_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_27_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_27_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_27_io_out_1; // @[Multiplier.scala 125:25]
  wire  c53_508_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_508_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_508_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_508_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_508_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_508_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_508_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_508_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_509_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_509_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_509_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_509_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_509_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_509_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_509_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_509_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_26_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_26_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_26_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_26_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_510_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_510_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_510_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_510_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_510_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_510_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_510_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_510_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_511_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_511_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_511_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_511_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_511_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_511_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_511_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_511_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_27_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_27_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_27_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_27_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_512_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_512_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_512_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_512_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_512_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_512_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_512_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_512_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_513_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_513_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_513_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_513_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_513_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_513_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_513_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_513_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_514_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_514_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_514_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_514_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_514_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_514_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_514_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_514_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_515_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_515_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_515_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_515_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_515_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_515_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_515_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_515_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_516_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_516_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_516_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_516_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_516_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_516_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_516_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_516_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_517_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_517_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_517_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_517_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_517_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_517_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_517_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_517_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_518_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_518_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_518_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_518_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_518_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_518_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_518_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_518_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_519_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_519_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_519_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_519_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_519_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_519_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_519_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_519_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_520_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_520_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_520_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_520_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_520_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_520_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_520_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_520_io_out_2; // @[Multiplier.scala 130:25]
  wire  c32_28_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_28_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_28_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_28_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_28_io_out_1; // @[Multiplier.scala 125:25]
  wire  c53_521_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_521_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_521_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_521_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_521_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_521_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_521_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_521_io_out_2; // @[Multiplier.scala 130:25]
  wire  c32_29_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_29_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_29_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_29_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_29_io_out_1; // @[Multiplier.scala 125:25]
  wire  c53_522_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_522_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_522_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_522_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_522_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_522_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_522_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_522_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_28_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_28_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_28_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_28_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_523_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_523_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_523_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_523_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_523_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_523_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_523_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_523_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_29_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_29_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_29_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_29_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_524_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_524_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_524_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_524_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_524_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_524_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_524_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_524_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_525_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_525_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_525_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_525_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_525_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_525_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_525_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_525_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_526_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_526_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_526_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_526_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_526_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_526_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_526_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_526_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_527_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_527_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_527_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_527_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_527_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_527_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_527_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_527_io_out_2; // @[Multiplier.scala 130:25]
  wire  c32_30_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_30_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_30_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_30_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_30_io_out_1; // @[Multiplier.scala 125:25]
  wire  c32_31_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_31_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_31_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_31_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_31_io_out_1; // @[Multiplier.scala 125:25]
  wire  c22_30_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_30_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_30_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_30_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_31_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_31_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_31_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_31_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_32_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_32_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_32_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_32_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_33_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_33_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_33_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_33_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_34_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_34_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_34_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_34_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_35_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_35_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_35_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_35_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_36_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_36_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_36_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_36_io_out_1; // @[Multiplier.scala 120:25]
  wire  c32_32_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_32_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_32_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_32_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_32_io_out_1; // @[Multiplier.scala 125:25]
  wire  c32_33_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_33_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_33_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_33_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_33_io_out_1; // @[Multiplier.scala 125:25]
  wire  c32_34_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_34_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_34_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_34_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_34_io_out_1; // @[Multiplier.scala 125:25]
  wire  c53_528_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_528_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_528_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_528_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_528_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_528_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_528_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_528_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_529_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_529_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_529_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_529_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_529_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_529_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_529_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_529_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_530_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_530_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_530_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_530_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_530_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_530_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_530_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_530_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_531_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_531_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_531_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_531_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_531_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_531_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_531_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_531_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_532_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_532_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_532_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_532_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_532_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_532_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_532_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_532_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_533_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_533_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_533_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_533_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_533_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_533_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_533_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_533_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_534_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_534_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_534_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_534_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_534_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_534_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_534_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_534_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_535_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_535_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_535_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_535_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_535_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_535_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_535_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_535_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_536_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_536_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_536_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_536_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_536_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_536_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_536_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_536_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_37_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_37_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_37_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_37_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_537_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_537_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_537_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_537_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_537_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_537_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_537_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_537_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_38_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_38_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_38_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_38_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_538_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_538_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_538_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_538_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_538_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_538_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_538_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_538_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_39_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_39_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_39_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_39_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_539_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_539_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_539_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_539_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_539_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_539_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_539_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_539_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_40_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_40_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_40_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_40_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_540_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_540_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_540_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_540_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_540_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_540_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_540_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_540_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_41_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_41_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_41_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_41_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_541_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_541_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_541_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_541_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_541_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_541_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_541_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_541_io_out_2; // @[Multiplier.scala 130:25]
  wire  c32_35_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_35_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_35_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_35_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_35_io_out_1; // @[Multiplier.scala 125:25]
  wire  c53_542_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_542_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_542_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_542_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_542_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_542_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_542_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_542_io_out_2; // @[Multiplier.scala 130:25]
  wire  c32_36_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_36_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_36_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_36_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_36_io_out_1; // @[Multiplier.scala 125:25]
  wire  c53_543_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_543_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_543_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_543_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_543_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_543_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_543_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_543_io_out_2; // @[Multiplier.scala 130:25]
  wire  c32_37_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_37_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_37_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_37_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_37_io_out_1; // @[Multiplier.scala 125:25]
  wire  c53_544_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_544_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_544_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_544_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_544_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_544_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_544_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_544_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_545_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_545_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_545_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_545_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_545_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_545_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_545_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_545_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_546_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_546_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_546_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_546_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_546_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_546_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_546_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_546_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_547_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_547_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_547_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_547_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_547_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_547_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_547_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_547_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_548_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_548_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_548_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_548_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_548_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_548_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_548_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_548_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_549_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_549_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_549_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_549_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_549_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_549_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_549_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_549_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_550_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_550_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_550_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_550_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_550_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_550_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_550_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_550_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_551_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_551_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_551_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_551_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_551_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_551_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_551_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_551_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_552_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_552_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_552_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_552_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_552_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_552_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_552_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_552_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_553_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_553_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_553_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_553_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_553_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_553_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_553_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_553_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_554_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_554_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_554_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_554_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_554_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_554_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_554_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_554_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_555_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_555_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_555_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_555_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_555_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_555_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_555_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_555_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_556_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_556_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_556_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_556_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_556_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_556_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_556_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_556_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_557_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_557_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_557_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_557_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_557_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_557_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_557_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_557_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_558_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_558_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_558_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_558_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_558_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_558_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_558_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_558_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_559_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_559_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_559_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_559_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_559_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_559_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_559_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_559_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_560_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_560_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_560_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_560_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_560_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_560_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_560_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_560_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_561_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_561_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_561_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_561_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_561_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_561_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_561_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_561_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_42_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_42_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_42_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_42_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_562_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_562_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_562_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_562_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_562_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_562_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_562_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_562_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_563_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_563_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_563_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_563_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_563_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_563_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_563_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_563_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_43_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_43_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_43_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_43_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_564_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_564_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_564_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_564_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_564_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_564_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_564_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_564_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_565_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_565_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_565_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_565_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_565_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_565_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_565_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_565_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_44_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_44_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_44_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_44_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_566_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_566_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_566_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_566_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_566_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_566_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_566_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_566_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_567_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_567_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_567_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_567_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_567_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_567_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_567_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_567_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_45_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_45_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_45_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_45_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_568_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_568_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_568_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_568_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_568_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_568_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_568_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_568_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_569_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_569_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_569_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_569_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_569_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_569_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_569_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_569_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_46_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_46_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_46_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_46_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_570_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_570_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_570_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_570_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_570_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_570_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_570_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_570_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_571_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_571_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_571_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_571_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_571_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_571_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_571_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_571_io_out_2; // @[Multiplier.scala 130:25]
  wire  c32_38_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_38_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_38_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_38_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_38_io_out_1; // @[Multiplier.scala 125:25]
  wire  c53_572_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_572_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_572_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_572_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_572_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_572_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_572_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_572_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_573_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_573_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_573_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_573_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_573_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_573_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_573_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_573_io_out_2; // @[Multiplier.scala 130:25]
  wire  c32_39_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_39_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_39_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_39_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_39_io_out_1; // @[Multiplier.scala 125:25]
  wire  c53_574_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_574_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_574_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_574_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_574_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_574_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_574_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_574_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_575_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_575_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_575_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_575_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_575_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_575_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_575_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_575_io_out_2; // @[Multiplier.scala 130:25]
  wire  c32_40_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_40_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_40_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_40_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_40_io_out_1; // @[Multiplier.scala 125:25]
  wire  c53_576_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_576_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_576_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_576_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_576_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_576_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_576_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_576_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_577_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_577_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_577_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_577_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_577_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_577_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_577_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_577_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_578_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_578_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_578_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_578_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_578_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_578_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_578_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_578_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_579_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_579_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_579_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_579_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_579_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_579_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_579_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_579_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_580_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_580_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_580_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_580_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_580_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_580_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_580_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_580_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_581_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_581_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_581_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_581_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_581_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_581_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_581_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_581_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_582_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_582_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_582_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_582_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_582_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_582_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_582_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_582_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_583_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_583_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_583_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_583_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_583_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_583_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_583_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_583_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_584_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_584_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_584_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_584_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_584_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_584_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_584_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_584_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_585_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_585_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_585_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_585_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_585_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_585_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_585_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_585_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_586_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_586_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_586_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_586_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_586_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_586_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_586_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_586_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_587_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_587_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_587_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_587_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_587_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_587_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_587_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_587_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_588_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_588_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_588_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_588_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_588_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_588_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_588_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_588_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_589_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_589_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_589_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_589_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_589_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_589_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_589_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_589_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_590_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_590_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_590_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_590_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_590_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_590_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_590_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_590_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_591_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_591_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_591_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_591_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_591_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_591_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_591_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_591_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_592_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_592_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_592_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_592_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_592_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_592_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_592_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_592_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_593_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_593_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_593_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_593_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_593_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_593_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_593_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_593_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_594_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_594_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_594_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_594_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_594_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_594_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_594_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_594_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_595_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_595_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_595_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_595_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_595_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_595_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_595_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_595_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_596_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_596_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_596_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_596_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_596_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_596_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_596_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_596_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_597_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_597_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_597_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_597_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_597_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_597_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_597_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_597_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_598_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_598_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_598_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_598_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_598_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_598_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_598_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_598_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_599_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_599_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_599_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_599_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_599_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_599_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_599_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_599_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_600_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_600_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_600_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_600_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_600_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_600_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_600_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_600_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_601_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_601_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_601_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_601_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_601_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_601_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_601_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_601_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_602_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_602_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_602_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_602_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_602_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_602_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_602_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_602_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_47_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_47_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_47_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_47_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_603_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_603_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_603_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_603_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_603_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_603_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_603_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_603_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_604_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_604_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_604_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_604_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_604_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_604_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_604_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_604_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_605_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_605_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_605_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_605_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_605_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_605_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_605_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_605_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_48_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_48_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_48_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_48_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_606_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_606_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_606_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_606_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_606_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_606_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_606_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_606_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_607_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_607_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_607_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_607_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_607_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_607_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_607_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_607_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_608_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_608_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_608_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_608_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_608_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_608_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_608_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_608_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_49_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_49_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_49_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_49_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_609_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_609_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_609_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_609_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_609_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_609_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_609_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_609_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_610_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_610_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_610_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_610_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_610_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_610_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_610_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_610_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_611_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_611_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_611_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_611_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_611_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_611_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_611_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_611_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_50_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_50_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_50_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_50_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_612_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_612_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_612_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_612_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_612_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_612_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_612_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_612_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_613_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_613_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_613_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_613_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_613_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_613_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_613_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_613_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_614_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_614_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_614_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_614_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_614_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_614_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_614_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_614_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_51_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_51_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_51_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_51_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_615_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_615_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_615_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_615_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_615_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_615_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_615_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_615_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_616_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_616_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_616_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_616_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_616_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_616_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_616_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_616_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_617_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_617_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_617_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_617_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_617_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_617_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_617_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_617_io_out_2; // @[Multiplier.scala 130:25]
  wire  c32_41_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_41_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_41_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_41_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_41_io_out_1; // @[Multiplier.scala 125:25]
  wire  c53_618_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_618_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_618_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_618_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_618_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_618_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_618_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_618_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_619_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_619_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_619_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_619_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_619_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_619_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_619_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_619_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_620_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_620_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_620_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_620_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_620_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_620_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_620_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_620_io_out_2; // @[Multiplier.scala 130:25]
  wire  c32_42_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_42_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_42_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_42_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_42_io_out_1; // @[Multiplier.scala 125:25]
  wire  c53_621_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_621_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_621_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_621_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_621_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_621_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_621_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_621_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_622_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_622_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_622_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_622_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_622_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_622_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_622_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_622_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_623_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_623_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_623_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_623_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_623_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_623_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_623_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_623_io_out_2; // @[Multiplier.scala 130:25]
  wire  c32_43_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_43_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_43_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_43_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_43_io_out_1; // @[Multiplier.scala 125:25]
  wire  c53_624_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_624_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_624_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_624_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_624_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_624_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_624_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_624_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_625_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_625_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_625_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_625_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_625_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_625_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_625_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_625_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_626_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_626_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_626_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_626_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_626_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_626_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_626_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_626_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_627_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_627_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_627_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_627_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_627_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_627_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_627_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_627_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_628_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_628_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_628_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_628_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_628_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_628_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_628_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_628_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_629_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_629_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_629_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_629_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_629_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_629_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_629_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_629_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_630_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_630_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_630_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_630_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_630_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_630_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_630_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_630_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_631_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_631_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_631_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_631_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_631_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_631_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_631_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_631_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_632_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_632_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_632_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_632_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_632_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_632_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_632_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_632_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_633_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_633_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_633_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_633_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_633_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_633_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_633_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_633_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_634_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_634_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_634_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_634_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_634_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_634_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_634_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_634_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_635_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_635_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_635_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_635_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_635_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_635_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_635_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_635_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_636_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_636_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_636_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_636_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_636_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_636_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_636_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_636_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_637_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_637_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_637_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_637_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_637_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_637_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_637_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_637_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_638_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_638_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_638_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_638_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_638_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_638_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_638_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_638_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_639_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_639_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_639_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_639_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_639_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_639_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_639_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_639_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_640_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_640_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_640_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_640_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_640_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_640_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_640_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_640_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_641_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_641_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_641_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_641_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_641_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_641_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_641_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_641_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_642_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_642_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_642_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_642_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_642_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_642_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_642_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_642_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_643_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_643_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_643_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_643_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_643_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_643_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_643_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_643_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_644_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_644_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_644_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_644_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_644_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_644_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_644_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_644_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_645_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_645_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_645_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_645_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_645_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_645_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_645_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_645_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_646_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_646_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_646_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_646_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_646_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_646_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_646_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_646_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_647_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_647_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_647_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_647_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_647_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_647_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_647_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_647_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_648_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_648_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_648_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_648_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_648_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_648_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_648_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_648_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_649_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_649_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_649_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_649_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_649_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_649_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_649_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_649_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_650_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_650_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_650_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_650_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_650_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_650_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_650_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_650_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_651_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_651_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_651_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_651_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_651_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_651_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_651_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_651_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_652_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_652_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_652_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_652_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_652_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_652_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_652_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_652_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_653_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_653_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_653_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_653_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_653_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_653_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_653_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_653_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_654_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_654_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_654_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_654_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_654_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_654_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_654_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_654_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_655_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_655_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_655_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_655_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_655_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_655_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_655_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_655_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_656_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_656_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_656_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_656_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_656_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_656_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_656_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_656_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_657_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_657_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_657_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_657_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_657_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_657_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_657_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_657_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_658_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_658_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_658_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_658_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_658_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_658_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_658_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_658_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_659_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_659_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_659_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_659_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_659_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_659_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_659_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_659_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_660_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_660_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_660_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_660_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_660_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_660_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_660_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_660_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_661_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_661_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_661_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_661_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_661_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_661_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_661_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_661_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_662_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_662_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_662_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_662_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_662_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_662_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_662_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_662_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_663_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_663_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_663_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_663_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_663_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_663_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_663_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_663_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_664_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_664_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_664_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_664_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_664_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_664_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_664_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_664_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_665_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_665_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_665_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_665_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_665_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_665_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_665_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_665_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_666_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_666_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_666_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_666_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_666_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_666_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_666_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_666_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_667_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_667_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_667_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_667_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_667_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_667_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_667_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_667_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_668_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_668_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_668_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_668_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_668_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_668_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_668_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_668_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_669_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_669_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_669_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_669_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_669_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_669_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_669_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_669_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_670_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_670_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_670_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_670_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_670_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_670_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_670_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_670_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_671_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_671_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_671_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_671_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_671_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_671_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_671_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_671_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_672_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_672_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_672_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_672_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_672_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_672_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_672_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_672_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_673_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_673_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_673_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_673_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_673_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_673_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_673_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_673_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_674_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_674_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_674_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_674_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_674_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_674_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_674_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_674_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_675_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_675_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_675_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_675_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_675_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_675_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_675_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_675_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_676_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_676_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_676_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_676_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_676_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_676_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_676_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_676_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_677_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_677_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_677_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_677_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_677_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_677_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_677_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_677_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_678_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_678_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_678_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_678_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_678_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_678_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_678_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_678_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_679_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_679_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_679_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_679_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_679_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_679_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_679_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_679_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_680_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_680_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_680_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_680_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_680_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_680_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_680_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_680_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_681_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_681_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_681_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_681_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_681_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_681_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_681_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_681_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_682_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_682_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_682_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_682_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_682_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_682_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_682_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_682_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_683_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_683_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_683_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_683_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_683_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_683_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_683_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_683_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_684_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_684_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_684_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_684_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_684_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_684_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_684_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_684_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_685_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_685_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_685_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_685_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_685_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_685_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_685_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_685_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_686_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_686_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_686_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_686_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_686_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_686_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_686_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_686_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_687_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_687_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_687_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_687_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_687_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_687_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_687_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_687_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_688_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_688_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_688_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_688_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_688_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_688_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_688_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_688_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_689_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_689_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_689_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_689_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_689_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_689_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_689_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_689_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_690_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_690_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_690_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_690_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_690_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_690_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_690_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_690_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_691_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_691_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_691_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_691_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_691_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_691_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_691_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_691_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_692_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_692_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_692_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_692_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_692_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_692_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_692_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_692_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_693_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_693_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_693_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_693_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_693_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_693_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_693_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_693_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_694_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_694_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_694_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_694_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_694_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_694_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_694_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_694_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_695_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_695_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_695_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_695_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_695_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_695_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_695_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_695_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_696_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_696_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_696_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_696_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_696_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_696_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_696_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_696_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_697_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_697_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_697_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_697_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_697_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_697_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_697_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_697_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_698_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_698_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_698_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_698_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_698_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_698_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_698_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_698_io_out_2; // @[Multiplier.scala 130:25]
  wire  c32_44_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_44_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_44_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_44_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_44_io_out_1; // @[Multiplier.scala 125:25]
  wire  c53_699_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_699_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_699_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_699_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_699_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_699_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_699_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_699_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_700_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_700_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_700_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_700_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_700_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_700_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_700_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_700_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_701_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_701_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_701_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_701_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_701_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_701_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_701_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_701_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_52_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_52_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_52_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_52_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_702_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_702_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_702_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_702_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_702_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_702_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_702_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_702_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_703_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_703_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_703_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_703_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_703_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_703_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_703_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_703_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_704_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_704_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_704_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_704_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_704_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_704_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_704_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_704_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_53_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_53_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_53_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_53_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_705_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_705_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_705_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_705_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_705_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_705_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_705_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_705_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_706_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_706_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_706_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_706_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_706_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_706_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_706_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_706_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_707_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_707_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_707_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_707_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_707_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_707_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_707_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_707_io_out_2; // @[Multiplier.scala 130:25]
  wire  c32_45_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_45_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_45_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_45_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_45_io_out_1; // @[Multiplier.scala 125:25]
  wire  c53_708_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_708_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_708_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_708_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_708_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_708_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_708_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_708_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_709_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_709_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_709_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_709_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_709_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_709_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_709_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_709_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_710_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_710_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_710_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_710_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_710_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_710_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_710_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_710_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_54_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_54_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_54_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_54_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_711_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_711_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_711_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_711_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_711_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_711_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_711_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_711_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_712_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_712_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_712_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_712_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_712_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_712_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_712_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_712_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_713_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_713_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_713_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_713_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_713_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_713_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_713_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_713_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_55_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_55_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_55_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_55_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_714_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_714_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_714_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_714_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_714_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_714_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_714_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_714_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_715_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_715_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_715_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_715_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_715_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_715_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_715_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_715_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_716_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_716_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_716_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_716_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_716_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_716_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_716_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_716_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_56_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_56_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_56_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_56_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_717_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_717_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_717_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_717_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_717_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_717_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_717_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_717_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_718_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_718_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_718_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_718_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_718_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_718_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_718_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_718_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_719_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_719_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_719_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_719_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_719_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_719_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_719_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_719_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_57_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_57_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_57_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_57_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_720_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_720_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_720_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_720_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_720_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_720_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_720_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_720_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_721_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_721_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_721_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_721_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_721_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_721_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_721_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_721_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_722_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_722_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_722_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_722_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_722_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_722_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_722_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_722_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_723_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_723_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_723_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_723_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_723_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_723_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_723_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_723_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_724_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_724_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_724_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_724_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_724_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_724_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_724_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_724_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_725_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_725_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_725_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_725_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_725_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_725_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_725_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_725_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_726_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_726_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_726_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_726_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_726_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_726_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_726_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_726_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_727_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_727_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_727_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_727_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_727_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_727_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_727_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_727_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_728_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_728_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_728_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_728_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_728_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_728_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_728_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_728_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_729_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_729_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_729_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_729_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_729_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_729_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_729_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_729_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_730_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_730_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_730_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_730_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_730_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_730_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_730_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_730_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_731_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_731_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_731_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_731_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_731_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_731_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_731_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_731_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_732_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_732_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_732_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_732_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_732_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_732_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_732_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_732_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_733_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_733_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_733_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_733_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_733_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_733_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_733_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_733_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_734_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_734_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_734_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_734_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_734_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_734_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_734_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_734_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_735_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_735_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_735_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_735_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_735_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_735_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_735_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_735_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_736_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_736_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_736_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_736_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_736_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_736_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_736_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_736_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_737_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_737_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_737_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_737_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_737_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_737_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_737_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_737_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_738_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_738_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_738_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_738_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_738_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_738_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_738_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_738_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_739_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_739_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_739_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_739_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_739_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_739_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_739_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_739_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_740_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_740_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_740_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_740_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_740_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_740_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_740_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_740_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_741_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_741_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_741_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_741_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_741_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_741_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_741_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_741_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_742_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_742_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_742_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_742_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_742_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_742_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_742_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_742_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_743_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_743_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_743_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_743_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_743_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_743_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_743_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_743_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_744_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_744_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_744_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_744_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_744_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_744_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_744_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_744_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_745_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_745_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_745_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_745_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_745_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_745_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_745_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_745_io_out_2; // @[Multiplier.scala 130:25]
  wire  c32_46_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_46_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_46_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_46_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_46_io_out_1; // @[Multiplier.scala 125:25]
  wire  c53_746_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_746_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_746_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_746_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_746_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_746_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_746_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_746_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_747_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_747_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_747_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_747_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_747_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_747_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_747_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_747_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_58_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_58_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_58_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_58_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_748_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_748_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_748_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_748_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_748_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_748_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_748_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_748_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_749_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_749_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_749_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_749_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_749_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_749_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_749_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_749_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_59_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_59_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_59_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_59_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_750_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_750_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_750_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_750_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_750_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_750_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_750_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_750_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_751_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_751_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_751_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_751_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_751_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_751_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_751_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_751_io_out_2; // @[Multiplier.scala 130:25]
  wire  c32_47_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_47_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_47_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_47_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_47_io_out_1; // @[Multiplier.scala 125:25]
  wire  c53_752_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_752_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_752_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_752_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_752_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_752_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_752_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_752_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_753_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_753_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_753_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_753_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_753_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_753_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_753_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_753_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_60_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_60_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_60_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_60_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_754_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_754_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_754_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_754_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_754_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_754_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_754_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_754_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_755_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_755_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_755_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_755_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_755_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_755_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_755_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_755_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_61_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_61_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_61_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_61_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_756_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_756_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_756_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_756_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_756_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_756_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_756_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_756_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_757_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_757_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_757_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_757_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_757_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_757_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_757_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_757_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_62_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_62_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_62_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_62_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_758_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_758_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_758_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_758_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_758_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_758_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_758_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_758_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_759_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_759_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_759_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_759_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_759_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_759_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_759_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_759_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_63_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_63_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_63_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_63_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_760_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_760_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_760_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_760_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_760_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_760_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_760_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_760_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_761_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_761_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_761_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_761_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_761_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_761_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_761_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_761_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_762_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_762_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_762_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_762_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_762_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_762_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_762_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_762_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_763_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_763_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_763_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_763_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_763_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_763_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_763_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_763_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_764_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_764_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_764_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_764_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_764_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_764_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_764_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_764_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_765_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_765_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_765_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_765_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_765_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_765_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_765_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_765_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_766_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_766_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_766_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_766_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_766_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_766_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_766_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_766_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_767_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_767_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_767_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_767_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_767_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_767_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_767_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_767_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_768_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_768_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_768_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_768_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_768_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_768_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_768_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_768_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_769_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_769_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_769_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_769_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_769_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_769_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_769_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_769_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_770_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_770_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_770_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_770_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_770_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_770_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_770_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_770_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_771_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_771_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_771_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_771_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_771_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_771_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_771_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_771_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_772_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_772_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_772_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_772_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_772_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_772_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_772_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_772_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_773_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_773_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_773_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_773_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_773_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_773_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_773_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_773_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_774_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_774_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_774_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_774_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_774_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_774_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_774_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_774_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_775_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_775_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_775_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_775_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_775_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_775_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_775_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_775_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_776_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_776_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_776_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_776_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_776_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_776_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_776_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_776_io_out_2; // @[Multiplier.scala 130:25]
  wire  c32_48_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_48_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_48_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_48_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_48_io_out_1; // @[Multiplier.scala 125:25]
  wire  c53_777_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_777_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_777_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_777_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_777_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_777_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_777_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_777_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_64_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_64_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_64_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_64_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_778_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_778_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_778_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_778_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_778_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_778_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_778_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_778_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_65_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_65_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_65_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_65_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_779_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_779_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_779_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_779_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_779_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_779_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_779_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_779_io_out_2; // @[Multiplier.scala 130:25]
  wire  c32_49_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_49_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_49_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_49_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_49_io_out_1; // @[Multiplier.scala 125:25]
  wire  c53_780_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_780_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_780_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_780_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_780_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_780_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_780_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_780_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_66_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_66_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_66_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_66_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_781_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_781_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_781_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_781_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_781_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_781_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_781_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_781_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_67_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_67_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_67_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_67_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_782_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_782_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_782_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_782_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_782_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_782_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_782_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_782_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_68_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_68_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_68_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_68_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_783_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_783_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_783_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_783_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_783_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_783_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_783_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_783_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_69_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_69_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_69_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_69_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_784_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_784_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_784_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_784_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_784_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_784_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_784_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_784_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_785_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_785_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_785_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_785_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_785_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_785_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_785_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_785_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_786_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_786_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_786_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_786_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_786_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_786_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_786_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_786_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_787_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_787_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_787_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_787_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_787_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_787_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_787_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_787_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_788_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_788_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_788_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_788_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_788_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_788_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_788_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_788_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_789_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_789_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_789_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_789_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_789_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_789_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_789_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_789_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_790_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_790_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_790_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_790_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_790_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_790_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_790_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_790_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_791_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_791_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_791_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_791_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_791_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_791_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_791_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_791_io_out_2; // @[Multiplier.scala 130:25]
  wire  c32_50_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_50_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_50_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_50_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_50_io_out_1; // @[Multiplier.scala 125:25]
  wire  c22_70_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_70_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_70_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_70_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_71_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_71_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_71_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_71_io_out_1; // @[Multiplier.scala 120:25]
  wire  c32_51_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_51_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_51_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_51_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_51_io_out_1; // @[Multiplier.scala 125:25]
  wire  c22_72_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_72_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_72_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_72_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_73_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_73_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_73_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_73_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_74_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_74_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_74_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_74_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_75_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_75_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_75_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_75_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_76_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_76_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_76_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_76_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_77_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_77_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_77_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_77_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_78_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_78_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_78_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_78_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_79_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_79_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_79_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_79_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_80_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_80_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_80_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_80_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_81_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_81_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_81_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_81_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_82_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_82_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_82_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_82_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_83_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_83_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_83_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_83_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_84_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_84_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_84_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_84_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_85_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_85_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_85_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_85_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_86_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_86_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_86_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_86_io_out_1; // @[Multiplier.scala 120:25]
  wire  c32_52_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_52_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_52_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_52_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_52_io_out_1; // @[Multiplier.scala 125:25]
  wire  c32_53_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_53_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_53_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_53_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_53_io_out_1; // @[Multiplier.scala 125:25]
  wire  c32_54_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_54_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_54_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_54_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_54_io_out_1; // @[Multiplier.scala 125:25]
  wire  c32_55_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_55_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_55_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_55_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_55_io_out_1; // @[Multiplier.scala 125:25]
  wire  c53_792_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_792_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_792_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_792_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_792_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_792_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_792_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_792_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_793_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_793_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_793_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_793_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_793_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_793_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_793_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_793_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_794_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_794_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_794_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_794_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_794_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_794_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_794_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_794_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_795_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_795_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_795_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_795_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_795_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_795_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_795_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_795_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_796_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_796_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_796_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_796_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_796_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_796_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_796_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_796_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_797_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_797_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_797_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_797_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_797_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_797_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_797_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_797_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_798_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_798_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_798_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_798_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_798_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_798_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_798_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_798_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_799_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_799_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_799_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_799_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_799_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_799_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_799_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_799_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_800_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_800_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_800_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_800_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_800_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_800_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_800_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_800_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_801_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_801_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_801_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_801_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_801_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_801_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_801_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_801_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_802_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_802_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_802_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_802_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_802_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_802_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_802_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_802_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_803_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_803_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_803_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_803_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_803_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_803_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_803_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_803_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_804_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_804_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_804_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_804_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_804_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_804_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_804_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_804_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_805_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_805_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_805_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_805_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_805_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_805_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_805_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_805_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_806_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_806_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_806_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_806_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_806_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_806_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_806_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_806_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_807_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_807_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_807_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_807_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_807_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_807_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_807_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_807_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_808_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_808_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_808_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_808_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_808_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_808_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_808_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_808_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_87_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_87_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_87_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_87_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_809_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_809_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_809_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_809_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_809_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_809_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_809_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_809_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_88_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_88_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_88_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_88_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_810_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_810_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_810_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_810_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_810_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_810_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_810_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_810_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_89_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_89_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_89_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_89_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_811_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_811_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_811_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_811_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_811_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_811_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_811_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_811_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_90_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_90_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_90_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_90_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_812_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_812_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_812_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_812_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_812_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_812_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_812_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_812_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_91_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_91_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_91_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_91_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_813_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_813_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_813_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_813_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_813_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_813_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_813_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_813_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_92_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_92_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_92_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_92_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_814_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_814_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_814_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_814_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_814_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_814_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_814_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_814_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_93_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_93_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_93_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_93_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_815_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_815_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_815_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_815_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_815_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_815_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_815_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_815_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_94_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_94_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_94_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_94_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_816_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_816_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_816_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_816_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_816_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_816_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_816_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_816_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_95_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_95_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_95_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_95_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_817_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_817_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_817_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_817_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_817_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_817_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_817_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_817_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_96_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_96_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_96_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_96_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_818_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_818_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_818_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_818_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_818_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_818_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_818_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_818_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_97_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_97_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_97_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_97_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_819_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_819_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_819_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_819_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_819_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_819_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_819_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_819_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_98_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_98_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_98_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_98_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_820_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_820_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_820_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_820_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_820_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_820_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_820_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_820_io_out_2; // @[Multiplier.scala 130:25]
  wire  c32_56_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_56_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_56_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_56_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_56_io_out_1; // @[Multiplier.scala 125:25]
  wire  c53_821_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_821_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_821_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_821_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_821_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_821_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_821_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_821_io_out_2; // @[Multiplier.scala 130:25]
  wire  c32_57_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_57_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_57_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_57_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_57_io_out_1; // @[Multiplier.scala 125:25]
  wire  c53_822_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_822_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_822_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_822_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_822_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_822_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_822_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_822_io_out_2; // @[Multiplier.scala 130:25]
  wire  c32_58_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_58_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_58_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_58_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_58_io_out_1; // @[Multiplier.scala 125:25]
  wire  c53_823_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_823_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_823_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_823_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_823_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_823_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_823_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_823_io_out_2; // @[Multiplier.scala 130:25]
  wire  c32_59_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_59_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_59_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_59_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_59_io_out_1; // @[Multiplier.scala 125:25]
  wire  c53_824_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_824_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_824_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_824_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_824_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_824_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_824_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_824_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_825_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_825_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_825_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_825_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_825_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_825_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_825_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_825_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_826_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_826_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_826_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_826_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_826_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_826_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_826_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_826_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_827_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_827_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_827_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_827_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_827_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_827_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_827_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_827_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_828_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_828_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_828_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_828_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_828_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_828_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_828_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_828_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_829_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_829_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_829_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_829_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_829_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_829_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_829_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_829_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_830_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_830_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_830_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_830_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_830_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_830_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_830_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_830_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_831_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_831_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_831_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_831_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_831_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_831_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_831_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_831_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_832_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_832_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_832_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_832_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_832_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_832_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_832_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_832_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_833_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_833_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_833_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_833_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_833_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_833_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_833_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_833_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_834_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_834_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_834_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_834_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_834_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_834_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_834_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_834_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_835_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_835_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_835_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_835_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_835_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_835_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_835_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_835_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_836_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_836_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_836_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_836_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_836_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_836_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_836_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_836_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_837_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_837_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_837_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_837_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_837_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_837_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_837_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_837_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_838_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_838_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_838_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_838_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_838_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_838_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_838_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_838_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_839_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_839_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_839_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_839_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_839_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_839_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_839_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_839_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_840_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_840_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_840_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_840_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_840_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_840_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_840_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_840_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_841_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_841_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_841_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_841_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_841_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_841_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_841_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_841_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_842_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_842_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_842_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_842_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_842_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_842_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_842_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_842_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_843_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_843_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_843_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_843_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_843_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_843_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_843_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_843_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_844_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_844_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_844_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_844_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_844_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_844_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_844_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_844_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_845_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_845_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_845_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_845_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_845_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_845_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_845_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_845_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_846_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_846_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_846_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_846_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_846_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_846_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_846_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_846_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_847_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_847_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_847_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_847_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_847_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_847_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_847_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_847_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_848_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_848_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_848_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_848_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_848_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_848_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_848_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_848_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_849_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_849_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_849_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_849_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_849_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_849_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_849_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_849_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_850_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_850_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_850_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_850_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_850_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_850_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_850_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_850_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_851_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_851_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_851_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_851_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_851_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_851_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_851_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_851_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_852_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_852_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_852_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_852_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_852_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_852_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_852_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_852_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_853_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_853_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_853_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_853_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_853_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_853_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_853_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_853_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_854_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_854_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_854_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_854_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_854_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_854_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_854_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_854_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_855_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_855_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_855_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_855_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_855_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_855_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_855_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_855_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_856_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_856_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_856_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_856_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_856_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_856_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_856_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_856_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_857_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_857_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_857_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_857_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_857_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_857_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_857_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_857_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_858_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_858_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_858_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_858_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_858_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_858_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_858_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_858_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_859_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_859_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_859_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_859_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_859_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_859_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_859_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_859_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_860_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_860_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_860_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_860_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_860_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_860_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_860_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_860_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_861_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_861_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_861_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_861_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_861_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_861_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_861_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_861_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_862_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_862_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_862_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_862_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_862_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_862_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_862_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_862_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_863_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_863_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_863_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_863_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_863_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_863_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_863_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_863_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_864_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_864_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_864_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_864_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_864_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_864_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_864_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_864_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_865_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_865_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_865_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_865_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_865_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_865_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_865_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_865_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_866_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_866_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_866_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_866_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_866_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_866_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_866_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_866_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_867_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_867_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_867_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_867_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_867_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_867_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_867_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_867_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_868_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_868_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_868_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_868_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_868_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_868_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_868_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_868_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_869_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_869_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_869_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_869_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_869_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_869_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_869_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_869_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_870_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_870_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_870_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_870_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_870_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_870_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_870_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_870_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_871_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_871_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_871_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_871_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_871_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_871_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_871_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_871_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_872_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_872_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_872_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_872_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_872_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_872_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_872_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_872_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_873_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_873_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_873_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_873_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_873_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_873_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_873_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_873_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_874_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_874_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_874_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_874_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_874_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_874_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_874_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_874_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_875_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_875_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_875_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_875_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_875_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_875_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_875_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_875_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_876_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_876_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_876_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_876_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_876_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_876_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_876_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_876_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_877_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_877_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_877_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_877_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_877_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_877_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_877_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_877_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_878_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_878_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_878_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_878_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_878_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_878_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_878_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_878_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_879_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_879_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_879_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_879_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_879_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_879_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_879_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_879_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_880_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_880_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_880_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_880_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_880_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_880_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_880_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_880_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_881_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_881_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_881_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_881_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_881_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_881_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_881_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_881_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_882_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_882_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_882_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_882_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_882_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_882_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_882_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_882_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_883_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_883_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_883_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_883_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_883_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_883_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_883_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_883_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_884_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_884_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_884_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_884_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_884_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_884_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_884_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_884_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_885_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_885_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_885_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_885_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_885_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_885_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_885_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_885_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_886_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_886_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_886_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_886_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_886_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_886_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_886_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_886_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_887_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_887_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_887_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_887_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_887_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_887_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_887_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_887_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_888_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_888_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_888_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_888_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_888_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_888_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_888_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_888_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_889_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_889_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_889_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_889_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_889_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_889_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_889_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_889_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_890_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_890_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_890_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_890_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_890_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_890_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_890_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_890_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_891_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_891_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_891_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_891_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_891_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_891_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_891_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_891_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_892_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_892_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_892_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_892_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_892_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_892_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_892_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_892_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_99_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_99_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_99_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_99_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_893_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_893_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_893_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_893_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_893_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_893_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_893_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_893_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_100_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_100_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_100_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_100_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_894_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_894_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_894_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_894_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_894_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_894_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_894_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_894_io_out_2; // @[Multiplier.scala 130:25]
  wire  c32_60_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_60_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_60_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_60_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_60_io_out_1; // @[Multiplier.scala 125:25]
  wire  c53_895_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_895_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_895_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_895_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_895_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_895_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_895_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_895_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_101_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_101_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_101_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_101_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_896_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_896_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_896_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_896_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_896_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_896_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_896_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_896_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_102_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_102_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_102_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_102_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_897_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_897_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_897_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_897_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_897_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_897_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_897_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_897_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_103_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_103_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_103_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_103_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_898_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_898_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_898_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_898_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_898_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_898_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_898_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_898_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_104_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_104_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_104_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_104_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_899_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_899_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_899_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_899_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_899_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_899_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_899_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_899_io_out_2; // @[Multiplier.scala 130:25]
  wire  c32_61_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_61_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_61_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_61_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_61_io_out_1; // @[Multiplier.scala 125:25]
  wire  c53_900_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_900_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_900_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_900_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_900_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_900_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_900_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_900_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_105_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_105_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_105_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_105_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_901_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_901_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_901_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_901_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_901_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_901_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_901_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_901_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_106_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_106_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_106_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_106_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_902_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_902_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_902_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_902_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_902_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_902_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_902_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_902_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_107_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_107_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_107_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_107_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_903_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_903_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_903_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_903_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_903_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_903_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_903_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_903_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_108_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_108_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_108_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_108_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_904_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_904_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_904_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_904_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_904_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_904_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_904_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_904_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_109_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_109_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_109_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_109_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_905_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_905_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_905_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_905_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_905_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_905_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_905_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_905_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_110_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_110_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_110_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_110_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_906_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_906_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_906_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_906_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_906_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_906_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_906_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_906_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_111_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_111_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_111_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_111_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_907_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_907_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_907_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_907_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_907_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_907_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_907_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_907_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_112_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_112_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_112_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_112_io_out_1; // @[Multiplier.scala 120:25]
  wire  c53_908_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_908_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_908_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_908_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_908_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_908_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_908_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_908_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_909_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_909_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_909_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_909_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_909_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_909_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_909_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_909_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_910_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_910_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_910_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_910_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_910_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_910_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_910_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_910_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_911_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_911_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_911_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_911_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_911_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_911_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_911_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_911_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_912_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_912_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_912_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_912_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_912_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_912_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_912_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_912_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_913_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_913_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_913_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_913_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_913_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_913_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_913_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_913_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_914_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_914_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_914_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_914_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_914_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_914_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_914_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_914_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_915_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_915_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_915_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_915_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_915_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_915_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_915_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_915_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_916_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_916_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_916_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_916_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_916_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_916_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_916_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_916_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_917_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_917_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_917_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_917_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_917_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_917_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_917_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_917_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_918_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_918_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_918_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_918_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_918_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_918_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_918_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_918_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_919_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_919_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_919_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_919_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_919_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_919_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_919_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_919_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_920_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_920_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_920_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_920_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_920_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_920_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_920_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_920_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_921_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_921_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_921_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_921_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_921_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_921_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_921_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_921_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_922_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_922_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_922_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_922_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_922_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_922_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_922_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_922_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_923_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_923_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_923_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_923_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_923_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_923_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_923_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_923_io_out_2; // @[Multiplier.scala 130:25]
  wire  c22_113_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_113_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_113_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_113_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_114_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_114_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_114_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_114_io_out_1; // @[Multiplier.scala 120:25]
  wire  c32_62_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_62_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_62_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_62_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_62_io_out_1; // @[Multiplier.scala 125:25]
  wire  c22_115_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_115_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_115_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_115_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_116_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_116_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_116_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_116_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_117_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_117_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_117_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_117_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_118_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_118_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_118_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_118_io_out_1; // @[Multiplier.scala 120:25]
  wire  c32_63_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_63_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_63_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_63_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_63_io_out_1; // @[Multiplier.scala 125:25]
  wire  c22_119_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_119_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_119_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_119_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_120_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_120_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_120_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_120_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_121_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_121_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_121_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_121_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_122_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_122_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_122_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_122_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_123_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_123_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_123_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_123_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_124_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_124_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_124_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_124_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_125_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_125_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_125_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_125_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_126_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_126_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_126_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_126_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_127_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_127_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_127_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_127_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_128_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_128_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_128_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_128_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_129_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_129_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_129_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_129_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_130_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_130_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_130_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_130_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_131_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_131_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_131_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_131_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_132_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_132_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_132_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_132_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_133_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_133_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_133_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_133_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_134_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_134_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_134_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_134_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_135_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_135_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_135_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_135_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_136_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_136_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_136_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_136_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_137_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_137_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_137_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_137_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_138_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_138_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_138_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_138_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_139_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_139_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_139_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_139_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_140_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_140_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_140_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_140_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_141_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_141_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_141_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_141_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_142_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_142_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_142_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_142_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_143_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_143_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_143_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_143_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_144_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_144_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_144_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_144_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_145_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_145_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_145_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_145_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_146_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_146_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_146_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_146_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_147_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_147_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_147_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_147_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_148_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_148_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_148_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_148_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_149_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_149_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_149_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_149_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_150_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_150_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_150_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_150_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_151_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_151_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_151_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_151_io_out_1; // @[Multiplier.scala 120:25]
  wire  c32_64_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_64_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_64_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_64_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_64_io_out_1; // @[Multiplier.scala 125:25]
  wire  c32_65_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_65_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_65_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_65_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_65_io_out_1; // @[Multiplier.scala 125:25]
  wire  c32_66_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_66_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_66_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_66_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_66_io_out_1; // @[Multiplier.scala 125:25]
  wire  c32_67_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_67_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_67_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_67_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_67_io_out_1; // @[Multiplier.scala 125:25]
  wire  c32_68_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_68_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_68_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_68_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_68_io_out_1; // @[Multiplier.scala 125:25]
  wire  c53_924_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_924_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_924_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_924_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_924_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_924_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_924_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_924_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_925_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_925_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_925_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_925_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_925_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_925_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_925_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_925_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_926_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_926_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_926_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_926_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_926_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_926_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_926_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_926_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_927_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_927_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_927_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_927_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_927_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_927_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_927_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_927_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_928_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_928_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_928_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_928_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_928_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_928_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_928_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_928_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_929_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_929_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_929_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_929_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_929_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_929_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_929_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_929_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_930_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_930_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_930_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_930_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_930_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_930_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_930_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_930_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_931_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_931_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_931_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_931_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_931_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_931_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_931_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_931_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_932_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_932_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_932_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_932_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_932_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_932_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_932_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_932_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_933_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_933_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_933_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_933_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_933_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_933_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_933_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_933_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_934_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_934_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_934_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_934_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_934_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_934_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_934_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_934_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_935_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_935_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_935_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_935_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_935_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_935_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_935_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_935_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_936_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_936_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_936_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_936_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_936_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_936_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_936_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_936_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_937_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_937_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_937_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_937_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_937_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_937_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_937_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_937_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_938_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_938_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_938_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_938_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_938_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_938_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_938_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_938_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_939_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_939_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_939_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_939_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_939_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_939_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_939_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_939_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_940_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_940_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_940_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_940_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_940_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_940_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_940_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_940_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_941_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_941_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_941_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_941_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_941_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_941_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_941_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_941_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_942_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_942_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_942_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_942_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_942_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_942_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_942_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_942_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_943_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_943_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_943_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_943_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_943_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_943_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_943_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_943_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_944_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_944_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_944_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_944_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_944_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_944_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_944_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_944_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_945_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_945_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_945_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_945_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_945_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_945_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_945_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_945_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_946_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_946_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_946_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_946_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_946_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_946_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_946_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_946_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_947_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_947_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_947_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_947_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_947_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_947_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_947_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_947_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_948_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_948_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_948_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_948_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_948_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_948_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_948_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_948_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_949_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_949_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_949_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_949_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_949_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_949_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_949_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_949_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_950_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_950_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_950_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_950_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_950_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_950_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_950_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_950_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_951_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_951_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_951_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_951_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_951_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_951_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_951_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_951_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_952_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_952_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_952_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_952_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_952_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_952_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_952_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_952_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_953_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_953_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_953_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_953_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_953_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_953_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_953_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_953_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_954_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_954_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_954_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_954_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_954_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_954_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_954_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_954_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_955_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_955_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_955_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_955_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_955_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_955_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_955_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_955_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_956_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_956_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_956_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_956_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_956_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_956_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_956_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_956_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_957_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_957_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_957_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_957_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_957_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_957_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_957_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_957_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_958_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_958_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_958_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_958_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_958_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_958_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_958_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_958_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_959_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_959_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_959_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_959_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_959_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_959_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_959_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_959_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_960_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_960_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_960_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_960_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_960_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_960_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_960_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_960_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_961_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_961_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_961_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_961_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_961_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_961_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_961_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_961_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_962_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_962_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_962_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_962_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_962_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_962_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_962_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_962_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_963_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_963_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_963_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_963_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_963_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_963_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_963_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_963_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_964_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_964_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_964_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_964_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_964_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_964_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_964_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_964_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_965_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_965_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_965_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_965_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_965_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_965_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_965_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_965_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_966_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_966_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_966_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_966_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_966_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_966_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_966_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_966_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_967_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_967_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_967_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_967_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_967_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_967_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_967_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_967_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_968_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_968_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_968_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_968_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_968_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_968_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_968_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_968_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_969_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_969_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_969_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_969_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_969_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_969_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_969_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_969_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_970_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_970_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_970_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_970_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_970_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_970_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_970_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_970_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_971_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_971_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_971_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_971_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_971_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_971_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_971_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_971_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_972_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_972_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_972_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_972_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_972_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_972_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_972_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_972_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_973_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_973_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_973_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_973_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_973_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_973_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_973_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_973_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_974_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_974_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_974_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_974_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_974_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_974_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_974_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_974_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_975_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_975_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_975_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_975_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_975_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_975_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_975_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_975_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_976_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_976_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_976_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_976_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_976_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_976_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_976_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_976_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_977_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_977_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_977_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_977_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_977_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_977_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_977_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_977_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_978_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_978_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_978_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_978_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_978_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_978_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_978_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_978_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_979_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_979_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_979_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_979_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_979_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_979_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_979_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_979_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_980_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_980_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_980_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_980_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_980_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_980_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_980_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_980_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_981_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_981_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_981_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_981_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_981_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_981_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_981_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_981_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_982_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_982_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_982_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_982_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_982_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_982_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_982_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_982_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_983_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_983_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_983_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_983_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_983_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_983_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_983_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_983_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_984_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_984_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_984_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_984_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_984_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_984_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_984_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_984_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_985_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_985_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_985_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_985_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_985_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_985_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_985_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_985_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_986_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_986_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_986_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_986_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_986_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_986_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_986_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_986_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_987_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_987_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_987_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_987_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_987_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_987_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_987_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_987_io_out_2; // @[Multiplier.scala 130:25]
  wire  c53_988_io_in_0; // @[Multiplier.scala 130:25]
  wire  c53_988_io_in_1; // @[Multiplier.scala 130:25]
  wire  c53_988_io_in_2; // @[Multiplier.scala 130:25]
  wire  c53_988_io_in_3; // @[Multiplier.scala 130:25]
  wire  c53_988_io_in_4; // @[Multiplier.scala 130:25]
  wire  c53_988_io_out_0; // @[Multiplier.scala 130:25]
  wire  c53_988_io_out_1; // @[Multiplier.scala 130:25]
  wire  c53_988_io_out_2; // @[Multiplier.scala 130:25]
  wire  c32_69_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_69_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_69_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_69_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_69_io_out_1; // @[Multiplier.scala 125:25]
  wire  c22_152_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_152_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_152_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_152_io_out_1; // @[Multiplier.scala 120:25]
  wire  c32_70_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_70_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_70_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_70_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_70_io_out_1; // @[Multiplier.scala 125:25]
  wire  c22_153_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_153_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_153_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_153_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_154_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_154_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_154_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_154_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_155_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_155_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_155_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_155_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_156_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_156_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_156_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_156_io_out_1; // @[Multiplier.scala 120:25]
  wire  c32_71_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_71_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_71_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_71_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_71_io_out_1; // @[Multiplier.scala 125:25]
  wire  c22_157_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_157_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_157_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_157_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_158_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_158_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_158_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_158_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_159_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_159_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_159_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_159_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_160_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_160_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_160_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_160_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_161_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_161_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_161_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_161_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_162_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_162_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_162_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_162_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_163_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_163_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_163_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_163_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_164_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_164_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_164_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_164_io_out_1; // @[Multiplier.scala 120:25]
  wire  c32_72_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_72_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_72_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_72_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_72_io_out_1; // @[Multiplier.scala 125:25]
  wire  c22_165_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_165_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_165_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_165_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_166_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_166_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_166_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_166_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_167_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_167_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_167_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_167_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_168_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_168_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_168_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_168_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_169_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_169_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_169_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_169_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_170_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_170_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_170_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_170_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_171_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_171_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_171_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_171_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_172_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_172_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_172_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_172_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_173_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_173_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_173_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_173_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_174_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_174_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_174_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_174_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_175_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_175_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_175_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_175_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_176_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_176_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_176_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_176_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_177_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_177_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_177_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_177_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_178_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_178_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_178_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_178_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_179_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_179_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_179_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_179_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_180_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_180_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_180_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_180_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_181_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_181_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_181_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_181_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_182_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_182_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_182_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_182_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_183_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_183_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_183_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_183_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_184_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_184_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_184_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_184_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_185_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_185_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_185_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_185_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_186_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_186_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_186_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_186_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_187_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_187_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_187_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_187_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_188_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_188_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_188_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_188_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_189_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_189_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_189_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_189_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_190_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_190_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_190_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_190_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_191_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_191_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_191_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_191_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_192_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_192_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_192_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_192_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_193_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_193_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_193_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_193_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_194_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_194_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_194_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_194_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_195_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_195_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_195_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_195_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_196_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_196_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_196_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_196_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_197_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_197_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_197_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_197_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_198_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_198_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_198_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_198_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_199_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_199_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_199_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_199_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_200_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_200_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_200_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_200_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_201_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_201_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_201_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_201_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_202_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_202_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_202_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_202_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_203_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_203_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_203_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_203_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_204_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_204_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_204_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_204_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_205_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_205_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_205_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_205_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_206_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_206_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_206_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_206_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_207_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_207_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_207_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_207_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_208_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_208_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_208_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_208_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_209_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_209_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_209_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_209_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_210_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_210_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_210_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_210_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_211_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_211_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_211_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_211_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_212_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_212_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_212_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_212_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_213_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_213_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_213_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_213_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_214_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_214_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_214_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_214_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_215_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_215_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_215_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_215_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_216_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_216_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_216_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_216_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_217_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_217_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_217_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_217_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_218_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_218_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_218_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_218_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_219_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_219_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_219_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_219_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_220_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_220_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_220_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_220_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_221_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_221_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_221_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_221_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_222_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_222_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_222_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_222_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_223_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_223_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_223_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_223_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_224_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_224_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_224_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_224_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_225_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_225_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_225_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_225_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_226_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_226_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_226_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_226_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_227_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_227_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_227_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_227_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_228_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_228_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_228_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_228_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_229_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_229_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_229_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_229_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_230_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_230_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_230_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_230_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_231_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_231_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_231_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_231_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_232_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_232_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_232_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_232_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_233_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_233_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_233_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_233_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_234_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_234_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_234_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_234_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_235_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_235_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_235_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_235_io_out_1; // @[Multiplier.scala 120:25]
  wire  c32_73_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_73_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_73_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_73_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_73_io_out_1; // @[Multiplier.scala 125:25]
  wire  c32_74_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_74_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_74_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_74_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_74_io_out_1; // @[Multiplier.scala 125:25]
  wire  c32_75_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_75_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_75_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_75_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_75_io_out_1; // @[Multiplier.scala 125:25]
  wire  c32_76_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_76_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_76_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_76_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_76_io_out_1; // @[Multiplier.scala 125:25]
  wire  c32_77_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_77_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_77_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_77_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_77_io_out_1; // @[Multiplier.scala 125:25]
  wire  c32_78_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_78_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_78_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_78_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_78_io_out_1; // @[Multiplier.scala 125:25]
  wire  c32_79_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_79_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_79_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_79_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_79_io_out_1; // @[Multiplier.scala 125:25]
  wire  c22_236_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_236_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_236_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_236_io_out_1; // @[Multiplier.scala 120:25]
  wire  c32_80_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_80_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_80_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_80_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_80_io_out_1; // @[Multiplier.scala 125:25]
  wire  c22_237_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_237_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_237_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_237_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_238_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_238_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_238_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_238_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_239_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_239_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_239_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_239_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_240_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_240_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_240_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_240_io_out_1; // @[Multiplier.scala 120:25]
  wire  c32_81_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_81_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_81_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_81_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_81_io_out_1; // @[Multiplier.scala 125:25]
  wire  c22_241_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_241_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_241_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_241_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_242_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_242_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_242_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_242_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_243_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_243_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_243_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_243_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_244_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_244_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_244_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_244_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_245_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_245_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_245_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_245_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_246_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_246_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_246_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_246_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_247_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_247_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_247_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_247_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_248_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_248_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_248_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_248_io_out_1; // @[Multiplier.scala 120:25]
  wire  c32_82_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_82_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_82_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_82_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_82_io_out_1; // @[Multiplier.scala 125:25]
  wire  c22_249_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_249_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_249_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_249_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_250_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_250_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_250_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_250_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_251_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_251_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_251_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_251_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_252_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_252_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_252_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_252_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_253_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_253_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_253_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_253_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_254_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_254_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_254_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_254_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_255_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_255_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_255_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_255_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_256_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_256_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_256_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_256_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_257_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_257_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_257_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_257_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_258_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_258_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_258_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_258_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_259_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_259_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_259_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_259_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_260_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_260_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_260_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_260_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_261_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_261_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_261_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_261_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_262_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_262_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_262_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_262_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_263_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_263_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_263_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_263_io_out_1; // @[Multiplier.scala 120:25]
  wire  c32_83_io_in_0; // @[Multiplier.scala 125:25]
  wire  c32_83_io_in_1; // @[Multiplier.scala 125:25]
  wire  c32_83_io_in_2; // @[Multiplier.scala 125:25]
  wire  c32_83_io_out_0; // @[Multiplier.scala 125:25]
  wire  c32_83_io_out_1; // @[Multiplier.scala 125:25]
  wire  c22_264_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_264_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_264_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_264_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_265_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_265_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_265_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_265_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_266_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_266_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_266_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_266_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_267_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_267_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_267_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_267_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_268_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_268_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_268_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_268_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_269_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_269_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_269_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_269_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_270_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_270_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_270_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_270_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_271_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_271_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_271_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_271_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_272_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_272_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_272_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_272_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_273_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_273_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_273_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_273_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_274_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_274_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_274_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_274_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_275_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_275_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_275_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_275_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_276_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_276_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_276_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_276_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_277_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_277_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_277_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_277_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_278_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_278_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_278_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_278_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_279_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_279_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_279_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_279_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_280_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_280_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_280_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_280_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_281_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_281_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_281_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_281_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_282_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_282_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_282_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_282_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_283_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_283_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_283_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_283_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_284_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_284_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_284_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_284_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_285_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_285_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_285_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_285_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_286_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_286_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_286_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_286_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_287_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_287_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_287_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_287_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_288_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_288_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_288_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_288_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_289_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_289_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_289_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_289_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_290_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_290_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_290_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_290_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_291_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_291_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_291_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_291_io_out_1; // @[Multiplier.scala 120:25]
  wire  c22_292_io_in_0; // @[Multiplier.scala 120:25]
  wire  c22_292_io_in_1; // @[Multiplier.scala 120:25]
  wire  c22_292_io_out_0; // @[Multiplier.scala 120:25]
  wire  c22_292_io_out_1; // @[Multiplier.scala 120:25]
  wire  b_sext_signBit = io_b[64]; // @[BitUtils.scala 80:20]
  wire [65:0] b_sext = {b_sext_signBit,io_b}; // @[Cat.scala 31:58]
  wire [66:0] _bx2_T = {b_sext, 1'h0}; // @[Multiplier.scala 73:17]
  wire [65:0] neg_b = ~b_sext; // @[Multiplier.scala 74:13]
  wire [66:0] _neg_bx2_T = {neg_b, 1'h0}; // @[Multiplier.scala 75:20]
  wire [2:0] x = {io_a[1:0],1'h0}; // @[Cat.scala 31:58]
  wire [65:0] _pp_temp_T_1 = 3'h1 == x ? b_sext : 66'h0; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_3 = 3'h2 == x ? b_sext : _pp_temp_T_1; // @[Mux.scala 81:58]
  wire [65:0] bx2 = _bx2_T[65:0]; // @[Multiplier.scala 71:41 73:7]
  wire [65:0] _pp_temp_T_5 = 3'h3 == x ? bx2 : _pp_temp_T_3; // @[Mux.scala 81:58]
  wire [65:0] neg_bx2 = _neg_bx2_T[65:0]; // @[Multiplier.scala 71:41 75:11]
  wire [65:0] _pp_temp_T_7 = 3'h4 == x ? neg_bx2 : _pp_temp_T_5; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_9 = 3'h5 == x ? neg_b : _pp_temp_T_7; // @[Mux.scala 81:58]
  wire [65:0] pp_temp = 3'h6 == x ? neg_b : _pp_temp_T_9; // @[Mux.scala 81:58]
  wire  s = pp_temp[65]; // @[Multiplier.scala 90:20]
  wire  _T = ~s; // @[Multiplier.scala 99:14]
  wire [68:0] pp = {_T,s,s,pp_temp}; // @[Cat.scala 31:58]
  wire [2:0] x_1 = io_a[3:1]; // @[Multiplier.scala 81:90]
  wire [65:0] _pp_temp_T_12 = 3'h1 == x_1 ? b_sext : 66'h0; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_14 = 3'h2 == x_1 ? b_sext : _pp_temp_T_12; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_16 = 3'h3 == x_1 ? bx2 : _pp_temp_T_14; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_18 = 3'h4 == x_1 ? neg_bx2 : _pp_temp_T_16; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_20 = 3'h5 == x_1 ? neg_b : _pp_temp_T_18; // @[Mux.scala 81:58]
  wire [65:0] pp_temp_1 = 3'h6 == x_1 ? neg_b : _pp_temp_T_20; // @[Mux.scala 81:58]
  wire  s_1 = pp_temp_1[65]; // @[Multiplier.scala 90:20]
  wire [1:0] _t_T_6 = 3'h4 == x ? 2'h2 : 2'h0; // @[Mux.scala 81:58]
  wire [1:0] _t_T_8 = 3'h5 == x ? 2'h1 : _t_T_6; // @[Mux.scala 81:58]
  wire [1:0] t_1 = 3'h6 == x ? 2'h1 : _t_T_8; // @[Mux.scala 81:58]
  wire  _T_70 = ~s_1; // @[Multiplier.scala 103:24]
  wire [69:0] pp_1 = {1'h1,_T_70,pp_temp_1,t_1}; // @[Cat.scala 31:58]
  wire [2:0] x_2 = io_a[5:3]; // @[Multiplier.scala 81:90]
  wire [65:0] _pp_temp_T_23 = 3'h1 == x_2 ? b_sext : 66'h0; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_25 = 3'h2 == x_2 ? b_sext : _pp_temp_T_23; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_27 = 3'h3 == x_2 ? bx2 : _pp_temp_T_25; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_29 = 3'h4 == x_2 ? neg_bx2 : _pp_temp_T_27; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_31 = 3'h5 == x_2 ? neg_b : _pp_temp_T_29; // @[Mux.scala 81:58]
  wire [65:0] pp_temp_2 = 3'h6 == x_2 ? neg_b : _pp_temp_T_31; // @[Mux.scala 81:58]
  wire  s_2 = pp_temp_2[65]; // @[Multiplier.scala 90:20]
  wire [1:0] _t_T_11 = 3'h4 == x_1 ? 2'h2 : 2'h0; // @[Mux.scala 81:58]
  wire [1:0] _t_T_13 = 3'h5 == x_1 ? 2'h1 : _t_T_11; // @[Mux.scala 81:58]
  wire [1:0] t_2 = 3'h6 == x_1 ? 2'h1 : _t_T_13; // @[Mux.scala 81:58]
  wire  _T_141 = ~s_2; // @[Multiplier.scala 103:24]
  wire [69:0] pp_2 = {1'h1,_T_141,pp_temp_2,t_2}; // @[Cat.scala 31:58]
  wire [2:0] x_3 = io_a[7:5]; // @[Multiplier.scala 81:90]
  wire [65:0] _pp_temp_T_34 = 3'h1 == x_3 ? b_sext : 66'h0; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_36 = 3'h2 == x_3 ? b_sext : _pp_temp_T_34; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_38 = 3'h3 == x_3 ? bx2 : _pp_temp_T_36; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_40 = 3'h4 == x_3 ? neg_bx2 : _pp_temp_T_38; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_42 = 3'h5 == x_3 ? neg_b : _pp_temp_T_40; // @[Mux.scala 81:58]
  wire [65:0] pp_temp_3 = 3'h6 == x_3 ? neg_b : _pp_temp_T_42; // @[Mux.scala 81:58]
  wire  s_3 = pp_temp_3[65]; // @[Multiplier.scala 90:20]
  wire [1:0] _t_T_16 = 3'h4 == x_2 ? 2'h2 : 2'h0; // @[Mux.scala 81:58]
  wire [1:0] _t_T_18 = 3'h5 == x_2 ? 2'h1 : _t_T_16; // @[Mux.scala 81:58]
  wire [1:0] t_3 = 3'h6 == x_2 ? 2'h1 : _t_T_18; // @[Mux.scala 81:58]
  wire  _T_212 = ~s_3; // @[Multiplier.scala 103:24]
  wire [69:0] pp_3 = {1'h1,_T_212,pp_temp_3,t_3}; // @[Cat.scala 31:58]
  wire [2:0] x_4 = io_a[9:7]; // @[Multiplier.scala 81:90]
  wire [65:0] _pp_temp_T_45 = 3'h1 == x_4 ? b_sext : 66'h0; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_47 = 3'h2 == x_4 ? b_sext : _pp_temp_T_45; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_49 = 3'h3 == x_4 ? bx2 : _pp_temp_T_47; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_51 = 3'h4 == x_4 ? neg_bx2 : _pp_temp_T_49; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_53 = 3'h5 == x_4 ? neg_b : _pp_temp_T_51; // @[Mux.scala 81:58]
  wire [65:0] pp_temp_4 = 3'h6 == x_4 ? neg_b : _pp_temp_T_53; // @[Mux.scala 81:58]
  wire  s_4 = pp_temp_4[65]; // @[Multiplier.scala 90:20]
  wire [1:0] _t_T_21 = 3'h4 == x_3 ? 2'h2 : 2'h0; // @[Mux.scala 81:58]
  wire [1:0] _t_T_23 = 3'h5 == x_3 ? 2'h1 : _t_T_21; // @[Mux.scala 81:58]
  wire [1:0] t_4 = 3'h6 == x_3 ? 2'h1 : _t_T_23; // @[Mux.scala 81:58]
  wire  _T_283 = ~s_4; // @[Multiplier.scala 103:24]
  wire [69:0] pp_4 = {1'h1,_T_283,pp_temp_4,t_4}; // @[Cat.scala 31:58]
  wire [2:0] x_5 = io_a[11:9]; // @[Multiplier.scala 81:90]
  wire [65:0] _pp_temp_T_56 = 3'h1 == x_5 ? b_sext : 66'h0; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_58 = 3'h2 == x_5 ? b_sext : _pp_temp_T_56; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_60 = 3'h3 == x_5 ? bx2 : _pp_temp_T_58; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_62 = 3'h4 == x_5 ? neg_bx2 : _pp_temp_T_60; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_64 = 3'h5 == x_5 ? neg_b : _pp_temp_T_62; // @[Mux.scala 81:58]
  wire [65:0] pp_temp_5 = 3'h6 == x_5 ? neg_b : _pp_temp_T_64; // @[Mux.scala 81:58]
  wire  s_5 = pp_temp_5[65]; // @[Multiplier.scala 90:20]
  wire [1:0] _t_T_26 = 3'h4 == x_4 ? 2'h2 : 2'h0; // @[Mux.scala 81:58]
  wire [1:0] _t_T_28 = 3'h5 == x_4 ? 2'h1 : _t_T_26; // @[Mux.scala 81:58]
  wire [1:0] t_5 = 3'h6 == x_4 ? 2'h1 : _t_T_28; // @[Mux.scala 81:58]
  wire  _T_354 = ~s_5; // @[Multiplier.scala 103:24]
  wire [69:0] pp_5 = {1'h1,_T_354,pp_temp_5,t_5}; // @[Cat.scala 31:58]
  wire [2:0] x_6 = io_a[13:11]; // @[Multiplier.scala 81:90]
  wire [65:0] _pp_temp_T_67 = 3'h1 == x_6 ? b_sext : 66'h0; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_69 = 3'h2 == x_6 ? b_sext : _pp_temp_T_67; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_71 = 3'h3 == x_6 ? bx2 : _pp_temp_T_69; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_73 = 3'h4 == x_6 ? neg_bx2 : _pp_temp_T_71; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_75 = 3'h5 == x_6 ? neg_b : _pp_temp_T_73; // @[Mux.scala 81:58]
  wire [65:0] pp_temp_6 = 3'h6 == x_6 ? neg_b : _pp_temp_T_75; // @[Mux.scala 81:58]
  wire  s_6 = pp_temp_6[65]; // @[Multiplier.scala 90:20]
  wire [1:0] _t_T_31 = 3'h4 == x_5 ? 2'h2 : 2'h0; // @[Mux.scala 81:58]
  wire [1:0] _t_T_33 = 3'h5 == x_5 ? 2'h1 : _t_T_31; // @[Mux.scala 81:58]
  wire [1:0] t_6 = 3'h6 == x_5 ? 2'h1 : _t_T_33; // @[Mux.scala 81:58]
  wire  _T_425 = ~s_6; // @[Multiplier.scala 103:24]
  wire [69:0] pp_6 = {1'h1,_T_425,pp_temp_6,t_6}; // @[Cat.scala 31:58]
  wire [2:0] x_7 = io_a[15:13]; // @[Multiplier.scala 81:90]
  wire [65:0] _pp_temp_T_78 = 3'h1 == x_7 ? b_sext : 66'h0; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_80 = 3'h2 == x_7 ? b_sext : _pp_temp_T_78; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_82 = 3'h3 == x_7 ? bx2 : _pp_temp_T_80; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_84 = 3'h4 == x_7 ? neg_bx2 : _pp_temp_T_82; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_86 = 3'h5 == x_7 ? neg_b : _pp_temp_T_84; // @[Mux.scala 81:58]
  wire [65:0] pp_temp_7 = 3'h6 == x_7 ? neg_b : _pp_temp_T_86; // @[Mux.scala 81:58]
  wire  s_7 = pp_temp_7[65]; // @[Multiplier.scala 90:20]
  wire [1:0] _t_T_36 = 3'h4 == x_6 ? 2'h2 : 2'h0; // @[Mux.scala 81:58]
  wire [1:0] _t_T_38 = 3'h5 == x_6 ? 2'h1 : _t_T_36; // @[Mux.scala 81:58]
  wire [1:0] t_7 = 3'h6 == x_6 ? 2'h1 : _t_T_38; // @[Mux.scala 81:58]
  wire  _T_496 = ~s_7; // @[Multiplier.scala 103:24]
  wire [69:0] pp_7 = {1'h1,_T_496,pp_temp_7,t_7}; // @[Cat.scala 31:58]
  wire [2:0] x_8 = io_a[17:15]; // @[Multiplier.scala 81:90]
  wire [65:0] _pp_temp_T_89 = 3'h1 == x_8 ? b_sext : 66'h0; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_91 = 3'h2 == x_8 ? b_sext : _pp_temp_T_89; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_93 = 3'h3 == x_8 ? bx2 : _pp_temp_T_91; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_95 = 3'h4 == x_8 ? neg_bx2 : _pp_temp_T_93; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_97 = 3'h5 == x_8 ? neg_b : _pp_temp_T_95; // @[Mux.scala 81:58]
  wire [65:0] pp_temp_8 = 3'h6 == x_8 ? neg_b : _pp_temp_T_97; // @[Mux.scala 81:58]
  wire  s_8 = pp_temp_8[65]; // @[Multiplier.scala 90:20]
  wire [1:0] _t_T_41 = 3'h4 == x_7 ? 2'h2 : 2'h0; // @[Mux.scala 81:58]
  wire [1:0] _t_T_43 = 3'h5 == x_7 ? 2'h1 : _t_T_41; // @[Mux.scala 81:58]
  wire [1:0] t_8 = 3'h6 == x_7 ? 2'h1 : _t_T_43; // @[Mux.scala 81:58]
  wire  _T_567 = ~s_8; // @[Multiplier.scala 103:24]
  wire [69:0] pp_8 = {1'h1,_T_567,pp_temp_8,t_8}; // @[Cat.scala 31:58]
  wire [2:0] x_9 = io_a[19:17]; // @[Multiplier.scala 81:90]
  wire [65:0] _pp_temp_T_100 = 3'h1 == x_9 ? b_sext : 66'h0; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_102 = 3'h2 == x_9 ? b_sext : _pp_temp_T_100; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_104 = 3'h3 == x_9 ? bx2 : _pp_temp_T_102; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_106 = 3'h4 == x_9 ? neg_bx2 : _pp_temp_T_104; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_108 = 3'h5 == x_9 ? neg_b : _pp_temp_T_106; // @[Mux.scala 81:58]
  wire [65:0] pp_temp_9 = 3'h6 == x_9 ? neg_b : _pp_temp_T_108; // @[Mux.scala 81:58]
  wire  s_9 = pp_temp_9[65]; // @[Multiplier.scala 90:20]
  wire [1:0] _t_T_46 = 3'h4 == x_8 ? 2'h2 : 2'h0; // @[Mux.scala 81:58]
  wire [1:0] _t_T_48 = 3'h5 == x_8 ? 2'h1 : _t_T_46; // @[Mux.scala 81:58]
  wire [1:0] t_9 = 3'h6 == x_8 ? 2'h1 : _t_T_48; // @[Mux.scala 81:58]
  wire  _T_638 = ~s_9; // @[Multiplier.scala 103:24]
  wire [69:0] pp_9 = {1'h1,_T_638,pp_temp_9,t_9}; // @[Cat.scala 31:58]
  wire [2:0] x_10 = io_a[21:19]; // @[Multiplier.scala 81:90]
  wire [65:0] _pp_temp_T_111 = 3'h1 == x_10 ? b_sext : 66'h0; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_113 = 3'h2 == x_10 ? b_sext : _pp_temp_T_111; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_115 = 3'h3 == x_10 ? bx2 : _pp_temp_T_113; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_117 = 3'h4 == x_10 ? neg_bx2 : _pp_temp_T_115; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_119 = 3'h5 == x_10 ? neg_b : _pp_temp_T_117; // @[Mux.scala 81:58]
  wire [65:0] pp_temp_10 = 3'h6 == x_10 ? neg_b : _pp_temp_T_119; // @[Mux.scala 81:58]
  wire  s_10 = pp_temp_10[65]; // @[Multiplier.scala 90:20]
  wire [1:0] _t_T_51 = 3'h4 == x_9 ? 2'h2 : 2'h0; // @[Mux.scala 81:58]
  wire [1:0] _t_T_53 = 3'h5 == x_9 ? 2'h1 : _t_T_51; // @[Mux.scala 81:58]
  wire [1:0] t_10 = 3'h6 == x_9 ? 2'h1 : _t_T_53; // @[Mux.scala 81:58]
  wire  _T_709 = ~s_10; // @[Multiplier.scala 103:24]
  wire [69:0] pp_10 = {1'h1,_T_709,pp_temp_10,t_10}; // @[Cat.scala 31:58]
  wire [2:0] x_11 = io_a[23:21]; // @[Multiplier.scala 81:90]
  wire [65:0] _pp_temp_T_122 = 3'h1 == x_11 ? b_sext : 66'h0; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_124 = 3'h2 == x_11 ? b_sext : _pp_temp_T_122; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_126 = 3'h3 == x_11 ? bx2 : _pp_temp_T_124; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_128 = 3'h4 == x_11 ? neg_bx2 : _pp_temp_T_126; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_130 = 3'h5 == x_11 ? neg_b : _pp_temp_T_128; // @[Mux.scala 81:58]
  wire [65:0] pp_temp_11 = 3'h6 == x_11 ? neg_b : _pp_temp_T_130; // @[Mux.scala 81:58]
  wire  s_11 = pp_temp_11[65]; // @[Multiplier.scala 90:20]
  wire [1:0] _t_T_56 = 3'h4 == x_10 ? 2'h2 : 2'h0; // @[Mux.scala 81:58]
  wire [1:0] _t_T_58 = 3'h5 == x_10 ? 2'h1 : _t_T_56; // @[Mux.scala 81:58]
  wire [1:0] t_11 = 3'h6 == x_10 ? 2'h1 : _t_T_58; // @[Mux.scala 81:58]
  wire  _T_780 = ~s_11; // @[Multiplier.scala 103:24]
  wire [69:0] pp_11 = {1'h1,_T_780,pp_temp_11,t_11}; // @[Cat.scala 31:58]
  wire [2:0] x_12 = io_a[25:23]; // @[Multiplier.scala 81:90]
  wire [65:0] _pp_temp_T_133 = 3'h1 == x_12 ? b_sext : 66'h0; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_135 = 3'h2 == x_12 ? b_sext : _pp_temp_T_133; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_137 = 3'h3 == x_12 ? bx2 : _pp_temp_T_135; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_139 = 3'h4 == x_12 ? neg_bx2 : _pp_temp_T_137; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_141 = 3'h5 == x_12 ? neg_b : _pp_temp_T_139; // @[Mux.scala 81:58]
  wire [65:0] pp_temp_12 = 3'h6 == x_12 ? neg_b : _pp_temp_T_141; // @[Mux.scala 81:58]
  wire  s_12 = pp_temp_12[65]; // @[Multiplier.scala 90:20]
  wire [1:0] _t_T_61 = 3'h4 == x_11 ? 2'h2 : 2'h0; // @[Mux.scala 81:58]
  wire [1:0] _t_T_63 = 3'h5 == x_11 ? 2'h1 : _t_T_61; // @[Mux.scala 81:58]
  wire [1:0] t_12 = 3'h6 == x_11 ? 2'h1 : _t_T_63; // @[Mux.scala 81:58]
  wire  _T_851 = ~s_12; // @[Multiplier.scala 103:24]
  wire [69:0] pp_12 = {1'h1,_T_851,pp_temp_12,t_12}; // @[Cat.scala 31:58]
  wire [2:0] x_13 = io_a[27:25]; // @[Multiplier.scala 81:90]
  wire [65:0] _pp_temp_T_144 = 3'h1 == x_13 ? b_sext : 66'h0; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_146 = 3'h2 == x_13 ? b_sext : _pp_temp_T_144; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_148 = 3'h3 == x_13 ? bx2 : _pp_temp_T_146; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_150 = 3'h4 == x_13 ? neg_bx2 : _pp_temp_T_148; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_152 = 3'h5 == x_13 ? neg_b : _pp_temp_T_150; // @[Mux.scala 81:58]
  wire [65:0] pp_temp_13 = 3'h6 == x_13 ? neg_b : _pp_temp_T_152; // @[Mux.scala 81:58]
  wire  s_13 = pp_temp_13[65]; // @[Multiplier.scala 90:20]
  wire [1:0] _t_T_66 = 3'h4 == x_12 ? 2'h2 : 2'h0; // @[Mux.scala 81:58]
  wire [1:0] _t_T_68 = 3'h5 == x_12 ? 2'h1 : _t_T_66; // @[Mux.scala 81:58]
  wire [1:0] t_13 = 3'h6 == x_12 ? 2'h1 : _t_T_68; // @[Mux.scala 81:58]
  wire  _T_922 = ~s_13; // @[Multiplier.scala 103:24]
  wire [69:0] pp_13 = {1'h1,_T_922,pp_temp_13,t_13}; // @[Cat.scala 31:58]
  wire [2:0] x_14 = io_a[29:27]; // @[Multiplier.scala 81:90]
  wire [65:0] _pp_temp_T_155 = 3'h1 == x_14 ? b_sext : 66'h0; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_157 = 3'h2 == x_14 ? b_sext : _pp_temp_T_155; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_159 = 3'h3 == x_14 ? bx2 : _pp_temp_T_157; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_161 = 3'h4 == x_14 ? neg_bx2 : _pp_temp_T_159; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_163 = 3'h5 == x_14 ? neg_b : _pp_temp_T_161; // @[Mux.scala 81:58]
  wire [65:0] pp_temp_14 = 3'h6 == x_14 ? neg_b : _pp_temp_T_163; // @[Mux.scala 81:58]
  wire  s_14 = pp_temp_14[65]; // @[Multiplier.scala 90:20]
  wire [1:0] _t_T_71 = 3'h4 == x_13 ? 2'h2 : 2'h0; // @[Mux.scala 81:58]
  wire [1:0] _t_T_73 = 3'h5 == x_13 ? 2'h1 : _t_T_71; // @[Mux.scala 81:58]
  wire [1:0] t_14 = 3'h6 == x_13 ? 2'h1 : _t_T_73; // @[Mux.scala 81:58]
  wire  _T_993 = ~s_14; // @[Multiplier.scala 103:24]
  wire [69:0] pp_14 = {1'h1,_T_993,pp_temp_14,t_14}; // @[Cat.scala 31:58]
  wire [2:0] x_15 = io_a[31:29]; // @[Multiplier.scala 81:90]
  wire [65:0] _pp_temp_T_166 = 3'h1 == x_15 ? b_sext : 66'h0; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_168 = 3'h2 == x_15 ? b_sext : _pp_temp_T_166; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_170 = 3'h3 == x_15 ? bx2 : _pp_temp_T_168; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_172 = 3'h4 == x_15 ? neg_bx2 : _pp_temp_T_170; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_174 = 3'h5 == x_15 ? neg_b : _pp_temp_T_172; // @[Mux.scala 81:58]
  wire [65:0] pp_temp_15 = 3'h6 == x_15 ? neg_b : _pp_temp_T_174; // @[Mux.scala 81:58]
  wire  s_15 = pp_temp_15[65]; // @[Multiplier.scala 90:20]
  wire [1:0] _t_T_76 = 3'h4 == x_14 ? 2'h2 : 2'h0; // @[Mux.scala 81:58]
  wire [1:0] _t_T_78 = 3'h5 == x_14 ? 2'h1 : _t_T_76; // @[Mux.scala 81:58]
  wire [1:0] t_15 = 3'h6 == x_14 ? 2'h1 : _t_T_78; // @[Mux.scala 81:58]
  wire  _T_1064 = ~s_15; // @[Multiplier.scala 103:24]
  wire [69:0] pp_15 = {1'h1,_T_1064,pp_temp_15,t_15}; // @[Cat.scala 31:58]
  wire [2:0] x_16 = io_a[33:31]; // @[Multiplier.scala 81:90]
  wire [65:0] _pp_temp_T_177 = 3'h1 == x_16 ? b_sext : 66'h0; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_179 = 3'h2 == x_16 ? b_sext : _pp_temp_T_177; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_181 = 3'h3 == x_16 ? bx2 : _pp_temp_T_179; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_183 = 3'h4 == x_16 ? neg_bx2 : _pp_temp_T_181; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_185 = 3'h5 == x_16 ? neg_b : _pp_temp_T_183; // @[Mux.scala 81:58]
  wire [65:0] pp_temp_16 = 3'h6 == x_16 ? neg_b : _pp_temp_T_185; // @[Mux.scala 81:58]
  wire  s_16 = pp_temp_16[65]; // @[Multiplier.scala 90:20]
  wire [1:0] _t_T_81 = 3'h4 == x_15 ? 2'h2 : 2'h0; // @[Mux.scala 81:58]
  wire [1:0] _t_T_83 = 3'h5 == x_15 ? 2'h1 : _t_T_81; // @[Mux.scala 81:58]
  wire [1:0] t_16 = 3'h6 == x_15 ? 2'h1 : _t_T_83; // @[Mux.scala 81:58]
  wire  _T_1135 = ~s_16; // @[Multiplier.scala 103:24]
  wire [69:0] pp_16 = {1'h1,_T_1135,pp_temp_16,t_16}; // @[Cat.scala 31:58]
  wire [2:0] x_17 = io_a[35:33]; // @[Multiplier.scala 81:90]
  wire [65:0] _pp_temp_T_188 = 3'h1 == x_17 ? b_sext : 66'h0; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_190 = 3'h2 == x_17 ? b_sext : _pp_temp_T_188; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_192 = 3'h3 == x_17 ? bx2 : _pp_temp_T_190; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_194 = 3'h4 == x_17 ? neg_bx2 : _pp_temp_T_192; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_196 = 3'h5 == x_17 ? neg_b : _pp_temp_T_194; // @[Mux.scala 81:58]
  wire [65:0] pp_temp_17 = 3'h6 == x_17 ? neg_b : _pp_temp_T_196; // @[Mux.scala 81:58]
  wire  s_17 = pp_temp_17[65]; // @[Multiplier.scala 90:20]
  wire [1:0] _t_T_86 = 3'h4 == x_16 ? 2'h2 : 2'h0; // @[Mux.scala 81:58]
  wire [1:0] _t_T_88 = 3'h5 == x_16 ? 2'h1 : _t_T_86; // @[Mux.scala 81:58]
  wire [1:0] t_17 = 3'h6 == x_16 ? 2'h1 : _t_T_88; // @[Mux.scala 81:58]
  wire  _T_1206 = ~s_17; // @[Multiplier.scala 103:24]
  wire [69:0] pp_17 = {1'h1,_T_1206,pp_temp_17,t_17}; // @[Cat.scala 31:58]
  wire [2:0] x_18 = io_a[37:35]; // @[Multiplier.scala 81:90]
  wire [65:0] _pp_temp_T_199 = 3'h1 == x_18 ? b_sext : 66'h0; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_201 = 3'h2 == x_18 ? b_sext : _pp_temp_T_199; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_203 = 3'h3 == x_18 ? bx2 : _pp_temp_T_201; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_205 = 3'h4 == x_18 ? neg_bx2 : _pp_temp_T_203; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_207 = 3'h5 == x_18 ? neg_b : _pp_temp_T_205; // @[Mux.scala 81:58]
  wire [65:0] pp_temp_18 = 3'h6 == x_18 ? neg_b : _pp_temp_T_207; // @[Mux.scala 81:58]
  wire  s_18 = pp_temp_18[65]; // @[Multiplier.scala 90:20]
  wire [1:0] _t_T_91 = 3'h4 == x_17 ? 2'h2 : 2'h0; // @[Mux.scala 81:58]
  wire [1:0] _t_T_93 = 3'h5 == x_17 ? 2'h1 : _t_T_91; // @[Mux.scala 81:58]
  wire [1:0] t_18 = 3'h6 == x_17 ? 2'h1 : _t_T_93; // @[Mux.scala 81:58]
  wire  _T_1277 = ~s_18; // @[Multiplier.scala 103:24]
  wire [69:0] pp_18 = {1'h1,_T_1277,pp_temp_18,t_18}; // @[Cat.scala 31:58]
  wire [2:0] x_19 = io_a[39:37]; // @[Multiplier.scala 81:90]
  wire [65:0] _pp_temp_T_210 = 3'h1 == x_19 ? b_sext : 66'h0; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_212 = 3'h2 == x_19 ? b_sext : _pp_temp_T_210; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_214 = 3'h3 == x_19 ? bx2 : _pp_temp_T_212; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_216 = 3'h4 == x_19 ? neg_bx2 : _pp_temp_T_214; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_218 = 3'h5 == x_19 ? neg_b : _pp_temp_T_216; // @[Mux.scala 81:58]
  wire [65:0] pp_temp_19 = 3'h6 == x_19 ? neg_b : _pp_temp_T_218; // @[Mux.scala 81:58]
  wire  s_19 = pp_temp_19[65]; // @[Multiplier.scala 90:20]
  wire [1:0] _t_T_96 = 3'h4 == x_18 ? 2'h2 : 2'h0; // @[Mux.scala 81:58]
  wire [1:0] _t_T_98 = 3'h5 == x_18 ? 2'h1 : _t_T_96; // @[Mux.scala 81:58]
  wire [1:0] t_19 = 3'h6 == x_18 ? 2'h1 : _t_T_98; // @[Mux.scala 81:58]
  wire  _T_1348 = ~s_19; // @[Multiplier.scala 103:24]
  wire [69:0] pp_19 = {1'h1,_T_1348,pp_temp_19,t_19}; // @[Cat.scala 31:58]
  wire [2:0] x_20 = io_a[41:39]; // @[Multiplier.scala 81:90]
  wire [65:0] _pp_temp_T_221 = 3'h1 == x_20 ? b_sext : 66'h0; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_223 = 3'h2 == x_20 ? b_sext : _pp_temp_T_221; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_225 = 3'h3 == x_20 ? bx2 : _pp_temp_T_223; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_227 = 3'h4 == x_20 ? neg_bx2 : _pp_temp_T_225; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_229 = 3'h5 == x_20 ? neg_b : _pp_temp_T_227; // @[Mux.scala 81:58]
  wire [65:0] pp_temp_20 = 3'h6 == x_20 ? neg_b : _pp_temp_T_229; // @[Mux.scala 81:58]
  wire  s_20 = pp_temp_20[65]; // @[Multiplier.scala 90:20]
  wire [1:0] _t_T_101 = 3'h4 == x_19 ? 2'h2 : 2'h0; // @[Mux.scala 81:58]
  wire [1:0] _t_T_103 = 3'h5 == x_19 ? 2'h1 : _t_T_101; // @[Mux.scala 81:58]
  wire [1:0] t_20 = 3'h6 == x_19 ? 2'h1 : _t_T_103; // @[Mux.scala 81:58]
  wire  _T_1419 = ~s_20; // @[Multiplier.scala 103:24]
  wire [69:0] pp_20 = {1'h1,_T_1419,pp_temp_20,t_20}; // @[Cat.scala 31:58]
  wire [2:0] x_21 = io_a[43:41]; // @[Multiplier.scala 81:90]
  wire [65:0] _pp_temp_T_232 = 3'h1 == x_21 ? b_sext : 66'h0; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_234 = 3'h2 == x_21 ? b_sext : _pp_temp_T_232; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_236 = 3'h3 == x_21 ? bx2 : _pp_temp_T_234; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_238 = 3'h4 == x_21 ? neg_bx2 : _pp_temp_T_236; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_240 = 3'h5 == x_21 ? neg_b : _pp_temp_T_238; // @[Mux.scala 81:58]
  wire [65:0] pp_temp_21 = 3'h6 == x_21 ? neg_b : _pp_temp_T_240; // @[Mux.scala 81:58]
  wire  s_21 = pp_temp_21[65]; // @[Multiplier.scala 90:20]
  wire [1:0] _t_T_106 = 3'h4 == x_20 ? 2'h2 : 2'h0; // @[Mux.scala 81:58]
  wire [1:0] _t_T_108 = 3'h5 == x_20 ? 2'h1 : _t_T_106; // @[Mux.scala 81:58]
  wire [1:0] t_21 = 3'h6 == x_20 ? 2'h1 : _t_T_108; // @[Mux.scala 81:58]
  wire  _T_1490 = ~s_21; // @[Multiplier.scala 103:24]
  wire [69:0] pp_21 = {1'h1,_T_1490,pp_temp_21,t_21}; // @[Cat.scala 31:58]
  wire [2:0] x_22 = io_a[45:43]; // @[Multiplier.scala 81:90]
  wire [65:0] _pp_temp_T_243 = 3'h1 == x_22 ? b_sext : 66'h0; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_245 = 3'h2 == x_22 ? b_sext : _pp_temp_T_243; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_247 = 3'h3 == x_22 ? bx2 : _pp_temp_T_245; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_249 = 3'h4 == x_22 ? neg_bx2 : _pp_temp_T_247; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_251 = 3'h5 == x_22 ? neg_b : _pp_temp_T_249; // @[Mux.scala 81:58]
  wire [65:0] pp_temp_22 = 3'h6 == x_22 ? neg_b : _pp_temp_T_251; // @[Mux.scala 81:58]
  wire  s_22 = pp_temp_22[65]; // @[Multiplier.scala 90:20]
  wire [1:0] _t_T_111 = 3'h4 == x_21 ? 2'h2 : 2'h0; // @[Mux.scala 81:58]
  wire [1:0] _t_T_113 = 3'h5 == x_21 ? 2'h1 : _t_T_111; // @[Mux.scala 81:58]
  wire [1:0] t_22 = 3'h6 == x_21 ? 2'h1 : _t_T_113; // @[Mux.scala 81:58]
  wire  _T_1561 = ~s_22; // @[Multiplier.scala 103:24]
  wire [69:0] pp_22 = {1'h1,_T_1561,pp_temp_22,t_22}; // @[Cat.scala 31:58]
  wire [2:0] x_23 = io_a[47:45]; // @[Multiplier.scala 81:90]
  wire [65:0] _pp_temp_T_254 = 3'h1 == x_23 ? b_sext : 66'h0; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_256 = 3'h2 == x_23 ? b_sext : _pp_temp_T_254; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_258 = 3'h3 == x_23 ? bx2 : _pp_temp_T_256; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_260 = 3'h4 == x_23 ? neg_bx2 : _pp_temp_T_258; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_262 = 3'h5 == x_23 ? neg_b : _pp_temp_T_260; // @[Mux.scala 81:58]
  wire [65:0] pp_temp_23 = 3'h6 == x_23 ? neg_b : _pp_temp_T_262; // @[Mux.scala 81:58]
  wire  s_23 = pp_temp_23[65]; // @[Multiplier.scala 90:20]
  wire [1:0] _t_T_116 = 3'h4 == x_22 ? 2'h2 : 2'h0; // @[Mux.scala 81:58]
  wire [1:0] _t_T_118 = 3'h5 == x_22 ? 2'h1 : _t_T_116; // @[Mux.scala 81:58]
  wire [1:0] t_23 = 3'h6 == x_22 ? 2'h1 : _t_T_118; // @[Mux.scala 81:58]
  wire  _T_1632 = ~s_23; // @[Multiplier.scala 103:24]
  wire [69:0] pp_23 = {1'h1,_T_1632,pp_temp_23,t_23}; // @[Cat.scala 31:58]
  wire [2:0] x_24 = io_a[49:47]; // @[Multiplier.scala 81:90]
  wire [65:0] _pp_temp_T_265 = 3'h1 == x_24 ? b_sext : 66'h0; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_267 = 3'h2 == x_24 ? b_sext : _pp_temp_T_265; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_269 = 3'h3 == x_24 ? bx2 : _pp_temp_T_267; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_271 = 3'h4 == x_24 ? neg_bx2 : _pp_temp_T_269; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_273 = 3'h5 == x_24 ? neg_b : _pp_temp_T_271; // @[Mux.scala 81:58]
  wire [65:0] pp_temp_24 = 3'h6 == x_24 ? neg_b : _pp_temp_T_273; // @[Mux.scala 81:58]
  wire  s_24 = pp_temp_24[65]; // @[Multiplier.scala 90:20]
  wire [1:0] _t_T_121 = 3'h4 == x_23 ? 2'h2 : 2'h0; // @[Mux.scala 81:58]
  wire [1:0] _t_T_123 = 3'h5 == x_23 ? 2'h1 : _t_T_121; // @[Mux.scala 81:58]
  wire [1:0] t_24 = 3'h6 == x_23 ? 2'h1 : _t_T_123; // @[Mux.scala 81:58]
  wire  _T_1703 = ~s_24; // @[Multiplier.scala 103:24]
  wire [69:0] pp_24 = {1'h1,_T_1703,pp_temp_24,t_24}; // @[Cat.scala 31:58]
  wire [2:0] x_25 = io_a[51:49]; // @[Multiplier.scala 81:90]
  wire [65:0] _pp_temp_T_276 = 3'h1 == x_25 ? b_sext : 66'h0; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_278 = 3'h2 == x_25 ? b_sext : _pp_temp_T_276; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_280 = 3'h3 == x_25 ? bx2 : _pp_temp_T_278; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_282 = 3'h4 == x_25 ? neg_bx2 : _pp_temp_T_280; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_284 = 3'h5 == x_25 ? neg_b : _pp_temp_T_282; // @[Mux.scala 81:58]
  wire [65:0] pp_temp_25 = 3'h6 == x_25 ? neg_b : _pp_temp_T_284; // @[Mux.scala 81:58]
  wire  s_25 = pp_temp_25[65]; // @[Multiplier.scala 90:20]
  wire [1:0] _t_T_126 = 3'h4 == x_24 ? 2'h2 : 2'h0; // @[Mux.scala 81:58]
  wire [1:0] _t_T_128 = 3'h5 == x_24 ? 2'h1 : _t_T_126; // @[Mux.scala 81:58]
  wire [1:0] t_25 = 3'h6 == x_24 ? 2'h1 : _t_T_128; // @[Mux.scala 81:58]
  wire  _T_1774 = ~s_25; // @[Multiplier.scala 103:24]
  wire [69:0] pp_25 = {1'h1,_T_1774,pp_temp_25,t_25}; // @[Cat.scala 31:58]
  wire [2:0] x_26 = io_a[53:51]; // @[Multiplier.scala 81:90]
  wire [65:0] _pp_temp_T_287 = 3'h1 == x_26 ? b_sext : 66'h0; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_289 = 3'h2 == x_26 ? b_sext : _pp_temp_T_287; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_291 = 3'h3 == x_26 ? bx2 : _pp_temp_T_289; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_293 = 3'h4 == x_26 ? neg_bx2 : _pp_temp_T_291; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_295 = 3'h5 == x_26 ? neg_b : _pp_temp_T_293; // @[Mux.scala 81:58]
  wire [65:0] pp_temp_26 = 3'h6 == x_26 ? neg_b : _pp_temp_T_295; // @[Mux.scala 81:58]
  wire  s_26 = pp_temp_26[65]; // @[Multiplier.scala 90:20]
  wire [1:0] _t_T_131 = 3'h4 == x_25 ? 2'h2 : 2'h0; // @[Mux.scala 81:58]
  wire [1:0] _t_T_133 = 3'h5 == x_25 ? 2'h1 : _t_T_131; // @[Mux.scala 81:58]
  wire [1:0] t_26 = 3'h6 == x_25 ? 2'h1 : _t_T_133; // @[Mux.scala 81:58]
  wire  _T_1845 = ~s_26; // @[Multiplier.scala 103:24]
  wire [69:0] pp_26 = {1'h1,_T_1845,pp_temp_26,t_26}; // @[Cat.scala 31:58]
  wire [2:0] x_27 = io_a[55:53]; // @[Multiplier.scala 81:90]
  wire [65:0] _pp_temp_T_298 = 3'h1 == x_27 ? b_sext : 66'h0; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_300 = 3'h2 == x_27 ? b_sext : _pp_temp_T_298; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_302 = 3'h3 == x_27 ? bx2 : _pp_temp_T_300; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_304 = 3'h4 == x_27 ? neg_bx2 : _pp_temp_T_302; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_306 = 3'h5 == x_27 ? neg_b : _pp_temp_T_304; // @[Mux.scala 81:58]
  wire [65:0] pp_temp_27 = 3'h6 == x_27 ? neg_b : _pp_temp_T_306; // @[Mux.scala 81:58]
  wire  s_27 = pp_temp_27[65]; // @[Multiplier.scala 90:20]
  wire [1:0] _t_T_136 = 3'h4 == x_26 ? 2'h2 : 2'h0; // @[Mux.scala 81:58]
  wire [1:0] _t_T_138 = 3'h5 == x_26 ? 2'h1 : _t_T_136; // @[Mux.scala 81:58]
  wire [1:0] t_27 = 3'h6 == x_26 ? 2'h1 : _t_T_138; // @[Mux.scala 81:58]
  wire  _T_1916 = ~s_27; // @[Multiplier.scala 103:24]
  wire [69:0] pp_27 = {1'h1,_T_1916,pp_temp_27,t_27}; // @[Cat.scala 31:58]
  wire [2:0] x_28 = io_a[57:55]; // @[Multiplier.scala 81:90]
  wire [65:0] _pp_temp_T_309 = 3'h1 == x_28 ? b_sext : 66'h0; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_311 = 3'h2 == x_28 ? b_sext : _pp_temp_T_309; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_313 = 3'h3 == x_28 ? bx2 : _pp_temp_T_311; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_315 = 3'h4 == x_28 ? neg_bx2 : _pp_temp_T_313; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_317 = 3'h5 == x_28 ? neg_b : _pp_temp_T_315; // @[Mux.scala 81:58]
  wire [65:0] pp_temp_28 = 3'h6 == x_28 ? neg_b : _pp_temp_T_317; // @[Mux.scala 81:58]
  wire  s_28 = pp_temp_28[65]; // @[Multiplier.scala 90:20]
  wire [1:0] _t_T_141 = 3'h4 == x_27 ? 2'h2 : 2'h0; // @[Mux.scala 81:58]
  wire [1:0] _t_T_143 = 3'h5 == x_27 ? 2'h1 : _t_T_141; // @[Mux.scala 81:58]
  wire [1:0] t_28 = 3'h6 == x_27 ? 2'h1 : _t_T_143; // @[Mux.scala 81:58]
  wire  _T_1987 = ~s_28; // @[Multiplier.scala 103:24]
  wire [69:0] pp_28 = {1'h1,_T_1987,pp_temp_28,t_28}; // @[Cat.scala 31:58]
  wire [2:0] x_29 = io_a[59:57]; // @[Multiplier.scala 81:90]
  wire [65:0] _pp_temp_T_320 = 3'h1 == x_29 ? b_sext : 66'h0; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_322 = 3'h2 == x_29 ? b_sext : _pp_temp_T_320; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_324 = 3'h3 == x_29 ? bx2 : _pp_temp_T_322; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_326 = 3'h4 == x_29 ? neg_bx2 : _pp_temp_T_324; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_328 = 3'h5 == x_29 ? neg_b : _pp_temp_T_326; // @[Mux.scala 81:58]
  wire [65:0] pp_temp_29 = 3'h6 == x_29 ? neg_b : _pp_temp_T_328; // @[Mux.scala 81:58]
  wire  s_29 = pp_temp_29[65]; // @[Multiplier.scala 90:20]
  wire [1:0] _t_T_146 = 3'h4 == x_28 ? 2'h2 : 2'h0; // @[Mux.scala 81:58]
  wire [1:0] _t_T_148 = 3'h5 == x_28 ? 2'h1 : _t_T_146; // @[Mux.scala 81:58]
  wire [1:0] t_29 = 3'h6 == x_28 ? 2'h1 : _t_T_148; // @[Mux.scala 81:58]
  wire  _T_2058 = ~s_29; // @[Multiplier.scala 103:24]
  wire [69:0] pp_29 = {1'h1,_T_2058,pp_temp_29,t_29}; // @[Cat.scala 31:58]
  wire [2:0] x_30 = io_a[61:59]; // @[Multiplier.scala 81:90]
  wire [65:0] _pp_temp_T_331 = 3'h1 == x_30 ? b_sext : 66'h0; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_333 = 3'h2 == x_30 ? b_sext : _pp_temp_T_331; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_335 = 3'h3 == x_30 ? bx2 : _pp_temp_T_333; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_337 = 3'h4 == x_30 ? neg_bx2 : _pp_temp_T_335; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_339 = 3'h5 == x_30 ? neg_b : _pp_temp_T_337; // @[Mux.scala 81:58]
  wire [65:0] pp_temp_30 = 3'h6 == x_30 ? neg_b : _pp_temp_T_339; // @[Mux.scala 81:58]
  wire  s_30 = pp_temp_30[65]; // @[Multiplier.scala 90:20]
  wire [1:0] _t_T_151 = 3'h4 == x_29 ? 2'h2 : 2'h0; // @[Mux.scala 81:58]
  wire [1:0] _t_T_153 = 3'h5 == x_29 ? 2'h1 : _t_T_151; // @[Mux.scala 81:58]
  wire [1:0] t_30 = 3'h6 == x_29 ? 2'h1 : _t_T_153; // @[Mux.scala 81:58]
  wire  _T_2129 = ~s_30; // @[Multiplier.scala 103:24]
  wire [69:0] pp_30 = {1'h1,_T_2129,pp_temp_30,t_30}; // @[Cat.scala 31:58]
  wire [2:0] x_31 = io_a[63:61]; // @[Multiplier.scala 81:90]
  wire [65:0] _pp_temp_T_342 = 3'h1 == x_31 ? b_sext : 66'h0; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_344 = 3'h2 == x_31 ? b_sext : _pp_temp_T_342; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_346 = 3'h3 == x_31 ? bx2 : _pp_temp_T_344; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_348 = 3'h4 == x_31 ? neg_bx2 : _pp_temp_T_346; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_350 = 3'h5 == x_31 ? neg_b : _pp_temp_T_348; // @[Mux.scala 81:58]
  wire [65:0] pp_temp_31 = 3'h6 == x_31 ? neg_b : _pp_temp_T_350; // @[Mux.scala 81:58]
  wire  s_31 = pp_temp_31[65]; // @[Multiplier.scala 90:20]
  wire [1:0] _t_T_156 = 3'h4 == x_30 ? 2'h2 : 2'h0; // @[Mux.scala 81:58]
  wire [1:0] _t_T_158 = 3'h5 == x_30 ? 2'h1 : _t_T_156; // @[Mux.scala 81:58]
  wire [1:0] t_31 = 3'h6 == x_30 ? 2'h1 : _t_T_158; // @[Mux.scala 81:58]
  wire  _T_2200 = ~s_31; // @[Multiplier.scala 103:24]
  wire [69:0] pp_31 = {1'h1,_T_2200,pp_temp_31,t_31}; // @[Cat.scala 31:58]
  wire  x_signBit = io_a[64]; // @[BitUtils.scala 80:20]
  wire [2:0] last_x_1 = {x_signBit,io_a[64:63]}; // @[Cat.scala 31:58]
  wire [65:0] _pp_temp_T_353 = 3'h1 == last_x_1 ? b_sext : 66'h0; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_355 = 3'h2 == last_x_1 ? b_sext : _pp_temp_T_353; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_357 = 3'h3 == last_x_1 ? bx2 : _pp_temp_T_355; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_359 = 3'h4 == last_x_1 ? neg_bx2 : _pp_temp_T_357; // @[Mux.scala 81:58]
  wire [65:0] _pp_temp_T_361 = 3'h5 == last_x_1 ? neg_b : _pp_temp_T_359; // @[Mux.scala 81:58]
  wire [65:0] pp_temp_32 = 3'h6 == last_x_1 ? neg_b : _pp_temp_T_361; // @[Mux.scala 81:58]
  wire  s_32 = pp_temp_32[65]; // @[Multiplier.scala 90:20]
  wire [1:0] _t_T_161 = 3'h4 == x_31 ? 2'h2 : 2'h0; // @[Mux.scala 81:58]
  wire [1:0] _t_T_163 = 3'h5 == x_31 ? 2'h1 : _t_T_161; // @[Mux.scala 81:58]
  wire [1:0] t_32 = 3'h6 == x_31 ? 2'h1 : _t_T_163; // @[Mux.scala 81:58]
  wire  _T_2271 = ~s_32; // @[Multiplier.scala 101:14]
  wire [68:0] pp_32 = {_T_2271,pp_temp_32,t_32}; // @[Cat.scala 31:58]
  reg  r; // @[Reg.scala 16:16]
  reg  r_1; // @[Reg.scala 16:16]
  reg  r_2; // @[Reg.scala 16:16]
  reg  r_3; // @[Reg.scala 16:16]
  reg  r_4; // @[Reg.scala 16:16]
  reg  r_5; // @[Reg.scala 16:16]
  reg  r_6; // @[Reg.scala 16:16]
  reg  r_7; // @[Reg.scala 16:16]
  reg  r_8; // @[Reg.scala 16:16]
  reg  r_9; // @[Reg.scala 16:16]
  reg  r_10; // @[Reg.scala 16:16]
  reg  r_11; // @[Reg.scala 16:16]
  reg  r_12; // @[Reg.scala 16:16]
  reg  r_13; // @[Reg.scala 16:16]
  reg  r_14; // @[Reg.scala 16:16]
  reg  r_15; // @[Reg.scala 16:16]
  reg  r_16; // @[Reg.scala 16:16]
  reg  r_17; // @[Reg.scala 16:16]
  reg  r_18; // @[Reg.scala 16:16]
  reg  r_19; // @[Reg.scala 16:16]
  reg  r_20; // @[Reg.scala 16:16]
  reg  r_21; // @[Reg.scala 16:16]
  reg  r_22; // @[Reg.scala 16:16]
  reg  r_23; // @[Reg.scala 16:16]
  reg  r_24; // @[Reg.scala 16:16]
  reg  r_25; // @[Reg.scala 16:16]
  reg  r_26; // @[Reg.scala 16:16]
  reg  r_27; // @[Reg.scala 16:16]
  reg  r_28; // @[Reg.scala 16:16]
  reg  r_29; // @[Reg.scala 16:16]
  reg  r_30; // @[Reg.scala 16:16]
  reg  r_31; // @[Reg.scala 16:16]
  reg  r_32; // @[Reg.scala 16:16]
  reg  r_33; // @[Reg.scala 16:16]
  reg  r_34; // @[Reg.scala 16:16]
  reg  r_35; // @[Reg.scala 16:16]
  reg  r_36; // @[Reg.scala 16:16]
  reg  r_37; // @[Reg.scala 16:16]
  reg  r_38; // @[Reg.scala 16:16]
  reg  r_39; // @[Reg.scala 16:16]
  reg  r_40; // @[Reg.scala 16:16]
  reg  r_41; // @[Reg.scala 16:16]
  reg  r_42; // @[Reg.scala 16:16]
  reg  r_43; // @[Reg.scala 16:16]
  reg  r_44; // @[Reg.scala 16:16]
  reg  r_45; // @[Reg.scala 16:16]
  reg  r_46; // @[Reg.scala 16:16]
  reg  r_47; // @[Reg.scala 16:16]
  reg  r_48; // @[Reg.scala 16:16]
  reg  r_49; // @[Reg.scala 16:16]
  reg  r_50; // @[Reg.scala 16:16]
  reg  r_51; // @[Reg.scala 16:16]
  reg  r_52; // @[Reg.scala 16:16]
  reg  r_53; // @[Reg.scala 16:16]
  reg  r_54; // @[Reg.scala 16:16]
  reg  r_55; // @[Reg.scala 16:16]
  reg  r_56; // @[Reg.scala 16:16]
  reg  r_57; // @[Reg.scala 16:16]
  reg  r_58; // @[Reg.scala 16:16]
  reg  r_59; // @[Reg.scala 16:16]
  reg  r_60; // @[Reg.scala 16:16]
  reg  r_61; // @[Reg.scala 16:16]
  reg  r_62; // @[Reg.scala 16:16]
  reg  r_63; // @[Reg.scala 16:16]
  reg  r_64; // @[Reg.scala 16:16]
  reg  r_65; // @[Reg.scala 16:16]
  reg  r_66; // @[Reg.scala 16:16]
  reg  r_67; // @[Reg.scala 16:16]
  reg  r_68; // @[Reg.scala 16:16]
  reg  r_69; // @[Reg.scala 16:16]
  reg  r_70; // @[Reg.scala 16:16]
  reg  r_71; // @[Reg.scala 16:16]
  reg  r_72; // @[Reg.scala 16:16]
  reg  r_73; // @[Reg.scala 16:16]
  reg  r_74; // @[Reg.scala 16:16]
  reg  r_75; // @[Reg.scala 16:16]
  reg  r_76; // @[Reg.scala 16:16]
  reg  r_77; // @[Reg.scala 16:16]
  reg  r_78; // @[Reg.scala 16:16]
  reg  r_79; // @[Reg.scala 16:16]
  reg  r_80; // @[Reg.scala 16:16]
  reg  r_81; // @[Reg.scala 16:16]
  reg  r_82; // @[Reg.scala 16:16]
  reg  r_83; // @[Reg.scala 16:16]
  reg  r_84; // @[Reg.scala 16:16]
  reg  r_85; // @[Reg.scala 16:16]
  reg  r_86; // @[Reg.scala 16:16]
  reg  r_87; // @[Reg.scala 16:16]
  reg  r_88; // @[Reg.scala 16:16]
  reg  r_89; // @[Reg.scala 16:16]
  reg  r_90; // @[Reg.scala 16:16]
  reg  r_91; // @[Reg.scala 16:16]
  reg  r_92; // @[Reg.scala 16:16]
  reg  r_93; // @[Reg.scala 16:16]
  reg  r_94; // @[Reg.scala 16:16]
  reg  r_95; // @[Reg.scala 16:16]
  reg  r_96; // @[Reg.scala 16:16]
  reg  r_97; // @[Reg.scala 16:16]
  reg  r_98; // @[Reg.scala 16:16]
  reg  r_99; // @[Reg.scala 16:16]
  reg  r_100; // @[Reg.scala 16:16]
  reg  r_101; // @[Reg.scala 16:16]
  reg  r_102; // @[Reg.scala 16:16]
  reg  r_103; // @[Reg.scala 16:16]
  reg  r_104; // @[Reg.scala 16:16]
  reg  r_105; // @[Reg.scala 16:16]
  reg  r_106; // @[Reg.scala 16:16]
  reg  r_107; // @[Reg.scala 16:16]
  reg  r_108; // @[Reg.scala 16:16]
  reg  r_109; // @[Reg.scala 16:16]
  reg  r_110; // @[Reg.scala 16:16]
  reg  r_111; // @[Reg.scala 16:16]
  reg  r_112; // @[Reg.scala 16:16]
  reg  r_113; // @[Reg.scala 16:16]
  reg  r_114; // @[Reg.scala 16:16]
  reg  r_115; // @[Reg.scala 16:16]
  reg  r_116; // @[Reg.scala 16:16]
  reg  r_117; // @[Reg.scala 16:16]
  reg  r_118; // @[Reg.scala 16:16]
  reg  r_119; // @[Reg.scala 16:16]
  reg  r_120; // @[Reg.scala 16:16]
  reg  r_121; // @[Reg.scala 16:16]
  reg  r_122; // @[Reg.scala 16:16]
  reg  r_123; // @[Reg.scala 16:16]
  reg  r_124; // @[Reg.scala 16:16]
  reg  r_125; // @[Reg.scala 16:16]
  reg  r_126; // @[Reg.scala 16:16]
  reg  r_127; // @[Reg.scala 16:16]
  reg  r_128; // @[Reg.scala 16:16]
  reg  r_129; // @[Reg.scala 16:16]
  reg  r_130; // @[Reg.scala 16:16]
  reg  r_131; // @[Reg.scala 16:16]
  reg  r_132; // @[Reg.scala 16:16]
  reg  r_133; // @[Reg.scala 16:16]
  reg  r_134; // @[Reg.scala 16:16]
  reg  r_135; // @[Reg.scala 16:16]
  reg  r_136; // @[Reg.scala 16:16]
  reg  r_137; // @[Reg.scala 16:16]
  reg  r_138; // @[Reg.scala 16:16]
  reg  r_139; // @[Reg.scala 16:16]
  reg  r_140; // @[Reg.scala 16:16]
  reg  r_141; // @[Reg.scala 16:16]
  reg  r_142; // @[Reg.scala 16:16]
  reg  r_143; // @[Reg.scala 16:16]
  reg  r_144; // @[Reg.scala 16:16]
  reg  r_145; // @[Reg.scala 16:16]
  reg  r_146; // @[Reg.scala 16:16]
  reg  r_147; // @[Reg.scala 16:16]
  reg  r_148; // @[Reg.scala 16:16]
  reg  r_149; // @[Reg.scala 16:16]
  reg  r_150; // @[Reg.scala 16:16]
  reg  r_151; // @[Reg.scala 16:16]
  reg  r_152; // @[Reg.scala 16:16]
  reg  r_153; // @[Reg.scala 16:16]
  reg  r_154; // @[Reg.scala 16:16]
  reg  r_155; // @[Reg.scala 16:16]
  reg  r_156; // @[Reg.scala 16:16]
  reg  r_157; // @[Reg.scala 16:16]
  reg  r_158; // @[Reg.scala 16:16]
  reg  r_159; // @[Reg.scala 16:16]
  reg  r_160; // @[Reg.scala 16:16]
  reg  r_161; // @[Reg.scala 16:16]
  reg  r_162; // @[Reg.scala 16:16]
  reg  r_163; // @[Reg.scala 16:16]
  reg  r_164; // @[Reg.scala 16:16]
  reg  r_165; // @[Reg.scala 16:16]
  reg  r_166; // @[Reg.scala 16:16]
  reg  r_167; // @[Reg.scala 16:16]
  reg  r_168; // @[Reg.scala 16:16]
  reg  r_169; // @[Reg.scala 16:16]
  reg  r_170; // @[Reg.scala 16:16]
  reg  r_171; // @[Reg.scala 16:16]
  reg  r_172; // @[Reg.scala 16:16]
  reg  r_173; // @[Reg.scala 16:16]
  reg  r_174; // @[Reg.scala 16:16]
  reg  r_175; // @[Reg.scala 16:16]
  reg  r_176; // @[Reg.scala 16:16]
  reg  r_177; // @[Reg.scala 16:16]
  reg  r_178; // @[Reg.scala 16:16]
  reg  r_179; // @[Reg.scala 16:16]
  reg  r_180; // @[Reg.scala 16:16]
  reg  r_181; // @[Reg.scala 16:16]
  reg  r_182; // @[Reg.scala 16:16]
  reg  r_183; // @[Reg.scala 16:16]
  reg  r_184; // @[Reg.scala 16:16]
  reg  r_185; // @[Reg.scala 16:16]
  reg  r_186; // @[Reg.scala 16:16]
  reg  r_187; // @[Reg.scala 16:16]
  reg  r_188; // @[Reg.scala 16:16]
  reg  r_189; // @[Reg.scala 16:16]
  reg  r_190; // @[Reg.scala 16:16]
  reg  r_191; // @[Reg.scala 16:16]
  reg  r_192; // @[Reg.scala 16:16]
  reg  r_193; // @[Reg.scala 16:16]
  reg  r_194; // @[Reg.scala 16:16]
  reg  r_195; // @[Reg.scala 16:16]
  reg  r_196; // @[Reg.scala 16:16]
  reg  r_197; // @[Reg.scala 16:16]
  reg  r_198; // @[Reg.scala 16:16]
  reg  r_199; // @[Reg.scala 16:16]
  reg  r_200; // @[Reg.scala 16:16]
  reg  r_201; // @[Reg.scala 16:16]
  reg  r_202; // @[Reg.scala 16:16]
  reg  r_203; // @[Reg.scala 16:16]
  reg  r_204; // @[Reg.scala 16:16]
  reg  r_205; // @[Reg.scala 16:16]
  reg  r_206; // @[Reg.scala 16:16]
  reg  r_207; // @[Reg.scala 16:16]
  reg  r_208; // @[Reg.scala 16:16]
  reg  r_209; // @[Reg.scala 16:16]
  reg  r_210; // @[Reg.scala 16:16]
  reg  r_211; // @[Reg.scala 16:16]
  reg  r_212; // @[Reg.scala 16:16]
  reg  r_213; // @[Reg.scala 16:16]
  reg  r_214; // @[Reg.scala 16:16]
  reg  r_215; // @[Reg.scala 16:16]
  reg  r_216; // @[Reg.scala 16:16]
  reg  r_217; // @[Reg.scala 16:16]
  reg  r_218; // @[Reg.scala 16:16]
  reg  r_219; // @[Reg.scala 16:16]
  reg  r_220; // @[Reg.scala 16:16]
  reg  r_221; // @[Reg.scala 16:16]
  reg  r_222; // @[Reg.scala 16:16]
  reg  r_223; // @[Reg.scala 16:16]
  reg  r_224; // @[Reg.scala 16:16]
  reg  r_225; // @[Reg.scala 16:16]
  reg  r_226; // @[Reg.scala 16:16]
  reg  r_227; // @[Reg.scala 16:16]
  reg  r_228; // @[Reg.scala 16:16]
  reg  r_229; // @[Reg.scala 16:16]
  reg  r_230; // @[Reg.scala 16:16]
  reg  r_231; // @[Reg.scala 16:16]
  reg  r_232; // @[Reg.scala 16:16]
  reg  r_233; // @[Reg.scala 16:16]
  reg  r_234; // @[Reg.scala 16:16]
  reg  r_235; // @[Reg.scala 16:16]
  reg  r_236; // @[Reg.scala 16:16]
  reg  r_237; // @[Reg.scala 16:16]
  reg  r_238; // @[Reg.scala 16:16]
  reg  r_239; // @[Reg.scala 16:16]
  reg  r_240; // @[Reg.scala 16:16]
  reg  r_241; // @[Reg.scala 16:16]
  reg  r_242; // @[Reg.scala 16:16]
  reg  r_243; // @[Reg.scala 16:16]
  reg  r_244; // @[Reg.scala 16:16]
  reg  r_245; // @[Reg.scala 16:16]
  reg  r_246; // @[Reg.scala 16:16]
  reg  r_247; // @[Reg.scala 16:16]
  reg  r_248; // @[Reg.scala 16:16]
  reg  r_249; // @[Reg.scala 16:16]
  reg  r_250; // @[Reg.scala 16:16]
  reg  r_251; // @[Reg.scala 16:16]
  reg  r_252; // @[Reg.scala 16:16]
  reg  r_253; // @[Reg.scala 16:16]
  reg  r_254; // @[Reg.scala 16:16]
  reg  r_255; // @[Reg.scala 16:16]
  reg  r_256; // @[Reg.scala 16:16]
  reg  r_257; // @[Reg.scala 16:16]
  reg  r_258; // @[Reg.scala 16:16]
  reg  r_259; // @[Reg.scala 16:16]
  reg  r_260; // @[Reg.scala 16:16]
  reg  r_261; // @[Reg.scala 16:16]
  reg  r_262; // @[Reg.scala 16:16]
  reg  r_263; // @[Reg.scala 16:16]
  reg  r_264; // @[Reg.scala 16:16]
  reg  r_265; // @[Reg.scala 16:16]
  reg  r_266; // @[Reg.scala 16:16]
  reg  r_267; // @[Reg.scala 16:16]
  reg  r_268; // @[Reg.scala 16:16]
  reg  r_269; // @[Reg.scala 16:16]
  reg  r_270; // @[Reg.scala 16:16]
  reg  r_271; // @[Reg.scala 16:16]
  reg  r_272; // @[Reg.scala 16:16]
  reg  r_273; // @[Reg.scala 16:16]
  reg  r_274; // @[Reg.scala 16:16]
  reg  r_275; // @[Reg.scala 16:16]
  reg  r_276; // @[Reg.scala 16:16]
  reg  r_277; // @[Reg.scala 16:16]
  reg  r_278; // @[Reg.scala 16:16]
  reg  r_279; // @[Reg.scala 16:16]
  reg  r_280; // @[Reg.scala 16:16]
  reg  r_281; // @[Reg.scala 16:16]
  reg  r_282; // @[Reg.scala 16:16]
  reg  r_283; // @[Reg.scala 16:16]
  reg  r_284; // @[Reg.scala 16:16]
  reg  r_285; // @[Reg.scala 16:16]
  reg  r_286; // @[Reg.scala 16:16]
  reg  r_287; // @[Reg.scala 16:16]
  reg  r_288; // @[Reg.scala 16:16]
  reg  r_289; // @[Reg.scala 16:16]
  reg  r_290; // @[Reg.scala 16:16]
  reg  r_291; // @[Reg.scala 16:16]
  reg  r_292; // @[Reg.scala 16:16]
  reg  r_293; // @[Reg.scala 16:16]
  reg  r_294; // @[Reg.scala 16:16]
  reg  r_295; // @[Reg.scala 16:16]
  reg  r_296; // @[Reg.scala 16:16]
  reg  r_297; // @[Reg.scala 16:16]
  reg  r_298; // @[Reg.scala 16:16]
  reg  r_299; // @[Reg.scala 16:16]
  reg  r_300; // @[Reg.scala 16:16]
  reg  r_301; // @[Reg.scala 16:16]
  reg  r_302; // @[Reg.scala 16:16]
  reg  r_303; // @[Reg.scala 16:16]
  reg  r_304; // @[Reg.scala 16:16]
  reg  r_305; // @[Reg.scala 16:16]
  reg  r_306; // @[Reg.scala 16:16]
  reg  r_307; // @[Reg.scala 16:16]
  reg  r_308; // @[Reg.scala 16:16]
  reg  r_309; // @[Reg.scala 16:16]
  reg  r_310; // @[Reg.scala 16:16]
  reg  r_311; // @[Reg.scala 16:16]
  reg  r_312; // @[Reg.scala 16:16]
  reg  r_313; // @[Reg.scala 16:16]
  reg  r_314; // @[Reg.scala 16:16]
  reg  r_315; // @[Reg.scala 16:16]
  reg  r_316; // @[Reg.scala 16:16]
  reg  r_317; // @[Reg.scala 16:16]
  reg  r_318; // @[Reg.scala 16:16]
  reg  r_319; // @[Reg.scala 16:16]
  reg  r_320; // @[Reg.scala 16:16]
  reg  r_321; // @[Reg.scala 16:16]
  reg  r_322; // @[Reg.scala 16:16]
  reg  r_323; // @[Reg.scala 16:16]
  reg  r_324; // @[Reg.scala 16:16]
  reg  r_325; // @[Reg.scala 16:16]
  reg  r_326; // @[Reg.scala 16:16]
  reg  r_327; // @[Reg.scala 16:16]
  reg  r_328; // @[Reg.scala 16:16]
  reg  r_329; // @[Reg.scala 16:16]
  reg  r_330; // @[Reg.scala 16:16]
  reg  r_331; // @[Reg.scala 16:16]
  reg  r_332; // @[Reg.scala 16:16]
  reg  r_333; // @[Reg.scala 16:16]
  reg  r_334; // @[Reg.scala 16:16]
  reg  r_335; // @[Reg.scala 16:16]
  reg  r_336; // @[Reg.scala 16:16]
  reg  r_337; // @[Reg.scala 16:16]
  reg  r_338; // @[Reg.scala 16:16]
  reg  r_339; // @[Reg.scala 16:16]
  reg  r_340; // @[Reg.scala 16:16]
  reg  r_341; // @[Reg.scala 16:16]
  reg  r_342; // @[Reg.scala 16:16]
  reg  r_343; // @[Reg.scala 16:16]
  reg  r_344; // @[Reg.scala 16:16]
  reg  r_345; // @[Reg.scala 16:16]
  reg  r_346; // @[Reg.scala 16:16]
  reg  r_347; // @[Reg.scala 16:16]
  reg  r_348; // @[Reg.scala 16:16]
  reg  r_349; // @[Reg.scala 16:16]
  reg  r_350; // @[Reg.scala 16:16]
  reg  r_351; // @[Reg.scala 16:16]
  reg  r_352; // @[Reg.scala 16:16]
  reg  r_353; // @[Reg.scala 16:16]
  reg  r_354; // @[Reg.scala 16:16]
  reg  r_355; // @[Reg.scala 16:16]
  reg  r_356; // @[Reg.scala 16:16]
  reg  r_357; // @[Reg.scala 16:16]
  reg  r_358; // @[Reg.scala 16:16]
  reg  r_359; // @[Reg.scala 16:16]
  reg  r_360; // @[Reg.scala 16:16]
  reg  r_361; // @[Reg.scala 16:16]
  reg  r_362; // @[Reg.scala 16:16]
  reg  r_363; // @[Reg.scala 16:16]
  reg  r_364; // @[Reg.scala 16:16]
  reg  r_365; // @[Reg.scala 16:16]
  reg  r_366; // @[Reg.scala 16:16]
  reg  r_367; // @[Reg.scala 16:16]
  reg  r_368; // @[Reg.scala 16:16]
  reg  r_369; // @[Reg.scala 16:16]
  reg  r_370; // @[Reg.scala 16:16]
  reg  r_371; // @[Reg.scala 16:16]
  reg  r_372; // @[Reg.scala 16:16]
  reg  r_373; // @[Reg.scala 16:16]
  reg  r_374; // @[Reg.scala 16:16]
  reg  r_375; // @[Reg.scala 16:16]
  reg  r_376; // @[Reg.scala 16:16]
  reg  r_377; // @[Reg.scala 16:16]
  reg  r_378; // @[Reg.scala 16:16]
  reg  r_379; // @[Reg.scala 16:16]
  reg  r_380; // @[Reg.scala 16:16]
  reg  r_381; // @[Reg.scala 16:16]
  reg  r_382; // @[Reg.scala 16:16]
  reg  r_383; // @[Reg.scala 16:16]
  reg  r_384; // @[Reg.scala 16:16]
  reg  r_385; // @[Reg.scala 16:16]
  reg  r_386; // @[Reg.scala 16:16]
  reg  r_387; // @[Reg.scala 16:16]
  reg  r_388; // @[Reg.scala 16:16]
  reg  r_389; // @[Reg.scala 16:16]
  reg  r_390; // @[Reg.scala 16:16]
  reg  r_391; // @[Reg.scala 16:16]
  reg  r_392; // @[Reg.scala 16:16]
  reg  r_393; // @[Reg.scala 16:16]
  reg  r_394; // @[Reg.scala 16:16]
  reg  r_395; // @[Reg.scala 16:16]
  reg  r_396; // @[Reg.scala 16:16]
  reg  r_397; // @[Reg.scala 16:16]
  reg  r_398; // @[Reg.scala 16:16]
  reg  r_399; // @[Reg.scala 16:16]
  reg  r_400; // @[Reg.scala 16:16]
  reg  r_401; // @[Reg.scala 16:16]
  reg  r_402; // @[Reg.scala 16:16]
  reg  r_403; // @[Reg.scala 16:16]
  reg  r_404; // @[Reg.scala 16:16]
  reg  r_405; // @[Reg.scala 16:16]
  reg  r_406; // @[Reg.scala 16:16]
  reg  r_407; // @[Reg.scala 16:16]
  reg  r_408; // @[Reg.scala 16:16]
  reg  r_409; // @[Reg.scala 16:16]
  reg  r_410; // @[Reg.scala 16:16]
  reg  r_411; // @[Reg.scala 16:16]
  reg  r_412; // @[Reg.scala 16:16]
  reg  r_413; // @[Reg.scala 16:16]
  reg  r_414; // @[Reg.scala 16:16]
  reg  r_415; // @[Reg.scala 16:16]
  reg  r_416; // @[Reg.scala 16:16]
  reg  r_417; // @[Reg.scala 16:16]
  reg  r_418; // @[Reg.scala 16:16]
  reg  r_419; // @[Reg.scala 16:16]
  reg  r_420; // @[Reg.scala 16:16]
  reg  r_421; // @[Reg.scala 16:16]
  reg  r_422; // @[Reg.scala 16:16]
  reg  r_423; // @[Reg.scala 16:16]
  reg  r_424; // @[Reg.scala 16:16]
  reg  r_425; // @[Reg.scala 16:16]
  reg  r_426; // @[Reg.scala 16:16]
  reg  r_427; // @[Reg.scala 16:16]
  reg  r_428; // @[Reg.scala 16:16]
  reg  r_429; // @[Reg.scala 16:16]
  reg  r_430; // @[Reg.scala 16:16]
  reg  r_431; // @[Reg.scala 16:16]
  reg  r_432; // @[Reg.scala 16:16]
  reg  r_433; // @[Reg.scala 16:16]
  reg  r_434; // @[Reg.scala 16:16]
  reg  r_435; // @[Reg.scala 16:16]
  reg  r_436; // @[Reg.scala 16:16]
  reg  r_437; // @[Reg.scala 16:16]
  reg  r_438; // @[Reg.scala 16:16]
  reg  r_439; // @[Reg.scala 16:16]
  reg  r_440; // @[Reg.scala 16:16]
  reg  r_441; // @[Reg.scala 16:16]
  reg  r_442; // @[Reg.scala 16:16]
  reg  r_443; // @[Reg.scala 16:16]
  reg  r_444; // @[Reg.scala 16:16]
  reg  r_445; // @[Reg.scala 16:16]
  reg  r_446; // @[Reg.scala 16:16]
  reg  r_447; // @[Reg.scala 16:16]
  reg  r_448; // @[Reg.scala 16:16]
  reg  r_449; // @[Reg.scala 16:16]
  reg  r_450; // @[Reg.scala 16:16]
  reg  r_451; // @[Reg.scala 16:16]
  reg  r_452; // @[Reg.scala 16:16]
  reg  r_453; // @[Reg.scala 16:16]
  reg  r_454; // @[Reg.scala 16:16]
  reg  r_455; // @[Reg.scala 16:16]
  reg  r_456; // @[Reg.scala 16:16]
  reg  r_457; // @[Reg.scala 16:16]
  reg  r_458; // @[Reg.scala 16:16]
  reg  r_459; // @[Reg.scala 16:16]
  reg  r_460; // @[Reg.scala 16:16]
  reg  r_461; // @[Reg.scala 16:16]
  reg  r_462; // @[Reg.scala 16:16]
  reg  r_463; // @[Reg.scala 16:16]
  reg  r_464; // @[Reg.scala 16:16]
  reg  r_465; // @[Reg.scala 16:16]
  reg  r_466; // @[Reg.scala 16:16]
  reg  r_467; // @[Reg.scala 16:16]
  reg  r_468; // @[Reg.scala 16:16]
  reg  r_469; // @[Reg.scala 16:16]
  reg  r_470; // @[Reg.scala 16:16]
  reg  r_471; // @[Reg.scala 16:16]
  reg  r_472; // @[Reg.scala 16:16]
  reg  r_473; // @[Reg.scala 16:16]
  reg  r_474; // @[Reg.scala 16:16]
  reg  r_475; // @[Reg.scala 16:16]
  reg  r_476; // @[Reg.scala 16:16]
  reg  r_477; // @[Reg.scala 16:16]
  reg  r_478; // @[Reg.scala 16:16]
  reg  r_479; // @[Reg.scala 16:16]
  reg  r_480; // @[Reg.scala 16:16]
  reg  r_481; // @[Reg.scala 16:16]
  reg  r_482; // @[Reg.scala 16:16]
  reg  r_483; // @[Reg.scala 16:16]
  reg  r_484; // @[Reg.scala 16:16]
  reg  r_485; // @[Reg.scala 16:16]
  reg  r_486; // @[Reg.scala 16:16]
  reg  r_487; // @[Reg.scala 16:16]
  reg  r_488; // @[Reg.scala 16:16]
  reg  r_489; // @[Reg.scala 16:16]
  reg  r_490; // @[Reg.scala 16:16]
  reg  r_491; // @[Reg.scala 16:16]
  reg  r_492; // @[Reg.scala 16:16]
  reg  r_493; // @[Reg.scala 16:16]
  reg  r_494; // @[Reg.scala 16:16]
  reg  r_495; // @[Reg.scala 16:16]
  reg  r_496; // @[Reg.scala 16:16]
  reg  r_497; // @[Reg.scala 16:16]
  reg  r_498; // @[Reg.scala 16:16]
  reg  r_499; // @[Reg.scala 16:16]
  reg  r_500; // @[Reg.scala 16:16]
  reg  r_501; // @[Reg.scala 16:16]
  reg  r_502; // @[Reg.scala 16:16]
  reg  r_503; // @[Reg.scala 16:16]
  reg  r_504; // @[Reg.scala 16:16]
  reg  r_505; // @[Reg.scala 16:16]
  reg  r_506; // @[Reg.scala 16:16]
  reg  r_507; // @[Reg.scala 16:16]
  reg  r_508; // @[Reg.scala 16:16]
  reg  r_509; // @[Reg.scala 16:16]
  reg  r_510; // @[Reg.scala 16:16]
  reg  r_511; // @[Reg.scala 16:16]
  reg  r_512; // @[Reg.scala 16:16]
  reg  r_513; // @[Reg.scala 16:16]
  reg  r_514; // @[Reg.scala 16:16]
  reg  r_515; // @[Reg.scala 16:16]
  reg  r_516; // @[Reg.scala 16:16]
  reg  r_517; // @[Reg.scala 16:16]
  reg  r_518; // @[Reg.scala 16:16]
  reg  r_519; // @[Reg.scala 16:16]
  reg  r_520; // @[Reg.scala 16:16]
  reg  r_521; // @[Reg.scala 16:16]
  reg  r_522; // @[Reg.scala 16:16]
  reg  r_523; // @[Reg.scala 16:16]
  reg  r_524; // @[Reg.scala 16:16]
  reg  r_525; // @[Reg.scala 16:16]
  reg  r_526; // @[Reg.scala 16:16]
  reg  r_527; // @[Reg.scala 16:16]
  reg  r_528; // @[Reg.scala 16:16]
  reg  r_529; // @[Reg.scala 16:16]
  reg  r_530; // @[Reg.scala 16:16]
  reg  r_531; // @[Reg.scala 16:16]
  reg  r_532; // @[Reg.scala 16:16]
  reg  r_533; // @[Reg.scala 16:16]
  reg  r_534; // @[Reg.scala 16:16]
  reg  r_535; // @[Reg.scala 16:16]
  reg  r_536; // @[Reg.scala 16:16]
  reg  r_537; // @[Reg.scala 16:16]
  reg  r_538; // @[Reg.scala 16:16]
  reg  r_539; // @[Reg.scala 16:16]
  reg  r_540; // @[Reg.scala 16:16]
  reg  r_541; // @[Reg.scala 16:16]
  reg  r_542; // @[Reg.scala 16:16]
  reg  r_543; // @[Reg.scala 16:16]
  reg  r_544; // @[Reg.scala 16:16]
  reg  r_545; // @[Reg.scala 16:16]
  reg  r_546; // @[Reg.scala 16:16]
  reg  r_547; // @[Reg.scala 16:16]
  reg  r_548; // @[Reg.scala 16:16]
  reg  r_549; // @[Reg.scala 16:16]
  reg  r_550; // @[Reg.scala 16:16]
  reg  r_551; // @[Reg.scala 16:16]
  reg  r_552; // @[Reg.scala 16:16]
  reg  r_553; // @[Reg.scala 16:16]
  reg  r_554; // @[Reg.scala 16:16]
  reg  r_555; // @[Reg.scala 16:16]
  reg  r_556; // @[Reg.scala 16:16]
  reg  r_557; // @[Reg.scala 16:16]
  reg  r_558; // @[Reg.scala 16:16]
  reg  r_559; // @[Reg.scala 16:16]
  reg  r_560; // @[Reg.scala 16:16]
  reg  r_561; // @[Reg.scala 16:16]
  reg  r_562; // @[Reg.scala 16:16]
  reg  r_563; // @[Reg.scala 16:16]
  reg  r_564; // @[Reg.scala 16:16]
  reg  r_565; // @[Reg.scala 16:16]
  reg  r_566; // @[Reg.scala 16:16]
  reg  r_567; // @[Reg.scala 16:16]
  reg  r_568; // @[Reg.scala 16:16]
  reg  r_569; // @[Reg.scala 16:16]
  reg  r_570; // @[Reg.scala 16:16]
  reg  r_571; // @[Reg.scala 16:16]
  reg  r_572; // @[Reg.scala 16:16]
  reg  r_573; // @[Reg.scala 16:16]
  reg  r_574; // @[Reg.scala 16:16]
  reg  r_575; // @[Reg.scala 16:16]
  reg  r_576; // @[Reg.scala 16:16]
  reg  r_577; // @[Reg.scala 16:16]
  reg  r_578; // @[Reg.scala 16:16]
  reg  r_579; // @[Reg.scala 16:16]
  reg  r_580; // @[Reg.scala 16:16]
  reg  r_581; // @[Reg.scala 16:16]
  reg  r_582; // @[Reg.scala 16:16]
  reg  r_583; // @[Reg.scala 16:16]
  reg  r_584; // @[Reg.scala 16:16]
  reg  r_585; // @[Reg.scala 16:16]
  reg  r_586; // @[Reg.scala 16:16]
  reg  r_587; // @[Reg.scala 16:16]
  reg  r_588; // @[Reg.scala 16:16]
  reg  r_589; // @[Reg.scala 16:16]
  reg  r_590; // @[Reg.scala 16:16]
  reg  r_591; // @[Reg.scala 16:16]
  reg  r_592; // @[Reg.scala 16:16]
  reg  r_593; // @[Reg.scala 16:16]
  reg  r_594; // @[Reg.scala 16:16]
  reg  r_595; // @[Reg.scala 16:16]
  reg  r_596; // @[Reg.scala 16:16]
  reg  r_597; // @[Reg.scala 16:16]
  reg  r_598; // @[Reg.scala 16:16]
  reg  r_599; // @[Reg.scala 16:16]
  reg  r_600; // @[Reg.scala 16:16]
  reg  r_601; // @[Reg.scala 16:16]
  reg  r_602; // @[Reg.scala 16:16]
  reg  r_603; // @[Reg.scala 16:16]
  reg  r_604; // @[Reg.scala 16:16]
  reg  r_605; // @[Reg.scala 16:16]
  reg  r_606; // @[Reg.scala 16:16]
  reg  r_607; // @[Reg.scala 16:16]
  reg  r_608; // @[Reg.scala 16:16]
  reg  r_609; // @[Reg.scala 16:16]
  reg  r_610; // @[Reg.scala 16:16]
  reg  r_611; // @[Reg.scala 16:16]
  reg  r_612; // @[Reg.scala 16:16]
  reg  r_613; // @[Reg.scala 16:16]
  reg  r_614; // @[Reg.scala 16:16]
  reg  r_615; // @[Reg.scala 16:16]
  reg  r_616; // @[Reg.scala 16:16]
  reg  r_617; // @[Reg.scala 16:16]
  reg  r_618; // @[Reg.scala 16:16]
  reg  r_619; // @[Reg.scala 16:16]
  reg  r_620; // @[Reg.scala 16:16]
  reg  r_621; // @[Reg.scala 16:16]
  reg  r_622; // @[Reg.scala 16:16]
  reg  r_623; // @[Reg.scala 16:16]
  reg  r_624; // @[Reg.scala 16:16]
  reg  r_625; // @[Reg.scala 16:16]
  reg  r_626; // @[Reg.scala 16:16]
  reg  r_627; // @[Reg.scala 16:16]
  reg  r_628; // @[Reg.scala 16:16]
  reg  r_629; // @[Reg.scala 16:16]
  reg  r_630; // @[Reg.scala 16:16]
  reg  r_631; // @[Reg.scala 16:16]
  reg  r_632; // @[Reg.scala 16:16]
  reg  r_633; // @[Reg.scala 16:16]
  reg  r_634; // @[Reg.scala 16:16]
  reg  r_635; // @[Reg.scala 16:16]
  reg  r_636; // @[Reg.scala 16:16]
  reg  r_637; // @[Reg.scala 16:16]
  reg  r_638; // @[Reg.scala 16:16]
  reg  r_639; // @[Reg.scala 16:16]
  reg  r_640; // @[Reg.scala 16:16]
  reg  r_641; // @[Reg.scala 16:16]
  reg  r_642; // @[Reg.scala 16:16]
  reg  r_643; // @[Reg.scala 16:16]
  reg  r_644; // @[Reg.scala 16:16]
  reg  r_645; // @[Reg.scala 16:16]
  reg  r_646; // @[Reg.scala 16:16]
  reg  r_647; // @[Reg.scala 16:16]
  reg  r_648; // @[Reg.scala 16:16]
  reg  r_649; // @[Reg.scala 16:16]
  reg  r_650; // @[Reg.scala 16:16]
  reg  r_651; // @[Reg.scala 16:16]
  reg  r_652; // @[Reg.scala 16:16]
  reg  r_653; // @[Reg.scala 16:16]
  reg  r_654; // @[Reg.scala 16:16]
  reg  r_655; // @[Reg.scala 16:16]
  reg  r_656; // @[Reg.scala 16:16]
  reg  r_657; // @[Reg.scala 16:16]
  reg  r_658; // @[Reg.scala 16:16]
  reg  r_659; // @[Reg.scala 16:16]
  reg  r_660; // @[Reg.scala 16:16]
  reg  r_661; // @[Reg.scala 16:16]
  reg  r_662; // @[Reg.scala 16:16]
  reg  r_663; // @[Reg.scala 16:16]
  reg  r_664; // @[Reg.scala 16:16]
  reg  r_665; // @[Reg.scala 16:16]
  reg  r_666; // @[Reg.scala 16:16]
  reg  r_667; // @[Reg.scala 16:16]
  reg  r_668; // @[Reg.scala 16:16]
  reg  r_669; // @[Reg.scala 16:16]
  reg  r_670; // @[Reg.scala 16:16]
  reg  r_671; // @[Reg.scala 16:16]
  reg  r_672; // @[Reg.scala 16:16]
  reg  r_673; // @[Reg.scala 16:16]
  reg  r_674; // @[Reg.scala 16:16]
  reg  r_675; // @[Reg.scala 16:16]
  reg  r_676; // @[Reg.scala 16:16]
  reg  r_677; // @[Reg.scala 16:16]
  reg  r_678; // @[Reg.scala 16:16]
  reg  r_679; // @[Reg.scala 16:16]
  reg  r_680; // @[Reg.scala 16:16]
  reg  r_681; // @[Reg.scala 16:16]
  reg  r_682; // @[Reg.scala 16:16]
  reg  r_683; // @[Reg.scala 16:16]
  reg  r_684; // @[Reg.scala 16:16]
  reg  r_685; // @[Reg.scala 16:16]
  reg  r_686; // @[Reg.scala 16:16]
  reg  r_687; // @[Reg.scala 16:16]
  reg  r_688; // @[Reg.scala 16:16]
  reg  r_689; // @[Reg.scala 16:16]
  reg  r_690; // @[Reg.scala 16:16]
  reg  r_691; // @[Reg.scala 16:16]
  reg  r_692; // @[Reg.scala 16:16]
  reg  r_693; // @[Reg.scala 16:16]
  reg  r_694; // @[Reg.scala 16:16]
  reg  r_695; // @[Reg.scala 16:16]
  reg  r_696; // @[Reg.scala 16:16]
  reg  r_697; // @[Reg.scala 16:16]
  reg  r_698; // @[Reg.scala 16:16]
  reg  r_699; // @[Reg.scala 16:16]
  reg  r_700; // @[Reg.scala 16:16]
  reg  r_701; // @[Reg.scala 16:16]
  reg  r_702; // @[Reg.scala 16:16]
  reg  r_703; // @[Reg.scala 16:16]
  reg  r_704; // @[Reg.scala 16:16]
  reg  r_705; // @[Reg.scala 16:16]
  reg  r_706; // @[Reg.scala 16:16]
  reg  r_707; // @[Reg.scala 16:16]
  reg  r_708; // @[Reg.scala 16:16]
  reg  r_709; // @[Reg.scala 16:16]
  reg  r_710; // @[Reg.scala 16:16]
  reg  r_711; // @[Reg.scala 16:16]
  reg  r_712; // @[Reg.scala 16:16]
  reg  r_713; // @[Reg.scala 16:16]
  reg  r_714; // @[Reg.scala 16:16]
  reg  r_715; // @[Reg.scala 16:16]
  reg  r_716; // @[Reg.scala 16:16]
  reg  r_717; // @[Reg.scala 16:16]
  reg  r_718; // @[Reg.scala 16:16]
  reg  r_719; // @[Reg.scala 16:16]
  reg  r_720; // @[Reg.scala 16:16]
  reg  r_721; // @[Reg.scala 16:16]
  reg  r_722; // @[Reg.scala 16:16]
  reg  r_723; // @[Reg.scala 16:16]
  reg  r_724; // @[Reg.scala 16:16]
  reg  r_725; // @[Reg.scala 16:16]
  reg  r_726; // @[Reg.scala 16:16]
  reg  r_727; // @[Reg.scala 16:16]
  reg  r_728; // @[Reg.scala 16:16]
  reg  r_729; // @[Reg.scala 16:16]
  reg  r_730; // @[Reg.scala 16:16]
  reg  r_731; // @[Reg.scala 16:16]
  reg  r_732; // @[Reg.scala 16:16]
  reg  r_733; // @[Reg.scala 16:16]
  reg  r_734; // @[Reg.scala 16:16]
  reg  r_735; // @[Reg.scala 16:16]
  reg  r_736; // @[Reg.scala 16:16]
  reg  r_737; // @[Reg.scala 16:16]
  reg  r_738; // @[Reg.scala 16:16]
  reg  r_739; // @[Reg.scala 16:16]
  reg  r_740; // @[Reg.scala 16:16]
  reg  r_741; // @[Reg.scala 16:16]
  reg  r_742; // @[Reg.scala 16:16]
  reg  r_743; // @[Reg.scala 16:16]
  reg  r_744; // @[Reg.scala 16:16]
  reg  r_745; // @[Reg.scala 16:16]
  reg  r_746; // @[Reg.scala 16:16]
  reg  r_747; // @[Reg.scala 16:16]
  reg  r_748; // @[Reg.scala 16:16]
  reg  r_749; // @[Reg.scala 16:16]
  reg  r_750; // @[Reg.scala 16:16]
  reg  r_751; // @[Reg.scala 16:16]
  reg  r_752; // @[Reg.scala 16:16]
  reg  r_753; // @[Reg.scala 16:16]
  reg  r_754; // @[Reg.scala 16:16]
  reg  r_755; // @[Reg.scala 16:16]
  reg  r_756; // @[Reg.scala 16:16]
  reg  r_757; // @[Reg.scala 16:16]
  reg  r_758; // @[Reg.scala 16:16]
  reg  r_759; // @[Reg.scala 16:16]
  reg  r_760; // @[Reg.scala 16:16]
  reg  r_761; // @[Reg.scala 16:16]
  reg  r_762; // @[Reg.scala 16:16]
  reg  r_763; // @[Reg.scala 16:16]
  reg  r_764; // @[Reg.scala 16:16]
  reg  r_765; // @[Reg.scala 16:16]
  reg  r_766; // @[Reg.scala 16:16]
  reg  r_767; // @[Reg.scala 16:16]
  reg  r_768; // @[Reg.scala 16:16]
  reg  r_769; // @[Reg.scala 16:16]
  reg  r_770; // @[Reg.scala 16:16]
  reg  r_771; // @[Reg.scala 16:16]
  reg  r_772; // @[Reg.scala 16:16]
  reg  r_773; // @[Reg.scala 16:16]
  reg  r_774; // @[Reg.scala 16:16]
  reg  r_775; // @[Reg.scala 16:16]
  reg  r_776; // @[Reg.scala 16:16]
  reg  r_777; // @[Reg.scala 16:16]
  reg  r_778; // @[Reg.scala 16:16]
  reg  r_779; // @[Reg.scala 16:16]
  reg  r_780; // @[Reg.scala 16:16]
  reg  r_781; // @[Reg.scala 16:16]
  reg  r_782; // @[Reg.scala 16:16]
  reg  r_783; // @[Reg.scala 16:16]
  reg  r_784; // @[Reg.scala 16:16]
  reg  r_785; // @[Reg.scala 16:16]
  reg  r_786; // @[Reg.scala 16:16]
  reg  r_787; // @[Reg.scala 16:16]
  reg  r_788; // @[Reg.scala 16:16]
  reg  r_789; // @[Reg.scala 16:16]
  reg  r_790; // @[Reg.scala 16:16]
  reg  r_791; // @[Reg.scala 16:16]
  reg  r_792; // @[Reg.scala 16:16]
  reg  r_793; // @[Reg.scala 16:16]
  reg  r_794; // @[Reg.scala 16:16]
  reg  r_795; // @[Reg.scala 16:16]
  reg  r_796; // @[Reg.scala 16:16]
  reg  r_797; // @[Reg.scala 16:16]
  reg  r_798; // @[Reg.scala 16:16]
  reg  r_799; // @[Reg.scala 16:16]
  reg  r_800; // @[Reg.scala 16:16]
  reg  r_801; // @[Reg.scala 16:16]
  reg  r_802; // @[Reg.scala 16:16]
  reg  r_803; // @[Reg.scala 16:16]
  reg  r_804; // @[Reg.scala 16:16]
  reg  r_805; // @[Reg.scala 16:16]
  reg  r_806; // @[Reg.scala 16:16]
  reg  r_807; // @[Reg.scala 16:16]
  reg  r_808; // @[Reg.scala 16:16]
  reg  r_809; // @[Reg.scala 16:16]
  reg  r_810; // @[Reg.scala 16:16]
  reg  r_811; // @[Reg.scala 16:16]
  reg  r_812; // @[Reg.scala 16:16]
  reg  r_813; // @[Reg.scala 16:16]
  reg  r_814; // @[Reg.scala 16:16]
  reg  r_815; // @[Reg.scala 16:16]
  reg  r_816; // @[Reg.scala 16:16]
  reg  r_817; // @[Reg.scala 16:16]
  reg  r_818; // @[Reg.scala 16:16]
  reg  r_819; // @[Reg.scala 16:16]
  reg  r_820; // @[Reg.scala 16:16]
  reg  r_821; // @[Reg.scala 16:16]
  reg  r_822; // @[Reg.scala 16:16]
  reg  r_823; // @[Reg.scala 16:16]
  reg  r_824; // @[Reg.scala 16:16]
  reg  r_825; // @[Reg.scala 16:16]
  reg  r_826; // @[Reg.scala 16:16]
  reg  r_827; // @[Reg.scala 16:16]
  reg  r_828; // @[Reg.scala 16:16]
  reg  r_829; // @[Reg.scala 16:16]
  reg  r_830; // @[Reg.scala 16:16]
  reg  r_831; // @[Reg.scala 16:16]
  reg  r_832; // @[Reg.scala 16:16]
  reg  r_833; // @[Reg.scala 16:16]
  reg  r_834; // @[Reg.scala 16:16]
  reg  r_835; // @[Reg.scala 16:16]
  reg  r_836; // @[Reg.scala 16:16]
  reg  r_837; // @[Reg.scala 16:16]
  reg  r_838; // @[Reg.scala 16:16]
  reg  r_839; // @[Reg.scala 16:16]
  reg  r_840; // @[Reg.scala 16:16]
  reg  r_841; // @[Reg.scala 16:16]
  reg  r_842; // @[Reg.scala 16:16]
  reg  r_843; // @[Reg.scala 16:16]
  reg  r_844; // @[Reg.scala 16:16]
  reg  r_845; // @[Reg.scala 16:16]
  reg  r_846; // @[Reg.scala 16:16]
  reg  r_847; // @[Reg.scala 16:16]
  reg  r_848; // @[Reg.scala 16:16]
  reg  r_849; // @[Reg.scala 16:16]
  reg  r_850; // @[Reg.scala 16:16]
  reg  r_851; // @[Reg.scala 16:16]
  reg  r_852; // @[Reg.scala 16:16]
  reg  r_853; // @[Reg.scala 16:16]
  reg  r_854; // @[Reg.scala 16:16]
  reg  r_855; // @[Reg.scala 16:16]
  reg  r_856; // @[Reg.scala 16:16]
  reg  r_857; // @[Reg.scala 16:16]
  reg  r_858; // @[Reg.scala 16:16]
  reg  r_859; // @[Reg.scala 16:16]
  reg  r_860; // @[Reg.scala 16:16]
  reg  r_861; // @[Reg.scala 16:16]
  reg  r_862; // @[Reg.scala 16:16]
  reg  r_863; // @[Reg.scala 16:16]
  reg  r_864; // @[Reg.scala 16:16]
  reg  r_865; // @[Reg.scala 16:16]
  reg  r_866; // @[Reg.scala 16:16]
  reg  r_867; // @[Reg.scala 16:16]
  reg  r_868; // @[Reg.scala 16:16]
  reg  r_869; // @[Reg.scala 16:16]
  reg  r_870; // @[Reg.scala 16:16]
  reg  r_871; // @[Reg.scala 16:16]
  reg  r_872; // @[Reg.scala 16:16]
  reg  r_873; // @[Reg.scala 16:16]
  reg  r_874; // @[Reg.scala 16:16]
  reg  r_875; // @[Reg.scala 16:16]
  reg  r_876; // @[Reg.scala 16:16]
  reg  r_877; // @[Reg.scala 16:16]
  reg  r_878; // @[Reg.scala 16:16]
  reg  r_879; // @[Reg.scala 16:16]
  reg  r_880; // @[Reg.scala 16:16]
  reg  r_881; // @[Reg.scala 16:16]
  reg  r_882; // @[Reg.scala 16:16]
  reg  r_883; // @[Reg.scala 16:16]
  reg  r_884; // @[Reg.scala 16:16]
  reg  r_885; // @[Reg.scala 16:16]
  reg  r_886; // @[Reg.scala 16:16]
  reg  r_887; // @[Reg.scala 16:16]
  reg  r_888; // @[Reg.scala 16:16]
  reg  r_889; // @[Reg.scala 16:16]
  reg  r_890; // @[Reg.scala 16:16]
  reg  r_891; // @[Reg.scala 16:16]
  reg  r_892; // @[Reg.scala 16:16]
  reg  r_893; // @[Reg.scala 16:16]
  reg  r_894; // @[Reg.scala 16:16]
  reg  r_895; // @[Reg.scala 16:16]
  reg  r_896; // @[Reg.scala 16:16]
  reg  r_897; // @[Reg.scala 16:16]
  reg  r_898; // @[Reg.scala 16:16]
  reg  r_899; // @[Reg.scala 16:16]
  reg  r_900; // @[Reg.scala 16:16]
  reg  r_901; // @[Reg.scala 16:16]
  reg  r_902; // @[Reg.scala 16:16]
  reg  r_903; // @[Reg.scala 16:16]
  reg  r_904; // @[Reg.scala 16:16]
  reg  r_905; // @[Reg.scala 16:16]
  reg  r_906; // @[Reg.scala 16:16]
  reg  r_907; // @[Reg.scala 16:16]
  reg  r_908; // @[Reg.scala 16:16]
  reg  r_909; // @[Reg.scala 16:16]
  reg  r_910; // @[Reg.scala 16:16]
  reg  r_911; // @[Reg.scala 16:16]
  reg  r_912; // @[Reg.scala 16:16]
  reg  r_913; // @[Reg.scala 16:16]
  reg  r_914; // @[Reg.scala 16:16]
  reg  r_915; // @[Reg.scala 16:16]
  reg  r_916; // @[Reg.scala 16:16]
  reg  r_917; // @[Reg.scala 16:16]
  reg  r_918; // @[Reg.scala 16:16]
  reg  r_919; // @[Reg.scala 16:16]
  reg  r_920; // @[Reg.scala 16:16]
  reg  r_921; // @[Reg.scala 16:16]
  reg  r_922; // @[Reg.scala 16:16]
  reg  r_923; // @[Reg.scala 16:16]
  reg  r_924; // @[Reg.scala 16:16]
  reg  r_925; // @[Reg.scala 16:16]
  reg  r_926; // @[Reg.scala 16:16]
  reg  r_927; // @[Reg.scala 16:16]
  reg  r_928; // @[Reg.scala 16:16]
  reg  r_929; // @[Reg.scala 16:16]
  reg  r_930; // @[Reg.scala 16:16]
  reg  r_931; // @[Reg.scala 16:16]
  reg  r_932; // @[Reg.scala 16:16]
  reg  r_933; // @[Reg.scala 16:16]
  reg  r_934; // @[Reg.scala 16:16]
  reg  r_935; // @[Reg.scala 16:16]
  reg  r_936; // @[Reg.scala 16:16]
  reg  r_937; // @[Reg.scala 16:16]
  reg  r_938; // @[Reg.scala 16:16]
  reg  r_939; // @[Reg.scala 16:16]
  reg  r_940; // @[Reg.scala 16:16]
  reg  r_941; // @[Reg.scala 16:16]
  reg  r_942; // @[Reg.scala 16:16]
  reg  r_943; // @[Reg.scala 16:16]
  reg  r_944; // @[Reg.scala 16:16]
  reg  r_945; // @[Reg.scala 16:16]
  reg  r_946; // @[Reg.scala 16:16]
  reg  r_947; // @[Reg.scala 16:16]
  reg  r_948; // @[Reg.scala 16:16]
  reg  r_949; // @[Reg.scala 16:16]
  reg  r_950; // @[Reg.scala 16:16]
  reg  r_951; // @[Reg.scala 16:16]
  reg  r_952; // @[Reg.scala 16:16]
  reg  r_953; // @[Reg.scala 16:16]
  reg  r_954; // @[Reg.scala 16:16]
  reg  r_955; // @[Reg.scala 16:16]
  reg  r_956; // @[Reg.scala 16:16]
  reg  r_957; // @[Reg.scala 16:16]
  reg  r_958; // @[Reg.scala 16:16]
  reg  r_959; // @[Reg.scala 16:16]
  reg  r_960; // @[Reg.scala 16:16]
  reg  r_961; // @[Reg.scala 16:16]
  reg  r_962; // @[Reg.scala 16:16]
  reg  r_963; // @[Reg.scala 16:16]
  reg  r_964; // @[Reg.scala 16:16]
  reg  r_965; // @[Reg.scala 16:16]
  reg  r_966; // @[Reg.scala 16:16]
  reg  r_967; // @[Reg.scala 16:16]
  reg  r_968; // @[Reg.scala 16:16]
  reg  r_969; // @[Reg.scala 16:16]
  reg  r_970; // @[Reg.scala 16:16]
  reg  r_971; // @[Reg.scala 16:16]
  reg  r_972; // @[Reg.scala 16:16]
  reg  r_973; // @[Reg.scala 16:16]
  reg  r_974; // @[Reg.scala 16:16]
  reg  r_975; // @[Reg.scala 16:16]
  reg  r_976; // @[Reg.scala 16:16]
  reg  r_977; // @[Reg.scala 16:16]
  reg  r_978; // @[Reg.scala 16:16]
  reg  r_979; // @[Reg.scala 16:16]
  reg  r_980; // @[Reg.scala 16:16]
  reg  r_981; // @[Reg.scala 16:16]
  reg  r_982; // @[Reg.scala 16:16]
  reg  r_983; // @[Reg.scala 16:16]
  reg  r_984; // @[Reg.scala 16:16]
  reg  r_985; // @[Reg.scala 16:16]
  reg  r_986; // @[Reg.scala 16:16]
  reg  r_987; // @[Reg.scala 16:16]
  reg  r_988; // @[Reg.scala 16:16]
  reg  r_989; // @[Reg.scala 16:16]
  reg  r_990; // @[Reg.scala 16:16]
  reg  r_991; // @[Reg.scala 16:16]
  reg  r_992; // @[Reg.scala 16:16]
  reg  r_993; // @[Reg.scala 16:16]
  reg  r_994; // @[Reg.scala 16:16]
  reg  r_995; // @[Reg.scala 16:16]
  reg  r_996; // @[Reg.scala 16:16]
  reg  r_997; // @[Reg.scala 16:16]
  reg  r_998; // @[Reg.scala 16:16]
  reg  r_999; // @[Reg.scala 16:16]
  reg  r_1000; // @[Reg.scala 16:16]
  reg  r_1001; // @[Reg.scala 16:16]
  reg  r_1002; // @[Reg.scala 16:16]
  reg  r_1003; // @[Reg.scala 16:16]
  reg  r_1004; // @[Reg.scala 16:16]
  reg  r_1005; // @[Reg.scala 16:16]
  reg  r_1006; // @[Reg.scala 16:16]
  reg  r_1007; // @[Reg.scala 16:16]
  reg  r_1008; // @[Reg.scala 16:16]
  reg  r_1009; // @[Reg.scala 16:16]
  reg  r_1010; // @[Reg.scala 16:16]
  reg  r_1011; // @[Reg.scala 16:16]
  reg  r_1012; // @[Reg.scala 16:16]
  reg  r_1013; // @[Reg.scala 16:16]
  reg  r_1014; // @[Reg.scala 16:16]
  reg  r_1015; // @[Reg.scala 16:16]
  reg  r_1016; // @[Reg.scala 16:16]
  reg  r_1017; // @[Reg.scala 16:16]
  reg  r_1018; // @[Reg.scala 16:16]
  reg  r_1019; // @[Reg.scala 16:16]
  reg  r_1020; // @[Reg.scala 16:16]
  reg  r_1021; // @[Reg.scala 16:16]
  reg  r_1022; // @[Reg.scala 16:16]
  reg  r_1023; // @[Reg.scala 16:16]
  reg  r_1024; // @[Reg.scala 16:16]
  reg  r_1025; // @[Reg.scala 16:16]
  reg  r_1026; // @[Reg.scala 16:16]
  reg  r_1027; // @[Reg.scala 16:16]
  reg  r_1028; // @[Reg.scala 16:16]
  reg  r_1029; // @[Reg.scala 16:16]
  reg  r_1030; // @[Reg.scala 16:16]
  reg  r_1031; // @[Reg.scala 16:16]
  reg  r_1032; // @[Reg.scala 16:16]
  reg  r_1033; // @[Reg.scala 16:16]
  reg  r_1034; // @[Reg.scala 16:16]
  reg  r_1035; // @[Reg.scala 16:16]
  reg  r_1036; // @[Reg.scala 16:16]
  reg  r_1037; // @[Reg.scala 16:16]
  reg  r_1038; // @[Reg.scala 16:16]
  reg  r_1039; // @[Reg.scala 16:16]
  reg  r_1040; // @[Reg.scala 16:16]
  reg  r_1041; // @[Reg.scala 16:16]
  reg  r_1042; // @[Reg.scala 16:16]
  reg  r_1043; // @[Reg.scala 16:16]
  reg  r_1044; // @[Reg.scala 16:16]
  reg  r_1045; // @[Reg.scala 16:16]
  reg  r_1046; // @[Reg.scala 16:16]
  reg  r_1047; // @[Reg.scala 16:16]
  reg  r_1048; // @[Reg.scala 16:16]
  reg  r_1049; // @[Reg.scala 16:16]
  reg  r_1050; // @[Reg.scala 16:16]
  reg  r_1051; // @[Reg.scala 16:16]
  reg  r_1052; // @[Reg.scala 16:16]
  reg  r_1053; // @[Reg.scala 16:16]
  reg  r_1054; // @[Reg.scala 16:16]
  reg  r_1055; // @[Reg.scala 16:16]
  reg  r_1056; // @[Reg.scala 16:16]
  reg  r_1057; // @[Reg.scala 16:16]
  reg  r_1058; // @[Reg.scala 16:16]
  reg  r_1059; // @[Reg.scala 16:16]
  reg  r_1060; // @[Reg.scala 16:16]
  reg  r_1061; // @[Reg.scala 16:16]
  reg  r_1062; // @[Reg.scala 16:16]
  reg  r_1063; // @[Reg.scala 16:16]
  reg  r_1064; // @[Reg.scala 16:16]
  reg  r_1065; // @[Reg.scala 16:16]
  reg  r_1066; // @[Reg.scala 16:16]
  reg  r_1067; // @[Reg.scala 16:16]
  reg  r_1068; // @[Reg.scala 16:16]
  reg  r_1069; // @[Reg.scala 16:16]
  reg  r_1070; // @[Reg.scala 16:16]
  reg  r_1071; // @[Reg.scala 16:16]
  reg  r_1072; // @[Reg.scala 16:16]
  reg  r_1073; // @[Reg.scala 16:16]
  reg  r_1074; // @[Reg.scala 16:16]
  reg  r_1075; // @[Reg.scala 16:16]
  reg  r_1076; // @[Reg.scala 16:16]
  reg  r_1077; // @[Reg.scala 16:16]
  reg  r_1078; // @[Reg.scala 16:16]
  reg  r_1079; // @[Reg.scala 16:16]
  reg  r_1080; // @[Reg.scala 16:16]
  reg  r_1081; // @[Reg.scala 16:16]
  reg  r_1082; // @[Reg.scala 16:16]
  reg  r_1083; // @[Reg.scala 16:16]
  reg  r_1084; // @[Reg.scala 16:16]
  reg  r_1085; // @[Reg.scala 16:16]
  reg  r_1086; // @[Reg.scala 16:16]
  reg  r_1087; // @[Reg.scala 16:16]
  reg  r_1088; // @[Reg.scala 16:16]
  reg  r_1089; // @[Reg.scala 16:16]
  reg  r_1090; // @[Reg.scala 16:16]
  reg  r_1091; // @[Reg.scala 16:16]
  reg  r_1092; // @[Reg.scala 16:16]
  reg  r_1093; // @[Reg.scala 16:16]
  reg  r_1094; // @[Reg.scala 16:16]
  reg  r_1095; // @[Reg.scala 16:16]
  reg  r_1096; // @[Reg.scala 16:16]
  reg  r_1097; // @[Reg.scala 16:16]
  reg  r_1098; // @[Reg.scala 16:16]
  reg  r_1099; // @[Reg.scala 16:16]
  reg  r_1100; // @[Reg.scala 16:16]
  reg  r_1101; // @[Reg.scala 16:16]
  reg  r_1102; // @[Reg.scala 16:16]
  reg  r_1103; // @[Reg.scala 16:16]
  reg  r_1104; // @[Reg.scala 16:16]
  reg  r_1105; // @[Reg.scala 16:16]
  reg  r_1106; // @[Reg.scala 16:16]
  reg  r_1107; // @[Reg.scala 16:16]
  reg  r_1108; // @[Reg.scala 16:16]
  reg  r_1109; // @[Reg.scala 16:16]
  reg  r_1110; // @[Reg.scala 16:16]
  reg  r_1111; // @[Reg.scala 16:16]
  reg  r_1112; // @[Reg.scala 16:16]
  reg  r_1113; // @[Reg.scala 16:16]
  reg  r_1114; // @[Reg.scala 16:16]
  reg  r_1115; // @[Reg.scala 16:16]
  reg  r_1116; // @[Reg.scala 16:16]
  reg  r_1117; // @[Reg.scala 16:16]
  reg  r_1118; // @[Reg.scala 16:16]
  reg  r_1119; // @[Reg.scala 16:16]
  reg  r_1120; // @[Reg.scala 16:16]
  reg  r_1121; // @[Reg.scala 16:16]
  reg  r_1122; // @[Reg.scala 16:16]
  reg  r_1123; // @[Reg.scala 16:16]
  reg  r_1124; // @[Reg.scala 16:16]
  reg  r_1125; // @[Reg.scala 16:16]
  reg  r_1126; // @[Reg.scala 16:16]
  reg  r_1127; // @[Reg.scala 16:16]
  reg  r_1128; // @[Reg.scala 16:16]
  reg  r_1129; // @[Reg.scala 16:16]
  reg  r_1130; // @[Reg.scala 16:16]
  reg  r_1131; // @[Reg.scala 16:16]
  reg  r_1132; // @[Reg.scala 16:16]
  reg  r_1133; // @[Reg.scala 16:16]
  reg  r_1134; // @[Reg.scala 16:16]
  reg  r_1135; // @[Reg.scala 16:16]
  reg  r_1136; // @[Reg.scala 16:16]
  reg  r_1137; // @[Reg.scala 16:16]
  reg  r_1138; // @[Reg.scala 16:16]
  reg  r_1139; // @[Reg.scala 16:16]
  reg  r_1140; // @[Reg.scala 16:16]
  reg  r_1141; // @[Reg.scala 16:16]
  reg  r_1142; // @[Reg.scala 16:16]
  reg  r_1143; // @[Reg.scala 16:16]
  reg  r_1144; // @[Reg.scala 16:16]
  reg  r_1145; // @[Reg.scala 16:16]
  reg  r_1146; // @[Reg.scala 16:16]
  reg  r_1147; // @[Reg.scala 16:16]
  reg  r_1148; // @[Reg.scala 16:16]
  reg  r_1149; // @[Reg.scala 16:16]
  reg  r_1150; // @[Reg.scala 16:16]
  reg  r_1151; // @[Reg.scala 16:16]
  reg  r_1152; // @[Reg.scala 16:16]
  reg  r_1153; // @[Reg.scala 16:16]
  reg  r_1154; // @[Reg.scala 16:16]
  reg  r_1155; // @[Reg.scala 16:16]
  reg  r_1156; // @[Reg.scala 16:16]
  reg  r_1157; // @[Reg.scala 16:16]
  reg  r_1158; // @[Reg.scala 16:16]
  reg  r_1159; // @[Reg.scala 16:16]
  reg  r_1160; // @[Reg.scala 16:16]
  reg  r_1161; // @[Reg.scala 16:16]
  reg  r_1162; // @[Reg.scala 16:16]
  reg  r_1163; // @[Reg.scala 16:16]
  reg  r_1164; // @[Reg.scala 16:16]
  reg  r_1165; // @[Reg.scala 16:16]
  reg  r_1166; // @[Reg.scala 16:16]
  reg  r_1167; // @[Reg.scala 16:16]
  reg  r_1168; // @[Reg.scala 16:16]
  reg  r_1169; // @[Reg.scala 16:16]
  reg  r_1170; // @[Reg.scala 16:16]
  reg  r_1171; // @[Reg.scala 16:16]
  reg  r_1172; // @[Reg.scala 16:16]
  reg  r_1173; // @[Reg.scala 16:16]
  reg  r_1174; // @[Reg.scala 16:16]
  reg  r_1175; // @[Reg.scala 16:16]
  reg  r_1176; // @[Reg.scala 16:16]
  reg  r_1177; // @[Reg.scala 16:16]
  reg  r_1178; // @[Reg.scala 16:16]
  reg  r_1179; // @[Reg.scala 16:16]
  reg  r_1180; // @[Reg.scala 16:16]
  reg  r_1181; // @[Reg.scala 16:16]
  reg  r_1182; // @[Reg.scala 16:16]
  reg  r_1183; // @[Reg.scala 16:16]
  reg  r_1184; // @[Reg.scala 16:16]
  reg  r_1185; // @[Reg.scala 16:16]
  reg  r_1186; // @[Reg.scala 16:16]
  reg  r_1187; // @[Reg.scala 16:16]
  reg  r_1188; // @[Reg.scala 16:16]
  reg  r_1189; // @[Reg.scala 16:16]
  reg  r_1190; // @[Reg.scala 16:16]
  reg  r_1191; // @[Reg.scala 16:16]
  reg  r_1192; // @[Reg.scala 16:16]
  reg  r_1193; // @[Reg.scala 16:16]
  reg  r_1194; // @[Reg.scala 16:16]
  reg  r_1195; // @[Reg.scala 16:16]
  reg  r_1196; // @[Reg.scala 16:16]
  reg  r_1197; // @[Reg.scala 16:16]
  reg  r_1198; // @[Reg.scala 16:16]
  reg  r_1199; // @[Reg.scala 16:16]
  reg  r_1200; // @[Reg.scala 16:16]
  reg  r_1201; // @[Reg.scala 16:16]
  reg  r_1202; // @[Reg.scala 16:16]
  reg  r_1203; // @[Reg.scala 16:16]
  reg  r_1204; // @[Reg.scala 16:16]
  reg  r_1205; // @[Reg.scala 16:16]
  reg  r_1206; // @[Reg.scala 16:16]
  reg  r_1207; // @[Reg.scala 16:16]
  reg  r_1208; // @[Reg.scala 16:16]
  reg  r_1209; // @[Reg.scala 16:16]
  reg  r_1210; // @[Reg.scala 16:16]
  reg  r_1211; // @[Reg.scala 16:16]
  reg  r_1212; // @[Reg.scala 16:16]
  reg  r_1213; // @[Reg.scala 16:16]
  reg  r_1214; // @[Reg.scala 16:16]
  reg  r_1215; // @[Reg.scala 16:16]
  reg  r_1216; // @[Reg.scala 16:16]
  reg  r_1217; // @[Reg.scala 16:16]
  reg  r_1218; // @[Reg.scala 16:16]
  reg  r_1219; // @[Reg.scala 16:16]
  reg  r_1220; // @[Reg.scala 16:16]
  reg  r_1221; // @[Reg.scala 16:16]
  reg  r_1222; // @[Reg.scala 16:16]
  reg  r_1223; // @[Reg.scala 16:16]
  reg  r_1224; // @[Reg.scala 16:16]
  reg  r_1225; // @[Reg.scala 16:16]
  reg  r_1226; // @[Reg.scala 16:16]
  reg  r_1227; // @[Reg.scala 16:16]
  reg  r_1228; // @[Reg.scala 16:16]
  reg  r_1229; // @[Reg.scala 16:16]
  reg  r_1230; // @[Reg.scala 16:16]
  reg  r_1231; // @[Reg.scala 16:16]
  reg  r_1232; // @[Reg.scala 16:16]
  reg  r_1233; // @[Reg.scala 16:16]
  reg  r_1234; // @[Reg.scala 16:16]
  reg  r_1235; // @[Reg.scala 16:16]
  reg  r_1236; // @[Reg.scala 16:16]
  reg  r_1237; // @[Reg.scala 16:16]
  reg  r_1238; // @[Reg.scala 16:16]
  reg  r_1239; // @[Reg.scala 16:16]
  reg  r_1240; // @[Reg.scala 16:16]
  reg  r_1241; // @[Reg.scala 16:16]
  reg  r_1242; // @[Reg.scala 16:16]
  reg  r_1243; // @[Reg.scala 16:16]
  reg  r_1244; // @[Reg.scala 16:16]
  reg  r_1245; // @[Reg.scala 16:16]
  reg  r_1246; // @[Reg.scala 16:16]
  reg  r_1247; // @[Reg.scala 16:16]
  reg  r_1248; // @[Reg.scala 16:16]
  reg  r_1249; // @[Reg.scala 16:16]
  reg  r_1250; // @[Reg.scala 16:16]
  reg  r_1251; // @[Reg.scala 16:16]
  reg  r_1252; // @[Reg.scala 16:16]
  reg  r_1253; // @[Reg.scala 16:16]
  reg  r_1254; // @[Reg.scala 16:16]
  reg  r_1255; // @[Reg.scala 16:16]
  reg  r_1256; // @[Reg.scala 16:16]
  reg  r_1257; // @[Reg.scala 16:16]
  reg  r_1258; // @[Reg.scala 16:16]
  reg  r_1259; // @[Reg.scala 16:16]
  reg  r_1260; // @[Reg.scala 16:16]
  reg  r_1261; // @[Reg.scala 16:16]
  reg  r_1262; // @[Reg.scala 16:16]
  reg  r_1263; // @[Reg.scala 16:16]
  reg  r_1264; // @[Reg.scala 16:16]
  reg  r_1265; // @[Reg.scala 16:16]
  reg  r_1266; // @[Reg.scala 16:16]
  reg  r_1267; // @[Reg.scala 16:16]
  reg  r_1268; // @[Reg.scala 16:16]
  reg  r_1269; // @[Reg.scala 16:16]
  reg  r_1270; // @[Reg.scala 16:16]
  reg  r_1271; // @[Reg.scala 16:16]
  reg  r_1272; // @[Reg.scala 16:16]
  reg  r_1273; // @[Reg.scala 16:16]
  reg  r_1274; // @[Reg.scala 16:16]
  reg  r_1275; // @[Reg.scala 16:16]
  reg  r_1276; // @[Reg.scala 16:16]
  reg  r_1277; // @[Reg.scala 16:16]
  reg  r_1278; // @[Reg.scala 16:16]
  reg  r_1279; // @[Reg.scala 16:16]
  reg  r_1280; // @[Reg.scala 16:16]
  reg  r_1281; // @[Reg.scala 16:16]
  reg  r_1282; // @[Reg.scala 16:16]
  reg  r_1283; // @[Reg.scala 16:16]
  reg  r_1284; // @[Reg.scala 16:16]
  reg  r_1285; // @[Reg.scala 16:16]
  reg  r_1286; // @[Reg.scala 16:16]
  reg  r_1287; // @[Reg.scala 16:16]
  reg  r_1288; // @[Reg.scala 16:16]
  reg  r_1289; // @[Reg.scala 16:16]
  reg  r_1290; // @[Reg.scala 16:16]
  reg  r_1291; // @[Reg.scala 16:16]
  reg  r_1292; // @[Reg.scala 16:16]
  reg  r_1293; // @[Reg.scala 16:16]
  reg  r_1294; // @[Reg.scala 16:16]
  reg  r_1295; // @[Reg.scala 16:16]
  reg  r_1296; // @[Reg.scala 16:16]
  reg  r_1297; // @[Reg.scala 16:16]
  reg  r_1298; // @[Reg.scala 16:16]
  reg  r_1299; // @[Reg.scala 16:16]
  reg  r_1300; // @[Reg.scala 16:16]
  reg  r_1301; // @[Reg.scala 16:16]
  reg  r_1302; // @[Reg.scala 16:16]
  reg  r_1303; // @[Reg.scala 16:16]
  reg  r_1304; // @[Reg.scala 16:16]
  reg  r_1305; // @[Reg.scala 16:16]
  reg  r_1306; // @[Reg.scala 16:16]
  reg  r_1307; // @[Reg.scala 16:16]
  reg  r_1308; // @[Reg.scala 16:16]
  reg  r_1309; // @[Reg.scala 16:16]
  reg  r_1310; // @[Reg.scala 16:16]
  reg  r_1311; // @[Reg.scala 16:16]
  reg  r_1312; // @[Reg.scala 16:16]
  reg  r_1313; // @[Reg.scala 16:16]
  reg  r_1314; // @[Reg.scala 16:16]
  reg  r_1315; // @[Reg.scala 16:16]
  reg  r_1316; // @[Reg.scala 16:16]
  reg  r_1317; // @[Reg.scala 16:16]
  reg  r_1318; // @[Reg.scala 16:16]
  reg  r_1319; // @[Reg.scala 16:16]
  reg  r_1320; // @[Reg.scala 16:16]
  reg  r_1321; // @[Reg.scala 16:16]
  reg  r_1322; // @[Reg.scala 16:16]
  reg  r_1323; // @[Reg.scala 16:16]
  reg  r_1324; // @[Reg.scala 16:16]
  reg  r_1325; // @[Reg.scala 16:16]
  reg  r_1326; // @[Reg.scala 16:16]
  reg  r_1327; // @[Reg.scala 16:16]
  reg  r_1328; // @[Reg.scala 16:16]
  reg  r_1329; // @[Reg.scala 16:16]
  reg  r_1330; // @[Reg.scala 16:16]
  reg  r_1331; // @[Reg.scala 16:16]
  reg  r_1332; // @[Reg.scala 16:16]
  reg  r_1333; // @[Reg.scala 16:16]
  reg  r_1334; // @[Reg.scala 16:16]
  reg  r_1335; // @[Reg.scala 16:16]
  reg  r_1336; // @[Reg.scala 16:16]
  reg  r_1337; // @[Reg.scala 16:16]
  reg  r_1338; // @[Reg.scala 16:16]
  reg  r_1339; // @[Reg.scala 16:16]
  reg  r_1340; // @[Reg.scala 16:16]
  reg  r_1341; // @[Reg.scala 16:16]
  reg  r_1342; // @[Reg.scala 16:16]
  reg  r_1343; // @[Reg.scala 16:16]
  reg  r_1344; // @[Reg.scala 16:16]
  reg  r_1345; // @[Reg.scala 16:16]
  reg  r_1346; // @[Reg.scala 16:16]
  reg  r_1347; // @[Reg.scala 16:16]
  reg  r_1348; // @[Reg.scala 16:16]
  reg  r_1349; // @[Reg.scala 16:16]
  reg  r_1350; // @[Reg.scala 16:16]
  reg  r_1351; // @[Reg.scala 16:16]
  reg  r_1352; // @[Reg.scala 16:16]
  reg  r_1353; // @[Reg.scala 16:16]
  reg  r_1354; // @[Reg.scala 16:16]
  reg  r_1355; // @[Reg.scala 16:16]
  reg  r_1356; // @[Reg.scala 16:16]
  reg  r_1357; // @[Reg.scala 16:16]
  reg  r_1358; // @[Reg.scala 16:16]
  reg  r_1359; // @[Reg.scala 16:16]
  reg  r_1360; // @[Reg.scala 16:16]
  reg  r_1361; // @[Reg.scala 16:16]
  reg  r_1362; // @[Reg.scala 16:16]
  reg  r_1363; // @[Reg.scala 16:16]
  reg  r_1364; // @[Reg.scala 16:16]
  reg  r_1365; // @[Reg.scala 16:16]
  reg  r_1366; // @[Reg.scala 16:16]
  reg  r_1367; // @[Reg.scala 16:16]
  reg  r_1368; // @[Reg.scala 16:16]
  reg  r_1369; // @[Reg.scala 16:16]
  reg  r_1370; // @[Reg.scala 16:16]
  reg  r_1371; // @[Reg.scala 16:16]
  reg  r_1372; // @[Reg.scala 16:16]
  reg  r_1373; // @[Reg.scala 16:16]
  reg  r_1374; // @[Reg.scala 16:16]
  reg  r_1375; // @[Reg.scala 16:16]
  reg  r_1376; // @[Reg.scala 16:16]
  reg  r_1377; // @[Reg.scala 16:16]
  reg  r_1378; // @[Reg.scala 16:16]
  reg  r_1379; // @[Reg.scala 16:16]
  reg  r_1380; // @[Reg.scala 16:16]
  reg  r_1381; // @[Reg.scala 16:16]
  reg  r_1382; // @[Reg.scala 16:16]
  reg  r_1383; // @[Reg.scala 16:16]
  reg  r_1384; // @[Reg.scala 16:16]
  reg  r_1385; // @[Reg.scala 16:16]
  reg  r_1386; // @[Reg.scala 16:16]
  reg  r_1387; // @[Reg.scala 16:16]
  reg  r_1388; // @[Reg.scala 16:16]
  reg  r_1389; // @[Reg.scala 16:16]
  reg  r_1390; // @[Reg.scala 16:16]
  reg  r_1391; // @[Reg.scala 16:16]
  reg  r_1392; // @[Reg.scala 16:16]
  reg  r_1393; // @[Reg.scala 16:16]
  reg  r_1394; // @[Reg.scala 16:16]
  reg  r_1395; // @[Reg.scala 16:16]
  reg  r_1396; // @[Reg.scala 16:16]
  reg  r_1397; // @[Reg.scala 16:16]
  reg  r_1398; // @[Reg.scala 16:16]
  reg  r_1399; // @[Reg.scala 16:16]
  reg  r_1400; // @[Reg.scala 16:16]
  reg  r_1401; // @[Reg.scala 16:16]
  reg  r_1402; // @[Reg.scala 16:16]
  reg  r_1403; // @[Reg.scala 16:16]
  reg  r_1404; // @[Reg.scala 16:16]
  reg  r_1405; // @[Reg.scala 16:16]
  reg  r_1406; // @[Reg.scala 16:16]
  reg  r_1407; // @[Reg.scala 16:16]
  reg  r_1408; // @[Reg.scala 16:16]
  reg  r_1409; // @[Reg.scala 16:16]
  reg  r_1410; // @[Reg.scala 16:16]
  reg  r_1411; // @[Reg.scala 16:16]
  reg  r_1412; // @[Reg.scala 16:16]
  reg  r_1413; // @[Reg.scala 16:16]
  reg  r_1414; // @[Reg.scala 16:16]
  reg  r_1415; // @[Reg.scala 16:16]
  reg  r_1416; // @[Reg.scala 16:16]
  reg  r_1417; // @[Reg.scala 16:16]
  reg  r_1418; // @[Reg.scala 16:16]
  reg  r_1419; // @[Reg.scala 16:16]
  reg  r_1420; // @[Reg.scala 16:16]
  reg  r_1421; // @[Reg.scala 16:16]
  reg  r_1422; // @[Reg.scala 16:16]
  reg  r_1423; // @[Reg.scala 16:16]
  reg  r_1424; // @[Reg.scala 16:16]
  reg  r_1425; // @[Reg.scala 16:16]
  reg  r_1426; // @[Reg.scala 16:16]
  reg  r_1427; // @[Reg.scala 16:16]
  reg  r_1428; // @[Reg.scala 16:16]
  reg  r_1429; // @[Reg.scala 16:16]
  reg  r_1430; // @[Reg.scala 16:16]
  reg  r_1431; // @[Reg.scala 16:16]
  reg  r_1432; // @[Reg.scala 16:16]
  reg  r_1433; // @[Reg.scala 16:16]
  reg  r_1434; // @[Reg.scala 16:16]
  reg  r_1435; // @[Reg.scala 16:16]
  reg  r_1436; // @[Reg.scala 16:16]
  reg  r_1437; // @[Reg.scala 16:16]
  reg  r_1438; // @[Reg.scala 16:16]
  reg  r_1439; // @[Reg.scala 16:16]
  reg  r_1440; // @[Reg.scala 16:16]
  reg  r_1441; // @[Reg.scala 16:16]
  reg  r_1442; // @[Reg.scala 16:16]
  reg  r_1443; // @[Reg.scala 16:16]
  reg  r_1444; // @[Reg.scala 16:16]
  reg  r_1445; // @[Reg.scala 16:16]
  reg  r_1446; // @[Reg.scala 16:16]
  reg  r_1447; // @[Reg.scala 16:16]
  reg  r_1448; // @[Reg.scala 16:16]
  reg  r_1449; // @[Reg.scala 16:16]
  reg  r_1450; // @[Reg.scala 16:16]
  reg  r_1451; // @[Reg.scala 16:16]
  reg  r_1452; // @[Reg.scala 16:16]
  reg  r_1453; // @[Reg.scala 16:16]
  reg  r_1454; // @[Reg.scala 16:16]
  reg  r_1455; // @[Reg.scala 16:16]
  reg  r_1456; // @[Reg.scala 16:16]
  reg  r_1457; // @[Reg.scala 16:16]
  reg  r_1458; // @[Reg.scala 16:16]
  reg  r_1459; // @[Reg.scala 16:16]
  reg  r_1460; // @[Reg.scala 16:16]
  reg  r_1461; // @[Reg.scala 16:16]
  reg  r_1462; // @[Reg.scala 16:16]
  reg  r_1463; // @[Reg.scala 16:16]
  reg  r_1464; // @[Reg.scala 16:16]
  reg  r_1465; // @[Reg.scala 16:16]
  reg  r_1466; // @[Reg.scala 16:16]
  reg  r_1467; // @[Reg.scala 16:16]
  reg  r_1468; // @[Reg.scala 16:16]
  reg  r_1469; // @[Reg.scala 16:16]
  reg  r_1470; // @[Reg.scala 16:16]
  reg  r_1471; // @[Reg.scala 16:16]
  reg  r_1472; // @[Reg.scala 16:16]
  reg  r_1473; // @[Reg.scala 16:16]
  reg  r_1474; // @[Reg.scala 16:16]
  reg  r_1475; // @[Reg.scala 16:16]
  reg  r_1476; // @[Reg.scala 16:16]
  reg  r_1477; // @[Reg.scala 16:16]
  reg  r_1478; // @[Reg.scala 16:16]
  reg  r_1479; // @[Reg.scala 16:16]
  reg  r_1480; // @[Reg.scala 16:16]
  reg  r_1481; // @[Reg.scala 16:16]
  reg  r_1482; // @[Reg.scala 16:16]
  reg  r_1483; // @[Reg.scala 16:16]
  reg  r_1484; // @[Reg.scala 16:16]
  reg  r_1485; // @[Reg.scala 16:16]
  reg  r_1486; // @[Reg.scala 16:16]
  reg  r_1487; // @[Reg.scala 16:16]
  reg  r_1488; // @[Reg.scala 16:16]
  reg  r_1489; // @[Reg.scala 16:16]
  reg  r_1490; // @[Reg.scala 16:16]
  reg  r_1491; // @[Reg.scala 16:16]
  reg  r_1492; // @[Reg.scala 16:16]
  reg  r_1493; // @[Reg.scala 16:16]
  reg  r_1494; // @[Reg.scala 16:16]
  reg  r_1495; // @[Reg.scala 16:16]
  reg  r_1496; // @[Reg.scala 16:16]
  reg  r_1497; // @[Reg.scala 16:16]
  reg  r_1498; // @[Reg.scala 16:16]
  reg  r_1499; // @[Reg.scala 16:16]
  reg  r_1500; // @[Reg.scala 16:16]
  reg  r_1501; // @[Reg.scala 16:16]
  reg  r_1502; // @[Reg.scala 16:16]
  reg  r_1503; // @[Reg.scala 16:16]
  reg  r_1504; // @[Reg.scala 16:16]
  reg  r_1505; // @[Reg.scala 16:16]
  reg  r_1506; // @[Reg.scala 16:16]
  reg  r_1507; // @[Reg.scala 16:16]
  reg  r_1508; // @[Reg.scala 16:16]
  reg  r_1509; // @[Reg.scala 16:16]
  reg  r_1510; // @[Reg.scala 16:16]
  reg  r_1511; // @[Reg.scala 16:16]
  reg  r_1512; // @[Reg.scala 16:16]
  reg  r_1513; // @[Reg.scala 16:16]
  reg  r_1514; // @[Reg.scala 16:16]
  reg  r_1515; // @[Reg.scala 16:16]
  reg  r_1516; // @[Reg.scala 16:16]
  reg  r_1517; // @[Reg.scala 16:16]
  reg  r_1518; // @[Reg.scala 16:16]
  reg  r_1519; // @[Reg.scala 16:16]
  reg  r_1520; // @[Reg.scala 16:16]
  reg  r_1521; // @[Reg.scala 16:16]
  reg  r_1522; // @[Reg.scala 16:16]
  reg  r_1523; // @[Reg.scala 16:16]
  reg  r_1524; // @[Reg.scala 16:16]
  reg  r_1525; // @[Reg.scala 16:16]
  reg  r_1526; // @[Reg.scala 16:16]
  reg  r_1527; // @[Reg.scala 16:16]
  reg  r_1528; // @[Reg.scala 16:16]
  reg  r_1529; // @[Reg.scala 16:16]
  reg  r_1530; // @[Reg.scala 16:16]
  reg  r_1531; // @[Reg.scala 16:16]
  reg  r_1532; // @[Reg.scala 16:16]
  reg  r_1533; // @[Reg.scala 16:16]
  reg  r_1534; // @[Reg.scala 16:16]
  reg  r_1535; // @[Reg.scala 16:16]
  reg  r_1536; // @[Reg.scala 16:16]
  reg  r_1537; // @[Reg.scala 16:16]
  reg  r_1538; // @[Reg.scala 16:16]
  reg  r_1539; // @[Reg.scala 16:16]
  reg  r_1540; // @[Reg.scala 16:16]
  reg  r_1541; // @[Reg.scala 16:16]
  reg  r_1542; // @[Reg.scala 16:16]
  reg  r_1543; // @[Reg.scala 16:16]
  reg  r_1544; // @[Reg.scala 16:16]
  reg  r_1545; // @[Reg.scala 16:16]
  reg  r_1546; // @[Reg.scala 16:16]
  reg  r_1547; // @[Reg.scala 16:16]
  reg  r_1548; // @[Reg.scala 16:16]
  reg  r_1549; // @[Reg.scala 16:16]
  reg  r_1550; // @[Reg.scala 16:16]
  reg  r_1551; // @[Reg.scala 16:16]
  reg  r_1552; // @[Reg.scala 16:16]
  reg  r_1553; // @[Reg.scala 16:16]
  reg  r_1554; // @[Reg.scala 16:16]
  reg  r_1555; // @[Reg.scala 16:16]
  reg  r_1556; // @[Reg.scala 16:16]
  reg  r_1557; // @[Reg.scala 16:16]
  reg  r_1558; // @[Reg.scala 16:16]
  reg  r_1559; // @[Reg.scala 16:16]
  reg  r_1560; // @[Reg.scala 16:16]
  reg  r_1561; // @[Reg.scala 16:16]
  reg  r_1562; // @[Reg.scala 16:16]
  reg  r_1563; // @[Reg.scala 16:16]
  reg  r_1564; // @[Reg.scala 16:16]
  reg  r_1565; // @[Reg.scala 16:16]
  reg  r_1566; // @[Reg.scala 16:16]
  reg  r_1567; // @[Reg.scala 16:16]
  reg  r_1568; // @[Reg.scala 16:16]
  reg  r_1569; // @[Reg.scala 16:16]
  reg  r_1570; // @[Reg.scala 16:16]
  reg  r_1571; // @[Reg.scala 16:16]
  reg  r_1572; // @[Reg.scala 16:16]
  reg  r_1573; // @[Reg.scala 16:16]
  reg  r_1574; // @[Reg.scala 16:16]
  reg  r_1575; // @[Reg.scala 16:16]
  reg  r_1576; // @[Reg.scala 16:16]
  reg  r_1577; // @[Reg.scala 16:16]
  reg  r_1578; // @[Reg.scala 16:16]
  reg  r_1579; // @[Reg.scala 16:16]
  reg  r_1580; // @[Reg.scala 16:16]
  reg  r_1581; // @[Reg.scala 16:16]
  reg  r_1582; // @[Reg.scala 16:16]
  reg  r_1583; // @[Reg.scala 16:16]
  reg  r_1584; // @[Reg.scala 16:16]
  reg  r_1585; // @[Reg.scala 16:16]
  reg  r_1586; // @[Reg.scala 16:16]
  reg  r_1587; // @[Reg.scala 16:16]
  reg  r_1588; // @[Reg.scala 16:16]
  reg  r_1589; // @[Reg.scala 16:16]
  reg  r_1590; // @[Reg.scala 16:16]
  reg  r_1591; // @[Reg.scala 16:16]
  reg  r_1592; // @[Reg.scala 16:16]
  reg  r_1593; // @[Reg.scala 16:16]
  reg  r_1594; // @[Reg.scala 16:16]
  reg  r_1595; // @[Reg.scala 16:16]
  reg  r_1596; // @[Reg.scala 16:16]
  reg  r_1597; // @[Reg.scala 16:16]
  reg  r_1598; // @[Reg.scala 16:16]
  reg  r_1599; // @[Reg.scala 16:16]
  reg  r_1600; // @[Reg.scala 16:16]
  reg  r_1601; // @[Reg.scala 16:16]
  reg  r_1602; // @[Reg.scala 16:16]
  reg  r_1603; // @[Reg.scala 16:16]
  reg  r_1604; // @[Reg.scala 16:16]
  reg  r_1605; // @[Reg.scala 16:16]
  reg  r_1606; // @[Reg.scala 16:16]
  reg  r_1607; // @[Reg.scala 16:16]
  reg  r_1608; // @[Reg.scala 16:16]
  reg  r_1609; // @[Reg.scala 16:16]
  reg  r_1610; // @[Reg.scala 16:16]
  reg  r_1611; // @[Reg.scala 16:16]
  reg  r_1612; // @[Reg.scala 16:16]
  reg  r_1613; // @[Reg.scala 16:16]
  reg  r_1614; // @[Reg.scala 16:16]
  reg  r_1615; // @[Reg.scala 16:16]
  reg  r_1616; // @[Reg.scala 16:16]
  reg  r_1617; // @[Reg.scala 16:16]
  reg  r_1618; // @[Reg.scala 16:16]
  reg  r_1619; // @[Reg.scala 16:16]
  reg  r_1620; // @[Reg.scala 16:16]
  reg  r_1621; // @[Reg.scala 16:16]
  reg  r_1622; // @[Reg.scala 16:16]
  reg  r_1623; // @[Reg.scala 16:16]
  reg  r_1624; // @[Reg.scala 16:16]
  reg  r_1625; // @[Reg.scala 16:16]
  reg  r_1626; // @[Reg.scala 16:16]
  reg  r_1627; // @[Reg.scala 16:16]
  reg  r_1628; // @[Reg.scala 16:16]
  reg  r_1629; // @[Reg.scala 16:16]
  reg  r_1630; // @[Reg.scala 16:16]
  reg  r_1631; // @[Reg.scala 16:16]
  reg  r_1632; // @[Reg.scala 16:16]
  reg  r_1633; // @[Reg.scala 16:16]
  reg  r_1634; // @[Reg.scala 16:16]
  reg  r_1635; // @[Reg.scala 16:16]
  reg  r_1636; // @[Reg.scala 16:16]
  reg  r_1637; // @[Reg.scala 16:16]
  reg  r_1638; // @[Reg.scala 16:16]
  reg  r_1639; // @[Reg.scala 16:16]
  reg  r_1640; // @[Reg.scala 16:16]
  reg  r_1641; // @[Reg.scala 16:16]
  reg  r_1642; // @[Reg.scala 16:16]
  reg  r_1643; // @[Reg.scala 16:16]
  reg  r_1644; // @[Reg.scala 16:16]
  reg  r_1645; // @[Reg.scala 16:16]
  reg  r_1646; // @[Reg.scala 16:16]
  reg  r_1647; // @[Reg.scala 16:16]
  reg  r_1648; // @[Reg.scala 16:16]
  reg  r_1649; // @[Reg.scala 16:16]
  reg  r_1650; // @[Reg.scala 16:16]
  reg  r_1651; // @[Reg.scala 16:16]
  reg  r_1652; // @[Reg.scala 16:16]
  reg  r_1653; // @[Reg.scala 16:16]
  reg  r_1654; // @[Reg.scala 16:16]
  reg  r_1655; // @[Reg.scala 16:16]
  reg  r_1656; // @[Reg.scala 16:16]
  reg  r_1657; // @[Reg.scala 16:16]
  reg  r_1658; // @[Reg.scala 16:16]
  reg  r_1659; // @[Reg.scala 16:16]
  reg  r_1660; // @[Reg.scala 16:16]
  reg  r_1661; // @[Reg.scala 16:16]
  reg  r_1662; // @[Reg.scala 16:16]
  reg  r_1663; // @[Reg.scala 16:16]
  reg  r_1664; // @[Reg.scala 16:16]
  reg  r_1665; // @[Reg.scala 16:16]
  reg  r_1666; // @[Reg.scala 16:16]
  reg  r_1667; // @[Reg.scala 16:16]
  reg  r_1668; // @[Reg.scala 16:16]
  reg  r_1669; // @[Reg.scala 16:16]
  reg  r_1670; // @[Reg.scala 16:16]
  reg  r_1671; // @[Reg.scala 16:16]
  reg  r_1672; // @[Reg.scala 16:16]
  reg  r_1673; // @[Reg.scala 16:16]
  reg  r_1674; // @[Reg.scala 16:16]
  reg  r_1675; // @[Reg.scala 16:16]
  reg  r_1676; // @[Reg.scala 16:16]
  reg  r_1677; // @[Reg.scala 16:16]
  reg  r_1678; // @[Reg.scala 16:16]
  reg  r_1679; // @[Reg.scala 16:16]
  reg  r_1680; // @[Reg.scala 16:16]
  reg  r_1681; // @[Reg.scala 16:16]
  reg  r_1682; // @[Reg.scala 16:16]
  reg  r_1683; // @[Reg.scala 16:16]
  reg  r_1684; // @[Reg.scala 16:16]
  reg  r_1685; // @[Reg.scala 16:16]
  reg  r_1686; // @[Reg.scala 16:16]
  reg  r_1687; // @[Reg.scala 16:16]
  reg  r_1688; // @[Reg.scala 16:16]
  reg  r_1689; // @[Reg.scala 16:16]
  reg  r_1690; // @[Reg.scala 16:16]
  reg  r_1691; // @[Reg.scala 16:16]
  reg  r_1692; // @[Reg.scala 16:16]
  reg  r_1693; // @[Reg.scala 16:16]
  reg  r_1694; // @[Reg.scala 16:16]
  reg  r_1695; // @[Reg.scala 16:16]
  reg  r_1696; // @[Reg.scala 16:16]
  reg  r_1697; // @[Reg.scala 16:16]
  reg  r_1698; // @[Reg.scala 16:16]
  reg  r_1699; // @[Reg.scala 16:16]
  reg  r_1700; // @[Reg.scala 16:16]
  reg  r_1701; // @[Reg.scala 16:16]
  reg  r_1702; // @[Reg.scala 16:16]
  reg  r_1703; // @[Reg.scala 16:16]
  reg  r_1704; // @[Reg.scala 16:16]
  reg  r_1705; // @[Reg.scala 16:16]
  reg  r_1706; // @[Reg.scala 16:16]
  reg  r_1707; // @[Reg.scala 16:16]
  reg  r_1708; // @[Reg.scala 16:16]
  reg  r_1709; // @[Reg.scala 16:16]
  reg  r_1710; // @[Reg.scala 16:16]
  reg  r_1711; // @[Reg.scala 16:16]
  reg  r_1712; // @[Reg.scala 16:16]
  reg  r_1713; // @[Reg.scala 16:16]
  reg  r_1714; // @[Reg.scala 16:16]
  reg  r_1715; // @[Reg.scala 16:16]
  reg  r_1716; // @[Reg.scala 16:16]
  reg  r_1717; // @[Reg.scala 16:16]
  reg  r_1718; // @[Reg.scala 16:16]
  reg  r_1719; // @[Reg.scala 16:16]
  reg  r_1720; // @[Reg.scala 16:16]
  reg  r_1721; // @[Reg.scala 16:16]
  reg  r_1722; // @[Reg.scala 16:16]
  reg  r_1723; // @[Reg.scala 16:16]
  reg  r_1724; // @[Reg.scala 16:16]
  reg  r_1725; // @[Reg.scala 16:16]
  reg  r_1726; // @[Reg.scala 16:16]
  reg  r_1727; // @[Reg.scala 16:16]
  reg  r_1728; // @[Reg.scala 16:16]
  reg  r_1729; // @[Reg.scala 16:16]
  reg  r_1730; // @[Reg.scala 16:16]
  reg  r_1731; // @[Reg.scala 16:16]
  reg  r_1732; // @[Reg.scala 16:16]
  reg  r_1733; // @[Reg.scala 16:16]
  reg  r_1734; // @[Reg.scala 16:16]
  reg  r_1735; // @[Reg.scala 16:16]
  reg  r_1736; // @[Reg.scala 16:16]
  reg  r_1737; // @[Reg.scala 16:16]
  reg  r_1738; // @[Reg.scala 16:16]
  reg  r_1739; // @[Reg.scala 16:16]
  reg  r_1740; // @[Reg.scala 16:16]
  reg  r_1741; // @[Reg.scala 16:16]
  reg  r_1742; // @[Reg.scala 16:16]
  reg  r_1743; // @[Reg.scala 16:16]
  reg  r_1744; // @[Reg.scala 16:16]
  reg  r_1745; // @[Reg.scala 16:16]
  reg  r_1746; // @[Reg.scala 16:16]
  reg  r_1747; // @[Reg.scala 16:16]
  reg  r_1748; // @[Reg.scala 16:16]
  reg  r_1749; // @[Reg.scala 16:16]
  reg  r_1750; // @[Reg.scala 16:16]
  reg  r_1751; // @[Reg.scala 16:16]
  reg  r_1752; // @[Reg.scala 16:16]
  reg  r_1753; // @[Reg.scala 16:16]
  reg  r_1754; // @[Reg.scala 16:16]
  reg  r_1755; // @[Reg.scala 16:16]
  reg  r_1756; // @[Reg.scala 16:16]
  reg  r_1757; // @[Reg.scala 16:16]
  reg  r_1758; // @[Reg.scala 16:16]
  reg  r_1759; // @[Reg.scala 16:16]
  reg  r_1760; // @[Reg.scala 16:16]
  reg  r_1761; // @[Reg.scala 16:16]
  reg  r_1762; // @[Reg.scala 16:16]
  reg  r_1763; // @[Reg.scala 16:16]
  reg  r_1764; // @[Reg.scala 16:16]
  reg  r_1765; // @[Reg.scala 16:16]
  reg  r_1766; // @[Reg.scala 16:16]
  reg  r_1767; // @[Reg.scala 16:16]
  reg  r_1768; // @[Reg.scala 16:16]
  reg  r_1769; // @[Reg.scala 16:16]
  reg  r_1770; // @[Reg.scala 16:16]
  reg  r_1771; // @[Reg.scala 16:16]
  reg  r_1772; // @[Reg.scala 16:16]
  reg  r_1773; // @[Reg.scala 16:16]
  reg  r_1774; // @[Reg.scala 16:16]
  reg  r_1775; // @[Reg.scala 16:16]
  reg  r_1776; // @[Reg.scala 16:16]
  reg  r_1777; // @[Reg.scala 16:16]
  reg  r_1778; // @[Reg.scala 16:16]
  reg  r_1779; // @[Reg.scala 16:16]
  reg  r_1780; // @[Reg.scala 16:16]
  reg  r_1781; // @[Reg.scala 16:16]
  reg  r_1782; // @[Reg.scala 16:16]
  reg  r_1783; // @[Reg.scala 16:16]
  reg  r_1784; // @[Reg.scala 16:16]
  reg  r_1785; // @[Reg.scala 16:16]
  reg  r_1786; // @[Reg.scala 16:16]
  reg  r_1787; // @[Reg.scala 16:16]
  reg  r_1788; // @[Reg.scala 16:16]
  reg  r_1789; // @[Reg.scala 16:16]
  reg  r_1790; // @[Reg.scala 16:16]
  reg  r_1791; // @[Reg.scala 16:16]
  reg  r_1792; // @[Reg.scala 16:16]
  reg  r_1793; // @[Reg.scala 16:16]
  reg  r_1794; // @[Reg.scala 16:16]
  reg  r_1795; // @[Reg.scala 16:16]
  reg  r_1796; // @[Reg.scala 16:16]
  reg  r_1797; // @[Reg.scala 16:16]
  reg  r_1798; // @[Reg.scala 16:16]
  reg  r_1799; // @[Reg.scala 16:16]
  reg  r_1800; // @[Reg.scala 16:16]
  reg  r_1801; // @[Reg.scala 16:16]
  reg  r_1802; // @[Reg.scala 16:16]
  reg  r_1803; // @[Reg.scala 16:16]
  reg  r_1804; // @[Reg.scala 16:16]
  reg  r_1805; // @[Reg.scala 16:16]
  reg  r_1806; // @[Reg.scala 16:16]
  reg  r_1807; // @[Reg.scala 16:16]
  reg  r_1808; // @[Reg.scala 16:16]
  reg  r_1809; // @[Reg.scala 16:16]
  reg  r_1810; // @[Reg.scala 16:16]
  reg  r_1811; // @[Reg.scala 16:16]
  reg  r_1812; // @[Reg.scala 16:16]
  reg  r_1813; // @[Reg.scala 16:16]
  reg  r_1814; // @[Reg.scala 16:16]
  reg  r_1815; // @[Reg.scala 16:16]
  reg  r_1816; // @[Reg.scala 16:16]
  reg  r_1817; // @[Reg.scala 16:16]
  reg  r_1818; // @[Reg.scala 16:16]
  reg  r_1819; // @[Reg.scala 16:16]
  reg  r_1820; // @[Reg.scala 16:16]
  reg  r_1821; // @[Reg.scala 16:16]
  reg  r_1822; // @[Reg.scala 16:16]
  reg  r_1823; // @[Reg.scala 16:16]
  reg  r_1824; // @[Reg.scala 16:16]
  reg  r_1825; // @[Reg.scala 16:16]
  reg  r_1826; // @[Reg.scala 16:16]
  reg  r_1827; // @[Reg.scala 16:16]
  reg  r_1828; // @[Reg.scala 16:16]
  reg  r_1829; // @[Reg.scala 16:16]
  reg  r_1830; // @[Reg.scala 16:16]
  reg  r_1831; // @[Reg.scala 16:16]
  reg  r_1832; // @[Reg.scala 16:16]
  reg  r_1833; // @[Reg.scala 16:16]
  reg  r_1834; // @[Reg.scala 16:16]
  reg  r_1835; // @[Reg.scala 16:16]
  reg  r_1836; // @[Reg.scala 16:16]
  reg  r_1837; // @[Reg.scala 16:16]
  reg  r_1838; // @[Reg.scala 16:16]
  reg  r_1839; // @[Reg.scala 16:16]
  reg  r_1840; // @[Reg.scala 16:16]
  reg  r_1841; // @[Reg.scala 16:16]
  reg  r_1842; // @[Reg.scala 16:16]
  reg  r_1843; // @[Reg.scala 16:16]
  reg  r_1844; // @[Reg.scala 16:16]
  reg  r_1845; // @[Reg.scala 16:16]
  reg  r_1846; // @[Reg.scala 16:16]
  reg  r_1847; // @[Reg.scala 16:16]
  reg  r_1848; // @[Reg.scala 16:16]
  reg  r_1849; // @[Reg.scala 16:16]
  reg  r_1850; // @[Reg.scala 16:16]
  reg  r_1851; // @[Reg.scala 16:16]
  reg  r_1852; // @[Reg.scala 16:16]
  reg  r_1853; // @[Reg.scala 16:16]
  reg  r_1854; // @[Reg.scala 16:16]
  reg  r_1855; // @[Reg.scala 16:16]
  reg  r_1856; // @[Reg.scala 16:16]
  reg  r_1857; // @[Reg.scala 16:16]
  reg  r_1858; // @[Reg.scala 16:16]
  reg  r_1859; // @[Reg.scala 16:16]
  reg  r_1860; // @[Reg.scala 16:16]
  reg  r_1861; // @[Reg.scala 16:16]
  reg  r_1862; // @[Reg.scala 16:16]
  reg  r_1863; // @[Reg.scala 16:16]
  reg  r_1864; // @[Reg.scala 16:16]
  reg  r_1865; // @[Reg.scala 16:16]
  reg  r_1866; // @[Reg.scala 16:16]
  reg  r_1867; // @[Reg.scala 16:16]
  reg  r_1868; // @[Reg.scala 16:16]
  reg  r_1869; // @[Reg.scala 16:16]
  reg  r_1870; // @[Reg.scala 16:16]
  reg  r_1871; // @[Reg.scala 16:16]
  reg  r_1872; // @[Reg.scala 16:16]
  reg  r_1873; // @[Reg.scala 16:16]
  reg  r_1874; // @[Reg.scala 16:16]
  reg  r_1875; // @[Reg.scala 16:16]
  reg  r_1876; // @[Reg.scala 16:16]
  reg  r_1877; // @[Reg.scala 16:16]
  reg  r_1878; // @[Reg.scala 16:16]
  reg  r_1879; // @[Reg.scala 16:16]
  reg  r_1880; // @[Reg.scala 16:16]
  reg  r_1881; // @[Reg.scala 16:16]
  reg  r_1882; // @[Reg.scala 16:16]
  reg  r_1883; // @[Reg.scala 16:16]
  reg  r_1884; // @[Reg.scala 16:16]
  reg  r_1885; // @[Reg.scala 16:16]
  reg  r_1886; // @[Reg.scala 16:16]
  reg  r_1887; // @[Reg.scala 16:16]
  reg  r_1888; // @[Reg.scala 16:16]
  reg  r_1889; // @[Reg.scala 16:16]
  reg  r_1890; // @[Reg.scala 16:16]
  reg  r_1891; // @[Reg.scala 16:16]
  reg  r_1892; // @[Reg.scala 16:16]
  reg  r_1893; // @[Reg.scala 16:16]
  reg  r_1894; // @[Reg.scala 16:16]
  reg  r_1895; // @[Reg.scala 16:16]
  reg  r_1896; // @[Reg.scala 16:16]
  reg  r_1897; // @[Reg.scala 16:16]
  reg  r_1898; // @[Reg.scala 16:16]
  reg  r_1899; // @[Reg.scala 16:16]
  reg  r_1900; // @[Reg.scala 16:16]
  reg  r_1901; // @[Reg.scala 16:16]
  reg  r_1902; // @[Reg.scala 16:16]
  reg  r_1903; // @[Reg.scala 16:16]
  reg  r_1904; // @[Reg.scala 16:16]
  reg  r_1905; // @[Reg.scala 16:16]
  reg  r_1906; // @[Reg.scala 16:16]
  reg  r_1907; // @[Reg.scala 16:16]
  reg  r_1908; // @[Reg.scala 16:16]
  reg  r_1909; // @[Reg.scala 16:16]
  reg  r_1910; // @[Reg.scala 16:16]
  reg  r_1911; // @[Reg.scala 16:16]
  reg  r_1912; // @[Reg.scala 16:16]
  reg  r_1913; // @[Reg.scala 16:16]
  reg  r_1914; // @[Reg.scala 16:16]
  reg  r_1915; // @[Reg.scala 16:16]
  reg  r_1916; // @[Reg.scala 16:16]
  reg  r_1917; // @[Reg.scala 16:16]
  reg  r_1918; // @[Reg.scala 16:16]
  reg  r_1919; // @[Reg.scala 16:16]
  reg  r_1920; // @[Reg.scala 16:16]
  reg  r_1921; // @[Reg.scala 16:16]
  reg  r_1922; // @[Reg.scala 16:16]
  reg  r_1923; // @[Reg.scala 16:16]
  reg  r_1924; // @[Reg.scala 16:16]
  reg  r_1925; // @[Reg.scala 16:16]
  reg  r_1926; // @[Reg.scala 16:16]
  reg  r_1927; // @[Reg.scala 16:16]
  reg  r_1928; // @[Reg.scala 16:16]
  reg  r_1929; // @[Reg.scala 16:16]
  reg  r_1930; // @[Reg.scala 16:16]
  reg  r_1931; // @[Reg.scala 16:16]
  reg  r_1932; // @[Reg.scala 16:16]
  reg  r_1933; // @[Reg.scala 16:16]
  reg  r_1934; // @[Reg.scala 16:16]
  reg  r_1935; // @[Reg.scala 16:16]
  reg  r_1936; // @[Reg.scala 16:16]
  reg  r_1937; // @[Reg.scala 16:16]
  reg  r_1938; // @[Reg.scala 16:16]
  reg  r_1939; // @[Reg.scala 16:16]
  reg  r_1940; // @[Reg.scala 16:16]
  reg  r_1941; // @[Reg.scala 16:16]
  reg  r_1942; // @[Reg.scala 16:16]
  reg  r_1943; // @[Reg.scala 16:16]
  reg  r_1944; // @[Reg.scala 16:16]
  reg  r_1945; // @[Reg.scala 16:16]
  reg  r_1946; // @[Reg.scala 16:16]
  reg  r_1947; // @[Reg.scala 16:16]
  reg  r_1948; // @[Reg.scala 16:16]
  reg  r_1949; // @[Reg.scala 16:16]
  reg  r_1950; // @[Reg.scala 16:16]
  reg  r_1951; // @[Reg.scala 16:16]
  reg  r_1952; // @[Reg.scala 16:16]
  reg  r_1953; // @[Reg.scala 16:16]
  reg  r_1954; // @[Reg.scala 16:16]
  reg  r_1955; // @[Reg.scala 16:16]
  reg  r_1956; // @[Reg.scala 16:16]
  reg  r_1957; // @[Reg.scala 16:16]
  reg  r_1958; // @[Reg.scala 16:16]
  reg  r_1959; // @[Reg.scala 16:16]
  reg  r_1960; // @[Reg.scala 16:16]
  reg  r_1961; // @[Reg.scala 16:16]
  reg  r_1962; // @[Reg.scala 16:16]
  reg  r_1963; // @[Reg.scala 16:16]
  reg  r_1964; // @[Reg.scala 16:16]
  reg  r_1965; // @[Reg.scala 16:16]
  reg  r_1966; // @[Reg.scala 16:16]
  reg  r_1967; // @[Reg.scala 16:16]
  reg  r_1968; // @[Reg.scala 16:16]
  reg  r_1969; // @[Reg.scala 16:16]
  reg  r_1970; // @[Reg.scala 16:16]
  reg  r_1971; // @[Reg.scala 16:16]
  reg  r_1972; // @[Reg.scala 16:16]
  reg  r_1973; // @[Reg.scala 16:16]
  reg  r_1974; // @[Reg.scala 16:16]
  reg  r_1975; // @[Reg.scala 16:16]
  reg  r_1976; // @[Reg.scala 16:16]
  reg  r_1977; // @[Reg.scala 16:16]
  reg  r_1978; // @[Reg.scala 16:16]
  reg  r_1979; // @[Reg.scala 16:16]
  reg  r_1980; // @[Reg.scala 16:16]
  reg  r_1981; // @[Reg.scala 16:16]
  reg  r_1982; // @[Reg.scala 16:16]
  reg  r_1983; // @[Reg.scala 16:16]
  reg  r_1984; // @[Reg.scala 16:16]
  reg  r_1985; // @[Reg.scala 16:16]
  reg  r_1986; // @[Reg.scala 16:16]
  reg  r_1987; // @[Reg.scala 16:16]
  reg  r_1988; // @[Reg.scala 16:16]
  reg  r_1989; // @[Reg.scala 16:16]
  reg  r_1990; // @[Reg.scala 16:16]
  reg  r_1991; // @[Reg.scala 16:16]
  reg  r_1992; // @[Reg.scala 16:16]
  reg  r_1993; // @[Reg.scala 16:16]
  reg  r_1994; // @[Reg.scala 16:16]
  reg  r_1995; // @[Reg.scala 16:16]
  reg  r_1996; // @[Reg.scala 16:16]
  reg  r_1997; // @[Reg.scala 16:16]
  reg  r_1998; // @[Reg.scala 16:16]
  reg  r_1999; // @[Reg.scala 16:16]
  reg  r_2000; // @[Reg.scala 16:16]
  reg  r_2001; // @[Reg.scala 16:16]
  reg  r_2002; // @[Reg.scala 16:16]
  reg  r_2003; // @[Reg.scala 16:16]
  reg  r_2004; // @[Reg.scala 16:16]
  reg  r_2005; // @[Reg.scala 16:16]
  reg  r_2006; // @[Reg.scala 16:16]
  reg  r_2007; // @[Reg.scala 16:16]
  reg  r_2008; // @[Reg.scala 16:16]
  reg  r_2009; // @[Reg.scala 16:16]
  reg  r_2010; // @[Reg.scala 16:16]
  reg  r_2011; // @[Reg.scala 16:16]
  reg  r_2012; // @[Reg.scala 16:16]
  reg  r_2013; // @[Reg.scala 16:16]
  reg  r_2014; // @[Reg.scala 16:16]
  reg  r_2015; // @[Reg.scala 16:16]
  reg  r_2016; // @[Reg.scala 16:16]
  reg  r_2017; // @[Reg.scala 16:16]
  reg  r_2018; // @[Reg.scala 16:16]
  reg  r_2019; // @[Reg.scala 16:16]
  reg  r_2020; // @[Reg.scala 16:16]
  reg  r_2021; // @[Reg.scala 16:16]
  reg  r_2022; // @[Reg.scala 16:16]
  reg  r_2023; // @[Reg.scala 16:16]
  reg  r_2024; // @[Reg.scala 16:16]
  reg  r_2025; // @[Reg.scala 16:16]
  reg  r_2026; // @[Reg.scala 16:16]
  reg  r_2027; // @[Reg.scala 16:16]
  reg  r_2028; // @[Reg.scala 16:16]
  reg  r_2029; // @[Reg.scala 16:16]
  reg  r_2030; // @[Reg.scala 16:16]
  reg  r_2031; // @[Reg.scala 16:16]
  reg  r_2032; // @[Reg.scala 16:16]
  reg  r_2033; // @[Reg.scala 16:16]
  reg  r_2034; // @[Reg.scala 16:16]
  reg  r_2035; // @[Reg.scala 16:16]
  reg  r_2036; // @[Reg.scala 16:16]
  reg  r_2037; // @[Reg.scala 16:16]
  reg  r_2038; // @[Reg.scala 16:16]
  reg  r_2039; // @[Reg.scala 16:16]
  reg  r_2040; // @[Reg.scala 16:16]
  reg  r_2041; // @[Reg.scala 16:16]
  reg  r_2042; // @[Reg.scala 16:16]
  reg  r_2043; // @[Reg.scala 16:16]
  reg  r_2044; // @[Reg.scala 16:16]
  reg  r_2045; // @[Reg.scala 16:16]
  reg  r_2046; // @[Reg.scala 16:16]
  reg  r_2047; // @[Reg.scala 16:16]
  reg  r_2048; // @[Reg.scala 16:16]
  reg  r_2049; // @[Reg.scala 16:16]
  reg  r_2050; // @[Reg.scala 16:16]
  reg  r_2051; // @[Reg.scala 16:16]
  reg  r_2052; // @[Reg.scala 16:16]
  reg  r_2053; // @[Reg.scala 16:16]
  reg  r_2054; // @[Reg.scala 16:16]
  reg  r_2055; // @[Reg.scala 16:16]
  reg  r_2056; // @[Reg.scala 16:16]
  reg  r_2057; // @[Reg.scala 16:16]
  reg  r_2058; // @[Reg.scala 16:16]
  reg  r_2059; // @[Reg.scala 16:16]
  reg  r_2060; // @[Reg.scala 16:16]
  reg  r_2061; // @[Reg.scala 16:16]
  reg  r_2062; // @[Reg.scala 16:16]
  reg  r_2063; // @[Reg.scala 16:16]
  reg  r_2064; // @[Reg.scala 16:16]
  reg  r_2065; // @[Reg.scala 16:16]
  reg  r_2066; // @[Reg.scala 16:16]
  reg  r_2067; // @[Reg.scala 16:16]
  reg  r_2068; // @[Reg.scala 16:16]
  reg  r_2069; // @[Reg.scala 16:16]
  reg  r_2070; // @[Reg.scala 16:16]
  reg  r_2071; // @[Reg.scala 16:16]
  reg  r_2072; // @[Reg.scala 16:16]
  reg  r_2073; // @[Reg.scala 16:16]
  reg  r_2074; // @[Reg.scala 16:16]
  reg  r_2075; // @[Reg.scala 16:16]
  reg  r_2076; // @[Reg.scala 16:16]
  reg  r_2077; // @[Reg.scala 16:16]
  reg  r_2078; // @[Reg.scala 16:16]
  reg  r_2079; // @[Reg.scala 16:16]
  reg  r_2080; // @[Reg.scala 16:16]
  reg  r_2081; // @[Reg.scala 16:16]
  reg  r_2082; // @[Reg.scala 16:16]
  reg  r_2083; // @[Reg.scala 16:16]
  reg  r_2084; // @[Reg.scala 16:16]
  reg  r_2085; // @[Reg.scala 16:16]
  reg  r_2086; // @[Reg.scala 16:16]
  reg  r_2087; // @[Reg.scala 16:16]
  reg  r_2088; // @[Reg.scala 16:16]
  reg  r_2089; // @[Reg.scala 16:16]
  reg  r_2090; // @[Reg.scala 16:16]
  reg  r_2091; // @[Reg.scala 16:16]
  reg  r_2092; // @[Reg.scala 16:16]
  reg  r_2093; // @[Reg.scala 16:16]
  reg  r_2094; // @[Reg.scala 16:16]
  reg  r_2095; // @[Reg.scala 16:16]
  reg  r_2096; // @[Reg.scala 16:16]
  reg  r_2097; // @[Reg.scala 16:16]
  reg  r_2098; // @[Reg.scala 16:16]
  reg  r_2099; // @[Reg.scala 16:16]
  reg  r_2100; // @[Reg.scala 16:16]
  reg  r_2101; // @[Reg.scala 16:16]
  reg  r_2102; // @[Reg.scala 16:16]
  reg  r_2103; // @[Reg.scala 16:16]
  reg  r_2104; // @[Reg.scala 16:16]
  reg  r_2105; // @[Reg.scala 16:16]
  reg  r_2106; // @[Reg.scala 16:16]
  reg  r_2107; // @[Reg.scala 16:16]
  reg  r_2108; // @[Reg.scala 16:16]
  reg  r_2109; // @[Reg.scala 16:16]
  reg  r_2110; // @[Reg.scala 16:16]
  reg  r_2111; // @[Reg.scala 16:16]
  reg  r_2112; // @[Reg.scala 16:16]
  reg  r_2113; // @[Reg.scala 16:16]
  reg  r_2114; // @[Reg.scala 16:16]
  reg  r_2115; // @[Reg.scala 16:16]
  reg  r_2116; // @[Reg.scala 16:16]
  reg  r_2117; // @[Reg.scala 16:16]
  reg  r_2118; // @[Reg.scala 16:16]
  reg  r_2119; // @[Reg.scala 16:16]
  reg  r_2120; // @[Reg.scala 16:16]
  reg  r_2121; // @[Reg.scala 16:16]
  reg  r_2122; // @[Reg.scala 16:16]
  reg  r_2123; // @[Reg.scala 16:16]
  reg  r_2124; // @[Reg.scala 16:16]
  reg  r_2125; // @[Reg.scala 16:16]
  reg  r_2126; // @[Reg.scala 16:16]
  reg  r_2127; // @[Reg.scala 16:16]
  reg  r_2128; // @[Reg.scala 16:16]
  reg  r_2129; // @[Reg.scala 16:16]
  reg  r_2130; // @[Reg.scala 16:16]
  reg  r_2131; // @[Reg.scala 16:16]
  reg  r_2132; // @[Reg.scala 16:16]
  reg  r_2133; // @[Reg.scala 16:16]
  reg  r_2134; // @[Reg.scala 16:16]
  reg  r_2135; // @[Reg.scala 16:16]
  reg  r_2136; // @[Reg.scala 16:16]
  reg  r_2137; // @[Reg.scala 16:16]
  reg  r_2138; // @[Reg.scala 16:16]
  reg  r_2139; // @[Reg.scala 16:16]
  reg  r_2140; // @[Reg.scala 16:16]
  reg  r_2141; // @[Reg.scala 16:16]
  reg  r_2142; // @[Reg.scala 16:16]
  reg  r_2143; // @[Reg.scala 16:16]
  reg  r_2144; // @[Reg.scala 16:16]
  reg  r_2145; // @[Reg.scala 16:16]
  reg  r_2146; // @[Reg.scala 16:16]
  reg  r_2147; // @[Reg.scala 16:16]
  reg  r_2148; // @[Reg.scala 16:16]
  reg  r_2149; // @[Reg.scala 16:16]
  reg  r_2150; // @[Reg.scala 16:16]
  reg  r_2151; // @[Reg.scala 16:16]
  reg  r_2152; // @[Reg.scala 16:16]
  reg  r_2153; // @[Reg.scala 16:16]
  reg  r_2154; // @[Reg.scala 16:16]
  reg  r_2155; // @[Reg.scala 16:16]
  reg  r_2156; // @[Reg.scala 16:16]
  reg  r_2157; // @[Reg.scala 16:16]
  reg  r_2158; // @[Reg.scala 16:16]
  reg  r_2159; // @[Reg.scala 16:16]
  reg  r_2160; // @[Reg.scala 16:16]
  reg  r_2161; // @[Reg.scala 16:16]
  reg  r_2162; // @[Reg.scala 16:16]
  reg  r_2163; // @[Reg.scala 16:16]
  reg  r_2164; // @[Reg.scala 16:16]
  reg  r_2165; // @[Reg.scala 16:16]
  reg  r_2166; // @[Reg.scala 16:16]
  reg  r_2167; // @[Reg.scala 16:16]
  reg  r_2168; // @[Reg.scala 16:16]
  reg  r_2169; // @[Reg.scala 16:16]
  reg  r_2170; // @[Reg.scala 16:16]
  reg  r_2171; // @[Reg.scala 16:16]
  reg  r_2172; // @[Reg.scala 16:16]
  reg  r_2173; // @[Reg.scala 16:16]
  reg  r_2174; // @[Reg.scala 16:16]
  reg  r_2175; // @[Reg.scala 16:16]
  reg  r_2176; // @[Reg.scala 16:16]
  reg  r_2177; // @[Reg.scala 16:16]
  reg  r_2178; // @[Reg.scala 16:16]
  reg  r_2179; // @[Reg.scala 16:16]
  reg  r_2180; // @[Reg.scala 16:16]
  reg  r_2181; // @[Reg.scala 16:16]
  reg  r_2182; // @[Reg.scala 16:16]
  reg  r_2183; // @[Reg.scala 16:16]
  reg  r_2184; // @[Reg.scala 16:16]
  reg  r_2185; // @[Reg.scala 16:16]
  reg  r_2186; // @[Reg.scala 16:16]
  reg  r_2187; // @[Reg.scala 16:16]
  reg  r_2188; // @[Reg.scala 16:16]
  reg  r_2189; // @[Reg.scala 16:16]
  reg  r_2190; // @[Reg.scala 16:16]
  reg  r_2191; // @[Reg.scala 16:16]
  reg  r_2192; // @[Reg.scala 16:16]
  reg  r_2193; // @[Reg.scala 16:16]
  reg  r_2194; // @[Reg.scala 16:16]
  reg  r_2195; // @[Reg.scala 16:16]
  reg  r_2196; // @[Reg.scala 16:16]
  reg  r_2197; // @[Reg.scala 16:16]
  reg  r_2198; // @[Reg.scala 16:16]
  reg  r_2199; // @[Reg.scala 16:16]
  reg  r_2200; // @[Reg.scala 16:16]
  reg  r_2201; // @[Reg.scala 16:16]
  reg  r_2202; // @[Reg.scala 16:16]
  reg  r_2203; // @[Reg.scala 16:16]
  reg  r_2204; // @[Reg.scala 16:16]
  reg  r_2205; // @[Reg.scala 16:16]
  reg  r_2206; // @[Reg.scala 16:16]
  reg  r_2207; // @[Reg.scala 16:16]
  reg  r_2208; // @[Reg.scala 16:16]
  reg  r_2209; // @[Reg.scala 16:16]
  reg  r_2210; // @[Reg.scala 16:16]
  reg  r_2211; // @[Reg.scala 16:16]
  reg  r_2212; // @[Reg.scala 16:16]
  reg  r_2213; // @[Reg.scala 16:16]
  reg  r_2214; // @[Reg.scala 16:16]
  reg  r_2215; // @[Reg.scala 16:16]
  reg  r_2216; // @[Reg.scala 16:16]
  reg  r_2217; // @[Reg.scala 16:16]
  reg  r_2218; // @[Reg.scala 16:16]
  reg  r_2219; // @[Reg.scala 16:16]
  reg  r_2220; // @[Reg.scala 16:16]
  reg  r_2221; // @[Reg.scala 16:16]
  reg  r_2222; // @[Reg.scala 16:16]
  reg  r_2223; // @[Reg.scala 16:16]
  reg  r_2224; // @[Reg.scala 16:16]
  reg  r_2225; // @[Reg.scala 16:16]
  reg  r_2226; // @[Reg.scala 16:16]
  reg  r_2227; // @[Reg.scala 16:16]
  reg  r_2228; // @[Reg.scala 16:16]
  reg  r_2229; // @[Reg.scala 16:16]
  reg  r_2230; // @[Reg.scala 16:16]
  reg  r_2231; // @[Reg.scala 16:16]
  reg  r_2232; // @[Reg.scala 16:16]
  reg  r_2233; // @[Reg.scala 16:16]
  reg  r_2234; // @[Reg.scala 16:16]
  reg  r_2235; // @[Reg.scala 16:16]
  reg  r_2236; // @[Reg.scala 16:16]
  reg  r_2237; // @[Reg.scala 16:16]
  reg  r_2238; // @[Reg.scala 16:16]
  reg  r_2239; // @[Reg.scala 16:16]
  reg  r_2240; // @[Reg.scala 16:16]
  reg  r_2241; // @[Reg.scala 16:16]
  reg  r_2242; // @[Reg.scala 16:16]
  reg  r_2243; // @[Reg.scala 16:16]
  reg  r_2244; // @[Reg.scala 16:16]
  reg  r_2245; // @[Reg.scala 16:16]
  reg  r_2246; // @[Reg.scala 16:16]
  reg  r_2247; // @[Reg.scala 16:16]
  reg  r_2248; // @[Reg.scala 16:16]
  reg  r_2249; // @[Reg.scala 16:16]
  reg  r_2250; // @[Reg.scala 16:16]
  reg  r_2251; // @[Reg.scala 16:16]
  reg  r_2252; // @[Reg.scala 16:16]
  reg  r_2253; // @[Reg.scala 16:16]
  reg  r_2254; // @[Reg.scala 16:16]
  reg  r_2255; // @[Reg.scala 16:16]
  reg  r_2256; // @[Reg.scala 16:16]
  reg  r_2257; // @[Reg.scala 16:16]
  reg  r_2258; // @[Reg.scala 16:16]
  reg  r_2259; // @[Reg.scala 16:16]
  reg  r_2260; // @[Reg.scala 16:16]
  reg  r_2261; // @[Reg.scala 16:16]
  reg  r_2262; // @[Reg.scala 16:16]
  reg  r_2263; // @[Reg.scala 16:16]
  reg  r_2264; // @[Reg.scala 16:16]
  reg  r_2265; // @[Reg.scala 16:16]
  reg  r_2266; // @[Reg.scala 16:16]
  reg  r_2267; // @[Reg.scala 16:16]
  reg  r_2268; // @[Reg.scala 16:16]
  reg  r_2269; // @[Reg.scala 16:16]
  reg  r_2270; // @[Reg.scala 16:16]
  reg  r_2271; // @[Reg.scala 16:16]
  reg  r_2272; // @[Reg.scala 16:16]
  reg  r_2273; // @[Reg.scala 16:16]
  reg  r_2274; // @[Reg.scala 16:16]
  reg  r_2275; // @[Reg.scala 16:16]
  reg  r_2276; // @[Reg.scala 16:16]
  reg  r_2277; // @[Reg.scala 16:16]
  reg  r_2278; // @[Reg.scala 16:16]
  reg  r_2279; // @[Reg.scala 16:16]
  reg  r_2280; // @[Reg.scala 16:16]
  reg  r_2281; // @[Reg.scala 16:16]
  reg  r_2282; // @[Reg.scala 16:16]
  reg  r_2283; // @[Reg.scala 16:16]
  reg  r_2284; // @[Reg.scala 16:16]
  reg  r_2285; // @[Reg.scala 16:16]
  reg  r_2286; // @[Reg.scala 16:16]
  reg  r_2287; // @[Reg.scala 16:16]
  reg  r_2288; // @[Reg.scala 16:16]
  reg  r_2289; // @[Reg.scala 16:16]
  reg  r_2290; // @[Reg.scala 16:16]
  reg  r_2291; // @[Reg.scala 16:16]
  reg  r_2292; // @[Reg.scala 16:16]
  reg  r_2293; // @[Reg.scala 16:16]
  reg  r_2294; // @[Reg.scala 16:16]
  reg  r_2295; // @[Reg.scala 16:16]
  reg  r_2296; // @[Reg.scala 16:16]
  reg  r_2297; // @[Reg.scala 16:16]
  reg  r_2298; // @[Reg.scala 16:16]
  reg  r_2299; // @[Reg.scala 16:16]
  reg  r_2300; // @[Reg.scala 16:16]
  reg  r_2301; // @[Reg.scala 16:16]
  reg  r_2302; // @[Reg.scala 16:16]
  reg  r_2303; // @[Reg.scala 16:16]
  reg  r_2304; // @[Reg.scala 16:16]
  reg  r_2305; // @[Reg.scala 16:16]
  reg  r_2306; // @[Reg.scala 16:16]
  wire  s_0 = c22_io_out_0; // @[Multiplier.scala 122:35]
  wire  s_0_130 = c22_32_io_out_0; // @[Multiplier.scala 122:35]
  wire  s_0_259 = c22_75_io_out_0; // @[Multiplier.scala 122:35]
  wire  s_0_387 = c22_125_io_out_0; // @[Multiplier.scala 122:35]
  wire  s_0_514 = c22_178_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_514 = c22_178_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_515 = c22_179_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_515 = c22_179_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_516 = c22_180_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_516 = c22_180_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_517 = c22_181_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_517 = c22_181_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_518 = c22_182_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_518 = c22_182_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_519 = c22_183_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_519 = c22_183_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_520 = c22_184_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_520 = c22_184_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_521 = c22_185_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_521 = c22_185_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_522 = c22_186_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_522 = c22_186_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_523 = c22_187_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_523 = c22_187_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_524 = c22_188_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_524 = c22_188_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_525 = c22_189_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_525 = c22_189_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_526 = c22_190_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_526 = c22_190_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_527 = c22_191_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_527 = c22_191_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_528 = c22_192_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_528 = c22_192_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_529 = c22_193_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_529 = c22_193_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_530 = c22_194_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_530 = c22_194_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_531 = c22_195_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_531 = c22_195_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_532 = c22_196_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_532 = c22_196_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_533 = c22_197_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_533 = c22_197_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_534 = c22_198_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_534 = c22_198_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_535 = c22_199_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_535 = c22_199_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_536 = c22_200_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_536 = c22_200_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_537 = c22_201_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_537 = c22_201_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_538 = c22_202_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_538 = c22_202_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_539 = c22_203_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_539 = c22_203_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_540 = c22_204_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_540 = c22_204_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_541 = c22_205_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_541 = c22_205_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_542 = c22_206_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_542 = c22_206_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_543 = c22_207_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_543 = c22_207_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_544 = c22_208_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_544 = c22_208_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_545 = c22_209_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_545 = c22_209_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_546 = c22_210_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_546 = c22_210_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_547 = c22_211_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_547 = c22_211_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_548 = c22_212_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_548 = c22_212_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_549 = c22_213_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_549 = c22_213_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_550 = c22_214_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_550 = c22_214_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_551 = c22_215_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_551 = c22_215_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_552 = c22_216_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_552 = c22_216_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_553 = c22_217_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_553 = c22_217_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_554 = c22_218_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_554 = c22_218_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_555 = c22_219_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_555 = c22_219_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_556 = c22_220_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_556 = c22_220_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_557 = c22_221_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_557 = c22_221_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_558 = c22_222_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_558 = c22_222_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_559 = c22_223_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_559 = c22_223_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_560 = c22_224_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_560 = c22_224_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_561 = c22_225_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_561 = c22_225_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_562 = c22_226_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_562 = c22_226_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_563 = c22_227_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_563 = c22_227_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_564 = c22_228_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_564 = c22_228_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_565 = c22_229_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_565 = c22_229_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_566 = c22_230_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_566 = c22_230_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_567 = c22_231_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_567 = c22_231_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_568 = c22_232_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_568 = c22_232_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_569 = c22_233_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_569 = c22_233_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_570 = c22_234_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_570 = c22_234_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_571 = c22_235_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_571 = c22_235_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_572 = c32_73_io_out_0; // @[Multiplier.scala 127:35]
  wire  c2_0_572 = c32_73_io_out_1; // @[Multiplier.scala 128:41]
  wire  s_0_573 = c32_74_io_out_0; // @[Multiplier.scala 127:35]
  wire  c2_0_573 = c32_74_io_out_1; // @[Multiplier.scala 128:41]
  wire  s_0_574 = c32_75_io_out_0; // @[Multiplier.scala 127:35]
  wire  c2_0_574 = c32_75_io_out_1; // @[Multiplier.scala 128:41]
  wire  s_0_575 = c32_76_io_out_0; // @[Multiplier.scala 127:35]
  wire  c2_0_575 = c32_76_io_out_1; // @[Multiplier.scala 128:41]
  wire  s_0_576 = c32_77_io_out_0; // @[Multiplier.scala 127:35]
  wire  c2_0_576 = c32_77_io_out_1; // @[Multiplier.scala 128:41]
  wire  s_0_577 = c32_78_io_out_0; // @[Multiplier.scala 127:35]
  wire  c2_0_577 = c32_78_io_out_1; // @[Multiplier.scala 128:41]
  wire  s_0_578 = c32_79_io_out_0; // @[Multiplier.scala 127:35]
  wire  c2_0_578 = c32_79_io_out_1; // @[Multiplier.scala 128:41]
  wire  s_0_579 = c22_236_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_579 = c22_236_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_580 = c32_80_io_out_0; // @[Multiplier.scala 127:35]
  wire  c2_0_580 = c32_80_io_out_1; // @[Multiplier.scala 128:41]
  wire  s_0_581 = c22_237_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_581 = c22_237_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_582 = c22_238_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_582 = c22_238_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_583 = c22_239_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_583 = c22_239_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_584 = c22_240_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_584 = c22_240_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_585 = c32_81_io_out_0; // @[Multiplier.scala 127:35]
  wire  c2_0_585 = c32_81_io_out_1; // @[Multiplier.scala 128:41]
  wire  s_0_586 = c22_241_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_586 = c22_241_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_587 = c22_242_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_587 = c22_242_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_588 = c22_243_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_588 = c22_243_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_589 = c22_244_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_589 = c22_244_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_590 = c22_245_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_590 = c22_245_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_591 = c22_246_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_591 = c22_246_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_592 = c22_247_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_592 = c22_247_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_593 = c22_248_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_593 = c22_248_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_594 = c32_82_io_out_0; // @[Multiplier.scala 127:35]
  wire  c2_0_594 = c32_82_io_out_1; // @[Multiplier.scala 128:41]
  wire  s_0_595 = c22_249_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_595 = c22_249_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_596 = c22_250_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_596 = c22_250_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_597 = c22_251_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_597 = c22_251_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_598 = c22_252_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_598 = c22_252_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_599 = c22_253_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_599 = c22_253_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_600 = c22_254_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_600 = c22_254_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_601 = c22_255_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_601 = c22_255_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_602 = c22_256_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_602 = c22_256_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_603 = c22_257_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_603 = c22_257_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_604 = c22_258_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_604 = c22_258_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_605 = c22_259_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_605 = c22_259_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_606 = c22_260_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_606 = c22_260_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_607 = c22_261_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_607 = c22_261_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_608 = c22_262_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_608 = c22_262_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_609 = c22_263_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_609 = c22_263_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_610 = c32_83_io_out_0; // @[Multiplier.scala 127:35]
  wire  c2_0_610 = c32_83_io_out_1; // @[Multiplier.scala 128:41]
  wire  s_0_611 = c22_264_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_611 = c22_264_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_612 = c22_265_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_612 = c22_265_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_613 = c22_266_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_613 = c22_266_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_614 = c22_267_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_614 = c22_267_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_615 = c22_268_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_615 = c22_268_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_616 = c22_269_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_616 = c22_269_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_617 = c22_270_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_617 = c22_270_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_618 = c22_271_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_618 = c22_271_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_619 = c22_272_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_619 = c22_272_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_620 = c22_273_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_620 = c22_273_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_621 = c22_274_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_621 = c22_274_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_622 = c22_275_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_622 = c22_275_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_623 = c22_276_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_623 = c22_276_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_624 = c22_277_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_624 = c22_277_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_625 = c22_278_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_625 = c22_278_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_626 = c22_279_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_626 = c22_279_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_627 = c22_280_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_627 = c22_280_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_628 = c22_281_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_628 = c22_281_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_629 = c22_282_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_629 = c22_282_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_630 = c22_283_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_630 = c22_283_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_631 = c22_284_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_631 = c22_284_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_632 = c22_285_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_632 = c22_285_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_633 = c22_286_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_633 = c22_286_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_634 = c22_287_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_634 = c22_287_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_635 = c22_288_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_635 = c22_288_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_636 = c22_289_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_636 = c22_289_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_637 = c22_290_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_637 = c22_290_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_638 = c22_291_io_out_0; // @[Multiplier.scala 122:35]
  wire  c2_0_638 = c22_291_io_out_1; // @[Multiplier.scala 123:41]
  wire  s_0_639 = c22_292_io_out_0; // @[Multiplier.scala 122:35]
  reg  r_2307; // @[Reg.scala 16:16]
  reg  r_2308; // @[Reg.scala 16:16]
  reg  r_2309; // @[Reg.scala 16:16]
  reg  r_2310; // @[Reg.scala 16:16]
  reg  r_2311; // @[Reg.scala 16:16]
  reg  r_2312; // @[Reg.scala 16:16]
  reg  r_2313; // @[Reg.scala 16:16]
  reg  r_2314; // @[Reg.scala 16:16]
  reg  r_2315; // @[Reg.scala 16:16]
  reg  r_2316; // @[Reg.scala 16:16]
  reg  r_2317; // @[Reg.scala 16:16]
  reg  r_2318; // @[Reg.scala 16:16]
  reg  r_2319; // @[Reg.scala 16:16]
  reg  r_2320; // @[Reg.scala 16:16]
  reg  r_2321; // @[Reg.scala 16:16]
  reg  r_2322; // @[Reg.scala 16:16]
  reg  r_2323; // @[Reg.scala 16:16]
  reg  r_2324; // @[Reg.scala 16:16]
  reg  r_2325; // @[Reg.scala 16:16]
  reg  r_2326; // @[Reg.scala 16:16]
  reg  r_2327; // @[Reg.scala 16:16]
  reg  r_2328; // @[Reg.scala 16:16]
  reg  r_2329; // @[Reg.scala 16:16]
  reg  r_2330; // @[Reg.scala 16:16]
  reg  r_2331; // @[Reg.scala 16:16]
  reg  r_2332; // @[Reg.scala 16:16]
  reg  r_2333; // @[Reg.scala 16:16]
  reg  r_2334; // @[Reg.scala 16:16]
  reg  r_2335; // @[Reg.scala 16:16]
  reg  r_2336; // @[Reg.scala 16:16]
  reg  r_2337; // @[Reg.scala 16:16]
  reg  r_2338; // @[Reg.scala 16:16]
  reg  r_2339; // @[Reg.scala 16:16]
  reg  r_2340; // @[Reg.scala 16:16]
  reg  r_2341; // @[Reg.scala 16:16]
  reg  r_2342; // @[Reg.scala 16:16]
  reg  r_2343; // @[Reg.scala 16:16]
  reg  r_2344; // @[Reg.scala 16:16]
  reg  r_2345; // @[Reg.scala 16:16]
  reg  r_2346; // @[Reg.scala 16:16]
  reg  r_2347; // @[Reg.scala 16:16]
  reg  r_2348; // @[Reg.scala 16:16]
  reg  r_2349; // @[Reg.scala 16:16]
  reg  r_2350; // @[Reg.scala 16:16]
  reg  r_2351; // @[Reg.scala 16:16]
  reg  r_2352; // @[Reg.scala 16:16]
  reg  r_2353; // @[Reg.scala 16:16]
  reg  r_2354; // @[Reg.scala 16:16]
  reg  r_2355; // @[Reg.scala 16:16]
  reg  r_2356; // @[Reg.scala 16:16]
  reg  r_2357; // @[Reg.scala 16:16]
  reg  r_2358; // @[Reg.scala 16:16]
  reg  r_2359; // @[Reg.scala 16:16]
  reg  r_2360; // @[Reg.scala 16:16]
  reg  r_2361; // @[Reg.scala 16:16]
  reg  r_2362; // @[Reg.scala 16:16]
  reg  r_2363; // @[Reg.scala 16:16]
  reg  r_2364; // @[Reg.scala 16:16]
  reg  r_2365; // @[Reg.scala 16:16]
  reg  r_2366; // @[Reg.scala 16:16]
  reg  r_2367; // @[Reg.scala 16:16]
  reg  r_2368; // @[Reg.scala 16:16]
  reg  r_2369; // @[Reg.scala 16:16]
  reg  r_2370; // @[Reg.scala 16:16]
  reg  r_2371; // @[Reg.scala 16:16]
  reg  r_2372; // @[Reg.scala 16:16]
  reg  r_2373; // @[Reg.scala 16:16]
  reg  r_2374; // @[Reg.scala 16:16]
  reg  r_2375; // @[Reg.scala 16:16]
  reg  r_2376; // @[Reg.scala 16:16]
  reg  r_2377; // @[Reg.scala 16:16]
  reg  r_2378; // @[Reg.scala 16:16]
  reg  r_2379; // @[Reg.scala 16:16]
  reg  r_2380; // @[Reg.scala 16:16]
  reg  r_2381; // @[Reg.scala 16:16]
  reg  r_2382; // @[Reg.scala 16:16]
  reg  r_2383; // @[Reg.scala 16:16]
  reg  r_2384; // @[Reg.scala 16:16]
  reg  r_2385; // @[Reg.scala 16:16]
  reg  r_2386; // @[Reg.scala 16:16]
  reg  r_2387; // @[Reg.scala 16:16]
  reg  r_2388; // @[Reg.scala 16:16]
  reg  r_2389; // @[Reg.scala 16:16]
  reg  r_2390; // @[Reg.scala 16:16]
  reg  r_2391; // @[Reg.scala 16:16]
  reg  r_2392; // @[Reg.scala 16:16]
  reg  r_2393; // @[Reg.scala 16:16]
  reg  r_2394; // @[Reg.scala 16:16]
  reg  r_2395; // @[Reg.scala 16:16]
  reg  r_2396; // @[Reg.scala 16:16]
  reg  r_2397; // @[Reg.scala 16:16]
  reg  r_2398; // @[Reg.scala 16:16]
  reg  r_2399; // @[Reg.scala 16:16]
  reg  r_2400; // @[Reg.scala 16:16]
  reg  r_2401; // @[Reg.scala 16:16]
  reg  r_2402; // @[Reg.scala 16:16]
  reg  r_2403; // @[Reg.scala 16:16]
  reg  r_2404; // @[Reg.scala 16:16]
  reg  r_2405; // @[Reg.scala 16:16]
  reg  r_2406; // @[Reg.scala 16:16]
  reg  r_2407; // @[Reg.scala 16:16]
  reg  r_2408; // @[Reg.scala 16:16]
  reg  r_2409; // @[Reg.scala 16:16]
  reg  r_2410; // @[Reg.scala 16:16]
  reg  r_2411; // @[Reg.scala 16:16]
  reg  r_2412; // @[Reg.scala 16:16]
  reg  r_2413; // @[Reg.scala 16:16]
  reg  r_2414; // @[Reg.scala 16:16]
  reg  r_2415; // @[Reg.scala 16:16]
  reg  r_2416; // @[Reg.scala 16:16]
  reg  r_2417; // @[Reg.scala 16:16]
  reg  r_2418; // @[Reg.scala 16:16]
  reg  r_2419; // @[Reg.scala 16:16]
  reg  r_2420; // @[Reg.scala 16:16]
  reg  r_2421; // @[Reg.scala 16:16]
  reg  r_2422; // @[Reg.scala 16:16]
  reg  r_2423; // @[Reg.scala 16:16]
  reg  r_2424; // @[Reg.scala 16:16]
  reg  r_2425; // @[Reg.scala 16:16]
  reg  r_2426; // @[Reg.scala 16:16]
  reg  r_2427; // @[Reg.scala 16:16]
  reg  r_2428; // @[Reg.scala 16:16]
  reg  r_2429; // @[Reg.scala 16:16]
  reg  r_2430; // @[Reg.scala 16:16]
  reg  r_2431; // @[Reg.scala 16:16]
  reg  r_2432; // @[Reg.scala 16:16]
  reg  r_2433; // @[Reg.scala 16:16]
  reg  r_2434; // @[Reg.scala 16:16]
  reg  r_2435; // @[Reg.scala 16:16]
  reg  r_2436; // @[Reg.scala 16:16]
  reg  r_2437; // @[Reg.scala 16:16]
  reg  r_2438; // @[Reg.scala 16:16]
  reg  r_2439; // @[Reg.scala 16:16]
  reg  r_2440; // @[Reg.scala 16:16]
  reg  r_2441; // @[Reg.scala 16:16]
  reg  r_2442; // @[Reg.scala 16:16]
  reg  r_2443; // @[Reg.scala 16:16]
  reg  r_2444; // @[Reg.scala 16:16]
  reg  r_2445; // @[Reg.scala 16:16]
  reg  r_2446; // @[Reg.scala 16:16]
  reg  r_2447; // @[Reg.scala 16:16]
  reg  r_2448; // @[Reg.scala 16:16]
  reg  r_2449; // @[Reg.scala 16:16]
  reg  r_2450; // @[Reg.scala 16:16]
  reg  r_2451; // @[Reg.scala 16:16]
  reg  r_2452; // @[Reg.scala 16:16]
  reg  r_2453; // @[Reg.scala 16:16]
  reg  r_2454; // @[Reg.scala 16:16]
  reg  r_2455; // @[Reg.scala 16:16]
  reg  r_2456; // @[Reg.scala 16:16]
  reg  r_2457; // @[Reg.scala 16:16]
  reg  r_2458; // @[Reg.scala 16:16]
  reg  r_2459; // @[Reg.scala 16:16]
  reg  r_2460; // @[Reg.scala 16:16]
  reg  r_2461; // @[Reg.scala 16:16]
  reg  r_2462; // @[Reg.scala 16:16]
  reg  r_2463; // @[Reg.scala 16:16]
  reg  r_2464; // @[Reg.scala 16:16]
  reg  r_2465; // @[Reg.scala 16:16]
  reg  r_2466; // @[Reg.scala 16:16]
  reg  r_2467; // @[Reg.scala 16:16]
  reg  r_2468; // @[Reg.scala 16:16]
  reg  r_2469; // @[Reg.scala 16:16]
  reg  r_2470; // @[Reg.scala 16:16]
  reg  r_2471; // @[Reg.scala 16:16]
  reg  r_2472; // @[Reg.scala 16:16]
  reg  r_2473; // @[Reg.scala 16:16]
  reg  r_2474; // @[Reg.scala 16:16]
  reg  r_2475; // @[Reg.scala 16:16]
  reg  r_2476; // @[Reg.scala 16:16]
  reg  r_2477; // @[Reg.scala 16:16]
  reg  r_2478; // @[Reg.scala 16:16]
  reg  r_2479; // @[Reg.scala 16:16]
  reg  r_2480; // @[Reg.scala 16:16]
  reg  r_2481; // @[Reg.scala 16:16]
  reg  r_2482; // @[Reg.scala 16:16]
  reg  r_2483; // @[Reg.scala 16:16]
  reg  r_2484; // @[Reg.scala 16:16]
  reg  r_2485; // @[Reg.scala 16:16]
  reg  r_2486; // @[Reg.scala 16:16]
  reg  r_2487; // @[Reg.scala 16:16]
  reg  r_2488; // @[Reg.scala 16:16]
  reg  r_2489; // @[Reg.scala 16:16]
  reg  r_2490; // @[Reg.scala 16:16]
  reg  r_2491; // @[Reg.scala 16:16]
  reg  r_2492; // @[Reg.scala 16:16]
  reg  r_2493; // @[Reg.scala 16:16]
  reg  r_2494; // @[Reg.scala 16:16]
  reg  r_2495; // @[Reg.scala 16:16]
  reg  r_2496; // @[Reg.scala 16:16]
  reg  r_2497; // @[Reg.scala 16:16]
  reg  r_2498; // @[Reg.scala 16:16]
  reg  r_2499; // @[Reg.scala 16:16]
  reg  r_2500; // @[Reg.scala 16:16]
  reg  r_2501; // @[Reg.scala 16:16]
  reg  r_2502; // @[Reg.scala 16:16]
  reg  r_2503; // @[Reg.scala 16:16]
  reg  r_2504; // @[Reg.scala 16:16]
  reg  r_2505; // @[Reg.scala 16:16]
  reg  r_2506; // @[Reg.scala 16:16]
  reg  r_2507; // @[Reg.scala 16:16]
  reg  r_2508; // @[Reg.scala 16:16]
  reg  r_2509; // @[Reg.scala 16:16]
  reg  r_2510; // @[Reg.scala 16:16]
  reg  r_2511; // @[Reg.scala 16:16]
  reg  r_2512; // @[Reg.scala 16:16]
  reg  r_2513; // @[Reg.scala 16:16]
  reg  r_2514; // @[Reg.scala 16:16]
  reg  r_2515; // @[Reg.scala 16:16]
  reg  r_2516; // @[Reg.scala 16:16]
  reg  r_2517; // @[Reg.scala 16:16]
  reg  r_2518; // @[Reg.scala 16:16]
  reg  r_2519; // @[Reg.scala 16:16]
  reg  r_2520; // @[Reg.scala 16:16]
  reg  r_2521; // @[Reg.scala 16:16]
  reg  r_2522; // @[Reg.scala 16:16]
  reg  r_2523; // @[Reg.scala 16:16]
  reg  r_2524; // @[Reg.scala 16:16]
  reg  r_2525; // @[Reg.scala 16:16]
  reg  r_2526; // @[Reg.scala 16:16]
  reg  r_2527; // @[Reg.scala 16:16]
  reg  r_2528; // @[Reg.scala 16:16]
  reg  r_2529; // @[Reg.scala 16:16]
  reg  r_2530; // @[Reg.scala 16:16]
  reg  r_2531; // @[Reg.scala 16:16]
  reg  r_2532; // @[Reg.scala 16:16]
  reg  r_2533; // @[Reg.scala 16:16]
  reg  r_2534; // @[Reg.scala 16:16]
  reg  r_2535; // @[Reg.scala 16:16]
  reg  r_2536; // @[Reg.scala 16:16]
  reg  r_2537; // @[Reg.scala 16:16]
  reg  r_2538; // @[Reg.scala 16:16]
  reg  r_2539; // @[Reg.scala 16:16]
  reg  r_2540; // @[Reg.scala 16:16]
  reg  r_2541; // @[Reg.scala 16:16]
  reg  r_2542; // @[Reg.scala 16:16]
  reg  r_2543; // @[Reg.scala 16:16]
  reg  r_2544; // @[Reg.scala 16:16]
  reg  r_2545; // @[Reg.scala 16:16]
  reg  r_2546; // @[Reg.scala 16:16]
  reg  r_2547; // @[Reg.scala 16:16]
  reg  r_2548; // @[Reg.scala 16:16]
  reg  r_2549; // @[Reg.scala 16:16]
  reg  r_2550; // @[Reg.scala 16:16]
  reg  r_2551; // @[Reg.scala 16:16]
  reg  r_2552; // @[Reg.scala 16:16]
  reg  r_2553; // @[Reg.scala 16:16]
  reg  r_2554; // @[Reg.scala 16:16]
  reg  r_2555; // @[Reg.scala 16:16]
  reg  r_2556; // @[Reg.scala 16:16]
  reg  r_2557; // @[Reg.scala 16:16]
  reg  r_2558; // @[Reg.scala 16:16]
  reg  r_2559; // @[Reg.scala 16:16]
  reg  r_2560; // @[Reg.scala 16:16]
  reg  r_2561; // @[Reg.scala 16:16]
  wire [7:0] sum_lo_lo_lo_lo = {r_2316,r_2314,r_2312,r_2311,r_2310,r_2309,r_2308,r_2307}; // @[Cat.scala 31:58]
  wire [15:0] sum_lo_lo_lo = {r_2332,r_2330,r_2328,r_2326,r_2324,r_2322,r_2320,r_2318,sum_lo_lo_lo_lo}; // @[Cat.scala 31:58]
  wire [7:0] sum_lo_lo_hi_lo = {r_2348,r_2346,r_2344,r_2342,r_2340,r_2338,r_2336,r_2334}; // @[Cat.scala 31:58]
  wire [31:0] sum_lo_lo = {r_2364,r_2362,r_2360,r_2358,r_2356,r_2354,r_2352,r_2350,sum_lo_lo_hi_lo,sum_lo_lo_lo}; // @[Cat.scala 31:58]
  wire [7:0] sum_lo_hi_lo_lo = {r_2380,r_2378,r_2376,r_2374,r_2372,r_2370,r_2368,r_2366}; // @[Cat.scala 31:58]
  wire [7:0] sum_lo_hi_hi_lo = {r_2412,r_2410,r_2408,r_2406,r_2404,r_2402,r_2400,r_2398}; // @[Cat.scala 31:58]
  wire [16:0] sum_lo_hi_hi = {r_2430,r_2428,r_2426,r_2424,r_2422,r_2420,r_2418,r_2416,r_2414,sum_lo_hi_hi_lo}; // @[Cat.scala 31:58]
  wire [32:0] sum_lo_hi = {sum_lo_hi_hi,r_2396,r_2394,r_2392,r_2390,r_2388,r_2386,r_2384,r_2382,sum_lo_hi_lo_lo}; // @[Cat.scala 31:58]
  wire [7:0] sum_hi_lo_lo_lo = {r_2446,r_2444,r_2442,r_2440,r_2438,r_2436,r_2434,r_2432}; // @[Cat.scala 31:58]
  wire [15:0] sum_hi_lo_lo = {r_2462,r_2460,r_2458,r_2456,r_2454,r_2452,r_2450,r_2448,sum_hi_lo_lo_lo}; // @[Cat.scala 31:58]
  wire [7:0] sum_hi_lo_hi_lo = {r_2478,r_2476,r_2474,r_2472,r_2470,r_2468,r_2466,r_2464}; // @[Cat.scala 31:58]
  wire [31:0] sum_hi_lo = {r_2494,r_2492,r_2490,r_2488,r_2486,r_2484,r_2482,r_2480,sum_hi_lo_hi_lo,sum_hi_lo_lo}; // @[Cat.scala 31:58]
  wire [7:0] sum_hi_hi_lo_lo = {r_2510,r_2508,r_2506,r_2504,r_2502,r_2500,r_2498,r_2496}; // @[Cat.scala 31:58]
  wire [7:0] sum_hi_hi_hi_lo = {r_2542,r_2540,r_2538,r_2536,r_2534,r_2532,r_2530,r_2528}; // @[Cat.scala 31:58]
  wire [16:0] sum_hi_hi_hi = {r_2560,r_2558,r_2556,r_2554,r_2552,r_2550,r_2548,r_2546,r_2544,sum_hi_hi_hi_lo}; // @[Cat.scala 31:58]
  wire [32:0] sum_hi_hi = {sum_hi_hi_hi,r_2526,r_2524,r_2522,r_2520,r_2518,r_2516,r_2514,r_2512,sum_hi_hi_lo_lo}; // @[Cat.scala 31:58]
  wire [129:0] sum = {sum_hi_hi,sum_hi_lo,sum_lo_hi,sum_lo_lo}; // @[Cat.scala 31:58]
  wire [6:0] carry_lo_lo_lo_lo = {r_2325,r_2323,r_2321,r_2319,r_2317,r_2315,r_2313}; // @[Cat.scala 31:58]
  wire [14:0] carry_lo_lo_lo = {r_2341,r_2339,r_2337,r_2335,r_2333,r_2331,r_2329,r_2327,carry_lo_lo_lo_lo}; // @[Cat.scala 31:58]
  wire [7:0] carry_lo_lo_hi_lo = {r_2357,r_2355,r_2353,r_2351,r_2349,r_2347,r_2345,r_2343}; // @[Cat.scala 31:58]
  wire [30:0] carry_lo_lo = {r_2373,r_2371,r_2369,r_2367,r_2365,r_2363,r_2361,r_2359,carry_lo_lo_hi_lo,carry_lo_lo_lo}; // @[Cat.scala 31:58]
  wire [6:0] carry_lo_hi_lo_lo = {r_2387,r_2385,r_2383,r_2381,r_2379,r_2377,r_2375}; // @[Cat.scala 31:58]
  wire [14:0] carry_lo_hi_lo = {r_2403,r_2401,r_2399,r_2397,r_2395,r_2393,r_2391,r_2389,carry_lo_hi_lo_lo}; // @[Cat.scala 31:58]
  wire [7:0] carry_lo_hi_hi_lo = {r_2419,r_2417,r_2415,r_2413,r_2411,r_2409,r_2407,r_2405}; // @[Cat.scala 31:58]
  wire [30:0] carry_lo_hi = {r_2435,r_2433,r_2431,r_2429,r_2427,r_2425,r_2423,r_2421,carry_lo_hi_hi_lo,carry_lo_hi_lo}; // @[Cat.scala 31:58]
  wire [6:0] carry_hi_lo_lo_lo = {r_2449,r_2447,r_2445,r_2443,r_2441,r_2439,r_2437}; // @[Cat.scala 31:58]
  wire [14:0] carry_hi_lo_lo = {r_2465,r_2463,r_2461,r_2459,r_2457,r_2455,r_2453,r_2451,carry_hi_lo_lo_lo}; // @[Cat.scala 31:58]
  wire [7:0] carry_hi_lo_hi_lo = {r_2481,r_2479,r_2477,r_2475,r_2473,r_2471,r_2469,r_2467}; // @[Cat.scala 31:58]
  wire [30:0] carry_hi_lo = {r_2497,r_2495,r_2493,r_2491,r_2489,r_2487,r_2485,r_2483,carry_hi_lo_hi_lo,carry_hi_lo_lo}; // @[Cat.scala 31:58]
  wire [7:0] carry_hi_hi_lo_lo = {r_2513,r_2511,r_2509,r_2507,r_2505,r_2503,r_2501,r_2499}; // @[Cat.scala 31:58]
  wire [15:0] carry_hi_hi_lo = {r_2529,r_2527,r_2525,r_2523,r_2521,r_2519,r_2517,r_2515,carry_hi_hi_lo_lo}; // @[Cat.scala 31:58]
  wire [7:0] carry_hi_hi_hi_lo = {r_2545,r_2543,r_2541,r_2539,r_2537,r_2535,r_2533,r_2531}; // @[Cat.scala 31:58]
  wire [31:0] carry_hi_hi = {r_2561,r_2559,r_2557,r_2555,r_2553,r_2551,r_2549,r_2547,carry_hi_hi_hi_lo,carry_hi_hi_lo}; // @[Cat.scala 31:58]
  wire [129:0] carry_1 = {carry_hi_hi,carry_hi_lo,carry_lo_hi,carry_lo_lo,5'h0}; // @[Cat.scala 31:58]
  C22 c22 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_io_in_0),
    .io_in_1(c22_io_in_1),
    .io_out_0(c22_io_out_0),
    .io_out_1(c22_io_out_1)
  );
  C22 c22_1 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_1_io_in_0),
    .io_in_1(c22_1_io_in_1),
    .io_out_0(c22_1_io_out_0),
    .io_out_1(c22_1_io_out_1)
  );
  C32 c32 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_io_in_0),
    .io_in_1(c32_io_in_1),
    .io_in_2(c32_io_in_2),
    .io_out_0(c32_io_out_0),
    .io_out_1(c32_io_out_1)
  );
  C32 c32_1 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_1_io_in_0),
    .io_in_1(c32_1_io_in_1),
    .io_in_2(c32_1_io_in_2),
    .io_out_0(c32_1_io_out_0),
    .io_out_1(c32_1_io_out_1)
  );
  C53 c53 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_io_in_0),
    .io_in_1(c53_io_in_1),
    .io_in_2(c53_io_in_2),
    .io_in_3(c53_io_in_3),
    .io_in_4(c53_io_in_4),
    .io_out_0(c53_io_out_0),
    .io_out_1(c53_io_out_1),
    .io_out_2(c53_io_out_2)
  );
  C53 c53_1 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_1_io_in_0),
    .io_in_1(c53_1_io_in_1),
    .io_in_2(c53_1_io_in_2),
    .io_in_3(c53_1_io_in_3),
    .io_in_4(c53_1_io_in_4),
    .io_out_0(c53_1_io_out_0),
    .io_out_1(c53_1_io_out_1),
    .io_out_2(c53_1_io_out_2)
  );
  C53 c53_2 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_2_io_in_0),
    .io_in_1(c53_2_io_in_1),
    .io_in_2(c53_2_io_in_2),
    .io_in_3(c53_2_io_in_3),
    .io_in_4(c53_2_io_in_4),
    .io_out_0(c53_2_io_out_0),
    .io_out_1(c53_2_io_out_1),
    .io_out_2(c53_2_io_out_2)
  );
  C53 c53_3 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_3_io_in_0),
    .io_in_1(c53_3_io_in_1),
    .io_in_2(c53_3_io_in_2),
    .io_in_3(c53_3_io_in_3),
    .io_in_4(c53_3_io_in_4),
    .io_out_0(c53_3_io_out_0),
    .io_out_1(c53_3_io_out_1),
    .io_out_2(c53_3_io_out_2)
  );
  C53 c53_4 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_4_io_in_0),
    .io_in_1(c53_4_io_in_1),
    .io_in_2(c53_4_io_in_2),
    .io_in_3(c53_4_io_in_3),
    .io_in_4(c53_4_io_in_4),
    .io_out_0(c53_4_io_out_0),
    .io_out_1(c53_4_io_out_1),
    .io_out_2(c53_4_io_out_2)
  );
  C22 c22_2 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_2_io_in_0),
    .io_in_1(c22_2_io_in_1),
    .io_out_0(c22_2_io_out_0),
    .io_out_1(c22_2_io_out_1)
  );
  C53 c53_5 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_5_io_in_0),
    .io_in_1(c53_5_io_in_1),
    .io_in_2(c53_5_io_in_2),
    .io_in_3(c53_5_io_in_3),
    .io_in_4(c53_5_io_in_4),
    .io_out_0(c53_5_io_out_0),
    .io_out_1(c53_5_io_out_1),
    .io_out_2(c53_5_io_out_2)
  );
  C22 c22_3 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_3_io_in_0),
    .io_in_1(c22_3_io_in_1),
    .io_out_0(c22_3_io_out_0),
    .io_out_1(c22_3_io_out_1)
  );
  C53 c53_6 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_6_io_in_0),
    .io_in_1(c53_6_io_in_1),
    .io_in_2(c53_6_io_in_2),
    .io_in_3(c53_6_io_in_3),
    .io_in_4(c53_6_io_in_4),
    .io_out_0(c53_6_io_out_0),
    .io_out_1(c53_6_io_out_1),
    .io_out_2(c53_6_io_out_2)
  );
  C32 c32_2 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_2_io_in_0),
    .io_in_1(c32_2_io_in_1),
    .io_in_2(c32_2_io_in_2),
    .io_out_0(c32_2_io_out_0),
    .io_out_1(c32_2_io_out_1)
  );
  C53 c53_7 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_7_io_in_0),
    .io_in_1(c53_7_io_in_1),
    .io_in_2(c53_7_io_in_2),
    .io_in_3(c53_7_io_in_3),
    .io_in_4(c53_7_io_in_4),
    .io_out_0(c53_7_io_out_0),
    .io_out_1(c53_7_io_out_1),
    .io_out_2(c53_7_io_out_2)
  );
  C32 c32_3 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_3_io_in_0),
    .io_in_1(c32_3_io_in_1),
    .io_in_2(c32_3_io_in_2),
    .io_out_0(c32_3_io_out_0),
    .io_out_1(c32_3_io_out_1)
  );
  C53 c53_8 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_8_io_in_0),
    .io_in_1(c53_8_io_in_1),
    .io_in_2(c53_8_io_in_2),
    .io_in_3(c53_8_io_in_3),
    .io_in_4(c53_8_io_in_4),
    .io_out_0(c53_8_io_out_0),
    .io_out_1(c53_8_io_out_1),
    .io_out_2(c53_8_io_out_2)
  );
  C53 c53_9 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_9_io_in_0),
    .io_in_1(c53_9_io_in_1),
    .io_in_2(c53_9_io_in_2),
    .io_in_3(c53_9_io_in_3),
    .io_in_4(c53_9_io_in_4),
    .io_out_0(c53_9_io_out_0),
    .io_out_1(c53_9_io_out_1),
    .io_out_2(c53_9_io_out_2)
  );
  C53 c53_10 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_10_io_in_0),
    .io_in_1(c53_10_io_in_1),
    .io_in_2(c53_10_io_in_2),
    .io_in_3(c53_10_io_in_3),
    .io_in_4(c53_10_io_in_4),
    .io_out_0(c53_10_io_out_0),
    .io_out_1(c53_10_io_out_1),
    .io_out_2(c53_10_io_out_2)
  );
  C53 c53_11 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_11_io_in_0),
    .io_in_1(c53_11_io_in_1),
    .io_in_2(c53_11_io_in_2),
    .io_in_3(c53_11_io_in_3),
    .io_in_4(c53_11_io_in_4),
    .io_out_0(c53_11_io_out_0),
    .io_out_1(c53_11_io_out_1),
    .io_out_2(c53_11_io_out_2)
  );
  C53 c53_12 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_12_io_in_0),
    .io_in_1(c53_12_io_in_1),
    .io_in_2(c53_12_io_in_2),
    .io_in_3(c53_12_io_in_3),
    .io_in_4(c53_12_io_in_4),
    .io_out_0(c53_12_io_out_0),
    .io_out_1(c53_12_io_out_1),
    .io_out_2(c53_12_io_out_2)
  );
  C53 c53_13 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_13_io_in_0),
    .io_in_1(c53_13_io_in_1),
    .io_in_2(c53_13_io_in_2),
    .io_in_3(c53_13_io_in_3),
    .io_in_4(c53_13_io_in_4),
    .io_out_0(c53_13_io_out_0),
    .io_out_1(c53_13_io_out_1),
    .io_out_2(c53_13_io_out_2)
  );
  C53 c53_14 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_14_io_in_0),
    .io_in_1(c53_14_io_in_1),
    .io_in_2(c53_14_io_in_2),
    .io_in_3(c53_14_io_in_3),
    .io_in_4(c53_14_io_in_4),
    .io_out_0(c53_14_io_out_0),
    .io_out_1(c53_14_io_out_1),
    .io_out_2(c53_14_io_out_2)
  );
  C53 c53_15 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_15_io_in_0),
    .io_in_1(c53_15_io_in_1),
    .io_in_2(c53_15_io_in_2),
    .io_in_3(c53_15_io_in_3),
    .io_in_4(c53_15_io_in_4),
    .io_out_0(c53_15_io_out_0),
    .io_out_1(c53_15_io_out_1),
    .io_out_2(c53_15_io_out_2)
  );
  C53 c53_16 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_16_io_in_0),
    .io_in_1(c53_16_io_in_1),
    .io_in_2(c53_16_io_in_2),
    .io_in_3(c53_16_io_in_3),
    .io_in_4(c53_16_io_in_4),
    .io_out_0(c53_16_io_out_0),
    .io_out_1(c53_16_io_out_1),
    .io_out_2(c53_16_io_out_2)
  );
  C53 c53_17 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_17_io_in_0),
    .io_in_1(c53_17_io_in_1),
    .io_in_2(c53_17_io_in_2),
    .io_in_3(c53_17_io_in_3),
    .io_in_4(c53_17_io_in_4),
    .io_out_0(c53_17_io_out_0),
    .io_out_1(c53_17_io_out_1),
    .io_out_2(c53_17_io_out_2)
  );
  C22 c22_4 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_4_io_in_0),
    .io_in_1(c22_4_io_in_1),
    .io_out_0(c22_4_io_out_0),
    .io_out_1(c22_4_io_out_1)
  );
  C53 c53_18 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_18_io_in_0),
    .io_in_1(c53_18_io_in_1),
    .io_in_2(c53_18_io_in_2),
    .io_in_3(c53_18_io_in_3),
    .io_in_4(c53_18_io_in_4),
    .io_out_0(c53_18_io_out_0),
    .io_out_1(c53_18_io_out_1),
    .io_out_2(c53_18_io_out_2)
  );
  C53 c53_19 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_19_io_in_0),
    .io_in_1(c53_19_io_in_1),
    .io_in_2(c53_19_io_in_2),
    .io_in_3(c53_19_io_in_3),
    .io_in_4(c53_19_io_in_4),
    .io_out_0(c53_19_io_out_0),
    .io_out_1(c53_19_io_out_1),
    .io_out_2(c53_19_io_out_2)
  );
  C22 c22_5 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_5_io_in_0),
    .io_in_1(c22_5_io_in_1),
    .io_out_0(c22_5_io_out_0),
    .io_out_1(c22_5_io_out_1)
  );
  C53 c53_20 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_20_io_in_0),
    .io_in_1(c53_20_io_in_1),
    .io_in_2(c53_20_io_in_2),
    .io_in_3(c53_20_io_in_3),
    .io_in_4(c53_20_io_in_4),
    .io_out_0(c53_20_io_out_0),
    .io_out_1(c53_20_io_out_1),
    .io_out_2(c53_20_io_out_2)
  );
  C53 c53_21 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_21_io_in_0),
    .io_in_1(c53_21_io_in_1),
    .io_in_2(c53_21_io_in_2),
    .io_in_3(c53_21_io_in_3),
    .io_in_4(c53_21_io_in_4),
    .io_out_0(c53_21_io_out_0),
    .io_out_1(c53_21_io_out_1),
    .io_out_2(c53_21_io_out_2)
  );
  C32 c32_4 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_4_io_in_0),
    .io_in_1(c32_4_io_in_1),
    .io_in_2(c32_4_io_in_2),
    .io_out_0(c32_4_io_out_0),
    .io_out_1(c32_4_io_out_1)
  );
  C53 c53_22 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_22_io_in_0),
    .io_in_1(c53_22_io_in_1),
    .io_in_2(c53_22_io_in_2),
    .io_in_3(c53_22_io_in_3),
    .io_in_4(c53_22_io_in_4),
    .io_out_0(c53_22_io_out_0),
    .io_out_1(c53_22_io_out_1),
    .io_out_2(c53_22_io_out_2)
  );
  C53 c53_23 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_23_io_in_0),
    .io_in_1(c53_23_io_in_1),
    .io_in_2(c53_23_io_in_2),
    .io_in_3(c53_23_io_in_3),
    .io_in_4(c53_23_io_in_4),
    .io_out_0(c53_23_io_out_0),
    .io_out_1(c53_23_io_out_1),
    .io_out_2(c53_23_io_out_2)
  );
  C32 c32_5 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_5_io_in_0),
    .io_in_1(c32_5_io_in_1),
    .io_in_2(c32_5_io_in_2),
    .io_out_0(c32_5_io_out_0),
    .io_out_1(c32_5_io_out_1)
  );
  C53 c53_24 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_24_io_in_0),
    .io_in_1(c53_24_io_in_1),
    .io_in_2(c53_24_io_in_2),
    .io_in_3(c53_24_io_in_3),
    .io_in_4(c53_24_io_in_4),
    .io_out_0(c53_24_io_out_0),
    .io_out_1(c53_24_io_out_1),
    .io_out_2(c53_24_io_out_2)
  );
  C53 c53_25 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_25_io_in_0),
    .io_in_1(c53_25_io_in_1),
    .io_in_2(c53_25_io_in_2),
    .io_in_3(c53_25_io_in_3),
    .io_in_4(c53_25_io_in_4),
    .io_out_0(c53_25_io_out_0),
    .io_out_1(c53_25_io_out_1),
    .io_out_2(c53_25_io_out_2)
  );
  C53 c53_26 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_26_io_in_0),
    .io_in_1(c53_26_io_in_1),
    .io_in_2(c53_26_io_in_2),
    .io_in_3(c53_26_io_in_3),
    .io_in_4(c53_26_io_in_4),
    .io_out_0(c53_26_io_out_0),
    .io_out_1(c53_26_io_out_1),
    .io_out_2(c53_26_io_out_2)
  );
  C53 c53_27 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_27_io_in_0),
    .io_in_1(c53_27_io_in_1),
    .io_in_2(c53_27_io_in_2),
    .io_in_3(c53_27_io_in_3),
    .io_in_4(c53_27_io_in_4),
    .io_out_0(c53_27_io_out_0),
    .io_out_1(c53_27_io_out_1),
    .io_out_2(c53_27_io_out_2)
  );
  C53 c53_28 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_28_io_in_0),
    .io_in_1(c53_28_io_in_1),
    .io_in_2(c53_28_io_in_2),
    .io_in_3(c53_28_io_in_3),
    .io_in_4(c53_28_io_in_4),
    .io_out_0(c53_28_io_out_0),
    .io_out_1(c53_28_io_out_1),
    .io_out_2(c53_28_io_out_2)
  );
  C53 c53_29 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_29_io_in_0),
    .io_in_1(c53_29_io_in_1),
    .io_in_2(c53_29_io_in_2),
    .io_in_3(c53_29_io_in_3),
    .io_in_4(c53_29_io_in_4),
    .io_out_0(c53_29_io_out_0),
    .io_out_1(c53_29_io_out_1),
    .io_out_2(c53_29_io_out_2)
  );
  C53 c53_30 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_30_io_in_0),
    .io_in_1(c53_30_io_in_1),
    .io_in_2(c53_30_io_in_2),
    .io_in_3(c53_30_io_in_3),
    .io_in_4(c53_30_io_in_4),
    .io_out_0(c53_30_io_out_0),
    .io_out_1(c53_30_io_out_1),
    .io_out_2(c53_30_io_out_2)
  );
  C53 c53_31 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_31_io_in_0),
    .io_in_1(c53_31_io_in_1),
    .io_in_2(c53_31_io_in_2),
    .io_in_3(c53_31_io_in_3),
    .io_in_4(c53_31_io_in_4),
    .io_out_0(c53_31_io_out_0),
    .io_out_1(c53_31_io_out_1),
    .io_out_2(c53_31_io_out_2)
  );
  C53 c53_32 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_32_io_in_0),
    .io_in_1(c53_32_io_in_1),
    .io_in_2(c53_32_io_in_2),
    .io_in_3(c53_32_io_in_3),
    .io_in_4(c53_32_io_in_4),
    .io_out_0(c53_32_io_out_0),
    .io_out_1(c53_32_io_out_1),
    .io_out_2(c53_32_io_out_2)
  );
  C53 c53_33 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_33_io_in_0),
    .io_in_1(c53_33_io_in_1),
    .io_in_2(c53_33_io_in_2),
    .io_in_3(c53_33_io_in_3),
    .io_in_4(c53_33_io_in_4),
    .io_out_0(c53_33_io_out_0),
    .io_out_1(c53_33_io_out_1),
    .io_out_2(c53_33_io_out_2)
  );
  C53 c53_34 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_34_io_in_0),
    .io_in_1(c53_34_io_in_1),
    .io_in_2(c53_34_io_in_2),
    .io_in_3(c53_34_io_in_3),
    .io_in_4(c53_34_io_in_4),
    .io_out_0(c53_34_io_out_0),
    .io_out_1(c53_34_io_out_1),
    .io_out_2(c53_34_io_out_2)
  );
  C53 c53_35 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_35_io_in_0),
    .io_in_1(c53_35_io_in_1),
    .io_in_2(c53_35_io_in_2),
    .io_in_3(c53_35_io_in_3),
    .io_in_4(c53_35_io_in_4),
    .io_out_0(c53_35_io_out_0),
    .io_out_1(c53_35_io_out_1),
    .io_out_2(c53_35_io_out_2)
  );
  C53 c53_36 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_36_io_in_0),
    .io_in_1(c53_36_io_in_1),
    .io_in_2(c53_36_io_in_2),
    .io_in_3(c53_36_io_in_3),
    .io_in_4(c53_36_io_in_4),
    .io_out_0(c53_36_io_out_0),
    .io_out_1(c53_36_io_out_1),
    .io_out_2(c53_36_io_out_2)
  );
  C53 c53_37 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_37_io_in_0),
    .io_in_1(c53_37_io_in_1),
    .io_in_2(c53_37_io_in_2),
    .io_in_3(c53_37_io_in_3),
    .io_in_4(c53_37_io_in_4),
    .io_out_0(c53_37_io_out_0),
    .io_out_1(c53_37_io_out_1),
    .io_out_2(c53_37_io_out_2)
  );
  C53 c53_38 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_38_io_in_0),
    .io_in_1(c53_38_io_in_1),
    .io_in_2(c53_38_io_in_2),
    .io_in_3(c53_38_io_in_3),
    .io_in_4(c53_38_io_in_4),
    .io_out_0(c53_38_io_out_0),
    .io_out_1(c53_38_io_out_1),
    .io_out_2(c53_38_io_out_2)
  );
  C22 c22_6 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_6_io_in_0),
    .io_in_1(c22_6_io_in_1),
    .io_out_0(c22_6_io_out_0),
    .io_out_1(c22_6_io_out_1)
  );
  C53 c53_39 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_39_io_in_0),
    .io_in_1(c53_39_io_in_1),
    .io_in_2(c53_39_io_in_2),
    .io_in_3(c53_39_io_in_3),
    .io_in_4(c53_39_io_in_4),
    .io_out_0(c53_39_io_out_0),
    .io_out_1(c53_39_io_out_1),
    .io_out_2(c53_39_io_out_2)
  );
  C53 c53_40 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_40_io_in_0),
    .io_in_1(c53_40_io_in_1),
    .io_in_2(c53_40_io_in_2),
    .io_in_3(c53_40_io_in_3),
    .io_in_4(c53_40_io_in_4),
    .io_out_0(c53_40_io_out_0),
    .io_out_1(c53_40_io_out_1),
    .io_out_2(c53_40_io_out_2)
  );
  C53 c53_41 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_41_io_in_0),
    .io_in_1(c53_41_io_in_1),
    .io_in_2(c53_41_io_in_2),
    .io_in_3(c53_41_io_in_3),
    .io_in_4(c53_41_io_in_4),
    .io_out_0(c53_41_io_out_0),
    .io_out_1(c53_41_io_out_1),
    .io_out_2(c53_41_io_out_2)
  );
  C22 c22_7 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_7_io_in_0),
    .io_in_1(c22_7_io_in_1),
    .io_out_0(c22_7_io_out_0),
    .io_out_1(c22_7_io_out_1)
  );
  C53 c53_42 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_42_io_in_0),
    .io_in_1(c53_42_io_in_1),
    .io_in_2(c53_42_io_in_2),
    .io_in_3(c53_42_io_in_3),
    .io_in_4(c53_42_io_in_4),
    .io_out_0(c53_42_io_out_0),
    .io_out_1(c53_42_io_out_1),
    .io_out_2(c53_42_io_out_2)
  );
  C53 c53_43 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_43_io_in_0),
    .io_in_1(c53_43_io_in_1),
    .io_in_2(c53_43_io_in_2),
    .io_in_3(c53_43_io_in_3),
    .io_in_4(c53_43_io_in_4),
    .io_out_0(c53_43_io_out_0),
    .io_out_1(c53_43_io_out_1),
    .io_out_2(c53_43_io_out_2)
  );
  C53 c53_44 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_44_io_in_0),
    .io_in_1(c53_44_io_in_1),
    .io_in_2(c53_44_io_in_2),
    .io_in_3(c53_44_io_in_3),
    .io_in_4(c53_44_io_in_4),
    .io_out_0(c53_44_io_out_0),
    .io_out_1(c53_44_io_out_1),
    .io_out_2(c53_44_io_out_2)
  );
  C32 c32_6 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_6_io_in_0),
    .io_in_1(c32_6_io_in_1),
    .io_in_2(c32_6_io_in_2),
    .io_out_0(c32_6_io_out_0),
    .io_out_1(c32_6_io_out_1)
  );
  C53 c53_45 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_45_io_in_0),
    .io_in_1(c53_45_io_in_1),
    .io_in_2(c53_45_io_in_2),
    .io_in_3(c53_45_io_in_3),
    .io_in_4(c53_45_io_in_4),
    .io_out_0(c53_45_io_out_0),
    .io_out_1(c53_45_io_out_1),
    .io_out_2(c53_45_io_out_2)
  );
  C53 c53_46 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_46_io_in_0),
    .io_in_1(c53_46_io_in_1),
    .io_in_2(c53_46_io_in_2),
    .io_in_3(c53_46_io_in_3),
    .io_in_4(c53_46_io_in_4),
    .io_out_0(c53_46_io_out_0),
    .io_out_1(c53_46_io_out_1),
    .io_out_2(c53_46_io_out_2)
  );
  C53 c53_47 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_47_io_in_0),
    .io_in_1(c53_47_io_in_1),
    .io_in_2(c53_47_io_in_2),
    .io_in_3(c53_47_io_in_3),
    .io_in_4(c53_47_io_in_4),
    .io_out_0(c53_47_io_out_0),
    .io_out_1(c53_47_io_out_1),
    .io_out_2(c53_47_io_out_2)
  );
  C32 c32_7 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_7_io_in_0),
    .io_in_1(c32_7_io_in_1),
    .io_in_2(c32_7_io_in_2),
    .io_out_0(c32_7_io_out_0),
    .io_out_1(c32_7_io_out_1)
  );
  C53 c53_48 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_48_io_in_0),
    .io_in_1(c53_48_io_in_1),
    .io_in_2(c53_48_io_in_2),
    .io_in_3(c53_48_io_in_3),
    .io_in_4(c53_48_io_in_4),
    .io_out_0(c53_48_io_out_0),
    .io_out_1(c53_48_io_out_1),
    .io_out_2(c53_48_io_out_2)
  );
  C53 c53_49 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_49_io_in_0),
    .io_in_1(c53_49_io_in_1),
    .io_in_2(c53_49_io_in_2),
    .io_in_3(c53_49_io_in_3),
    .io_in_4(c53_49_io_in_4),
    .io_out_0(c53_49_io_out_0),
    .io_out_1(c53_49_io_out_1),
    .io_out_2(c53_49_io_out_2)
  );
  C53 c53_50 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_50_io_in_0),
    .io_in_1(c53_50_io_in_1),
    .io_in_2(c53_50_io_in_2),
    .io_in_3(c53_50_io_in_3),
    .io_in_4(c53_50_io_in_4),
    .io_out_0(c53_50_io_out_0),
    .io_out_1(c53_50_io_out_1),
    .io_out_2(c53_50_io_out_2)
  );
  C53 c53_51 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_51_io_in_0),
    .io_in_1(c53_51_io_in_1),
    .io_in_2(c53_51_io_in_2),
    .io_in_3(c53_51_io_in_3),
    .io_in_4(c53_51_io_in_4),
    .io_out_0(c53_51_io_out_0),
    .io_out_1(c53_51_io_out_1),
    .io_out_2(c53_51_io_out_2)
  );
  C53 c53_52 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_52_io_in_0),
    .io_in_1(c53_52_io_in_1),
    .io_in_2(c53_52_io_in_2),
    .io_in_3(c53_52_io_in_3),
    .io_in_4(c53_52_io_in_4),
    .io_out_0(c53_52_io_out_0),
    .io_out_1(c53_52_io_out_1),
    .io_out_2(c53_52_io_out_2)
  );
  C53 c53_53 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_53_io_in_0),
    .io_in_1(c53_53_io_in_1),
    .io_in_2(c53_53_io_in_2),
    .io_in_3(c53_53_io_in_3),
    .io_in_4(c53_53_io_in_4),
    .io_out_0(c53_53_io_out_0),
    .io_out_1(c53_53_io_out_1),
    .io_out_2(c53_53_io_out_2)
  );
  C53 c53_54 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_54_io_in_0),
    .io_in_1(c53_54_io_in_1),
    .io_in_2(c53_54_io_in_2),
    .io_in_3(c53_54_io_in_3),
    .io_in_4(c53_54_io_in_4),
    .io_out_0(c53_54_io_out_0),
    .io_out_1(c53_54_io_out_1),
    .io_out_2(c53_54_io_out_2)
  );
  C53 c53_55 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_55_io_in_0),
    .io_in_1(c53_55_io_in_1),
    .io_in_2(c53_55_io_in_2),
    .io_in_3(c53_55_io_in_3),
    .io_in_4(c53_55_io_in_4),
    .io_out_0(c53_55_io_out_0),
    .io_out_1(c53_55_io_out_1),
    .io_out_2(c53_55_io_out_2)
  );
  C53 c53_56 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_56_io_in_0),
    .io_in_1(c53_56_io_in_1),
    .io_in_2(c53_56_io_in_2),
    .io_in_3(c53_56_io_in_3),
    .io_in_4(c53_56_io_in_4),
    .io_out_0(c53_56_io_out_0),
    .io_out_1(c53_56_io_out_1),
    .io_out_2(c53_56_io_out_2)
  );
  C53 c53_57 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_57_io_in_0),
    .io_in_1(c53_57_io_in_1),
    .io_in_2(c53_57_io_in_2),
    .io_in_3(c53_57_io_in_3),
    .io_in_4(c53_57_io_in_4),
    .io_out_0(c53_57_io_out_0),
    .io_out_1(c53_57_io_out_1),
    .io_out_2(c53_57_io_out_2)
  );
  C53 c53_58 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_58_io_in_0),
    .io_in_1(c53_58_io_in_1),
    .io_in_2(c53_58_io_in_2),
    .io_in_3(c53_58_io_in_3),
    .io_in_4(c53_58_io_in_4),
    .io_out_0(c53_58_io_out_0),
    .io_out_1(c53_58_io_out_1),
    .io_out_2(c53_58_io_out_2)
  );
  C53 c53_59 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_59_io_in_0),
    .io_in_1(c53_59_io_in_1),
    .io_in_2(c53_59_io_in_2),
    .io_in_3(c53_59_io_in_3),
    .io_in_4(c53_59_io_in_4),
    .io_out_0(c53_59_io_out_0),
    .io_out_1(c53_59_io_out_1),
    .io_out_2(c53_59_io_out_2)
  );
  C53 c53_60 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_60_io_in_0),
    .io_in_1(c53_60_io_in_1),
    .io_in_2(c53_60_io_in_2),
    .io_in_3(c53_60_io_in_3),
    .io_in_4(c53_60_io_in_4),
    .io_out_0(c53_60_io_out_0),
    .io_out_1(c53_60_io_out_1),
    .io_out_2(c53_60_io_out_2)
  );
  C53 c53_61 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_61_io_in_0),
    .io_in_1(c53_61_io_in_1),
    .io_in_2(c53_61_io_in_2),
    .io_in_3(c53_61_io_in_3),
    .io_in_4(c53_61_io_in_4),
    .io_out_0(c53_61_io_out_0),
    .io_out_1(c53_61_io_out_1),
    .io_out_2(c53_61_io_out_2)
  );
  C53 c53_62 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_62_io_in_0),
    .io_in_1(c53_62_io_in_1),
    .io_in_2(c53_62_io_in_2),
    .io_in_3(c53_62_io_in_3),
    .io_in_4(c53_62_io_in_4),
    .io_out_0(c53_62_io_out_0),
    .io_out_1(c53_62_io_out_1),
    .io_out_2(c53_62_io_out_2)
  );
  C53 c53_63 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_63_io_in_0),
    .io_in_1(c53_63_io_in_1),
    .io_in_2(c53_63_io_in_2),
    .io_in_3(c53_63_io_in_3),
    .io_in_4(c53_63_io_in_4),
    .io_out_0(c53_63_io_out_0),
    .io_out_1(c53_63_io_out_1),
    .io_out_2(c53_63_io_out_2)
  );
  C53 c53_64 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_64_io_in_0),
    .io_in_1(c53_64_io_in_1),
    .io_in_2(c53_64_io_in_2),
    .io_in_3(c53_64_io_in_3),
    .io_in_4(c53_64_io_in_4),
    .io_out_0(c53_64_io_out_0),
    .io_out_1(c53_64_io_out_1),
    .io_out_2(c53_64_io_out_2)
  );
  C53 c53_65 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_65_io_in_0),
    .io_in_1(c53_65_io_in_1),
    .io_in_2(c53_65_io_in_2),
    .io_in_3(c53_65_io_in_3),
    .io_in_4(c53_65_io_in_4),
    .io_out_0(c53_65_io_out_0),
    .io_out_1(c53_65_io_out_1),
    .io_out_2(c53_65_io_out_2)
  );
  C53 c53_66 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_66_io_in_0),
    .io_in_1(c53_66_io_in_1),
    .io_in_2(c53_66_io_in_2),
    .io_in_3(c53_66_io_in_3),
    .io_in_4(c53_66_io_in_4),
    .io_out_0(c53_66_io_out_0),
    .io_out_1(c53_66_io_out_1),
    .io_out_2(c53_66_io_out_2)
  );
  C53 c53_67 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_67_io_in_0),
    .io_in_1(c53_67_io_in_1),
    .io_in_2(c53_67_io_in_2),
    .io_in_3(c53_67_io_in_3),
    .io_in_4(c53_67_io_in_4),
    .io_out_0(c53_67_io_out_0),
    .io_out_1(c53_67_io_out_1),
    .io_out_2(c53_67_io_out_2)
  );
  C22 c22_8 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_8_io_in_0),
    .io_in_1(c22_8_io_in_1),
    .io_out_0(c22_8_io_out_0),
    .io_out_1(c22_8_io_out_1)
  );
  C53 c53_68 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_68_io_in_0),
    .io_in_1(c53_68_io_in_1),
    .io_in_2(c53_68_io_in_2),
    .io_in_3(c53_68_io_in_3),
    .io_in_4(c53_68_io_in_4),
    .io_out_0(c53_68_io_out_0),
    .io_out_1(c53_68_io_out_1),
    .io_out_2(c53_68_io_out_2)
  );
  C53 c53_69 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_69_io_in_0),
    .io_in_1(c53_69_io_in_1),
    .io_in_2(c53_69_io_in_2),
    .io_in_3(c53_69_io_in_3),
    .io_in_4(c53_69_io_in_4),
    .io_out_0(c53_69_io_out_0),
    .io_out_1(c53_69_io_out_1),
    .io_out_2(c53_69_io_out_2)
  );
  C53 c53_70 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_70_io_in_0),
    .io_in_1(c53_70_io_in_1),
    .io_in_2(c53_70_io_in_2),
    .io_in_3(c53_70_io_in_3),
    .io_in_4(c53_70_io_in_4),
    .io_out_0(c53_70_io_out_0),
    .io_out_1(c53_70_io_out_1),
    .io_out_2(c53_70_io_out_2)
  );
  C53 c53_71 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_71_io_in_0),
    .io_in_1(c53_71_io_in_1),
    .io_in_2(c53_71_io_in_2),
    .io_in_3(c53_71_io_in_3),
    .io_in_4(c53_71_io_in_4),
    .io_out_0(c53_71_io_out_0),
    .io_out_1(c53_71_io_out_1),
    .io_out_2(c53_71_io_out_2)
  );
  C22 c22_9 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_9_io_in_0),
    .io_in_1(c22_9_io_in_1),
    .io_out_0(c22_9_io_out_0),
    .io_out_1(c22_9_io_out_1)
  );
  C53 c53_72 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_72_io_in_0),
    .io_in_1(c53_72_io_in_1),
    .io_in_2(c53_72_io_in_2),
    .io_in_3(c53_72_io_in_3),
    .io_in_4(c53_72_io_in_4),
    .io_out_0(c53_72_io_out_0),
    .io_out_1(c53_72_io_out_1),
    .io_out_2(c53_72_io_out_2)
  );
  C53 c53_73 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_73_io_in_0),
    .io_in_1(c53_73_io_in_1),
    .io_in_2(c53_73_io_in_2),
    .io_in_3(c53_73_io_in_3),
    .io_in_4(c53_73_io_in_4),
    .io_out_0(c53_73_io_out_0),
    .io_out_1(c53_73_io_out_1),
    .io_out_2(c53_73_io_out_2)
  );
  C53 c53_74 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_74_io_in_0),
    .io_in_1(c53_74_io_in_1),
    .io_in_2(c53_74_io_in_2),
    .io_in_3(c53_74_io_in_3),
    .io_in_4(c53_74_io_in_4),
    .io_out_0(c53_74_io_out_0),
    .io_out_1(c53_74_io_out_1),
    .io_out_2(c53_74_io_out_2)
  );
  C53 c53_75 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_75_io_in_0),
    .io_in_1(c53_75_io_in_1),
    .io_in_2(c53_75_io_in_2),
    .io_in_3(c53_75_io_in_3),
    .io_in_4(c53_75_io_in_4),
    .io_out_0(c53_75_io_out_0),
    .io_out_1(c53_75_io_out_1),
    .io_out_2(c53_75_io_out_2)
  );
  C32 c32_8 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_8_io_in_0),
    .io_in_1(c32_8_io_in_1),
    .io_in_2(c32_8_io_in_2),
    .io_out_0(c32_8_io_out_0),
    .io_out_1(c32_8_io_out_1)
  );
  C53 c53_76 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_76_io_in_0),
    .io_in_1(c53_76_io_in_1),
    .io_in_2(c53_76_io_in_2),
    .io_in_3(c53_76_io_in_3),
    .io_in_4(c53_76_io_in_4),
    .io_out_0(c53_76_io_out_0),
    .io_out_1(c53_76_io_out_1),
    .io_out_2(c53_76_io_out_2)
  );
  C53 c53_77 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_77_io_in_0),
    .io_in_1(c53_77_io_in_1),
    .io_in_2(c53_77_io_in_2),
    .io_in_3(c53_77_io_in_3),
    .io_in_4(c53_77_io_in_4),
    .io_out_0(c53_77_io_out_0),
    .io_out_1(c53_77_io_out_1),
    .io_out_2(c53_77_io_out_2)
  );
  C53 c53_78 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_78_io_in_0),
    .io_in_1(c53_78_io_in_1),
    .io_in_2(c53_78_io_in_2),
    .io_in_3(c53_78_io_in_3),
    .io_in_4(c53_78_io_in_4),
    .io_out_0(c53_78_io_out_0),
    .io_out_1(c53_78_io_out_1),
    .io_out_2(c53_78_io_out_2)
  );
  C53 c53_79 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_79_io_in_0),
    .io_in_1(c53_79_io_in_1),
    .io_in_2(c53_79_io_in_2),
    .io_in_3(c53_79_io_in_3),
    .io_in_4(c53_79_io_in_4),
    .io_out_0(c53_79_io_out_0),
    .io_out_1(c53_79_io_out_1),
    .io_out_2(c53_79_io_out_2)
  );
  C32 c32_9 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_9_io_in_0),
    .io_in_1(c32_9_io_in_1),
    .io_in_2(c32_9_io_in_2),
    .io_out_0(c32_9_io_out_0),
    .io_out_1(c32_9_io_out_1)
  );
  C53 c53_80 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_80_io_in_0),
    .io_in_1(c53_80_io_in_1),
    .io_in_2(c53_80_io_in_2),
    .io_in_3(c53_80_io_in_3),
    .io_in_4(c53_80_io_in_4),
    .io_out_0(c53_80_io_out_0),
    .io_out_1(c53_80_io_out_1),
    .io_out_2(c53_80_io_out_2)
  );
  C53 c53_81 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_81_io_in_0),
    .io_in_1(c53_81_io_in_1),
    .io_in_2(c53_81_io_in_2),
    .io_in_3(c53_81_io_in_3),
    .io_in_4(c53_81_io_in_4),
    .io_out_0(c53_81_io_out_0),
    .io_out_1(c53_81_io_out_1),
    .io_out_2(c53_81_io_out_2)
  );
  C53 c53_82 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_82_io_in_0),
    .io_in_1(c53_82_io_in_1),
    .io_in_2(c53_82_io_in_2),
    .io_in_3(c53_82_io_in_3),
    .io_in_4(c53_82_io_in_4),
    .io_out_0(c53_82_io_out_0),
    .io_out_1(c53_82_io_out_1),
    .io_out_2(c53_82_io_out_2)
  );
  C53 c53_83 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_83_io_in_0),
    .io_in_1(c53_83_io_in_1),
    .io_in_2(c53_83_io_in_2),
    .io_in_3(c53_83_io_in_3),
    .io_in_4(c53_83_io_in_4),
    .io_out_0(c53_83_io_out_0),
    .io_out_1(c53_83_io_out_1),
    .io_out_2(c53_83_io_out_2)
  );
  C53 c53_84 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_84_io_in_0),
    .io_in_1(c53_84_io_in_1),
    .io_in_2(c53_84_io_in_2),
    .io_in_3(c53_84_io_in_3),
    .io_in_4(c53_84_io_in_4),
    .io_out_0(c53_84_io_out_0),
    .io_out_1(c53_84_io_out_1),
    .io_out_2(c53_84_io_out_2)
  );
  C53 c53_85 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_85_io_in_0),
    .io_in_1(c53_85_io_in_1),
    .io_in_2(c53_85_io_in_2),
    .io_in_3(c53_85_io_in_3),
    .io_in_4(c53_85_io_in_4),
    .io_out_0(c53_85_io_out_0),
    .io_out_1(c53_85_io_out_1),
    .io_out_2(c53_85_io_out_2)
  );
  C53 c53_86 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_86_io_in_0),
    .io_in_1(c53_86_io_in_1),
    .io_in_2(c53_86_io_in_2),
    .io_in_3(c53_86_io_in_3),
    .io_in_4(c53_86_io_in_4),
    .io_out_0(c53_86_io_out_0),
    .io_out_1(c53_86_io_out_1),
    .io_out_2(c53_86_io_out_2)
  );
  C53 c53_87 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_87_io_in_0),
    .io_in_1(c53_87_io_in_1),
    .io_in_2(c53_87_io_in_2),
    .io_in_3(c53_87_io_in_3),
    .io_in_4(c53_87_io_in_4),
    .io_out_0(c53_87_io_out_0),
    .io_out_1(c53_87_io_out_1),
    .io_out_2(c53_87_io_out_2)
  );
  C53 c53_88 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_88_io_in_0),
    .io_in_1(c53_88_io_in_1),
    .io_in_2(c53_88_io_in_2),
    .io_in_3(c53_88_io_in_3),
    .io_in_4(c53_88_io_in_4),
    .io_out_0(c53_88_io_out_0),
    .io_out_1(c53_88_io_out_1),
    .io_out_2(c53_88_io_out_2)
  );
  C53 c53_89 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_89_io_in_0),
    .io_in_1(c53_89_io_in_1),
    .io_in_2(c53_89_io_in_2),
    .io_in_3(c53_89_io_in_3),
    .io_in_4(c53_89_io_in_4),
    .io_out_0(c53_89_io_out_0),
    .io_out_1(c53_89_io_out_1),
    .io_out_2(c53_89_io_out_2)
  );
  C53 c53_90 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_90_io_in_0),
    .io_in_1(c53_90_io_in_1),
    .io_in_2(c53_90_io_in_2),
    .io_in_3(c53_90_io_in_3),
    .io_in_4(c53_90_io_in_4),
    .io_out_0(c53_90_io_out_0),
    .io_out_1(c53_90_io_out_1),
    .io_out_2(c53_90_io_out_2)
  );
  C53 c53_91 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_91_io_in_0),
    .io_in_1(c53_91_io_in_1),
    .io_in_2(c53_91_io_in_2),
    .io_in_3(c53_91_io_in_3),
    .io_in_4(c53_91_io_in_4),
    .io_out_0(c53_91_io_out_0),
    .io_out_1(c53_91_io_out_1),
    .io_out_2(c53_91_io_out_2)
  );
  C53 c53_92 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_92_io_in_0),
    .io_in_1(c53_92_io_in_1),
    .io_in_2(c53_92_io_in_2),
    .io_in_3(c53_92_io_in_3),
    .io_in_4(c53_92_io_in_4),
    .io_out_0(c53_92_io_out_0),
    .io_out_1(c53_92_io_out_1),
    .io_out_2(c53_92_io_out_2)
  );
  C53 c53_93 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_93_io_in_0),
    .io_in_1(c53_93_io_in_1),
    .io_in_2(c53_93_io_in_2),
    .io_in_3(c53_93_io_in_3),
    .io_in_4(c53_93_io_in_4),
    .io_out_0(c53_93_io_out_0),
    .io_out_1(c53_93_io_out_1),
    .io_out_2(c53_93_io_out_2)
  );
  C53 c53_94 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_94_io_in_0),
    .io_in_1(c53_94_io_in_1),
    .io_in_2(c53_94_io_in_2),
    .io_in_3(c53_94_io_in_3),
    .io_in_4(c53_94_io_in_4),
    .io_out_0(c53_94_io_out_0),
    .io_out_1(c53_94_io_out_1),
    .io_out_2(c53_94_io_out_2)
  );
  C53 c53_95 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_95_io_in_0),
    .io_in_1(c53_95_io_in_1),
    .io_in_2(c53_95_io_in_2),
    .io_in_3(c53_95_io_in_3),
    .io_in_4(c53_95_io_in_4),
    .io_out_0(c53_95_io_out_0),
    .io_out_1(c53_95_io_out_1),
    .io_out_2(c53_95_io_out_2)
  );
  C53 c53_96 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_96_io_in_0),
    .io_in_1(c53_96_io_in_1),
    .io_in_2(c53_96_io_in_2),
    .io_in_3(c53_96_io_in_3),
    .io_in_4(c53_96_io_in_4),
    .io_out_0(c53_96_io_out_0),
    .io_out_1(c53_96_io_out_1),
    .io_out_2(c53_96_io_out_2)
  );
  C53 c53_97 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_97_io_in_0),
    .io_in_1(c53_97_io_in_1),
    .io_in_2(c53_97_io_in_2),
    .io_in_3(c53_97_io_in_3),
    .io_in_4(c53_97_io_in_4),
    .io_out_0(c53_97_io_out_0),
    .io_out_1(c53_97_io_out_1),
    .io_out_2(c53_97_io_out_2)
  );
  C53 c53_98 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_98_io_in_0),
    .io_in_1(c53_98_io_in_1),
    .io_in_2(c53_98_io_in_2),
    .io_in_3(c53_98_io_in_3),
    .io_in_4(c53_98_io_in_4),
    .io_out_0(c53_98_io_out_0),
    .io_out_1(c53_98_io_out_1),
    .io_out_2(c53_98_io_out_2)
  );
  C53 c53_99 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_99_io_in_0),
    .io_in_1(c53_99_io_in_1),
    .io_in_2(c53_99_io_in_2),
    .io_in_3(c53_99_io_in_3),
    .io_in_4(c53_99_io_in_4),
    .io_out_0(c53_99_io_out_0),
    .io_out_1(c53_99_io_out_1),
    .io_out_2(c53_99_io_out_2)
  );
  C53 c53_100 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_100_io_in_0),
    .io_in_1(c53_100_io_in_1),
    .io_in_2(c53_100_io_in_2),
    .io_in_3(c53_100_io_in_3),
    .io_in_4(c53_100_io_in_4),
    .io_out_0(c53_100_io_out_0),
    .io_out_1(c53_100_io_out_1),
    .io_out_2(c53_100_io_out_2)
  );
  C53 c53_101 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_101_io_in_0),
    .io_in_1(c53_101_io_in_1),
    .io_in_2(c53_101_io_in_2),
    .io_in_3(c53_101_io_in_3),
    .io_in_4(c53_101_io_in_4),
    .io_out_0(c53_101_io_out_0),
    .io_out_1(c53_101_io_out_1),
    .io_out_2(c53_101_io_out_2)
  );
  C53 c53_102 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_102_io_in_0),
    .io_in_1(c53_102_io_in_1),
    .io_in_2(c53_102_io_in_2),
    .io_in_3(c53_102_io_in_3),
    .io_in_4(c53_102_io_in_4),
    .io_out_0(c53_102_io_out_0),
    .io_out_1(c53_102_io_out_1),
    .io_out_2(c53_102_io_out_2)
  );
  C53 c53_103 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_103_io_in_0),
    .io_in_1(c53_103_io_in_1),
    .io_in_2(c53_103_io_in_2),
    .io_in_3(c53_103_io_in_3),
    .io_in_4(c53_103_io_in_4),
    .io_out_0(c53_103_io_out_0),
    .io_out_1(c53_103_io_out_1),
    .io_out_2(c53_103_io_out_2)
  );
  C53 c53_104 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_104_io_in_0),
    .io_in_1(c53_104_io_in_1),
    .io_in_2(c53_104_io_in_2),
    .io_in_3(c53_104_io_in_3),
    .io_in_4(c53_104_io_in_4),
    .io_out_0(c53_104_io_out_0),
    .io_out_1(c53_104_io_out_1),
    .io_out_2(c53_104_io_out_2)
  );
  C22 c22_10 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_10_io_in_0),
    .io_in_1(c22_10_io_in_1),
    .io_out_0(c22_10_io_out_0),
    .io_out_1(c22_10_io_out_1)
  );
  C53 c53_105 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_105_io_in_0),
    .io_in_1(c53_105_io_in_1),
    .io_in_2(c53_105_io_in_2),
    .io_in_3(c53_105_io_in_3),
    .io_in_4(c53_105_io_in_4),
    .io_out_0(c53_105_io_out_0),
    .io_out_1(c53_105_io_out_1),
    .io_out_2(c53_105_io_out_2)
  );
  C53 c53_106 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_106_io_in_0),
    .io_in_1(c53_106_io_in_1),
    .io_in_2(c53_106_io_in_2),
    .io_in_3(c53_106_io_in_3),
    .io_in_4(c53_106_io_in_4),
    .io_out_0(c53_106_io_out_0),
    .io_out_1(c53_106_io_out_1),
    .io_out_2(c53_106_io_out_2)
  );
  C53 c53_107 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_107_io_in_0),
    .io_in_1(c53_107_io_in_1),
    .io_in_2(c53_107_io_in_2),
    .io_in_3(c53_107_io_in_3),
    .io_in_4(c53_107_io_in_4),
    .io_out_0(c53_107_io_out_0),
    .io_out_1(c53_107_io_out_1),
    .io_out_2(c53_107_io_out_2)
  );
  C53 c53_108 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_108_io_in_0),
    .io_in_1(c53_108_io_in_1),
    .io_in_2(c53_108_io_in_2),
    .io_in_3(c53_108_io_in_3),
    .io_in_4(c53_108_io_in_4),
    .io_out_0(c53_108_io_out_0),
    .io_out_1(c53_108_io_out_1),
    .io_out_2(c53_108_io_out_2)
  );
  C53 c53_109 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_109_io_in_0),
    .io_in_1(c53_109_io_in_1),
    .io_in_2(c53_109_io_in_2),
    .io_in_3(c53_109_io_in_3),
    .io_in_4(c53_109_io_in_4),
    .io_out_0(c53_109_io_out_0),
    .io_out_1(c53_109_io_out_1),
    .io_out_2(c53_109_io_out_2)
  );
  C22 c22_11 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_11_io_in_0),
    .io_in_1(c22_11_io_in_1),
    .io_out_0(c22_11_io_out_0),
    .io_out_1(c22_11_io_out_1)
  );
  C53 c53_110 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_110_io_in_0),
    .io_in_1(c53_110_io_in_1),
    .io_in_2(c53_110_io_in_2),
    .io_in_3(c53_110_io_in_3),
    .io_in_4(c53_110_io_in_4),
    .io_out_0(c53_110_io_out_0),
    .io_out_1(c53_110_io_out_1),
    .io_out_2(c53_110_io_out_2)
  );
  C53 c53_111 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_111_io_in_0),
    .io_in_1(c53_111_io_in_1),
    .io_in_2(c53_111_io_in_2),
    .io_in_3(c53_111_io_in_3),
    .io_in_4(c53_111_io_in_4),
    .io_out_0(c53_111_io_out_0),
    .io_out_1(c53_111_io_out_1),
    .io_out_2(c53_111_io_out_2)
  );
  C53 c53_112 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_112_io_in_0),
    .io_in_1(c53_112_io_in_1),
    .io_in_2(c53_112_io_in_2),
    .io_in_3(c53_112_io_in_3),
    .io_in_4(c53_112_io_in_4),
    .io_out_0(c53_112_io_out_0),
    .io_out_1(c53_112_io_out_1),
    .io_out_2(c53_112_io_out_2)
  );
  C53 c53_113 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_113_io_in_0),
    .io_in_1(c53_113_io_in_1),
    .io_in_2(c53_113_io_in_2),
    .io_in_3(c53_113_io_in_3),
    .io_in_4(c53_113_io_in_4),
    .io_out_0(c53_113_io_out_0),
    .io_out_1(c53_113_io_out_1),
    .io_out_2(c53_113_io_out_2)
  );
  C53 c53_114 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_114_io_in_0),
    .io_in_1(c53_114_io_in_1),
    .io_in_2(c53_114_io_in_2),
    .io_in_3(c53_114_io_in_3),
    .io_in_4(c53_114_io_in_4),
    .io_out_0(c53_114_io_out_0),
    .io_out_1(c53_114_io_out_1),
    .io_out_2(c53_114_io_out_2)
  );
  C32 c32_10 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_10_io_in_0),
    .io_in_1(c32_10_io_in_1),
    .io_in_2(c32_10_io_in_2),
    .io_out_0(c32_10_io_out_0),
    .io_out_1(c32_10_io_out_1)
  );
  C53 c53_115 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_115_io_in_0),
    .io_in_1(c53_115_io_in_1),
    .io_in_2(c53_115_io_in_2),
    .io_in_3(c53_115_io_in_3),
    .io_in_4(c53_115_io_in_4),
    .io_out_0(c53_115_io_out_0),
    .io_out_1(c53_115_io_out_1),
    .io_out_2(c53_115_io_out_2)
  );
  C53 c53_116 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_116_io_in_0),
    .io_in_1(c53_116_io_in_1),
    .io_in_2(c53_116_io_in_2),
    .io_in_3(c53_116_io_in_3),
    .io_in_4(c53_116_io_in_4),
    .io_out_0(c53_116_io_out_0),
    .io_out_1(c53_116_io_out_1),
    .io_out_2(c53_116_io_out_2)
  );
  C53 c53_117 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_117_io_in_0),
    .io_in_1(c53_117_io_in_1),
    .io_in_2(c53_117_io_in_2),
    .io_in_3(c53_117_io_in_3),
    .io_in_4(c53_117_io_in_4),
    .io_out_0(c53_117_io_out_0),
    .io_out_1(c53_117_io_out_1),
    .io_out_2(c53_117_io_out_2)
  );
  C53 c53_118 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_118_io_in_0),
    .io_in_1(c53_118_io_in_1),
    .io_in_2(c53_118_io_in_2),
    .io_in_3(c53_118_io_in_3),
    .io_in_4(c53_118_io_in_4),
    .io_out_0(c53_118_io_out_0),
    .io_out_1(c53_118_io_out_1),
    .io_out_2(c53_118_io_out_2)
  );
  C53 c53_119 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_119_io_in_0),
    .io_in_1(c53_119_io_in_1),
    .io_in_2(c53_119_io_in_2),
    .io_in_3(c53_119_io_in_3),
    .io_in_4(c53_119_io_in_4),
    .io_out_0(c53_119_io_out_0),
    .io_out_1(c53_119_io_out_1),
    .io_out_2(c53_119_io_out_2)
  );
  C32 c32_11 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_11_io_in_0),
    .io_in_1(c32_11_io_in_1),
    .io_in_2(c32_11_io_in_2),
    .io_out_0(c32_11_io_out_0),
    .io_out_1(c32_11_io_out_1)
  );
  C53 c53_120 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_120_io_in_0),
    .io_in_1(c53_120_io_in_1),
    .io_in_2(c53_120_io_in_2),
    .io_in_3(c53_120_io_in_3),
    .io_in_4(c53_120_io_in_4),
    .io_out_0(c53_120_io_out_0),
    .io_out_1(c53_120_io_out_1),
    .io_out_2(c53_120_io_out_2)
  );
  C53 c53_121 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_121_io_in_0),
    .io_in_1(c53_121_io_in_1),
    .io_in_2(c53_121_io_in_2),
    .io_in_3(c53_121_io_in_3),
    .io_in_4(c53_121_io_in_4),
    .io_out_0(c53_121_io_out_0),
    .io_out_1(c53_121_io_out_1),
    .io_out_2(c53_121_io_out_2)
  );
  C53 c53_122 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_122_io_in_0),
    .io_in_1(c53_122_io_in_1),
    .io_in_2(c53_122_io_in_2),
    .io_in_3(c53_122_io_in_3),
    .io_in_4(c53_122_io_in_4),
    .io_out_0(c53_122_io_out_0),
    .io_out_1(c53_122_io_out_1),
    .io_out_2(c53_122_io_out_2)
  );
  C53 c53_123 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_123_io_in_0),
    .io_in_1(c53_123_io_in_1),
    .io_in_2(c53_123_io_in_2),
    .io_in_3(c53_123_io_in_3),
    .io_in_4(c53_123_io_in_4),
    .io_out_0(c53_123_io_out_0),
    .io_out_1(c53_123_io_out_1),
    .io_out_2(c53_123_io_out_2)
  );
  C53 c53_124 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_124_io_in_0),
    .io_in_1(c53_124_io_in_1),
    .io_in_2(c53_124_io_in_2),
    .io_in_3(c53_124_io_in_3),
    .io_in_4(c53_124_io_in_4),
    .io_out_0(c53_124_io_out_0),
    .io_out_1(c53_124_io_out_1),
    .io_out_2(c53_124_io_out_2)
  );
  C53 c53_125 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_125_io_in_0),
    .io_in_1(c53_125_io_in_1),
    .io_in_2(c53_125_io_in_2),
    .io_in_3(c53_125_io_in_3),
    .io_in_4(c53_125_io_in_4),
    .io_out_0(c53_125_io_out_0),
    .io_out_1(c53_125_io_out_1),
    .io_out_2(c53_125_io_out_2)
  );
  C53 c53_126 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_126_io_in_0),
    .io_in_1(c53_126_io_in_1),
    .io_in_2(c53_126_io_in_2),
    .io_in_3(c53_126_io_in_3),
    .io_in_4(c53_126_io_in_4),
    .io_out_0(c53_126_io_out_0),
    .io_out_1(c53_126_io_out_1),
    .io_out_2(c53_126_io_out_2)
  );
  C53 c53_127 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_127_io_in_0),
    .io_in_1(c53_127_io_in_1),
    .io_in_2(c53_127_io_in_2),
    .io_in_3(c53_127_io_in_3),
    .io_in_4(c53_127_io_in_4),
    .io_out_0(c53_127_io_out_0),
    .io_out_1(c53_127_io_out_1),
    .io_out_2(c53_127_io_out_2)
  );
  C53 c53_128 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_128_io_in_0),
    .io_in_1(c53_128_io_in_1),
    .io_in_2(c53_128_io_in_2),
    .io_in_3(c53_128_io_in_3),
    .io_in_4(c53_128_io_in_4),
    .io_out_0(c53_128_io_out_0),
    .io_out_1(c53_128_io_out_1),
    .io_out_2(c53_128_io_out_2)
  );
  C53 c53_129 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_129_io_in_0),
    .io_in_1(c53_129_io_in_1),
    .io_in_2(c53_129_io_in_2),
    .io_in_3(c53_129_io_in_3),
    .io_in_4(c53_129_io_in_4),
    .io_out_0(c53_129_io_out_0),
    .io_out_1(c53_129_io_out_1),
    .io_out_2(c53_129_io_out_2)
  );
  C53 c53_130 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_130_io_in_0),
    .io_in_1(c53_130_io_in_1),
    .io_in_2(c53_130_io_in_2),
    .io_in_3(c53_130_io_in_3),
    .io_in_4(c53_130_io_in_4),
    .io_out_0(c53_130_io_out_0),
    .io_out_1(c53_130_io_out_1),
    .io_out_2(c53_130_io_out_2)
  );
  C53 c53_131 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_131_io_in_0),
    .io_in_1(c53_131_io_in_1),
    .io_in_2(c53_131_io_in_2),
    .io_in_3(c53_131_io_in_3),
    .io_in_4(c53_131_io_in_4),
    .io_out_0(c53_131_io_out_0),
    .io_out_1(c53_131_io_out_1),
    .io_out_2(c53_131_io_out_2)
  );
  C53 c53_132 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_132_io_in_0),
    .io_in_1(c53_132_io_in_1),
    .io_in_2(c53_132_io_in_2),
    .io_in_3(c53_132_io_in_3),
    .io_in_4(c53_132_io_in_4),
    .io_out_0(c53_132_io_out_0),
    .io_out_1(c53_132_io_out_1),
    .io_out_2(c53_132_io_out_2)
  );
  C53 c53_133 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_133_io_in_0),
    .io_in_1(c53_133_io_in_1),
    .io_in_2(c53_133_io_in_2),
    .io_in_3(c53_133_io_in_3),
    .io_in_4(c53_133_io_in_4),
    .io_out_0(c53_133_io_out_0),
    .io_out_1(c53_133_io_out_1),
    .io_out_2(c53_133_io_out_2)
  );
  C53 c53_134 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_134_io_in_0),
    .io_in_1(c53_134_io_in_1),
    .io_in_2(c53_134_io_in_2),
    .io_in_3(c53_134_io_in_3),
    .io_in_4(c53_134_io_in_4),
    .io_out_0(c53_134_io_out_0),
    .io_out_1(c53_134_io_out_1),
    .io_out_2(c53_134_io_out_2)
  );
  C53 c53_135 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_135_io_in_0),
    .io_in_1(c53_135_io_in_1),
    .io_in_2(c53_135_io_in_2),
    .io_in_3(c53_135_io_in_3),
    .io_in_4(c53_135_io_in_4),
    .io_out_0(c53_135_io_out_0),
    .io_out_1(c53_135_io_out_1),
    .io_out_2(c53_135_io_out_2)
  );
  C53 c53_136 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_136_io_in_0),
    .io_in_1(c53_136_io_in_1),
    .io_in_2(c53_136_io_in_2),
    .io_in_3(c53_136_io_in_3),
    .io_in_4(c53_136_io_in_4),
    .io_out_0(c53_136_io_out_0),
    .io_out_1(c53_136_io_out_1),
    .io_out_2(c53_136_io_out_2)
  );
  C53 c53_137 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_137_io_in_0),
    .io_in_1(c53_137_io_in_1),
    .io_in_2(c53_137_io_in_2),
    .io_in_3(c53_137_io_in_3),
    .io_in_4(c53_137_io_in_4),
    .io_out_0(c53_137_io_out_0),
    .io_out_1(c53_137_io_out_1),
    .io_out_2(c53_137_io_out_2)
  );
  C53 c53_138 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_138_io_in_0),
    .io_in_1(c53_138_io_in_1),
    .io_in_2(c53_138_io_in_2),
    .io_in_3(c53_138_io_in_3),
    .io_in_4(c53_138_io_in_4),
    .io_out_0(c53_138_io_out_0),
    .io_out_1(c53_138_io_out_1),
    .io_out_2(c53_138_io_out_2)
  );
  C53 c53_139 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_139_io_in_0),
    .io_in_1(c53_139_io_in_1),
    .io_in_2(c53_139_io_in_2),
    .io_in_3(c53_139_io_in_3),
    .io_in_4(c53_139_io_in_4),
    .io_out_0(c53_139_io_out_0),
    .io_out_1(c53_139_io_out_1),
    .io_out_2(c53_139_io_out_2)
  );
  C53 c53_140 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_140_io_in_0),
    .io_in_1(c53_140_io_in_1),
    .io_in_2(c53_140_io_in_2),
    .io_in_3(c53_140_io_in_3),
    .io_in_4(c53_140_io_in_4),
    .io_out_0(c53_140_io_out_0),
    .io_out_1(c53_140_io_out_1),
    .io_out_2(c53_140_io_out_2)
  );
  C53 c53_141 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_141_io_in_0),
    .io_in_1(c53_141_io_in_1),
    .io_in_2(c53_141_io_in_2),
    .io_in_3(c53_141_io_in_3),
    .io_in_4(c53_141_io_in_4),
    .io_out_0(c53_141_io_out_0),
    .io_out_1(c53_141_io_out_1),
    .io_out_2(c53_141_io_out_2)
  );
  C53 c53_142 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_142_io_in_0),
    .io_in_1(c53_142_io_in_1),
    .io_in_2(c53_142_io_in_2),
    .io_in_3(c53_142_io_in_3),
    .io_in_4(c53_142_io_in_4),
    .io_out_0(c53_142_io_out_0),
    .io_out_1(c53_142_io_out_1),
    .io_out_2(c53_142_io_out_2)
  );
  C53 c53_143 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_143_io_in_0),
    .io_in_1(c53_143_io_in_1),
    .io_in_2(c53_143_io_in_2),
    .io_in_3(c53_143_io_in_3),
    .io_in_4(c53_143_io_in_4),
    .io_out_0(c53_143_io_out_0),
    .io_out_1(c53_143_io_out_1),
    .io_out_2(c53_143_io_out_2)
  );
  C53 c53_144 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_144_io_in_0),
    .io_in_1(c53_144_io_in_1),
    .io_in_2(c53_144_io_in_2),
    .io_in_3(c53_144_io_in_3),
    .io_in_4(c53_144_io_in_4),
    .io_out_0(c53_144_io_out_0),
    .io_out_1(c53_144_io_out_1),
    .io_out_2(c53_144_io_out_2)
  );
  C53 c53_145 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_145_io_in_0),
    .io_in_1(c53_145_io_in_1),
    .io_in_2(c53_145_io_in_2),
    .io_in_3(c53_145_io_in_3),
    .io_in_4(c53_145_io_in_4),
    .io_out_0(c53_145_io_out_0),
    .io_out_1(c53_145_io_out_1),
    .io_out_2(c53_145_io_out_2)
  );
  C53 c53_146 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_146_io_in_0),
    .io_in_1(c53_146_io_in_1),
    .io_in_2(c53_146_io_in_2),
    .io_in_3(c53_146_io_in_3),
    .io_in_4(c53_146_io_in_4),
    .io_out_0(c53_146_io_out_0),
    .io_out_1(c53_146_io_out_1),
    .io_out_2(c53_146_io_out_2)
  );
  C53 c53_147 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_147_io_in_0),
    .io_in_1(c53_147_io_in_1),
    .io_in_2(c53_147_io_in_2),
    .io_in_3(c53_147_io_in_3),
    .io_in_4(c53_147_io_in_4),
    .io_out_0(c53_147_io_out_0),
    .io_out_1(c53_147_io_out_1),
    .io_out_2(c53_147_io_out_2)
  );
  C53 c53_148 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_148_io_in_0),
    .io_in_1(c53_148_io_in_1),
    .io_in_2(c53_148_io_in_2),
    .io_in_3(c53_148_io_in_3),
    .io_in_4(c53_148_io_in_4),
    .io_out_0(c53_148_io_out_0),
    .io_out_1(c53_148_io_out_1),
    .io_out_2(c53_148_io_out_2)
  );
  C53 c53_149 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_149_io_in_0),
    .io_in_1(c53_149_io_in_1),
    .io_in_2(c53_149_io_in_2),
    .io_in_3(c53_149_io_in_3),
    .io_in_4(c53_149_io_in_4),
    .io_out_0(c53_149_io_out_0),
    .io_out_1(c53_149_io_out_1),
    .io_out_2(c53_149_io_out_2)
  );
  C22 c22_12 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_12_io_in_0),
    .io_in_1(c22_12_io_in_1),
    .io_out_0(c22_12_io_out_0),
    .io_out_1(c22_12_io_out_1)
  );
  C53 c53_150 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_150_io_in_0),
    .io_in_1(c53_150_io_in_1),
    .io_in_2(c53_150_io_in_2),
    .io_in_3(c53_150_io_in_3),
    .io_in_4(c53_150_io_in_4),
    .io_out_0(c53_150_io_out_0),
    .io_out_1(c53_150_io_out_1),
    .io_out_2(c53_150_io_out_2)
  );
  C53 c53_151 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_151_io_in_0),
    .io_in_1(c53_151_io_in_1),
    .io_in_2(c53_151_io_in_2),
    .io_in_3(c53_151_io_in_3),
    .io_in_4(c53_151_io_in_4),
    .io_out_0(c53_151_io_out_0),
    .io_out_1(c53_151_io_out_1),
    .io_out_2(c53_151_io_out_2)
  );
  C53 c53_152 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_152_io_in_0),
    .io_in_1(c53_152_io_in_1),
    .io_in_2(c53_152_io_in_2),
    .io_in_3(c53_152_io_in_3),
    .io_in_4(c53_152_io_in_4),
    .io_out_0(c53_152_io_out_0),
    .io_out_1(c53_152_io_out_1),
    .io_out_2(c53_152_io_out_2)
  );
  C53 c53_153 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_153_io_in_0),
    .io_in_1(c53_153_io_in_1),
    .io_in_2(c53_153_io_in_2),
    .io_in_3(c53_153_io_in_3),
    .io_in_4(c53_153_io_in_4),
    .io_out_0(c53_153_io_out_0),
    .io_out_1(c53_153_io_out_1),
    .io_out_2(c53_153_io_out_2)
  );
  C53 c53_154 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_154_io_in_0),
    .io_in_1(c53_154_io_in_1),
    .io_in_2(c53_154_io_in_2),
    .io_in_3(c53_154_io_in_3),
    .io_in_4(c53_154_io_in_4),
    .io_out_0(c53_154_io_out_0),
    .io_out_1(c53_154_io_out_1),
    .io_out_2(c53_154_io_out_2)
  );
  C53 c53_155 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_155_io_in_0),
    .io_in_1(c53_155_io_in_1),
    .io_in_2(c53_155_io_in_2),
    .io_in_3(c53_155_io_in_3),
    .io_in_4(c53_155_io_in_4),
    .io_out_0(c53_155_io_out_0),
    .io_out_1(c53_155_io_out_1),
    .io_out_2(c53_155_io_out_2)
  );
  C22 c22_13 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_13_io_in_0),
    .io_in_1(c22_13_io_in_1),
    .io_out_0(c22_13_io_out_0),
    .io_out_1(c22_13_io_out_1)
  );
  C53 c53_156 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_156_io_in_0),
    .io_in_1(c53_156_io_in_1),
    .io_in_2(c53_156_io_in_2),
    .io_in_3(c53_156_io_in_3),
    .io_in_4(c53_156_io_in_4),
    .io_out_0(c53_156_io_out_0),
    .io_out_1(c53_156_io_out_1),
    .io_out_2(c53_156_io_out_2)
  );
  C53 c53_157 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_157_io_in_0),
    .io_in_1(c53_157_io_in_1),
    .io_in_2(c53_157_io_in_2),
    .io_in_3(c53_157_io_in_3),
    .io_in_4(c53_157_io_in_4),
    .io_out_0(c53_157_io_out_0),
    .io_out_1(c53_157_io_out_1),
    .io_out_2(c53_157_io_out_2)
  );
  C53 c53_158 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_158_io_in_0),
    .io_in_1(c53_158_io_in_1),
    .io_in_2(c53_158_io_in_2),
    .io_in_3(c53_158_io_in_3),
    .io_in_4(c53_158_io_in_4),
    .io_out_0(c53_158_io_out_0),
    .io_out_1(c53_158_io_out_1),
    .io_out_2(c53_158_io_out_2)
  );
  C53 c53_159 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_159_io_in_0),
    .io_in_1(c53_159_io_in_1),
    .io_in_2(c53_159_io_in_2),
    .io_in_3(c53_159_io_in_3),
    .io_in_4(c53_159_io_in_4),
    .io_out_0(c53_159_io_out_0),
    .io_out_1(c53_159_io_out_1),
    .io_out_2(c53_159_io_out_2)
  );
  C53 c53_160 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_160_io_in_0),
    .io_in_1(c53_160_io_in_1),
    .io_in_2(c53_160_io_in_2),
    .io_in_3(c53_160_io_in_3),
    .io_in_4(c53_160_io_in_4),
    .io_out_0(c53_160_io_out_0),
    .io_out_1(c53_160_io_out_1),
    .io_out_2(c53_160_io_out_2)
  );
  C53 c53_161 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_161_io_in_0),
    .io_in_1(c53_161_io_in_1),
    .io_in_2(c53_161_io_in_2),
    .io_in_3(c53_161_io_in_3),
    .io_in_4(c53_161_io_in_4),
    .io_out_0(c53_161_io_out_0),
    .io_out_1(c53_161_io_out_1),
    .io_out_2(c53_161_io_out_2)
  );
  C32 c32_12 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_12_io_in_0),
    .io_in_1(c32_12_io_in_1),
    .io_in_2(c32_12_io_in_2),
    .io_out_0(c32_12_io_out_0),
    .io_out_1(c32_12_io_out_1)
  );
  C53 c53_162 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_162_io_in_0),
    .io_in_1(c53_162_io_in_1),
    .io_in_2(c53_162_io_in_2),
    .io_in_3(c53_162_io_in_3),
    .io_in_4(c53_162_io_in_4),
    .io_out_0(c53_162_io_out_0),
    .io_out_1(c53_162_io_out_1),
    .io_out_2(c53_162_io_out_2)
  );
  C53 c53_163 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_163_io_in_0),
    .io_in_1(c53_163_io_in_1),
    .io_in_2(c53_163_io_in_2),
    .io_in_3(c53_163_io_in_3),
    .io_in_4(c53_163_io_in_4),
    .io_out_0(c53_163_io_out_0),
    .io_out_1(c53_163_io_out_1),
    .io_out_2(c53_163_io_out_2)
  );
  C53 c53_164 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_164_io_in_0),
    .io_in_1(c53_164_io_in_1),
    .io_in_2(c53_164_io_in_2),
    .io_in_3(c53_164_io_in_3),
    .io_in_4(c53_164_io_in_4),
    .io_out_0(c53_164_io_out_0),
    .io_out_1(c53_164_io_out_1),
    .io_out_2(c53_164_io_out_2)
  );
  C53 c53_165 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_165_io_in_0),
    .io_in_1(c53_165_io_in_1),
    .io_in_2(c53_165_io_in_2),
    .io_in_3(c53_165_io_in_3),
    .io_in_4(c53_165_io_in_4),
    .io_out_0(c53_165_io_out_0),
    .io_out_1(c53_165_io_out_1),
    .io_out_2(c53_165_io_out_2)
  );
  C53 c53_166 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_166_io_in_0),
    .io_in_1(c53_166_io_in_1),
    .io_in_2(c53_166_io_in_2),
    .io_in_3(c53_166_io_in_3),
    .io_in_4(c53_166_io_in_4),
    .io_out_0(c53_166_io_out_0),
    .io_out_1(c53_166_io_out_1),
    .io_out_2(c53_166_io_out_2)
  );
  C53 c53_167 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_167_io_in_0),
    .io_in_1(c53_167_io_in_1),
    .io_in_2(c53_167_io_in_2),
    .io_in_3(c53_167_io_in_3),
    .io_in_4(c53_167_io_in_4),
    .io_out_0(c53_167_io_out_0),
    .io_out_1(c53_167_io_out_1),
    .io_out_2(c53_167_io_out_2)
  );
  C32 c32_13 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_13_io_in_0),
    .io_in_1(c32_13_io_in_1),
    .io_in_2(c32_13_io_in_2),
    .io_out_0(c32_13_io_out_0),
    .io_out_1(c32_13_io_out_1)
  );
  C53 c53_168 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_168_io_in_0),
    .io_in_1(c53_168_io_in_1),
    .io_in_2(c53_168_io_in_2),
    .io_in_3(c53_168_io_in_3),
    .io_in_4(c53_168_io_in_4),
    .io_out_0(c53_168_io_out_0),
    .io_out_1(c53_168_io_out_1),
    .io_out_2(c53_168_io_out_2)
  );
  C53 c53_169 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_169_io_in_0),
    .io_in_1(c53_169_io_in_1),
    .io_in_2(c53_169_io_in_2),
    .io_in_3(c53_169_io_in_3),
    .io_in_4(c53_169_io_in_4),
    .io_out_0(c53_169_io_out_0),
    .io_out_1(c53_169_io_out_1),
    .io_out_2(c53_169_io_out_2)
  );
  C53 c53_170 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_170_io_in_0),
    .io_in_1(c53_170_io_in_1),
    .io_in_2(c53_170_io_in_2),
    .io_in_3(c53_170_io_in_3),
    .io_in_4(c53_170_io_in_4),
    .io_out_0(c53_170_io_out_0),
    .io_out_1(c53_170_io_out_1),
    .io_out_2(c53_170_io_out_2)
  );
  C53 c53_171 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_171_io_in_0),
    .io_in_1(c53_171_io_in_1),
    .io_in_2(c53_171_io_in_2),
    .io_in_3(c53_171_io_in_3),
    .io_in_4(c53_171_io_in_4),
    .io_out_0(c53_171_io_out_0),
    .io_out_1(c53_171_io_out_1),
    .io_out_2(c53_171_io_out_2)
  );
  C53 c53_172 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_172_io_in_0),
    .io_in_1(c53_172_io_in_1),
    .io_in_2(c53_172_io_in_2),
    .io_in_3(c53_172_io_in_3),
    .io_in_4(c53_172_io_in_4),
    .io_out_0(c53_172_io_out_0),
    .io_out_1(c53_172_io_out_1),
    .io_out_2(c53_172_io_out_2)
  );
  C53 c53_173 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_173_io_in_0),
    .io_in_1(c53_173_io_in_1),
    .io_in_2(c53_173_io_in_2),
    .io_in_3(c53_173_io_in_3),
    .io_in_4(c53_173_io_in_4),
    .io_out_0(c53_173_io_out_0),
    .io_out_1(c53_173_io_out_1),
    .io_out_2(c53_173_io_out_2)
  );
  C53 c53_174 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_174_io_in_0),
    .io_in_1(c53_174_io_in_1),
    .io_in_2(c53_174_io_in_2),
    .io_in_3(c53_174_io_in_3),
    .io_in_4(c53_174_io_in_4),
    .io_out_0(c53_174_io_out_0),
    .io_out_1(c53_174_io_out_1),
    .io_out_2(c53_174_io_out_2)
  );
  C53 c53_175 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_175_io_in_0),
    .io_in_1(c53_175_io_in_1),
    .io_in_2(c53_175_io_in_2),
    .io_in_3(c53_175_io_in_3),
    .io_in_4(c53_175_io_in_4),
    .io_out_0(c53_175_io_out_0),
    .io_out_1(c53_175_io_out_1),
    .io_out_2(c53_175_io_out_2)
  );
  C53 c53_176 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_176_io_in_0),
    .io_in_1(c53_176_io_in_1),
    .io_in_2(c53_176_io_in_2),
    .io_in_3(c53_176_io_in_3),
    .io_in_4(c53_176_io_in_4),
    .io_out_0(c53_176_io_out_0),
    .io_out_1(c53_176_io_out_1),
    .io_out_2(c53_176_io_out_2)
  );
  C53 c53_177 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_177_io_in_0),
    .io_in_1(c53_177_io_in_1),
    .io_in_2(c53_177_io_in_2),
    .io_in_3(c53_177_io_in_3),
    .io_in_4(c53_177_io_in_4),
    .io_out_0(c53_177_io_out_0),
    .io_out_1(c53_177_io_out_1),
    .io_out_2(c53_177_io_out_2)
  );
  C53 c53_178 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_178_io_in_0),
    .io_in_1(c53_178_io_in_1),
    .io_in_2(c53_178_io_in_2),
    .io_in_3(c53_178_io_in_3),
    .io_in_4(c53_178_io_in_4),
    .io_out_0(c53_178_io_out_0),
    .io_out_1(c53_178_io_out_1),
    .io_out_2(c53_178_io_out_2)
  );
  C53 c53_179 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_179_io_in_0),
    .io_in_1(c53_179_io_in_1),
    .io_in_2(c53_179_io_in_2),
    .io_in_3(c53_179_io_in_3),
    .io_in_4(c53_179_io_in_4),
    .io_out_0(c53_179_io_out_0),
    .io_out_1(c53_179_io_out_1),
    .io_out_2(c53_179_io_out_2)
  );
  C53 c53_180 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_180_io_in_0),
    .io_in_1(c53_180_io_in_1),
    .io_in_2(c53_180_io_in_2),
    .io_in_3(c53_180_io_in_3),
    .io_in_4(c53_180_io_in_4),
    .io_out_0(c53_180_io_out_0),
    .io_out_1(c53_180_io_out_1),
    .io_out_2(c53_180_io_out_2)
  );
  C53 c53_181 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_181_io_in_0),
    .io_in_1(c53_181_io_in_1),
    .io_in_2(c53_181_io_in_2),
    .io_in_3(c53_181_io_in_3),
    .io_in_4(c53_181_io_in_4),
    .io_out_0(c53_181_io_out_0),
    .io_out_1(c53_181_io_out_1),
    .io_out_2(c53_181_io_out_2)
  );
  C53 c53_182 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_182_io_in_0),
    .io_in_1(c53_182_io_in_1),
    .io_in_2(c53_182_io_in_2),
    .io_in_3(c53_182_io_in_3),
    .io_in_4(c53_182_io_in_4),
    .io_out_0(c53_182_io_out_0),
    .io_out_1(c53_182_io_out_1),
    .io_out_2(c53_182_io_out_2)
  );
  C53 c53_183 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_183_io_in_0),
    .io_in_1(c53_183_io_in_1),
    .io_in_2(c53_183_io_in_2),
    .io_in_3(c53_183_io_in_3),
    .io_in_4(c53_183_io_in_4),
    .io_out_0(c53_183_io_out_0),
    .io_out_1(c53_183_io_out_1),
    .io_out_2(c53_183_io_out_2)
  );
  C53 c53_184 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_184_io_in_0),
    .io_in_1(c53_184_io_in_1),
    .io_in_2(c53_184_io_in_2),
    .io_in_3(c53_184_io_in_3),
    .io_in_4(c53_184_io_in_4),
    .io_out_0(c53_184_io_out_0),
    .io_out_1(c53_184_io_out_1),
    .io_out_2(c53_184_io_out_2)
  );
  C53 c53_185 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_185_io_in_0),
    .io_in_1(c53_185_io_in_1),
    .io_in_2(c53_185_io_in_2),
    .io_in_3(c53_185_io_in_3),
    .io_in_4(c53_185_io_in_4),
    .io_out_0(c53_185_io_out_0),
    .io_out_1(c53_185_io_out_1),
    .io_out_2(c53_185_io_out_2)
  );
  C53 c53_186 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_186_io_in_0),
    .io_in_1(c53_186_io_in_1),
    .io_in_2(c53_186_io_in_2),
    .io_in_3(c53_186_io_in_3),
    .io_in_4(c53_186_io_in_4),
    .io_out_0(c53_186_io_out_0),
    .io_out_1(c53_186_io_out_1),
    .io_out_2(c53_186_io_out_2)
  );
  C53 c53_187 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_187_io_in_0),
    .io_in_1(c53_187_io_in_1),
    .io_in_2(c53_187_io_in_2),
    .io_in_3(c53_187_io_in_3),
    .io_in_4(c53_187_io_in_4),
    .io_out_0(c53_187_io_out_0),
    .io_out_1(c53_187_io_out_1),
    .io_out_2(c53_187_io_out_2)
  );
  C53 c53_188 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_188_io_in_0),
    .io_in_1(c53_188_io_in_1),
    .io_in_2(c53_188_io_in_2),
    .io_in_3(c53_188_io_in_3),
    .io_in_4(c53_188_io_in_4),
    .io_out_0(c53_188_io_out_0),
    .io_out_1(c53_188_io_out_1),
    .io_out_2(c53_188_io_out_2)
  );
  C53 c53_189 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_189_io_in_0),
    .io_in_1(c53_189_io_in_1),
    .io_in_2(c53_189_io_in_2),
    .io_in_3(c53_189_io_in_3),
    .io_in_4(c53_189_io_in_4),
    .io_out_0(c53_189_io_out_0),
    .io_out_1(c53_189_io_out_1),
    .io_out_2(c53_189_io_out_2)
  );
  C53 c53_190 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_190_io_in_0),
    .io_in_1(c53_190_io_in_1),
    .io_in_2(c53_190_io_in_2),
    .io_in_3(c53_190_io_in_3),
    .io_in_4(c53_190_io_in_4),
    .io_out_0(c53_190_io_out_0),
    .io_out_1(c53_190_io_out_1),
    .io_out_2(c53_190_io_out_2)
  );
  C53 c53_191 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_191_io_in_0),
    .io_in_1(c53_191_io_in_1),
    .io_in_2(c53_191_io_in_2),
    .io_in_3(c53_191_io_in_3),
    .io_in_4(c53_191_io_in_4),
    .io_out_0(c53_191_io_out_0),
    .io_out_1(c53_191_io_out_1),
    .io_out_2(c53_191_io_out_2)
  );
  C53 c53_192 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_192_io_in_0),
    .io_in_1(c53_192_io_in_1),
    .io_in_2(c53_192_io_in_2),
    .io_in_3(c53_192_io_in_3),
    .io_in_4(c53_192_io_in_4),
    .io_out_0(c53_192_io_out_0),
    .io_out_1(c53_192_io_out_1),
    .io_out_2(c53_192_io_out_2)
  );
  C53 c53_193 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_193_io_in_0),
    .io_in_1(c53_193_io_in_1),
    .io_in_2(c53_193_io_in_2),
    .io_in_3(c53_193_io_in_3),
    .io_in_4(c53_193_io_in_4),
    .io_out_0(c53_193_io_out_0),
    .io_out_1(c53_193_io_out_1),
    .io_out_2(c53_193_io_out_2)
  );
  C53 c53_194 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_194_io_in_0),
    .io_in_1(c53_194_io_in_1),
    .io_in_2(c53_194_io_in_2),
    .io_in_3(c53_194_io_in_3),
    .io_in_4(c53_194_io_in_4),
    .io_out_0(c53_194_io_out_0),
    .io_out_1(c53_194_io_out_1),
    .io_out_2(c53_194_io_out_2)
  );
  C53 c53_195 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_195_io_in_0),
    .io_in_1(c53_195_io_in_1),
    .io_in_2(c53_195_io_in_2),
    .io_in_3(c53_195_io_in_3),
    .io_in_4(c53_195_io_in_4),
    .io_out_0(c53_195_io_out_0),
    .io_out_1(c53_195_io_out_1),
    .io_out_2(c53_195_io_out_2)
  );
  C53 c53_196 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_196_io_in_0),
    .io_in_1(c53_196_io_in_1),
    .io_in_2(c53_196_io_in_2),
    .io_in_3(c53_196_io_in_3),
    .io_in_4(c53_196_io_in_4),
    .io_out_0(c53_196_io_out_0),
    .io_out_1(c53_196_io_out_1),
    .io_out_2(c53_196_io_out_2)
  );
  C53 c53_197 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_197_io_in_0),
    .io_in_1(c53_197_io_in_1),
    .io_in_2(c53_197_io_in_2),
    .io_in_3(c53_197_io_in_3),
    .io_in_4(c53_197_io_in_4),
    .io_out_0(c53_197_io_out_0),
    .io_out_1(c53_197_io_out_1),
    .io_out_2(c53_197_io_out_2)
  );
  C53 c53_198 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_198_io_in_0),
    .io_in_1(c53_198_io_in_1),
    .io_in_2(c53_198_io_in_2),
    .io_in_3(c53_198_io_in_3),
    .io_in_4(c53_198_io_in_4),
    .io_out_0(c53_198_io_out_0),
    .io_out_1(c53_198_io_out_1),
    .io_out_2(c53_198_io_out_2)
  );
  C53 c53_199 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_199_io_in_0),
    .io_in_1(c53_199_io_in_1),
    .io_in_2(c53_199_io_in_2),
    .io_in_3(c53_199_io_in_3),
    .io_in_4(c53_199_io_in_4),
    .io_out_0(c53_199_io_out_0),
    .io_out_1(c53_199_io_out_1),
    .io_out_2(c53_199_io_out_2)
  );
  C53 c53_200 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_200_io_in_0),
    .io_in_1(c53_200_io_in_1),
    .io_in_2(c53_200_io_in_2),
    .io_in_3(c53_200_io_in_3),
    .io_in_4(c53_200_io_in_4),
    .io_out_0(c53_200_io_out_0),
    .io_out_1(c53_200_io_out_1),
    .io_out_2(c53_200_io_out_2)
  );
  C53 c53_201 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_201_io_in_0),
    .io_in_1(c53_201_io_in_1),
    .io_in_2(c53_201_io_in_2),
    .io_in_3(c53_201_io_in_3),
    .io_in_4(c53_201_io_in_4),
    .io_out_0(c53_201_io_out_0),
    .io_out_1(c53_201_io_out_1),
    .io_out_2(c53_201_io_out_2)
  );
  C53 c53_202 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_202_io_in_0),
    .io_in_1(c53_202_io_in_1),
    .io_in_2(c53_202_io_in_2),
    .io_in_3(c53_202_io_in_3),
    .io_in_4(c53_202_io_in_4),
    .io_out_0(c53_202_io_out_0),
    .io_out_1(c53_202_io_out_1),
    .io_out_2(c53_202_io_out_2)
  );
  C22 c22_14 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_14_io_in_0),
    .io_in_1(c22_14_io_in_1),
    .io_out_0(c22_14_io_out_0),
    .io_out_1(c22_14_io_out_1)
  );
  C53 c53_203 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_203_io_in_0),
    .io_in_1(c53_203_io_in_1),
    .io_in_2(c53_203_io_in_2),
    .io_in_3(c53_203_io_in_3),
    .io_in_4(c53_203_io_in_4),
    .io_out_0(c53_203_io_out_0),
    .io_out_1(c53_203_io_out_1),
    .io_out_2(c53_203_io_out_2)
  );
  C53 c53_204 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_204_io_in_0),
    .io_in_1(c53_204_io_in_1),
    .io_in_2(c53_204_io_in_2),
    .io_in_3(c53_204_io_in_3),
    .io_in_4(c53_204_io_in_4),
    .io_out_0(c53_204_io_out_0),
    .io_out_1(c53_204_io_out_1),
    .io_out_2(c53_204_io_out_2)
  );
  C53 c53_205 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_205_io_in_0),
    .io_in_1(c53_205_io_in_1),
    .io_in_2(c53_205_io_in_2),
    .io_in_3(c53_205_io_in_3),
    .io_in_4(c53_205_io_in_4),
    .io_out_0(c53_205_io_out_0),
    .io_out_1(c53_205_io_out_1),
    .io_out_2(c53_205_io_out_2)
  );
  C53 c53_206 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_206_io_in_0),
    .io_in_1(c53_206_io_in_1),
    .io_in_2(c53_206_io_in_2),
    .io_in_3(c53_206_io_in_3),
    .io_in_4(c53_206_io_in_4),
    .io_out_0(c53_206_io_out_0),
    .io_out_1(c53_206_io_out_1),
    .io_out_2(c53_206_io_out_2)
  );
  C53 c53_207 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_207_io_in_0),
    .io_in_1(c53_207_io_in_1),
    .io_in_2(c53_207_io_in_2),
    .io_in_3(c53_207_io_in_3),
    .io_in_4(c53_207_io_in_4),
    .io_out_0(c53_207_io_out_0),
    .io_out_1(c53_207_io_out_1),
    .io_out_2(c53_207_io_out_2)
  );
  C53 c53_208 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_208_io_in_0),
    .io_in_1(c53_208_io_in_1),
    .io_in_2(c53_208_io_in_2),
    .io_in_3(c53_208_io_in_3),
    .io_in_4(c53_208_io_in_4),
    .io_out_0(c53_208_io_out_0),
    .io_out_1(c53_208_io_out_1),
    .io_out_2(c53_208_io_out_2)
  );
  C53 c53_209 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_209_io_in_0),
    .io_in_1(c53_209_io_in_1),
    .io_in_2(c53_209_io_in_2),
    .io_in_3(c53_209_io_in_3),
    .io_in_4(c53_209_io_in_4),
    .io_out_0(c53_209_io_out_0),
    .io_out_1(c53_209_io_out_1),
    .io_out_2(c53_209_io_out_2)
  );
  C22 c22_15 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_15_io_in_0),
    .io_in_1(c22_15_io_in_1),
    .io_out_0(c22_15_io_out_0),
    .io_out_1(c22_15_io_out_1)
  );
  C53 c53_210 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_210_io_in_0),
    .io_in_1(c53_210_io_in_1),
    .io_in_2(c53_210_io_in_2),
    .io_in_3(c53_210_io_in_3),
    .io_in_4(c53_210_io_in_4),
    .io_out_0(c53_210_io_out_0),
    .io_out_1(c53_210_io_out_1),
    .io_out_2(c53_210_io_out_2)
  );
  C53 c53_211 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_211_io_in_0),
    .io_in_1(c53_211_io_in_1),
    .io_in_2(c53_211_io_in_2),
    .io_in_3(c53_211_io_in_3),
    .io_in_4(c53_211_io_in_4),
    .io_out_0(c53_211_io_out_0),
    .io_out_1(c53_211_io_out_1),
    .io_out_2(c53_211_io_out_2)
  );
  C53 c53_212 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_212_io_in_0),
    .io_in_1(c53_212_io_in_1),
    .io_in_2(c53_212_io_in_2),
    .io_in_3(c53_212_io_in_3),
    .io_in_4(c53_212_io_in_4),
    .io_out_0(c53_212_io_out_0),
    .io_out_1(c53_212_io_out_1),
    .io_out_2(c53_212_io_out_2)
  );
  C53 c53_213 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_213_io_in_0),
    .io_in_1(c53_213_io_in_1),
    .io_in_2(c53_213_io_in_2),
    .io_in_3(c53_213_io_in_3),
    .io_in_4(c53_213_io_in_4),
    .io_out_0(c53_213_io_out_0),
    .io_out_1(c53_213_io_out_1),
    .io_out_2(c53_213_io_out_2)
  );
  C53 c53_214 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_214_io_in_0),
    .io_in_1(c53_214_io_in_1),
    .io_in_2(c53_214_io_in_2),
    .io_in_3(c53_214_io_in_3),
    .io_in_4(c53_214_io_in_4),
    .io_out_0(c53_214_io_out_0),
    .io_out_1(c53_214_io_out_1),
    .io_out_2(c53_214_io_out_2)
  );
  C53 c53_215 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_215_io_in_0),
    .io_in_1(c53_215_io_in_1),
    .io_in_2(c53_215_io_in_2),
    .io_in_3(c53_215_io_in_3),
    .io_in_4(c53_215_io_in_4),
    .io_out_0(c53_215_io_out_0),
    .io_out_1(c53_215_io_out_1),
    .io_out_2(c53_215_io_out_2)
  );
  C53 c53_216 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_216_io_in_0),
    .io_in_1(c53_216_io_in_1),
    .io_in_2(c53_216_io_in_2),
    .io_in_3(c53_216_io_in_3),
    .io_in_4(c53_216_io_in_4),
    .io_out_0(c53_216_io_out_0),
    .io_out_1(c53_216_io_out_1),
    .io_out_2(c53_216_io_out_2)
  );
  C32 c32_14 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_14_io_in_0),
    .io_in_1(c32_14_io_in_1),
    .io_in_2(c32_14_io_in_2),
    .io_out_0(c32_14_io_out_0),
    .io_out_1(c32_14_io_out_1)
  );
  C53 c53_217 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_217_io_in_0),
    .io_in_1(c53_217_io_in_1),
    .io_in_2(c53_217_io_in_2),
    .io_in_3(c53_217_io_in_3),
    .io_in_4(c53_217_io_in_4),
    .io_out_0(c53_217_io_out_0),
    .io_out_1(c53_217_io_out_1),
    .io_out_2(c53_217_io_out_2)
  );
  C53 c53_218 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_218_io_in_0),
    .io_in_1(c53_218_io_in_1),
    .io_in_2(c53_218_io_in_2),
    .io_in_3(c53_218_io_in_3),
    .io_in_4(c53_218_io_in_4),
    .io_out_0(c53_218_io_out_0),
    .io_out_1(c53_218_io_out_1),
    .io_out_2(c53_218_io_out_2)
  );
  C53 c53_219 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_219_io_in_0),
    .io_in_1(c53_219_io_in_1),
    .io_in_2(c53_219_io_in_2),
    .io_in_3(c53_219_io_in_3),
    .io_in_4(c53_219_io_in_4),
    .io_out_0(c53_219_io_out_0),
    .io_out_1(c53_219_io_out_1),
    .io_out_2(c53_219_io_out_2)
  );
  C53 c53_220 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_220_io_in_0),
    .io_in_1(c53_220_io_in_1),
    .io_in_2(c53_220_io_in_2),
    .io_in_3(c53_220_io_in_3),
    .io_in_4(c53_220_io_in_4),
    .io_out_0(c53_220_io_out_0),
    .io_out_1(c53_220_io_out_1),
    .io_out_2(c53_220_io_out_2)
  );
  C53 c53_221 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_221_io_in_0),
    .io_in_1(c53_221_io_in_1),
    .io_in_2(c53_221_io_in_2),
    .io_in_3(c53_221_io_in_3),
    .io_in_4(c53_221_io_in_4),
    .io_out_0(c53_221_io_out_0),
    .io_out_1(c53_221_io_out_1),
    .io_out_2(c53_221_io_out_2)
  );
  C53 c53_222 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_222_io_in_0),
    .io_in_1(c53_222_io_in_1),
    .io_in_2(c53_222_io_in_2),
    .io_in_3(c53_222_io_in_3),
    .io_in_4(c53_222_io_in_4),
    .io_out_0(c53_222_io_out_0),
    .io_out_1(c53_222_io_out_1),
    .io_out_2(c53_222_io_out_2)
  );
  C53 c53_223 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_223_io_in_0),
    .io_in_1(c53_223_io_in_1),
    .io_in_2(c53_223_io_in_2),
    .io_in_3(c53_223_io_in_3),
    .io_in_4(c53_223_io_in_4),
    .io_out_0(c53_223_io_out_0),
    .io_out_1(c53_223_io_out_1),
    .io_out_2(c53_223_io_out_2)
  );
  C32 c32_15 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_15_io_in_0),
    .io_in_1(c32_15_io_in_1),
    .io_in_2(c32_15_io_in_2),
    .io_out_0(c32_15_io_out_0),
    .io_out_1(c32_15_io_out_1)
  );
  C53 c53_224 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_224_io_in_0),
    .io_in_1(c53_224_io_in_1),
    .io_in_2(c53_224_io_in_2),
    .io_in_3(c53_224_io_in_3),
    .io_in_4(c53_224_io_in_4),
    .io_out_0(c53_224_io_out_0),
    .io_out_1(c53_224_io_out_1),
    .io_out_2(c53_224_io_out_2)
  );
  C53 c53_225 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_225_io_in_0),
    .io_in_1(c53_225_io_in_1),
    .io_in_2(c53_225_io_in_2),
    .io_in_3(c53_225_io_in_3),
    .io_in_4(c53_225_io_in_4),
    .io_out_0(c53_225_io_out_0),
    .io_out_1(c53_225_io_out_1),
    .io_out_2(c53_225_io_out_2)
  );
  C53 c53_226 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_226_io_in_0),
    .io_in_1(c53_226_io_in_1),
    .io_in_2(c53_226_io_in_2),
    .io_in_3(c53_226_io_in_3),
    .io_in_4(c53_226_io_in_4),
    .io_out_0(c53_226_io_out_0),
    .io_out_1(c53_226_io_out_1),
    .io_out_2(c53_226_io_out_2)
  );
  C53 c53_227 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_227_io_in_0),
    .io_in_1(c53_227_io_in_1),
    .io_in_2(c53_227_io_in_2),
    .io_in_3(c53_227_io_in_3),
    .io_in_4(c53_227_io_in_4),
    .io_out_0(c53_227_io_out_0),
    .io_out_1(c53_227_io_out_1),
    .io_out_2(c53_227_io_out_2)
  );
  C53 c53_228 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_228_io_in_0),
    .io_in_1(c53_228_io_in_1),
    .io_in_2(c53_228_io_in_2),
    .io_in_3(c53_228_io_in_3),
    .io_in_4(c53_228_io_in_4),
    .io_out_0(c53_228_io_out_0),
    .io_out_1(c53_228_io_out_1),
    .io_out_2(c53_228_io_out_2)
  );
  C53 c53_229 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_229_io_in_0),
    .io_in_1(c53_229_io_in_1),
    .io_in_2(c53_229_io_in_2),
    .io_in_3(c53_229_io_in_3),
    .io_in_4(c53_229_io_in_4),
    .io_out_0(c53_229_io_out_0),
    .io_out_1(c53_229_io_out_1),
    .io_out_2(c53_229_io_out_2)
  );
  C53 c53_230 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_230_io_in_0),
    .io_in_1(c53_230_io_in_1),
    .io_in_2(c53_230_io_in_2),
    .io_in_3(c53_230_io_in_3),
    .io_in_4(c53_230_io_in_4),
    .io_out_0(c53_230_io_out_0),
    .io_out_1(c53_230_io_out_1),
    .io_out_2(c53_230_io_out_2)
  );
  C53 c53_231 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_231_io_in_0),
    .io_in_1(c53_231_io_in_1),
    .io_in_2(c53_231_io_in_2),
    .io_in_3(c53_231_io_in_3),
    .io_in_4(c53_231_io_in_4),
    .io_out_0(c53_231_io_out_0),
    .io_out_1(c53_231_io_out_1),
    .io_out_2(c53_231_io_out_2)
  );
  C53 c53_232 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_232_io_in_0),
    .io_in_1(c53_232_io_in_1),
    .io_in_2(c53_232_io_in_2),
    .io_in_3(c53_232_io_in_3),
    .io_in_4(c53_232_io_in_4),
    .io_out_0(c53_232_io_out_0),
    .io_out_1(c53_232_io_out_1),
    .io_out_2(c53_232_io_out_2)
  );
  C53 c53_233 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_233_io_in_0),
    .io_in_1(c53_233_io_in_1),
    .io_in_2(c53_233_io_in_2),
    .io_in_3(c53_233_io_in_3),
    .io_in_4(c53_233_io_in_4),
    .io_out_0(c53_233_io_out_0),
    .io_out_1(c53_233_io_out_1),
    .io_out_2(c53_233_io_out_2)
  );
  C53 c53_234 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_234_io_in_0),
    .io_in_1(c53_234_io_in_1),
    .io_in_2(c53_234_io_in_2),
    .io_in_3(c53_234_io_in_3),
    .io_in_4(c53_234_io_in_4),
    .io_out_0(c53_234_io_out_0),
    .io_out_1(c53_234_io_out_1),
    .io_out_2(c53_234_io_out_2)
  );
  C53 c53_235 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_235_io_in_0),
    .io_in_1(c53_235_io_in_1),
    .io_in_2(c53_235_io_in_2),
    .io_in_3(c53_235_io_in_3),
    .io_in_4(c53_235_io_in_4),
    .io_out_0(c53_235_io_out_0),
    .io_out_1(c53_235_io_out_1),
    .io_out_2(c53_235_io_out_2)
  );
  C53 c53_236 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_236_io_in_0),
    .io_in_1(c53_236_io_in_1),
    .io_in_2(c53_236_io_in_2),
    .io_in_3(c53_236_io_in_3),
    .io_in_4(c53_236_io_in_4),
    .io_out_0(c53_236_io_out_0),
    .io_out_1(c53_236_io_out_1),
    .io_out_2(c53_236_io_out_2)
  );
  C53 c53_237 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_237_io_in_0),
    .io_in_1(c53_237_io_in_1),
    .io_in_2(c53_237_io_in_2),
    .io_in_3(c53_237_io_in_3),
    .io_in_4(c53_237_io_in_4),
    .io_out_0(c53_237_io_out_0),
    .io_out_1(c53_237_io_out_1),
    .io_out_2(c53_237_io_out_2)
  );
  C53 c53_238 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_238_io_in_0),
    .io_in_1(c53_238_io_in_1),
    .io_in_2(c53_238_io_in_2),
    .io_in_3(c53_238_io_in_3),
    .io_in_4(c53_238_io_in_4),
    .io_out_0(c53_238_io_out_0),
    .io_out_1(c53_238_io_out_1),
    .io_out_2(c53_238_io_out_2)
  );
  C53 c53_239 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_239_io_in_0),
    .io_in_1(c53_239_io_in_1),
    .io_in_2(c53_239_io_in_2),
    .io_in_3(c53_239_io_in_3),
    .io_in_4(c53_239_io_in_4),
    .io_out_0(c53_239_io_out_0),
    .io_out_1(c53_239_io_out_1),
    .io_out_2(c53_239_io_out_2)
  );
  C53 c53_240 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_240_io_in_0),
    .io_in_1(c53_240_io_in_1),
    .io_in_2(c53_240_io_in_2),
    .io_in_3(c53_240_io_in_3),
    .io_in_4(c53_240_io_in_4),
    .io_out_0(c53_240_io_out_0),
    .io_out_1(c53_240_io_out_1),
    .io_out_2(c53_240_io_out_2)
  );
  C53 c53_241 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_241_io_in_0),
    .io_in_1(c53_241_io_in_1),
    .io_in_2(c53_241_io_in_2),
    .io_in_3(c53_241_io_in_3),
    .io_in_4(c53_241_io_in_4),
    .io_out_0(c53_241_io_out_0),
    .io_out_1(c53_241_io_out_1),
    .io_out_2(c53_241_io_out_2)
  );
  C53 c53_242 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_242_io_in_0),
    .io_in_1(c53_242_io_in_1),
    .io_in_2(c53_242_io_in_2),
    .io_in_3(c53_242_io_in_3),
    .io_in_4(c53_242_io_in_4),
    .io_out_0(c53_242_io_out_0),
    .io_out_1(c53_242_io_out_1),
    .io_out_2(c53_242_io_out_2)
  );
  C53 c53_243 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_243_io_in_0),
    .io_in_1(c53_243_io_in_1),
    .io_in_2(c53_243_io_in_2),
    .io_in_3(c53_243_io_in_3),
    .io_in_4(c53_243_io_in_4),
    .io_out_0(c53_243_io_out_0),
    .io_out_1(c53_243_io_out_1),
    .io_out_2(c53_243_io_out_2)
  );
  C53 c53_244 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_244_io_in_0),
    .io_in_1(c53_244_io_in_1),
    .io_in_2(c53_244_io_in_2),
    .io_in_3(c53_244_io_in_3),
    .io_in_4(c53_244_io_in_4),
    .io_out_0(c53_244_io_out_0),
    .io_out_1(c53_244_io_out_1),
    .io_out_2(c53_244_io_out_2)
  );
  C53 c53_245 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_245_io_in_0),
    .io_in_1(c53_245_io_in_1),
    .io_in_2(c53_245_io_in_2),
    .io_in_3(c53_245_io_in_3),
    .io_in_4(c53_245_io_in_4),
    .io_out_0(c53_245_io_out_0),
    .io_out_1(c53_245_io_out_1),
    .io_out_2(c53_245_io_out_2)
  );
  C53 c53_246 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_246_io_in_0),
    .io_in_1(c53_246_io_in_1),
    .io_in_2(c53_246_io_in_2),
    .io_in_3(c53_246_io_in_3),
    .io_in_4(c53_246_io_in_4),
    .io_out_0(c53_246_io_out_0),
    .io_out_1(c53_246_io_out_1),
    .io_out_2(c53_246_io_out_2)
  );
  C53 c53_247 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_247_io_in_0),
    .io_in_1(c53_247_io_in_1),
    .io_in_2(c53_247_io_in_2),
    .io_in_3(c53_247_io_in_3),
    .io_in_4(c53_247_io_in_4),
    .io_out_0(c53_247_io_out_0),
    .io_out_1(c53_247_io_out_1),
    .io_out_2(c53_247_io_out_2)
  );
  C53 c53_248 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_248_io_in_0),
    .io_in_1(c53_248_io_in_1),
    .io_in_2(c53_248_io_in_2),
    .io_in_3(c53_248_io_in_3),
    .io_in_4(c53_248_io_in_4),
    .io_out_0(c53_248_io_out_0),
    .io_out_1(c53_248_io_out_1),
    .io_out_2(c53_248_io_out_2)
  );
  C53 c53_249 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_249_io_in_0),
    .io_in_1(c53_249_io_in_1),
    .io_in_2(c53_249_io_in_2),
    .io_in_3(c53_249_io_in_3),
    .io_in_4(c53_249_io_in_4),
    .io_out_0(c53_249_io_out_0),
    .io_out_1(c53_249_io_out_1),
    .io_out_2(c53_249_io_out_2)
  );
  C53 c53_250 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_250_io_in_0),
    .io_in_1(c53_250_io_in_1),
    .io_in_2(c53_250_io_in_2),
    .io_in_3(c53_250_io_in_3),
    .io_in_4(c53_250_io_in_4),
    .io_out_0(c53_250_io_out_0),
    .io_out_1(c53_250_io_out_1),
    .io_out_2(c53_250_io_out_2)
  );
  C53 c53_251 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_251_io_in_0),
    .io_in_1(c53_251_io_in_1),
    .io_in_2(c53_251_io_in_2),
    .io_in_3(c53_251_io_in_3),
    .io_in_4(c53_251_io_in_4),
    .io_out_0(c53_251_io_out_0),
    .io_out_1(c53_251_io_out_1),
    .io_out_2(c53_251_io_out_2)
  );
  C53 c53_252 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_252_io_in_0),
    .io_in_1(c53_252_io_in_1),
    .io_in_2(c53_252_io_in_2),
    .io_in_3(c53_252_io_in_3),
    .io_in_4(c53_252_io_in_4),
    .io_out_0(c53_252_io_out_0),
    .io_out_1(c53_252_io_out_1),
    .io_out_2(c53_252_io_out_2)
  );
  C53 c53_253 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_253_io_in_0),
    .io_in_1(c53_253_io_in_1),
    .io_in_2(c53_253_io_in_2),
    .io_in_3(c53_253_io_in_3),
    .io_in_4(c53_253_io_in_4),
    .io_out_0(c53_253_io_out_0),
    .io_out_1(c53_253_io_out_1),
    .io_out_2(c53_253_io_out_2)
  );
  C53 c53_254 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_254_io_in_0),
    .io_in_1(c53_254_io_in_1),
    .io_in_2(c53_254_io_in_2),
    .io_in_3(c53_254_io_in_3),
    .io_in_4(c53_254_io_in_4),
    .io_out_0(c53_254_io_out_0),
    .io_out_1(c53_254_io_out_1),
    .io_out_2(c53_254_io_out_2)
  );
  C53 c53_255 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_255_io_in_0),
    .io_in_1(c53_255_io_in_1),
    .io_in_2(c53_255_io_in_2),
    .io_in_3(c53_255_io_in_3),
    .io_in_4(c53_255_io_in_4),
    .io_out_0(c53_255_io_out_0),
    .io_out_1(c53_255_io_out_1),
    .io_out_2(c53_255_io_out_2)
  );
  C53 c53_256 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_256_io_in_0),
    .io_in_1(c53_256_io_in_1),
    .io_in_2(c53_256_io_in_2),
    .io_in_3(c53_256_io_in_3),
    .io_in_4(c53_256_io_in_4),
    .io_out_0(c53_256_io_out_0),
    .io_out_1(c53_256_io_out_1),
    .io_out_2(c53_256_io_out_2)
  );
  C53 c53_257 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_257_io_in_0),
    .io_in_1(c53_257_io_in_1),
    .io_in_2(c53_257_io_in_2),
    .io_in_3(c53_257_io_in_3),
    .io_in_4(c53_257_io_in_4),
    .io_out_0(c53_257_io_out_0),
    .io_out_1(c53_257_io_out_1),
    .io_out_2(c53_257_io_out_2)
  );
  C53 c53_258 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_258_io_in_0),
    .io_in_1(c53_258_io_in_1),
    .io_in_2(c53_258_io_in_2),
    .io_in_3(c53_258_io_in_3),
    .io_in_4(c53_258_io_in_4),
    .io_out_0(c53_258_io_out_0),
    .io_out_1(c53_258_io_out_1),
    .io_out_2(c53_258_io_out_2)
  );
  C53 c53_259 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_259_io_in_0),
    .io_in_1(c53_259_io_in_1),
    .io_in_2(c53_259_io_in_2),
    .io_in_3(c53_259_io_in_3),
    .io_in_4(c53_259_io_in_4),
    .io_out_0(c53_259_io_out_0),
    .io_out_1(c53_259_io_out_1),
    .io_out_2(c53_259_io_out_2)
  );
  C53 c53_260 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_260_io_in_0),
    .io_in_1(c53_260_io_in_1),
    .io_in_2(c53_260_io_in_2),
    .io_in_3(c53_260_io_in_3),
    .io_in_4(c53_260_io_in_4),
    .io_out_0(c53_260_io_out_0),
    .io_out_1(c53_260_io_out_1),
    .io_out_2(c53_260_io_out_2)
  );
  C53 c53_261 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_261_io_in_0),
    .io_in_1(c53_261_io_in_1),
    .io_in_2(c53_261_io_in_2),
    .io_in_3(c53_261_io_in_3),
    .io_in_4(c53_261_io_in_4),
    .io_out_0(c53_261_io_out_0),
    .io_out_1(c53_261_io_out_1),
    .io_out_2(c53_261_io_out_2)
  );
  C53 c53_262 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_262_io_in_0),
    .io_in_1(c53_262_io_in_1),
    .io_in_2(c53_262_io_in_2),
    .io_in_3(c53_262_io_in_3),
    .io_in_4(c53_262_io_in_4),
    .io_out_0(c53_262_io_out_0),
    .io_out_1(c53_262_io_out_1),
    .io_out_2(c53_262_io_out_2)
  );
  C53 c53_263 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_263_io_in_0),
    .io_in_1(c53_263_io_in_1),
    .io_in_2(c53_263_io_in_2),
    .io_in_3(c53_263_io_in_3),
    .io_in_4(c53_263_io_in_4),
    .io_out_0(c53_263_io_out_0),
    .io_out_1(c53_263_io_out_1),
    .io_out_2(c53_263_io_out_2)
  );
  C53 c53_264 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_264_io_in_0),
    .io_in_1(c53_264_io_in_1),
    .io_in_2(c53_264_io_in_2),
    .io_in_3(c53_264_io_in_3),
    .io_in_4(c53_264_io_in_4),
    .io_out_0(c53_264_io_out_0),
    .io_out_1(c53_264_io_out_1),
    .io_out_2(c53_264_io_out_2)
  );
  C53 c53_265 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_265_io_in_0),
    .io_in_1(c53_265_io_in_1),
    .io_in_2(c53_265_io_in_2),
    .io_in_3(c53_265_io_in_3),
    .io_in_4(c53_265_io_in_4),
    .io_out_0(c53_265_io_out_0),
    .io_out_1(c53_265_io_out_1),
    .io_out_2(c53_265_io_out_2)
  );
  C53 c53_266 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_266_io_in_0),
    .io_in_1(c53_266_io_in_1),
    .io_in_2(c53_266_io_in_2),
    .io_in_3(c53_266_io_in_3),
    .io_in_4(c53_266_io_in_4),
    .io_out_0(c53_266_io_out_0),
    .io_out_1(c53_266_io_out_1),
    .io_out_2(c53_266_io_out_2)
  );
  C53 c53_267 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_267_io_in_0),
    .io_in_1(c53_267_io_in_1),
    .io_in_2(c53_267_io_in_2),
    .io_in_3(c53_267_io_in_3),
    .io_in_4(c53_267_io_in_4),
    .io_out_0(c53_267_io_out_0),
    .io_out_1(c53_267_io_out_1),
    .io_out_2(c53_267_io_out_2)
  );
  C53 c53_268 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_268_io_in_0),
    .io_in_1(c53_268_io_in_1),
    .io_in_2(c53_268_io_in_2),
    .io_in_3(c53_268_io_in_3),
    .io_in_4(c53_268_io_in_4),
    .io_out_0(c53_268_io_out_0),
    .io_out_1(c53_268_io_out_1),
    .io_out_2(c53_268_io_out_2)
  );
  C53 c53_269 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_269_io_in_0),
    .io_in_1(c53_269_io_in_1),
    .io_in_2(c53_269_io_in_2),
    .io_in_3(c53_269_io_in_3),
    .io_in_4(c53_269_io_in_4),
    .io_out_0(c53_269_io_out_0),
    .io_out_1(c53_269_io_out_1),
    .io_out_2(c53_269_io_out_2)
  );
  C53 c53_270 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_270_io_in_0),
    .io_in_1(c53_270_io_in_1),
    .io_in_2(c53_270_io_in_2),
    .io_in_3(c53_270_io_in_3),
    .io_in_4(c53_270_io_in_4),
    .io_out_0(c53_270_io_out_0),
    .io_out_1(c53_270_io_out_1),
    .io_out_2(c53_270_io_out_2)
  );
  C53 c53_271 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_271_io_in_0),
    .io_in_1(c53_271_io_in_1),
    .io_in_2(c53_271_io_in_2),
    .io_in_3(c53_271_io_in_3),
    .io_in_4(c53_271_io_in_4),
    .io_out_0(c53_271_io_out_0),
    .io_out_1(c53_271_io_out_1),
    .io_out_2(c53_271_io_out_2)
  );
  C53 c53_272 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_272_io_in_0),
    .io_in_1(c53_272_io_in_1),
    .io_in_2(c53_272_io_in_2),
    .io_in_3(c53_272_io_in_3),
    .io_in_4(c53_272_io_in_4),
    .io_out_0(c53_272_io_out_0),
    .io_out_1(c53_272_io_out_1),
    .io_out_2(c53_272_io_out_2)
  );
  C53 c53_273 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_273_io_in_0),
    .io_in_1(c53_273_io_in_1),
    .io_in_2(c53_273_io_in_2),
    .io_in_3(c53_273_io_in_3),
    .io_in_4(c53_273_io_in_4),
    .io_out_0(c53_273_io_out_0),
    .io_out_1(c53_273_io_out_1),
    .io_out_2(c53_273_io_out_2)
  );
  C53 c53_274 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_274_io_in_0),
    .io_in_1(c53_274_io_in_1),
    .io_in_2(c53_274_io_in_2),
    .io_in_3(c53_274_io_in_3),
    .io_in_4(c53_274_io_in_4),
    .io_out_0(c53_274_io_out_0),
    .io_out_1(c53_274_io_out_1),
    .io_out_2(c53_274_io_out_2)
  );
  C53 c53_275 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_275_io_in_0),
    .io_in_1(c53_275_io_in_1),
    .io_in_2(c53_275_io_in_2),
    .io_in_3(c53_275_io_in_3),
    .io_in_4(c53_275_io_in_4),
    .io_out_0(c53_275_io_out_0),
    .io_out_1(c53_275_io_out_1),
    .io_out_2(c53_275_io_out_2)
  );
  C53 c53_276 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_276_io_in_0),
    .io_in_1(c53_276_io_in_1),
    .io_in_2(c53_276_io_in_2),
    .io_in_3(c53_276_io_in_3),
    .io_in_4(c53_276_io_in_4),
    .io_out_0(c53_276_io_out_0),
    .io_out_1(c53_276_io_out_1),
    .io_out_2(c53_276_io_out_2)
  );
  C53 c53_277 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_277_io_in_0),
    .io_in_1(c53_277_io_in_1),
    .io_in_2(c53_277_io_in_2),
    .io_in_3(c53_277_io_in_3),
    .io_in_4(c53_277_io_in_4),
    .io_out_0(c53_277_io_out_0),
    .io_out_1(c53_277_io_out_1),
    .io_out_2(c53_277_io_out_2)
  );
  C53 c53_278 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_278_io_in_0),
    .io_in_1(c53_278_io_in_1),
    .io_in_2(c53_278_io_in_2),
    .io_in_3(c53_278_io_in_3),
    .io_in_4(c53_278_io_in_4),
    .io_out_0(c53_278_io_out_0),
    .io_out_1(c53_278_io_out_1),
    .io_out_2(c53_278_io_out_2)
  );
  C53 c53_279 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_279_io_in_0),
    .io_in_1(c53_279_io_in_1),
    .io_in_2(c53_279_io_in_2),
    .io_in_3(c53_279_io_in_3),
    .io_in_4(c53_279_io_in_4),
    .io_out_0(c53_279_io_out_0),
    .io_out_1(c53_279_io_out_1),
    .io_out_2(c53_279_io_out_2)
  );
  C53 c53_280 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_280_io_in_0),
    .io_in_1(c53_280_io_in_1),
    .io_in_2(c53_280_io_in_2),
    .io_in_3(c53_280_io_in_3),
    .io_in_4(c53_280_io_in_4),
    .io_out_0(c53_280_io_out_0),
    .io_out_1(c53_280_io_out_1),
    .io_out_2(c53_280_io_out_2)
  );
  C53 c53_281 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_281_io_in_0),
    .io_in_1(c53_281_io_in_1),
    .io_in_2(c53_281_io_in_2),
    .io_in_3(c53_281_io_in_3),
    .io_in_4(c53_281_io_in_4),
    .io_out_0(c53_281_io_out_0),
    .io_out_1(c53_281_io_out_1),
    .io_out_2(c53_281_io_out_2)
  );
  C53 c53_282 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_282_io_in_0),
    .io_in_1(c53_282_io_in_1),
    .io_in_2(c53_282_io_in_2),
    .io_in_3(c53_282_io_in_3),
    .io_in_4(c53_282_io_in_4),
    .io_out_0(c53_282_io_out_0),
    .io_out_1(c53_282_io_out_1),
    .io_out_2(c53_282_io_out_2)
  );
  C53 c53_283 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_283_io_in_0),
    .io_in_1(c53_283_io_in_1),
    .io_in_2(c53_283_io_in_2),
    .io_in_3(c53_283_io_in_3),
    .io_in_4(c53_283_io_in_4),
    .io_out_0(c53_283_io_out_0),
    .io_out_1(c53_283_io_out_1),
    .io_out_2(c53_283_io_out_2)
  );
  C53 c53_284 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_284_io_in_0),
    .io_in_1(c53_284_io_in_1),
    .io_in_2(c53_284_io_in_2),
    .io_in_3(c53_284_io_in_3),
    .io_in_4(c53_284_io_in_4),
    .io_out_0(c53_284_io_out_0),
    .io_out_1(c53_284_io_out_1),
    .io_out_2(c53_284_io_out_2)
  );
  C53 c53_285 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_285_io_in_0),
    .io_in_1(c53_285_io_in_1),
    .io_in_2(c53_285_io_in_2),
    .io_in_3(c53_285_io_in_3),
    .io_in_4(c53_285_io_in_4),
    .io_out_0(c53_285_io_out_0),
    .io_out_1(c53_285_io_out_1),
    .io_out_2(c53_285_io_out_2)
  );
  C53 c53_286 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_286_io_in_0),
    .io_in_1(c53_286_io_in_1),
    .io_in_2(c53_286_io_in_2),
    .io_in_3(c53_286_io_in_3),
    .io_in_4(c53_286_io_in_4),
    .io_out_0(c53_286_io_out_0),
    .io_out_1(c53_286_io_out_1),
    .io_out_2(c53_286_io_out_2)
  );
  C53 c53_287 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_287_io_in_0),
    .io_in_1(c53_287_io_in_1),
    .io_in_2(c53_287_io_in_2),
    .io_in_3(c53_287_io_in_3),
    .io_in_4(c53_287_io_in_4),
    .io_out_0(c53_287_io_out_0),
    .io_out_1(c53_287_io_out_1),
    .io_out_2(c53_287_io_out_2)
  );
  C53 c53_288 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_288_io_in_0),
    .io_in_1(c53_288_io_in_1),
    .io_in_2(c53_288_io_in_2),
    .io_in_3(c53_288_io_in_3),
    .io_in_4(c53_288_io_in_4),
    .io_out_0(c53_288_io_out_0),
    .io_out_1(c53_288_io_out_1),
    .io_out_2(c53_288_io_out_2)
  );
  C53 c53_289 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_289_io_in_0),
    .io_in_1(c53_289_io_in_1),
    .io_in_2(c53_289_io_in_2),
    .io_in_3(c53_289_io_in_3),
    .io_in_4(c53_289_io_in_4),
    .io_out_0(c53_289_io_out_0),
    .io_out_1(c53_289_io_out_1),
    .io_out_2(c53_289_io_out_2)
  );
  C53 c53_290 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_290_io_in_0),
    .io_in_1(c53_290_io_in_1),
    .io_in_2(c53_290_io_in_2),
    .io_in_3(c53_290_io_in_3),
    .io_in_4(c53_290_io_in_4),
    .io_out_0(c53_290_io_out_0),
    .io_out_1(c53_290_io_out_1),
    .io_out_2(c53_290_io_out_2)
  );
  C53 c53_291 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_291_io_in_0),
    .io_in_1(c53_291_io_in_1),
    .io_in_2(c53_291_io_in_2),
    .io_in_3(c53_291_io_in_3),
    .io_in_4(c53_291_io_in_4),
    .io_out_0(c53_291_io_out_0),
    .io_out_1(c53_291_io_out_1),
    .io_out_2(c53_291_io_out_2)
  );
  C53 c53_292 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_292_io_in_0),
    .io_in_1(c53_292_io_in_1),
    .io_in_2(c53_292_io_in_2),
    .io_in_3(c53_292_io_in_3),
    .io_in_4(c53_292_io_in_4),
    .io_out_0(c53_292_io_out_0),
    .io_out_1(c53_292_io_out_1),
    .io_out_2(c53_292_io_out_2)
  );
  C53 c53_293 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_293_io_in_0),
    .io_in_1(c53_293_io_in_1),
    .io_in_2(c53_293_io_in_2),
    .io_in_3(c53_293_io_in_3),
    .io_in_4(c53_293_io_in_4),
    .io_out_0(c53_293_io_out_0),
    .io_out_1(c53_293_io_out_1),
    .io_out_2(c53_293_io_out_2)
  );
  C53 c53_294 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_294_io_in_0),
    .io_in_1(c53_294_io_in_1),
    .io_in_2(c53_294_io_in_2),
    .io_in_3(c53_294_io_in_3),
    .io_in_4(c53_294_io_in_4),
    .io_out_0(c53_294_io_out_0),
    .io_out_1(c53_294_io_out_1),
    .io_out_2(c53_294_io_out_2)
  );
  C53 c53_295 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_295_io_in_0),
    .io_in_1(c53_295_io_in_1),
    .io_in_2(c53_295_io_in_2),
    .io_in_3(c53_295_io_in_3),
    .io_in_4(c53_295_io_in_4),
    .io_out_0(c53_295_io_out_0),
    .io_out_1(c53_295_io_out_1),
    .io_out_2(c53_295_io_out_2)
  );
  C53 c53_296 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_296_io_in_0),
    .io_in_1(c53_296_io_in_1),
    .io_in_2(c53_296_io_in_2),
    .io_in_3(c53_296_io_in_3),
    .io_in_4(c53_296_io_in_4),
    .io_out_0(c53_296_io_out_0),
    .io_out_1(c53_296_io_out_1),
    .io_out_2(c53_296_io_out_2)
  );
  C53 c53_297 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_297_io_in_0),
    .io_in_1(c53_297_io_in_1),
    .io_in_2(c53_297_io_in_2),
    .io_in_3(c53_297_io_in_3),
    .io_in_4(c53_297_io_in_4),
    .io_out_0(c53_297_io_out_0),
    .io_out_1(c53_297_io_out_1),
    .io_out_2(c53_297_io_out_2)
  );
  C53 c53_298 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_298_io_in_0),
    .io_in_1(c53_298_io_in_1),
    .io_in_2(c53_298_io_in_2),
    .io_in_3(c53_298_io_in_3),
    .io_in_4(c53_298_io_in_4),
    .io_out_0(c53_298_io_out_0),
    .io_out_1(c53_298_io_out_1),
    .io_out_2(c53_298_io_out_2)
  );
  C53 c53_299 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_299_io_in_0),
    .io_in_1(c53_299_io_in_1),
    .io_in_2(c53_299_io_in_2),
    .io_in_3(c53_299_io_in_3),
    .io_in_4(c53_299_io_in_4),
    .io_out_0(c53_299_io_out_0),
    .io_out_1(c53_299_io_out_1),
    .io_out_2(c53_299_io_out_2)
  );
  C53 c53_300 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_300_io_in_0),
    .io_in_1(c53_300_io_in_1),
    .io_in_2(c53_300_io_in_2),
    .io_in_3(c53_300_io_in_3),
    .io_in_4(c53_300_io_in_4),
    .io_out_0(c53_300_io_out_0),
    .io_out_1(c53_300_io_out_1),
    .io_out_2(c53_300_io_out_2)
  );
  C53 c53_301 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_301_io_in_0),
    .io_in_1(c53_301_io_in_1),
    .io_in_2(c53_301_io_in_2),
    .io_in_3(c53_301_io_in_3),
    .io_in_4(c53_301_io_in_4),
    .io_out_0(c53_301_io_out_0),
    .io_out_1(c53_301_io_out_1),
    .io_out_2(c53_301_io_out_2)
  );
  C53 c53_302 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_302_io_in_0),
    .io_in_1(c53_302_io_in_1),
    .io_in_2(c53_302_io_in_2),
    .io_in_3(c53_302_io_in_3),
    .io_in_4(c53_302_io_in_4),
    .io_out_0(c53_302_io_out_0),
    .io_out_1(c53_302_io_out_1),
    .io_out_2(c53_302_io_out_2)
  );
  C53 c53_303 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_303_io_in_0),
    .io_in_1(c53_303_io_in_1),
    .io_in_2(c53_303_io_in_2),
    .io_in_3(c53_303_io_in_3),
    .io_in_4(c53_303_io_in_4),
    .io_out_0(c53_303_io_out_0),
    .io_out_1(c53_303_io_out_1),
    .io_out_2(c53_303_io_out_2)
  );
  C53 c53_304 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_304_io_in_0),
    .io_in_1(c53_304_io_in_1),
    .io_in_2(c53_304_io_in_2),
    .io_in_3(c53_304_io_in_3),
    .io_in_4(c53_304_io_in_4),
    .io_out_0(c53_304_io_out_0),
    .io_out_1(c53_304_io_out_1),
    .io_out_2(c53_304_io_out_2)
  );
  C53 c53_305 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_305_io_in_0),
    .io_in_1(c53_305_io_in_1),
    .io_in_2(c53_305_io_in_2),
    .io_in_3(c53_305_io_in_3),
    .io_in_4(c53_305_io_in_4),
    .io_out_0(c53_305_io_out_0),
    .io_out_1(c53_305_io_out_1),
    .io_out_2(c53_305_io_out_2)
  );
  C53 c53_306 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_306_io_in_0),
    .io_in_1(c53_306_io_in_1),
    .io_in_2(c53_306_io_in_2),
    .io_in_3(c53_306_io_in_3),
    .io_in_4(c53_306_io_in_4),
    .io_out_0(c53_306_io_out_0),
    .io_out_1(c53_306_io_out_1),
    .io_out_2(c53_306_io_out_2)
  );
  C53 c53_307 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_307_io_in_0),
    .io_in_1(c53_307_io_in_1),
    .io_in_2(c53_307_io_in_2),
    .io_in_3(c53_307_io_in_3),
    .io_in_4(c53_307_io_in_4),
    .io_out_0(c53_307_io_out_0),
    .io_out_1(c53_307_io_out_1),
    .io_out_2(c53_307_io_out_2)
  );
  C53 c53_308 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_308_io_in_0),
    .io_in_1(c53_308_io_in_1),
    .io_in_2(c53_308_io_in_2),
    .io_in_3(c53_308_io_in_3),
    .io_in_4(c53_308_io_in_4),
    .io_out_0(c53_308_io_out_0),
    .io_out_1(c53_308_io_out_1),
    .io_out_2(c53_308_io_out_2)
  );
  C53 c53_309 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_309_io_in_0),
    .io_in_1(c53_309_io_in_1),
    .io_in_2(c53_309_io_in_2),
    .io_in_3(c53_309_io_in_3),
    .io_in_4(c53_309_io_in_4),
    .io_out_0(c53_309_io_out_0),
    .io_out_1(c53_309_io_out_1),
    .io_out_2(c53_309_io_out_2)
  );
  C53 c53_310 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_310_io_in_0),
    .io_in_1(c53_310_io_in_1),
    .io_in_2(c53_310_io_in_2),
    .io_in_3(c53_310_io_in_3),
    .io_in_4(c53_310_io_in_4),
    .io_out_0(c53_310_io_out_0),
    .io_out_1(c53_310_io_out_1),
    .io_out_2(c53_310_io_out_2)
  );
  C32 c32_16 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_16_io_in_0),
    .io_in_1(c32_16_io_in_1),
    .io_in_2(c32_16_io_in_2),
    .io_out_0(c32_16_io_out_0),
    .io_out_1(c32_16_io_out_1)
  );
  C53 c53_311 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_311_io_in_0),
    .io_in_1(c53_311_io_in_1),
    .io_in_2(c53_311_io_in_2),
    .io_in_3(c53_311_io_in_3),
    .io_in_4(c53_311_io_in_4),
    .io_out_0(c53_311_io_out_0),
    .io_out_1(c53_311_io_out_1),
    .io_out_2(c53_311_io_out_2)
  );
  C53 c53_312 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_312_io_in_0),
    .io_in_1(c53_312_io_in_1),
    .io_in_2(c53_312_io_in_2),
    .io_in_3(c53_312_io_in_3),
    .io_in_4(c53_312_io_in_4),
    .io_out_0(c53_312_io_out_0),
    .io_out_1(c53_312_io_out_1),
    .io_out_2(c53_312_io_out_2)
  );
  C53 c53_313 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_313_io_in_0),
    .io_in_1(c53_313_io_in_1),
    .io_in_2(c53_313_io_in_2),
    .io_in_3(c53_313_io_in_3),
    .io_in_4(c53_313_io_in_4),
    .io_out_0(c53_313_io_out_0),
    .io_out_1(c53_313_io_out_1),
    .io_out_2(c53_313_io_out_2)
  );
  C53 c53_314 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_314_io_in_0),
    .io_in_1(c53_314_io_in_1),
    .io_in_2(c53_314_io_in_2),
    .io_in_3(c53_314_io_in_3),
    .io_in_4(c53_314_io_in_4),
    .io_out_0(c53_314_io_out_0),
    .io_out_1(c53_314_io_out_1),
    .io_out_2(c53_314_io_out_2)
  );
  C53 c53_315 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_315_io_in_0),
    .io_in_1(c53_315_io_in_1),
    .io_in_2(c53_315_io_in_2),
    .io_in_3(c53_315_io_in_3),
    .io_in_4(c53_315_io_in_4),
    .io_out_0(c53_315_io_out_0),
    .io_out_1(c53_315_io_out_1),
    .io_out_2(c53_315_io_out_2)
  );
  C53 c53_316 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_316_io_in_0),
    .io_in_1(c53_316_io_in_1),
    .io_in_2(c53_316_io_in_2),
    .io_in_3(c53_316_io_in_3),
    .io_in_4(c53_316_io_in_4),
    .io_out_0(c53_316_io_out_0),
    .io_out_1(c53_316_io_out_1),
    .io_out_2(c53_316_io_out_2)
  );
  C53 c53_317 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_317_io_in_0),
    .io_in_1(c53_317_io_in_1),
    .io_in_2(c53_317_io_in_2),
    .io_in_3(c53_317_io_in_3),
    .io_in_4(c53_317_io_in_4),
    .io_out_0(c53_317_io_out_0),
    .io_out_1(c53_317_io_out_1),
    .io_out_2(c53_317_io_out_2)
  );
  C32 c32_17 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_17_io_in_0),
    .io_in_1(c32_17_io_in_1),
    .io_in_2(c32_17_io_in_2),
    .io_out_0(c32_17_io_out_0),
    .io_out_1(c32_17_io_out_1)
  );
  C53 c53_318 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_318_io_in_0),
    .io_in_1(c53_318_io_in_1),
    .io_in_2(c53_318_io_in_2),
    .io_in_3(c53_318_io_in_3),
    .io_in_4(c53_318_io_in_4),
    .io_out_0(c53_318_io_out_0),
    .io_out_1(c53_318_io_out_1),
    .io_out_2(c53_318_io_out_2)
  );
  C53 c53_319 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_319_io_in_0),
    .io_in_1(c53_319_io_in_1),
    .io_in_2(c53_319_io_in_2),
    .io_in_3(c53_319_io_in_3),
    .io_in_4(c53_319_io_in_4),
    .io_out_0(c53_319_io_out_0),
    .io_out_1(c53_319_io_out_1),
    .io_out_2(c53_319_io_out_2)
  );
  C53 c53_320 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_320_io_in_0),
    .io_in_1(c53_320_io_in_1),
    .io_in_2(c53_320_io_in_2),
    .io_in_3(c53_320_io_in_3),
    .io_in_4(c53_320_io_in_4),
    .io_out_0(c53_320_io_out_0),
    .io_out_1(c53_320_io_out_1),
    .io_out_2(c53_320_io_out_2)
  );
  C53 c53_321 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_321_io_in_0),
    .io_in_1(c53_321_io_in_1),
    .io_in_2(c53_321_io_in_2),
    .io_in_3(c53_321_io_in_3),
    .io_in_4(c53_321_io_in_4),
    .io_out_0(c53_321_io_out_0),
    .io_out_1(c53_321_io_out_1),
    .io_out_2(c53_321_io_out_2)
  );
  C53 c53_322 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_322_io_in_0),
    .io_in_1(c53_322_io_in_1),
    .io_in_2(c53_322_io_in_2),
    .io_in_3(c53_322_io_in_3),
    .io_in_4(c53_322_io_in_4),
    .io_out_0(c53_322_io_out_0),
    .io_out_1(c53_322_io_out_1),
    .io_out_2(c53_322_io_out_2)
  );
  C53 c53_323 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_323_io_in_0),
    .io_in_1(c53_323_io_in_1),
    .io_in_2(c53_323_io_in_2),
    .io_in_3(c53_323_io_in_3),
    .io_in_4(c53_323_io_in_4),
    .io_out_0(c53_323_io_out_0),
    .io_out_1(c53_323_io_out_1),
    .io_out_2(c53_323_io_out_2)
  );
  C53 c53_324 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_324_io_in_0),
    .io_in_1(c53_324_io_in_1),
    .io_in_2(c53_324_io_in_2),
    .io_in_3(c53_324_io_in_3),
    .io_in_4(c53_324_io_in_4),
    .io_out_0(c53_324_io_out_0),
    .io_out_1(c53_324_io_out_1),
    .io_out_2(c53_324_io_out_2)
  );
  C22 c22_16 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_16_io_in_0),
    .io_in_1(c22_16_io_in_1),
    .io_out_0(c22_16_io_out_0),
    .io_out_1(c22_16_io_out_1)
  );
  C53 c53_325 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_325_io_in_0),
    .io_in_1(c53_325_io_in_1),
    .io_in_2(c53_325_io_in_2),
    .io_in_3(c53_325_io_in_3),
    .io_in_4(c53_325_io_in_4),
    .io_out_0(c53_325_io_out_0),
    .io_out_1(c53_325_io_out_1),
    .io_out_2(c53_325_io_out_2)
  );
  C53 c53_326 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_326_io_in_0),
    .io_in_1(c53_326_io_in_1),
    .io_in_2(c53_326_io_in_2),
    .io_in_3(c53_326_io_in_3),
    .io_in_4(c53_326_io_in_4),
    .io_out_0(c53_326_io_out_0),
    .io_out_1(c53_326_io_out_1),
    .io_out_2(c53_326_io_out_2)
  );
  C53 c53_327 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_327_io_in_0),
    .io_in_1(c53_327_io_in_1),
    .io_in_2(c53_327_io_in_2),
    .io_in_3(c53_327_io_in_3),
    .io_in_4(c53_327_io_in_4),
    .io_out_0(c53_327_io_out_0),
    .io_out_1(c53_327_io_out_1),
    .io_out_2(c53_327_io_out_2)
  );
  C53 c53_328 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_328_io_in_0),
    .io_in_1(c53_328_io_in_1),
    .io_in_2(c53_328_io_in_2),
    .io_in_3(c53_328_io_in_3),
    .io_in_4(c53_328_io_in_4),
    .io_out_0(c53_328_io_out_0),
    .io_out_1(c53_328_io_out_1),
    .io_out_2(c53_328_io_out_2)
  );
  C53 c53_329 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_329_io_in_0),
    .io_in_1(c53_329_io_in_1),
    .io_in_2(c53_329_io_in_2),
    .io_in_3(c53_329_io_in_3),
    .io_in_4(c53_329_io_in_4),
    .io_out_0(c53_329_io_out_0),
    .io_out_1(c53_329_io_out_1),
    .io_out_2(c53_329_io_out_2)
  );
  C53 c53_330 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_330_io_in_0),
    .io_in_1(c53_330_io_in_1),
    .io_in_2(c53_330_io_in_2),
    .io_in_3(c53_330_io_in_3),
    .io_in_4(c53_330_io_in_4),
    .io_out_0(c53_330_io_out_0),
    .io_out_1(c53_330_io_out_1),
    .io_out_2(c53_330_io_out_2)
  );
  C53 c53_331 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_331_io_in_0),
    .io_in_1(c53_331_io_in_1),
    .io_in_2(c53_331_io_in_2),
    .io_in_3(c53_331_io_in_3),
    .io_in_4(c53_331_io_in_4),
    .io_out_0(c53_331_io_out_0),
    .io_out_1(c53_331_io_out_1),
    .io_out_2(c53_331_io_out_2)
  );
  C22 c22_17 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_17_io_in_0),
    .io_in_1(c22_17_io_in_1),
    .io_out_0(c22_17_io_out_0),
    .io_out_1(c22_17_io_out_1)
  );
  C53 c53_332 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_332_io_in_0),
    .io_in_1(c53_332_io_in_1),
    .io_in_2(c53_332_io_in_2),
    .io_in_3(c53_332_io_in_3),
    .io_in_4(c53_332_io_in_4),
    .io_out_0(c53_332_io_out_0),
    .io_out_1(c53_332_io_out_1),
    .io_out_2(c53_332_io_out_2)
  );
  C53 c53_333 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_333_io_in_0),
    .io_in_1(c53_333_io_in_1),
    .io_in_2(c53_333_io_in_2),
    .io_in_3(c53_333_io_in_3),
    .io_in_4(c53_333_io_in_4),
    .io_out_0(c53_333_io_out_0),
    .io_out_1(c53_333_io_out_1),
    .io_out_2(c53_333_io_out_2)
  );
  C53 c53_334 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_334_io_in_0),
    .io_in_1(c53_334_io_in_1),
    .io_in_2(c53_334_io_in_2),
    .io_in_3(c53_334_io_in_3),
    .io_in_4(c53_334_io_in_4),
    .io_out_0(c53_334_io_out_0),
    .io_out_1(c53_334_io_out_1),
    .io_out_2(c53_334_io_out_2)
  );
  C53 c53_335 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_335_io_in_0),
    .io_in_1(c53_335_io_in_1),
    .io_in_2(c53_335_io_in_2),
    .io_in_3(c53_335_io_in_3),
    .io_in_4(c53_335_io_in_4),
    .io_out_0(c53_335_io_out_0),
    .io_out_1(c53_335_io_out_1),
    .io_out_2(c53_335_io_out_2)
  );
  C53 c53_336 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_336_io_in_0),
    .io_in_1(c53_336_io_in_1),
    .io_in_2(c53_336_io_in_2),
    .io_in_3(c53_336_io_in_3),
    .io_in_4(c53_336_io_in_4),
    .io_out_0(c53_336_io_out_0),
    .io_out_1(c53_336_io_out_1),
    .io_out_2(c53_336_io_out_2)
  );
  C53 c53_337 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_337_io_in_0),
    .io_in_1(c53_337_io_in_1),
    .io_in_2(c53_337_io_in_2),
    .io_in_3(c53_337_io_in_3),
    .io_in_4(c53_337_io_in_4),
    .io_out_0(c53_337_io_out_0),
    .io_out_1(c53_337_io_out_1),
    .io_out_2(c53_337_io_out_2)
  );
  C53 c53_338 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_338_io_in_0),
    .io_in_1(c53_338_io_in_1),
    .io_in_2(c53_338_io_in_2),
    .io_in_3(c53_338_io_in_3),
    .io_in_4(c53_338_io_in_4),
    .io_out_0(c53_338_io_out_0),
    .io_out_1(c53_338_io_out_1),
    .io_out_2(c53_338_io_out_2)
  );
  C53 c53_339 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_339_io_in_0),
    .io_in_1(c53_339_io_in_1),
    .io_in_2(c53_339_io_in_2),
    .io_in_3(c53_339_io_in_3),
    .io_in_4(c53_339_io_in_4),
    .io_out_0(c53_339_io_out_0),
    .io_out_1(c53_339_io_out_1),
    .io_out_2(c53_339_io_out_2)
  );
  C53 c53_340 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_340_io_in_0),
    .io_in_1(c53_340_io_in_1),
    .io_in_2(c53_340_io_in_2),
    .io_in_3(c53_340_io_in_3),
    .io_in_4(c53_340_io_in_4),
    .io_out_0(c53_340_io_out_0),
    .io_out_1(c53_340_io_out_1),
    .io_out_2(c53_340_io_out_2)
  );
  C53 c53_341 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_341_io_in_0),
    .io_in_1(c53_341_io_in_1),
    .io_in_2(c53_341_io_in_2),
    .io_in_3(c53_341_io_in_3),
    .io_in_4(c53_341_io_in_4),
    .io_out_0(c53_341_io_out_0),
    .io_out_1(c53_341_io_out_1),
    .io_out_2(c53_341_io_out_2)
  );
  C53 c53_342 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_342_io_in_0),
    .io_in_1(c53_342_io_in_1),
    .io_in_2(c53_342_io_in_2),
    .io_in_3(c53_342_io_in_3),
    .io_in_4(c53_342_io_in_4),
    .io_out_0(c53_342_io_out_0),
    .io_out_1(c53_342_io_out_1),
    .io_out_2(c53_342_io_out_2)
  );
  C53 c53_343 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_343_io_in_0),
    .io_in_1(c53_343_io_in_1),
    .io_in_2(c53_343_io_in_2),
    .io_in_3(c53_343_io_in_3),
    .io_in_4(c53_343_io_in_4),
    .io_out_0(c53_343_io_out_0),
    .io_out_1(c53_343_io_out_1),
    .io_out_2(c53_343_io_out_2)
  );
  C53 c53_344 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_344_io_in_0),
    .io_in_1(c53_344_io_in_1),
    .io_in_2(c53_344_io_in_2),
    .io_in_3(c53_344_io_in_3),
    .io_in_4(c53_344_io_in_4),
    .io_out_0(c53_344_io_out_0),
    .io_out_1(c53_344_io_out_1),
    .io_out_2(c53_344_io_out_2)
  );
  C53 c53_345 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_345_io_in_0),
    .io_in_1(c53_345_io_in_1),
    .io_in_2(c53_345_io_in_2),
    .io_in_3(c53_345_io_in_3),
    .io_in_4(c53_345_io_in_4),
    .io_out_0(c53_345_io_out_0),
    .io_out_1(c53_345_io_out_1),
    .io_out_2(c53_345_io_out_2)
  );
  C53 c53_346 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_346_io_in_0),
    .io_in_1(c53_346_io_in_1),
    .io_in_2(c53_346_io_in_2),
    .io_in_3(c53_346_io_in_3),
    .io_in_4(c53_346_io_in_4),
    .io_out_0(c53_346_io_out_0),
    .io_out_1(c53_346_io_out_1),
    .io_out_2(c53_346_io_out_2)
  );
  C53 c53_347 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_347_io_in_0),
    .io_in_1(c53_347_io_in_1),
    .io_in_2(c53_347_io_in_2),
    .io_in_3(c53_347_io_in_3),
    .io_in_4(c53_347_io_in_4),
    .io_out_0(c53_347_io_out_0),
    .io_out_1(c53_347_io_out_1),
    .io_out_2(c53_347_io_out_2)
  );
  C53 c53_348 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_348_io_in_0),
    .io_in_1(c53_348_io_in_1),
    .io_in_2(c53_348_io_in_2),
    .io_in_3(c53_348_io_in_3),
    .io_in_4(c53_348_io_in_4),
    .io_out_0(c53_348_io_out_0),
    .io_out_1(c53_348_io_out_1),
    .io_out_2(c53_348_io_out_2)
  );
  C53 c53_349 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_349_io_in_0),
    .io_in_1(c53_349_io_in_1),
    .io_in_2(c53_349_io_in_2),
    .io_in_3(c53_349_io_in_3),
    .io_in_4(c53_349_io_in_4),
    .io_out_0(c53_349_io_out_0),
    .io_out_1(c53_349_io_out_1),
    .io_out_2(c53_349_io_out_2)
  );
  C53 c53_350 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_350_io_in_0),
    .io_in_1(c53_350_io_in_1),
    .io_in_2(c53_350_io_in_2),
    .io_in_3(c53_350_io_in_3),
    .io_in_4(c53_350_io_in_4),
    .io_out_0(c53_350_io_out_0),
    .io_out_1(c53_350_io_out_1),
    .io_out_2(c53_350_io_out_2)
  );
  C53 c53_351 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_351_io_in_0),
    .io_in_1(c53_351_io_in_1),
    .io_in_2(c53_351_io_in_2),
    .io_in_3(c53_351_io_in_3),
    .io_in_4(c53_351_io_in_4),
    .io_out_0(c53_351_io_out_0),
    .io_out_1(c53_351_io_out_1),
    .io_out_2(c53_351_io_out_2)
  );
  C53 c53_352 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_352_io_in_0),
    .io_in_1(c53_352_io_in_1),
    .io_in_2(c53_352_io_in_2),
    .io_in_3(c53_352_io_in_3),
    .io_in_4(c53_352_io_in_4),
    .io_out_0(c53_352_io_out_0),
    .io_out_1(c53_352_io_out_1),
    .io_out_2(c53_352_io_out_2)
  );
  C53 c53_353 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_353_io_in_0),
    .io_in_1(c53_353_io_in_1),
    .io_in_2(c53_353_io_in_2),
    .io_in_3(c53_353_io_in_3),
    .io_in_4(c53_353_io_in_4),
    .io_out_0(c53_353_io_out_0),
    .io_out_1(c53_353_io_out_1),
    .io_out_2(c53_353_io_out_2)
  );
  C53 c53_354 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_354_io_in_0),
    .io_in_1(c53_354_io_in_1),
    .io_in_2(c53_354_io_in_2),
    .io_in_3(c53_354_io_in_3),
    .io_in_4(c53_354_io_in_4),
    .io_out_0(c53_354_io_out_0),
    .io_out_1(c53_354_io_out_1),
    .io_out_2(c53_354_io_out_2)
  );
  C53 c53_355 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_355_io_in_0),
    .io_in_1(c53_355_io_in_1),
    .io_in_2(c53_355_io_in_2),
    .io_in_3(c53_355_io_in_3),
    .io_in_4(c53_355_io_in_4),
    .io_out_0(c53_355_io_out_0),
    .io_out_1(c53_355_io_out_1),
    .io_out_2(c53_355_io_out_2)
  );
  C53 c53_356 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_356_io_in_0),
    .io_in_1(c53_356_io_in_1),
    .io_in_2(c53_356_io_in_2),
    .io_in_3(c53_356_io_in_3),
    .io_in_4(c53_356_io_in_4),
    .io_out_0(c53_356_io_out_0),
    .io_out_1(c53_356_io_out_1),
    .io_out_2(c53_356_io_out_2)
  );
  C53 c53_357 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_357_io_in_0),
    .io_in_1(c53_357_io_in_1),
    .io_in_2(c53_357_io_in_2),
    .io_in_3(c53_357_io_in_3),
    .io_in_4(c53_357_io_in_4),
    .io_out_0(c53_357_io_out_0),
    .io_out_1(c53_357_io_out_1),
    .io_out_2(c53_357_io_out_2)
  );
  C53 c53_358 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_358_io_in_0),
    .io_in_1(c53_358_io_in_1),
    .io_in_2(c53_358_io_in_2),
    .io_in_3(c53_358_io_in_3),
    .io_in_4(c53_358_io_in_4),
    .io_out_0(c53_358_io_out_0),
    .io_out_1(c53_358_io_out_1),
    .io_out_2(c53_358_io_out_2)
  );
  C53 c53_359 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_359_io_in_0),
    .io_in_1(c53_359_io_in_1),
    .io_in_2(c53_359_io_in_2),
    .io_in_3(c53_359_io_in_3),
    .io_in_4(c53_359_io_in_4),
    .io_out_0(c53_359_io_out_0),
    .io_out_1(c53_359_io_out_1),
    .io_out_2(c53_359_io_out_2)
  );
  C53 c53_360 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_360_io_in_0),
    .io_in_1(c53_360_io_in_1),
    .io_in_2(c53_360_io_in_2),
    .io_in_3(c53_360_io_in_3),
    .io_in_4(c53_360_io_in_4),
    .io_out_0(c53_360_io_out_0),
    .io_out_1(c53_360_io_out_1),
    .io_out_2(c53_360_io_out_2)
  );
  C53 c53_361 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_361_io_in_0),
    .io_in_1(c53_361_io_in_1),
    .io_in_2(c53_361_io_in_2),
    .io_in_3(c53_361_io_in_3),
    .io_in_4(c53_361_io_in_4),
    .io_out_0(c53_361_io_out_0),
    .io_out_1(c53_361_io_out_1),
    .io_out_2(c53_361_io_out_2)
  );
  C53 c53_362 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_362_io_in_0),
    .io_in_1(c53_362_io_in_1),
    .io_in_2(c53_362_io_in_2),
    .io_in_3(c53_362_io_in_3),
    .io_in_4(c53_362_io_in_4),
    .io_out_0(c53_362_io_out_0),
    .io_out_1(c53_362_io_out_1),
    .io_out_2(c53_362_io_out_2)
  );
  C53 c53_363 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_363_io_in_0),
    .io_in_1(c53_363_io_in_1),
    .io_in_2(c53_363_io_in_2),
    .io_in_3(c53_363_io_in_3),
    .io_in_4(c53_363_io_in_4),
    .io_out_0(c53_363_io_out_0),
    .io_out_1(c53_363_io_out_1),
    .io_out_2(c53_363_io_out_2)
  );
  C53 c53_364 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_364_io_in_0),
    .io_in_1(c53_364_io_in_1),
    .io_in_2(c53_364_io_in_2),
    .io_in_3(c53_364_io_in_3),
    .io_in_4(c53_364_io_in_4),
    .io_out_0(c53_364_io_out_0),
    .io_out_1(c53_364_io_out_1),
    .io_out_2(c53_364_io_out_2)
  );
  C53 c53_365 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_365_io_in_0),
    .io_in_1(c53_365_io_in_1),
    .io_in_2(c53_365_io_in_2),
    .io_in_3(c53_365_io_in_3),
    .io_in_4(c53_365_io_in_4),
    .io_out_0(c53_365_io_out_0),
    .io_out_1(c53_365_io_out_1),
    .io_out_2(c53_365_io_out_2)
  );
  C32 c32_18 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_18_io_in_0),
    .io_in_1(c32_18_io_in_1),
    .io_in_2(c32_18_io_in_2),
    .io_out_0(c32_18_io_out_0),
    .io_out_1(c32_18_io_out_1)
  );
  C53 c53_366 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_366_io_in_0),
    .io_in_1(c53_366_io_in_1),
    .io_in_2(c53_366_io_in_2),
    .io_in_3(c53_366_io_in_3),
    .io_in_4(c53_366_io_in_4),
    .io_out_0(c53_366_io_out_0),
    .io_out_1(c53_366_io_out_1),
    .io_out_2(c53_366_io_out_2)
  );
  C53 c53_367 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_367_io_in_0),
    .io_in_1(c53_367_io_in_1),
    .io_in_2(c53_367_io_in_2),
    .io_in_3(c53_367_io_in_3),
    .io_in_4(c53_367_io_in_4),
    .io_out_0(c53_367_io_out_0),
    .io_out_1(c53_367_io_out_1),
    .io_out_2(c53_367_io_out_2)
  );
  C53 c53_368 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_368_io_in_0),
    .io_in_1(c53_368_io_in_1),
    .io_in_2(c53_368_io_in_2),
    .io_in_3(c53_368_io_in_3),
    .io_in_4(c53_368_io_in_4),
    .io_out_0(c53_368_io_out_0),
    .io_out_1(c53_368_io_out_1),
    .io_out_2(c53_368_io_out_2)
  );
  C53 c53_369 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_369_io_in_0),
    .io_in_1(c53_369_io_in_1),
    .io_in_2(c53_369_io_in_2),
    .io_in_3(c53_369_io_in_3),
    .io_in_4(c53_369_io_in_4),
    .io_out_0(c53_369_io_out_0),
    .io_out_1(c53_369_io_out_1),
    .io_out_2(c53_369_io_out_2)
  );
  C53 c53_370 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_370_io_in_0),
    .io_in_1(c53_370_io_in_1),
    .io_in_2(c53_370_io_in_2),
    .io_in_3(c53_370_io_in_3),
    .io_in_4(c53_370_io_in_4),
    .io_out_0(c53_370_io_out_0),
    .io_out_1(c53_370_io_out_1),
    .io_out_2(c53_370_io_out_2)
  );
  C53 c53_371 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_371_io_in_0),
    .io_in_1(c53_371_io_in_1),
    .io_in_2(c53_371_io_in_2),
    .io_in_3(c53_371_io_in_3),
    .io_in_4(c53_371_io_in_4),
    .io_out_0(c53_371_io_out_0),
    .io_out_1(c53_371_io_out_1),
    .io_out_2(c53_371_io_out_2)
  );
  C32 c32_19 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_19_io_in_0),
    .io_in_1(c32_19_io_in_1),
    .io_in_2(c32_19_io_in_2),
    .io_out_0(c32_19_io_out_0),
    .io_out_1(c32_19_io_out_1)
  );
  C53 c53_372 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_372_io_in_0),
    .io_in_1(c53_372_io_in_1),
    .io_in_2(c53_372_io_in_2),
    .io_in_3(c53_372_io_in_3),
    .io_in_4(c53_372_io_in_4),
    .io_out_0(c53_372_io_out_0),
    .io_out_1(c53_372_io_out_1),
    .io_out_2(c53_372_io_out_2)
  );
  C53 c53_373 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_373_io_in_0),
    .io_in_1(c53_373_io_in_1),
    .io_in_2(c53_373_io_in_2),
    .io_in_3(c53_373_io_in_3),
    .io_in_4(c53_373_io_in_4),
    .io_out_0(c53_373_io_out_0),
    .io_out_1(c53_373_io_out_1),
    .io_out_2(c53_373_io_out_2)
  );
  C53 c53_374 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_374_io_in_0),
    .io_in_1(c53_374_io_in_1),
    .io_in_2(c53_374_io_in_2),
    .io_in_3(c53_374_io_in_3),
    .io_in_4(c53_374_io_in_4),
    .io_out_0(c53_374_io_out_0),
    .io_out_1(c53_374_io_out_1),
    .io_out_2(c53_374_io_out_2)
  );
  C53 c53_375 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_375_io_in_0),
    .io_in_1(c53_375_io_in_1),
    .io_in_2(c53_375_io_in_2),
    .io_in_3(c53_375_io_in_3),
    .io_in_4(c53_375_io_in_4),
    .io_out_0(c53_375_io_out_0),
    .io_out_1(c53_375_io_out_1),
    .io_out_2(c53_375_io_out_2)
  );
  C53 c53_376 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_376_io_in_0),
    .io_in_1(c53_376_io_in_1),
    .io_in_2(c53_376_io_in_2),
    .io_in_3(c53_376_io_in_3),
    .io_in_4(c53_376_io_in_4),
    .io_out_0(c53_376_io_out_0),
    .io_out_1(c53_376_io_out_1),
    .io_out_2(c53_376_io_out_2)
  );
  C53 c53_377 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_377_io_in_0),
    .io_in_1(c53_377_io_in_1),
    .io_in_2(c53_377_io_in_2),
    .io_in_3(c53_377_io_in_3),
    .io_in_4(c53_377_io_in_4),
    .io_out_0(c53_377_io_out_0),
    .io_out_1(c53_377_io_out_1),
    .io_out_2(c53_377_io_out_2)
  );
  C22 c22_18 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_18_io_in_0),
    .io_in_1(c22_18_io_in_1),
    .io_out_0(c22_18_io_out_0),
    .io_out_1(c22_18_io_out_1)
  );
  C53 c53_378 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_378_io_in_0),
    .io_in_1(c53_378_io_in_1),
    .io_in_2(c53_378_io_in_2),
    .io_in_3(c53_378_io_in_3),
    .io_in_4(c53_378_io_in_4),
    .io_out_0(c53_378_io_out_0),
    .io_out_1(c53_378_io_out_1),
    .io_out_2(c53_378_io_out_2)
  );
  C53 c53_379 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_379_io_in_0),
    .io_in_1(c53_379_io_in_1),
    .io_in_2(c53_379_io_in_2),
    .io_in_3(c53_379_io_in_3),
    .io_in_4(c53_379_io_in_4),
    .io_out_0(c53_379_io_out_0),
    .io_out_1(c53_379_io_out_1),
    .io_out_2(c53_379_io_out_2)
  );
  C53 c53_380 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_380_io_in_0),
    .io_in_1(c53_380_io_in_1),
    .io_in_2(c53_380_io_in_2),
    .io_in_3(c53_380_io_in_3),
    .io_in_4(c53_380_io_in_4),
    .io_out_0(c53_380_io_out_0),
    .io_out_1(c53_380_io_out_1),
    .io_out_2(c53_380_io_out_2)
  );
  C53 c53_381 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_381_io_in_0),
    .io_in_1(c53_381_io_in_1),
    .io_in_2(c53_381_io_in_2),
    .io_in_3(c53_381_io_in_3),
    .io_in_4(c53_381_io_in_4),
    .io_out_0(c53_381_io_out_0),
    .io_out_1(c53_381_io_out_1),
    .io_out_2(c53_381_io_out_2)
  );
  C53 c53_382 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_382_io_in_0),
    .io_in_1(c53_382_io_in_1),
    .io_in_2(c53_382_io_in_2),
    .io_in_3(c53_382_io_in_3),
    .io_in_4(c53_382_io_in_4),
    .io_out_0(c53_382_io_out_0),
    .io_out_1(c53_382_io_out_1),
    .io_out_2(c53_382_io_out_2)
  );
  C53 c53_383 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_383_io_in_0),
    .io_in_1(c53_383_io_in_1),
    .io_in_2(c53_383_io_in_2),
    .io_in_3(c53_383_io_in_3),
    .io_in_4(c53_383_io_in_4),
    .io_out_0(c53_383_io_out_0),
    .io_out_1(c53_383_io_out_1),
    .io_out_2(c53_383_io_out_2)
  );
  C22 c22_19 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_19_io_in_0),
    .io_in_1(c22_19_io_in_1),
    .io_out_0(c22_19_io_out_0),
    .io_out_1(c22_19_io_out_1)
  );
  C53 c53_384 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_384_io_in_0),
    .io_in_1(c53_384_io_in_1),
    .io_in_2(c53_384_io_in_2),
    .io_in_3(c53_384_io_in_3),
    .io_in_4(c53_384_io_in_4),
    .io_out_0(c53_384_io_out_0),
    .io_out_1(c53_384_io_out_1),
    .io_out_2(c53_384_io_out_2)
  );
  C53 c53_385 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_385_io_in_0),
    .io_in_1(c53_385_io_in_1),
    .io_in_2(c53_385_io_in_2),
    .io_in_3(c53_385_io_in_3),
    .io_in_4(c53_385_io_in_4),
    .io_out_0(c53_385_io_out_0),
    .io_out_1(c53_385_io_out_1),
    .io_out_2(c53_385_io_out_2)
  );
  C53 c53_386 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_386_io_in_0),
    .io_in_1(c53_386_io_in_1),
    .io_in_2(c53_386_io_in_2),
    .io_in_3(c53_386_io_in_3),
    .io_in_4(c53_386_io_in_4),
    .io_out_0(c53_386_io_out_0),
    .io_out_1(c53_386_io_out_1),
    .io_out_2(c53_386_io_out_2)
  );
  C53 c53_387 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_387_io_in_0),
    .io_in_1(c53_387_io_in_1),
    .io_in_2(c53_387_io_in_2),
    .io_in_3(c53_387_io_in_3),
    .io_in_4(c53_387_io_in_4),
    .io_out_0(c53_387_io_out_0),
    .io_out_1(c53_387_io_out_1),
    .io_out_2(c53_387_io_out_2)
  );
  C53 c53_388 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_388_io_in_0),
    .io_in_1(c53_388_io_in_1),
    .io_in_2(c53_388_io_in_2),
    .io_in_3(c53_388_io_in_3),
    .io_in_4(c53_388_io_in_4),
    .io_out_0(c53_388_io_out_0),
    .io_out_1(c53_388_io_out_1),
    .io_out_2(c53_388_io_out_2)
  );
  C53 c53_389 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_389_io_in_0),
    .io_in_1(c53_389_io_in_1),
    .io_in_2(c53_389_io_in_2),
    .io_in_3(c53_389_io_in_3),
    .io_in_4(c53_389_io_in_4),
    .io_out_0(c53_389_io_out_0),
    .io_out_1(c53_389_io_out_1),
    .io_out_2(c53_389_io_out_2)
  );
  C53 c53_390 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_390_io_in_0),
    .io_in_1(c53_390_io_in_1),
    .io_in_2(c53_390_io_in_2),
    .io_in_3(c53_390_io_in_3),
    .io_in_4(c53_390_io_in_4),
    .io_out_0(c53_390_io_out_0),
    .io_out_1(c53_390_io_out_1),
    .io_out_2(c53_390_io_out_2)
  );
  C53 c53_391 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_391_io_in_0),
    .io_in_1(c53_391_io_in_1),
    .io_in_2(c53_391_io_in_2),
    .io_in_3(c53_391_io_in_3),
    .io_in_4(c53_391_io_in_4),
    .io_out_0(c53_391_io_out_0),
    .io_out_1(c53_391_io_out_1),
    .io_out_2(c53_391_io_out_2)
  );
  C53 c53_392 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_392_io_in_0),
    .io_in_1(c53_392_io_in_1),
    .io_in_2(c53_392_io_in_2),
    .io_in_3(c53_392_io_in_3),
    .io_in_4(c53_392_io_in_4),
    .io_out_0(c53_392_io_out_0),
    .io_out_1(c53_392_io_out_1),
    .io_out_2(c53_392_io_out_2)
  );
  C53 c53_393 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_393_io_in_0),
    .io_in_1(c53_393_io_in_1),
    .io_in_2(c53_393_io_in_2),
    .io_in_3(c53_393_io_in_3),
    .io_in_4(c53_393_io_in_4),
    .io_out_0(c53_393_io_out_0),
    .io_out_1(c53_393_io_out_1),
    .io_out_2(c53_393_io_out_2)
  );
  C53 c53_394 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_394_io_in_0),
    .io_in_1(c53_394_io_in_1),
    .io_in_2(c53_394_io_in_2),
    .io_in_3(c53_394_io_in_3),
    .io_in_4(c53_394_io_in_4),
    .io_out_0(c53_394_io_out_0),
    .io_out_1(c53_394_io_out_1),
    .io_out_2(c53_394_io_out_2)
  );
  C53 c53_395 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_395_io_in_0),
    .io_in_1(c53_395_io_in_1),
    .io_in_2(c53_395_io_in_2),
    .io_in_3(c53_395_io_in_3),
    .io_in_4(c53_395_io_in_4),
    .io_out_0(c53_395_io_out_0),
    .io_out_1(c53_395_io_out_1),
    .io_out_2(c53_395_io_out_2)
  );
  C53 c53_396 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_396_io_in_0),
    .io_in_1(c53_396_io_in_1),
    .io_in_2(c53_396_io_in_2),
    .io_in_3(c53_396_io_in_3),
    .io_in_4(c53_396_io_in_4),
    .io_out_0(c53_396_io_out_0),
    .io_out_1(c53_396_io_out_1),
    .io_out_2(c53_396_io_out_2)
  );
  C53 c53_397 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_397_io_in_0),
    .io_in_1(c53_397_io_in_1),
    .io_in_2(c53_397_io_in_2),
    .io_in_3(c53_397_io_in_3),
    .io_in_4(c53_397_io_in_4),
    .io_out_0(c53_397_io_out_0),
    .io_out_1(c53_397_io_out_1),
    .io_out_2(c53_397_io_out_2)
  );
  C53 c53_398 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_398_io_in_0),
    .io_in_1(c53_398_io_in_1),
    .io_in_2(c53_398_io_in_2),
    .io_in_3(c53_398_io_in_3),
    .io_in_4(c53_398_io_in_4),
    .io_out_0(c53_398_io_out_0),
    .io_out_1(c53_398_io_out_1),
    .io_out_2(c53_398_io_out_2)
  );
  C53 c53_399 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_399_io_in_0),
    .io_in_1(c53_399_io_in_1),
    .io_in_2(c53_399_io_in_2),
    .io_in_3(c53_399_io_in_3),
    .io_in_4(c53_399_io_in_4),
    .io_out_0(c53_399_io_out_0),
    .io_out_1(c53_399_io_out_1),
    .io_out_2(c53_399_io_out_2)
  );
  C53 c53_400 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_400_io_in_0),
    .io_in_1(c53_400_io_in_1),
    .io_in_2(c53_400_io_in_2),
    .io_in_3(c53_400_io_in_3),
    .io_in_4(c53_400_io_in_4),
    .io_out_0(c53_400_io_out_0),
    .io_out_1(c53_400_io_out_1),
    .io_out_2(c53_400_io_out_2)
  );
  C53 c53_401 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_401_io_in_0),
    .io_in_1(c53_401_io_in_1),
    .io_in_2(c53_401_io_in_2),
    .io_in_3(c53_401_io_in_3),
    .io_in_4(c53_401_io_in_4),
    .io_out_0(c53_401_io_out_0),
    .io_out_1(c53_401_io_out_1),
    .io_out_2(c53_401_io_out_2)
  );
  C53 c53_402 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_402_io_in_0),
    .io_in_1(c53_402_io_in_1),
    .io_in_2(c53_402_io_in_2),
    .io_in_3(c53_402_io_in_3),
    .io_in_4(c53_402_io_in_4),
    .io_out_0(c53_402_io_out_0),
    .io_out_1(c53_402_io_out_1),
    .io_out_2(c53_402_io_out_2)
  );
  C53 c53_403 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_403_io_in_0),
    .io_in_1(c53_403_io_in_1),
    .io_in_2(c53_403_io_in_2),
    .io_in_3(c53_403_io_in_3),
    .io_in_4(c53_403_io_in_4),
    .io_out_0(c53_403_io_out_0),
    .io_out_1(c53_403_io_out_1),
    .io_out_2(c53_403_io_out_2)
  );
  C53 c53_404 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_404_io_in_0),
    .io_in_1(c53_404_io_in_1),
    .io_in_2(c53_404_io_in_2),
    .io_in_3(c53_404_io_in_3),
    .io_in_4(c53_404_io_in_4),
    .io_out_0(c53_404_io_out_0),
    .io_out_1(c53_404_io_out_1),
    .io_out_2(c53_404_io_out_2)
  );
  C53 c53_405 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_405_io_in_0),
    .io_in_1(c53_405_io_in_1),
    .io_in_2(c53_405_io_in_2),
    .io_in_3(c53_405_io_in_3),
    .io_in_4(c53_405_io_in_4),
    .io_out_0(c53_405_io_out_0),
    .io_out_1(c53_405_io_out_1),
    .io_out_2(c53_405_io_out_2)
  );
  C53 c53_406 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_406_io_in_0),
    .io_in_1(c53_406_io_in_1),
    .io_in_2(c53_406_io_in_2),
    .io_in_3(c53_406_io_in_3),
    .io_in_4(c53_406_io_in_4),
    .io_out_0(c53_406_io_out_0),
    .io_out_1(c53_406_io_out_1),
    .io_out_2(c53_406_io_out_2)
  );
  C53 c53_407 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_407_io_in_0),
    .io_in_1(c53_407_io_in_1),
    .io_in_2(c53_407_io_in_2),
    .io_in_3(c53_407_io_in_3),
    .io_in_4(c53_407_io_in_4),
    .io_out_0(c53_407_io_out_0),
    .io_out_1(c53_407_io_out_1),
    .io_out_2(c53_407_io_out_2)
  );
  C53 c53_408 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_408_io_in_0),
    .io_in_1(c53_408_io_in_1),
    .io_in_2(c53_408_io_in_2),
    .io_in_3(c53_408_io_in_3),
    .io_in_4(c53_408_io_in_4),
    .io_out_0(c53_408_io_out_0),
    .io_out_1(c53_408_io_out_1),
    .io_out_2(c53_408_io_out_2)
  );
  C53 c53_409 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_409_io_in_0),
    .io_in_1(c53_409_io_in_1),
    .io_in_2(c53_409_io_in_2),
    .io_in_3(c53_409_io_in_3),
    .io_in_4(c53_409_io_in_4),
    .io_out_0(c53_409_io_out_0),
    .io_out_1(c53_409_io_out_1),
    .io_out_2(c53_409_io_out_2)
  );
  C53 c53_410 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_410_io_in_0),
    .io_in_1(c53_410_io_in_1),
    .io_in_2(c53_410_io_in_2),
    .io_in_3(c53_410_io_in_3),
    .io_in_4(c53_410_io_in_4),
    .io_out_0(c53_410_io_out_0),
    .io_out_1(c53_410_io_out_1),
    .io_out_2(c53_410_io_out_2)
  );
  C53 c53_411 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_411_io_in_0),
    .io_in_1(c53_411_io_in_1),
    .io_in_2(c53_411_io_in_2),
    .io_in_3(c53_411_io_in_3),
    .io_in_4(c53_411_io_in_4),
    .io_out_0(c53_411_io_out_0),
    .io_out_1(c53_411_io_out_1),
    .io_out_2(c53_411_io_out_2)
  );
  C53 c53_412 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_412_io_in_0),
    .io_in_1(c53_412_io_in_1),
    .io_in_2(c53_412_io_in_2),
    .io_in_3(c53_412_io_in_3),
    .io_in_4(c53_412_io_in_4),
    .io_out_0(c53_412_io_out_0),
    .io_out_1(c53_412_io_out_1),
    .io_out_2(c53_412_io_out_2)
  );
  C32 c32_20 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_20_io_in_0),
    .io_in_1(c32_20_io_in_1),
    .io_in_2(c32_20_io_in_2),
    .io_out_0(c32_20_io_out_0),
    .io_out_1(c32_20_io_out_1)
  );
  C53 c53_413 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_413_io_in_0),
    .io_in_1(c53_413_io_in_1),
    .io_in_2(c53_413_io_in_2),
    .io_in_3(c53_413_io_in_3),
    .io_in_4(c53_413_io_in_4),
    .io_out_0(c53_413_io_out_0),
    .io_out_1(c53_413_io_out_1),
    .io_out_2(c53_413_io_out_2)
  );
  C53 c53_414 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_414_io_in_0),
    .io_in_1(c53_414_io_in_1),
    .io_in_2(c53_414_io_in_2),
    .io_in_3(c53_414_io_in_3),
    .io_in_4(c53_414_io_in_4),
    .io_out_0(c53_414_io_out_0),
    .io_out_1(c53_414_io_out_1),
    .io_out_2(c53_414_io_out_2)
  );
  C53 c53_415 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_415_io_in_0),
    .io_in_1(c53_415_io_in_1),
    .io_in_2(c53_415_io_in_2),
    .io_in_3(c53_415_io_in_3),
    .io_in_4(c53_415_io_in_4),
    .io_out_0(c53_415_io_out_0),
    .io_out_1(c53_415_io_out_1),
    .io_out_2(c53_415_io_out_2)
  );
  C53 c53_416 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_416_io_in_0),
    .io_in_1(c53_416_io_in_1),
    .io_in_2(c53_416_io_in_2),
    .io_in_3(c53_416_io_in_3),
    .io_in_4(c53_416_io_in_4),
    .io_out_0(c53_416_io_out_0),
    .io_out_1(c53_416_io_out_1),
    .io_out_2(c53_416_io_out_2)
  );
  C53 c53_417 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_417_io_in_0),
    .io_in_1(c53_417_io_in_1),
    .io_in_2(c53_417_io_in_2),
    .io_in_3(c53_417_io_in_3),
    .io_in_4(c53_417_io_in_4),
    .io_out_0(c53_417_io_out_0),
    .io_out_1(c53_417_io_out_1),
    .io_out_2(c53_417_io_out_2)
  );
  C32 c32_21 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_21_io_in_0),
    .io_in_1(c32_21_io_in_1),
    .io_in_2(c32_21_io_in_2),
    .io_out_0(c32_21_io_out_0),
    .io_out_1(c32_21_io_out_1)
  );
  C53 c53_418 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_418_io_in_0),
    .io_in_1(c53_418_io_in_1),
    .io_in_2(c53_418_io_in_2),
    .io_in_3(c53_418_io_in_3),
    .io_in_4(c53_418_io_in_4),
    .io_out_0(c53_418_io_out_0),
    .io_out_1(c53_418_io_out_1),
    .io_out_2(c53_418_io_out_2)
  );
  C53 c53_419 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_419_io_in_0),
    .io_in_1(c53_419_io_in_1),
    .io_in_2(c53_419_io_in_2),
    .io_in_3(c53_419_io_in_3),
    .io_in_4(c53_419_io_in_4),
    .io_out_0(c53_419_io_out_0),
    .io_out_1(c53_419_io_out_1),
    .io_out_2(c53_419_io_out_2)
  );
  C53 c53_420 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_420_io_in_0),
    .io_in_1(c53_420_io_in_1),
    .io_in_2(c53_420_io_in_2),
    .io_in_3(c53_420_io_in_3),
    .io_in_4(c53_420_io_in_4),
    .io_out_0(c53_420_io_out_0),
    .io_out_1(c53_420_io_out_1),
    .io_out_2(c53_420_io_out_2)
  );
  C53 c53_421 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_421_io_in_0),
    .io_in_1(c53_421_io_in_1),
    .io_in_2(c53_421_io_in_2),
    .io_in_3(c53_421_io_in_3),
    .io_in_4(c53_421_io_in_4),
    .io_out_0(c53_421_io_out_0),
    .io_out_1(c53_421_io_out_1),
    .io_out_2(c53_421_io_out_2)
  );
  C53 c53_422 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_422_io_in_0),
    .io_in_1(c53_422_io_in_1),
    .io_in_2(c53_422_io_in_2),
    .io_in_3(c53_422_io_in_3),
    .io_in_4(c53_422_io_in_4),
    .io_out_0(c53_422_io_out_0),
    .io_out_1(c53_422_io_out_1),
    .io_out_2(c53_422_io_out_2)
  );
  C22 c22_20 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_20_io_in_0),
    .io_in_1(c22_20_io_in_1),
    .io_out_0(c22_20_io_out_0),
    .io_out_1(c22_20_io_out_1)
  );
  C53 c53_423 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_423_io_in_0),
    .io_in_1(c53_423_io_in_1),
    .io_in_2(c53_423_io_in_2),
    .io_in_3(c53_423_io_in_3),
    .io_in_4(c53_423_io_in_4),
    .io_out_0(c53_423_io_out_0),
    .io_out_1(c53_423_io_out_1),
    .io_out_2(c53_423_io_out_2)
  );
  C53 c53_424 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_424_io_in_0),
    .io_in_1(c53_424_io_in_1),
    .io_in_2(c53_424_io_in_2),
    .io_in_3(c53_424_io_in_3),
    .io_in_4(c53_424_io_in_4),
    .io_out_0(c53_424_io_out_0),
    .io_out_1(c53_424_io_out_1),
    .io_out_2(c53_424_io_out_2)
  );
  C53 c53_425 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_425_io_in_0),
    .io_in_1(c53_425_io_in_1),
    .io_in_2(c53_425_io_in_2),
    .io_in_3(c53_425_io_in_3),
    .io_in_4(c53_425_io_in_4),
    .io_out_0(c53_425_io_out_0),
    .io_out_1(c53_425_io_out_1),
    .io_out_2(c53_425_io_out_2)
  );
  C53 c53_426 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_426_io_in_0),
    .io_in_1(c53_426_io_in_1),
    .io_in_2(c53_426_io_in_2),
    .io_in_3(c53_426_io_in_3),
    .io_in_4(c53_426_io_in_4),
    .io_out_0(c53_426_io_out_0),
    .io_out_1(c53_426_io_out_1),
    .io_out_2(c53_426_io_out_2)
  );
  C53 c53_427 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_427_io_in_0),
    .io_in_1(c53_427_io_in_1),
    .io_in_2(c53_427_io_in_2),
    .io_in_3(c53_427_io_in_3),
    .io_in_4(c53_427_io_in_4),
    .io_out_0(c53_427_io_out_0),
    .io_out_1(c53_427_io_out_1),
    .io_out_2(c53_427_io_out_2)
  );
  C22 c22_21 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_21_io_in_0),
    .io_in_1(c22_21_io_in_1),
    .io_out_0(c22_21_io_out_0),
    .io_out_1(c22_21_io_out_1)
  );
  C53 c53_428 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_428_io_in_0),
    .io_in_1(c53_428_io_in_1),
    .io_in_2(c53_428_io_in_2),
    .io_in_3(c53_428_io_in_3),
    .io_in_4(c53_428_io_in_4),
    .io_out_0(c53_428_io_out_0),
    .io_out_1(c53_428_io_out_1),
    .io_out_2(c53_428_io_out_2)
  );
  C53 c53_429 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_429_io_in_0),
    .io_in_1(c53_429_io_in_1),
    .io_in_2(c53_429_io_in_2),
    .io_in_3(c53_429_io_in_3),
    .io_in_4(c53_429_io_in_4),
    .io_out_0(c53_429_io_out_0),
    .io_out_1(c53_429_io_out_1),
    .io_out_2(c53_429_io_out_2)
  );
  C53 c53_430 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_430_io_in_0),
    .io_in_1(c53_430_io_in_1),
    .io_in_2(c53_430_io_in_2),
    .io_in_3(c53_430_io_in_3),
    .io_in_4(c53_430_io_in_4),
    .io_out_0(c53_430_io_out_0),
    .io_out_1(c53_430_io_out_1),
    .io_out_2(c53_430_io_out_2)
  );
  C53 c53_431 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_431_io_in_0),
    .io_in_1(c53_431_io_in_1),
    .io_in_2(c53_431_io_in_2),
    .io_in_3(c53_431_io_in_3),
    .io_in_4(c53_431_io_in_4),
    .io_out_0(c53_431_io_out_0),
    .io_out_1(c53_431_io_out_1),
    .io_out_2(c53_431_io_out_2)
  );
  C53 c53_432 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_432_io_in_0),
    .io_in_1(c53_432_io_in_1),
    .io_in_2(c53_432_io_in_2),
    .io_in_3(c53_432_io_in_3),
    .io_in_4(c53_432_io_in_4),
    .io_out_0(c53_432_io_out_0),
    .io_out_1(c53_432_io_out_1),
    .io_out_2(c53_432_io_out_2)
  );
  C53 c53_433 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_433_io_in_0),
    .io_in_1(c53_433_io_in_1),
    .io_in_2(c53_433_io_in_2),
    .io_in_3(c53_433_io_in_3),
    .io_in_4(c53_433_io_in_4),
    .io_out_0(c53_433_io_out_0),
    .io_out_1(c53_433_io_out_1),
    .io_out_2(c53_433_io_out_2)
  );
  C53 c53_434 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_434_io_in_0),
    .io_in_1(c53_434_io_in_1),
    .io_in_2(c53_434_io_in_2),
    .io_in_3(c53_434_io_in_3),
    .io_in_4(c53_434_io_in_4),
    .io_out_0(c53_434_io_out_0),
    .io_out_1(c53_434_io_out_1),
    .io_out_2(c53_434_io_out_2)
  );
  C53 c53_435 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_435_io_in_0),
    .io_in_1(c53_435_io_in_1),
    .io_in_2(c53_435_io_in_2),
    .io_in_3(c53_435_io_in_3),
    .io_in_4(c53_435_io_in_4),
    .io_out_0(c53_435_io_out_0),
    .io_out_1(c53_435_io_out_1),
    .io_out_2(c53_435_io_out_2)
  );
  C53 c53_436 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_436_io_in_0),
    .io_in_1(c53_436_io_in_1),
    .io_in_2(c53_436_io_in_2),
    .io_in_3(c53_436_io_in_3),
    .io_in_4(c53_436_io_in_4),
    .io_out_0(c53_436_io_out_0),
    .io_out_1(c53_436_io_out_1),
    .io_out_2(c53_436_io_out_2)
  );
  C53 c53_437 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_437_io_in_0),
    .io_in_1(c53_437_io_in_1),
    .io_in_2(c53_437_io_in_2),
    .io_in_3(c53_437_io_in_3),
    .io_in_4(c53_437_io_in_4),
    .io_out_0(c53_437_io_out_0),
    .io_out_1(c53_437_io_out_1),
    .io_out_2(c53_437_io_out_2)
  );
  C53 c53_438 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_438_io_in_0),
    .io_in_1(c53_438_io_in_1),
    .io_in_2(c53_438_io_in_2),
    .io_in_3(c53_438_io_in_3),
    .io_in_4(c53_438_io_in_4),
    .io_out_0(c53_438_io_out_0),
    .io_out_1(c53_438_io_out_1),
    .io_out_2(c53_438_io_out_2)
  );
  C53 c53_439 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_439_io_in_0),
    .io_in_1(c53_439_io_in_1),
    .io_in_2(c53_439_io_in_2),
    .io_in_3(c53_439_io_in_3),
    .io_in_4(c53_439_io_in_4),
    .io_out_0(c53_439_io_out_0),
    .io_out_1(c53_439_io_out_1),
    .io_out_2(c53_439_io_out_2)
  );
  C53 c53_440 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_440_io_in_0),
    .io_in_1(c53_440_io_in_1),
    .io_in_2(c53_440_io_in_2),
    .io_in_3(c53_440_io_in_3),
    .io_in_4(c53_440_io_in_4),
    .io_out_0(c53_440_io_out_0),
    .io_out_1(c53_440_io_out_1),
    .io_out_2(c53_440_io_out_2)
  );
  C53 c53_441 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_441_io_in_0),
    .io_in_1(c53_441_io_in_1),
    .io_in_2(c53_441_io_in_2),
    .io_in_3(c53_441_io_in_3),
    .io_in_4(c53_441_io_in_4),
    .io_out_0(c53_441_io_out_0),
    .io_out_1(c53_441_io_out_1),
    .io_out_2(c53_441_io_out_2)
  );
  C53 c53_442 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_442_io_in_0),
    .io_in_1(c53_442_io_in_1),
    .io_in_2(c53_442_io_in_2),
    .io_in_3(c53_442_io_in_3),
    .io_in_4(c53_442_io_in_4),
    .io_out_0(c53_442_io_out_0),
    .io_out_1(c53_442_io_out_1),
    .io_out_2(c53_442_io_out_2)
  );
  C53 c53_443 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_443_io_in_0),
    .io_in_1(c53_443_io_in_1),
    .io_in_2(c53_443_io_in_2),
    .io_in_3(c53_443_io_in_3),
    .io_in_4(c53_443_io_in_4),
    .io_out_0(c53_443_io_out_0),
    .io_out_1(c53_443_io_out_1),
    .io_out_2(c53_443_io_out_2)
  );
  C53 c53_444 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_444_io_in_0),
    .io_in_1(c53_444_io_in_1),
    .io_in_2(c53_444_io_in_2),
    .io_in_3(c53_444_io_in_3),
    .io_in_4(c53_444_io_in_4),
    .io_out_0(c53_444_io_out_0),
    .io_out_1(c53_444_io_out_1),
    .io_out_2(c53_444_io_out_2)
  );
  C53 c53_445 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_445_io_in_0),
    .io_in_1(c53_445_io_in_1),
    .io_in_2(c53_445_io_in_2),
    .io_in_3(c53_445_io_in_3),
    .io_in_4(c53_445_io_in_4),
    .io_out_0(c53_445_io_out_0),
    .io_out_1(c53_445_io_out_1),
    .io_out_2(c53_445_io_out_2)
  );
  C53 c53_446 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_446_io_in_0),
    .io_in_1(c53_446_io_in_1),
    .io_in_2(c53_446_io_in_2),
    .io_in_3(c53_446_io_in_3),
    .io_in_4(c53_446_io_in_4),
    .io_out_0(c53_446_io_out_0),
    .io_out_1(c53_446_io_out_1),
    .io_out_2(c53_446_io_out_2)
  );
  C53 c53_447 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_447_io_in_0),
    .io_in_1(c53_447_io_in_1),
    .io_in_2(c53_447_io_in_2),
    .io_in_3(c53_447_io_in_3),
    .io_in_4(c53_447_io_in_4),
    .io_out_0(c53_447_io_out_0),
    .io_out_1(c53_447_io_out_1),
    .io_out_2(c53_447_io_out_2)
  );
  C53 c53_448 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_448_io_in_0),
    .io_in_1(c53_448_io_in_1),
    .io_in_2(c53_448_io_in_2),
    .io_in_3(c53_448_io_in_3),
    .io_in_4(c53_448_io_in_4),
    .io_out_0(c53_448_io_out_0),
    .io_out_1(c53_448_io_out_1),
    .io_out_2(c53_448_io_out_2)
  );
  C53 c53_449 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_449_io_in_0),
    .io_in_1(c53_449_io_in_1),
    .io_in_2(c53_449_io_in_2),
    .io_in_3(c53_449_io_in_3),
    .io_in_4(c53_449_io_in_4),
    .io_out_0(c53_449_io_out_0),
    .io_out_1(c53_449_io_out_1),
    .io_out_2(c53_449_io_out_2)
  );
  C53 c53_450 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_450_io_in_0),
    .io_in_1(c53_450_io_in_1),
    .io_in_2(c53_450_io_in_2),
    .io_in_3(c53_450_io_in_3),
    .io_in_4(c53_450_io_in_4),
    .io_out_0(c53_450_io_out_0),
    .io_out_1(c53_450_io_out_1),
    .io_out_2(c53_450_io_out_2)
  );
  C53 c53_451 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_451_io_in_0),
    .io_in_1(c53_451_io_in_1),
    .io_in_2(c53_451_io_in_2),
    .io_in_3(c53_451_io_in_3),
    .io_in_4(c53_451_io_in_4),
    .io_out_0(c53_451_io_out_0),
    .io_out_1(c53_451_io_out_1),
    .io_out_2(c53_451_io_out_2)
  );
  C32 c32_22 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_22_io_in_0),
    .io_in_1(c32_22_io_in_1),
    .io_in_2(c32_22_io_in_2),
    .io_out_0(c32_22_io_out_0),
    .io_out_1(c32_22_io_out_1)
  );
  C53 c53_452 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_452_io_in_0),
    .io_in_1(c53_452_io_in_1),
    .io_in_2(c53_452_io_in_2),
    .io_in_3(c53_452_io_in_3),
    .io_in_4(c53_452_io_in_4),
    .io_out_0(c53_452_io_out_0),
    .io_out_1(c53_452_io_out_1),
    .io_out_2(c53_452_io_out_2)
  );
  C53 c53_453 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_453_io_in_0),
    .io_in_1(c53_453_io_in_1),
    .io_in_2(c53_453_io_in_2),
    .io_in_3(c53_453_io_in_3),
    .io_in_4(c53_453_io_in_4),
    .io_out_0(c53_453_io_out_0),
    .io_out_1(c53_453_io_out_1),
    .io_out_2(c53_453_io_out_2)
  );
  C53 c53_454 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_454_io_in_0),
    .io_in_1(c53_454_io_in_1),
    .io_in_2(c53_454_io_in_2),
    .io_in_3(c53_454_io_in_3),
    .io_in_4(c53_454_io_in_4),
    .io_out_0(c53_454_io_out_0),
    .io_out_1(c53_454_io_out_1),
    .io_out_2(c53_454_io_out_2)
  );
  C53 c53_455 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_455_io_in_0),
    .io_in_1(c53_455_io_in_1),
    .io_in_2(c53_455_io_in_2),
    .io_in_3(c53_455_io_in_3),
    .io_in_4(c53_455_io_in_4),
    .io_out_0(c53_455_io_out_0),
    .io_out_1(c53_455_io_out_1),
    .io_out_2(c53_455_io_out_2)
  );
  C32 c32_23 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_23_io_in_0),
    .io_in_1(c32_23_io_in_1),
    .io_in_2(c32_23_io_in_2),
    .io_out_0(c32_23_io_out_0),
    .io_out_1(c32_23_io_out_1)
  );
  C53 c53_456 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_456_io_in_0),
    .io_in_1(c53_456_io_in_1),
    .io_in_2(c53_456_io_in_2),
    .io_in_3(c53_456_io_in_3),
    .io_in_4(c53_456_io_in_4),
    .io_out_0(c53_456_io_out_0),
    .io_out_1(c53_456_io_out_1),
    .io_out_2(c53_456_io_out_2)
  );
  C53 c53_457 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_457_io_in_0),
    .io_in_1(c53_457_io_in_1),
    .io_in_2(c53_457_io_in_2),
    .io_in_3(c53_457_io_in_3),
    .io_in_4(c53_457_io_in_4),
    .io_out_0(c53_457_io_out_0),
    .io_out_1(c53_457_io_out_1),
    .io_out_2(c53_457_io_out_2)
  );
  C53 c53_458 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_458_io_in_0),
    .io_in_1(c53_458_io_in_1),
    .io_in_2(c53_458_io_in_2),
    .io_in_3(c53_458_io_in_3),
    .io_in_4(c53_458_io_in_4),
    .io_out_0(c53_458_io_out_0),
    .io_out_1(c53_458_io_out_1),
    .io_out_2(c53_458_io_out_2)
  );
  C53 c53_459 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_459_io_in_0),
    .io_in_1(c53_459_io_in_1),
    .io_in_2(c53_459_io_in_2),
    .io_in_3(c53_459_io_in_3),
    .io_in_4(c53_459_io_in_4),
    .io_out_0(c53_459_io_out_0),
    .io_out_1(c53_459_io_out_1),
    .io_out_2(c53_459_io_out_2)
  );
  C22 c22_22 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_22_io_in_0),
    .io_in_1(c22_22_io_in_1),
    .io_out_0(c22_22_io_out_0),
    .io_out_1(c22_22_io_out_1)
  );
  C53 c53_460 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_460_io_in_0),
    .io_in_1(c53_460_io_in_1),
    .io_in_2(c53_460_io_in_2),
    .io_in_3(c53_460_io_in_3),
    .io_in_4(c53_460_io_in_4),
    .io_out_0(c53_460_io_out_0),
    .io_out_1(c53_460_io_out_1),
    .io_out_2(c53_460_io_out_2)
  );
  C53 c53_461 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_461_io_in_0),
    .io_in_1(c53_461_io_in_1),
    .io_in_2(c53_461_io_in_2),
    .io_in_3(c53_461_io_in_3),
    .io_in_4(c53_461_io_in_4),
    .io_out_0(c53_461_io_out_0),
    .io_out_1(c53_461_io_out_1),
    .io_out_2(c53_461_io_out_2)
  );
  C53 c53_462 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_462_io_in_0),
    .io_in_1(c53_462_io_in_1),
    .io_in_2(c53_462_io_in_2),
    .io_in_3(c53_462_io_in_3),
    .io_in_4(c53_462_io_in_4),
    .io_out_0(c53_462_io_out_0),
    .io_out_1(c53_462_io_out_1),
    .io_out_2(c53_462_io_out_2)
  );
  C53 c53_463 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_463_io_in_0),
    .io_in_1(c53_463_io_in_1),
    .io_in_2(c53_463_io_in_2),
    .io_in_3(c53_463_io_in_3),
    .io_in_4(c53_463_io_in_4),
    .io_out_0(c53_463_io_out_0),
    .io_out_1(c53_463_io_out_1),
    .io_out_2(c53_463_io_out_2)
  );
  C22 c22_23 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_23_io_in_0),
    .io_in_1(c22_23_io_in_1),
    .io_out_0(c22_23_io_out_0),
    .io_out_1(c22_23_io_out_1)
  );
  C53 c53_464 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_464_io_in_0),
    .io_in_1(c53_464_io_in_1),
    .io_in_2(c53_464_io_in_2),
    .io_in_3(c53_464_io_in_3),
    .io_in_4(c53_464_io_in_4),
    .io_out_0(c53_464_io_out_0),
    .io_out_1(c53_464_io_out_1),
    .io_out_2(c53_464_io_out_2)
  );
  C53 c53_465 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_465_io_in_0),
    .io_in_1(c53_465_io_in_1),
    .io_in_2(c53_465_io_in_2),
    .io_in_3(c53_465_io_in_3),
    .io_in_4(c53_465_io_in_4),
    .io_out_0(c53_465_io_out_0),
    .io_out_1(c53_465_io_out_1),
    .io_out_2(c53_465_io_out_2)
  );
  C53 c53_466 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_466_io_in_0),
    .io_in_1(c53_466_io_in_1),
    .io_in_2(c53_466_io_in_2),
    .io_in_3(c53_466_io_in_3),
    .io_in_4(c53_466_io_in_4),
    .io_out_0(c53_466_io_out_0),
    .io_out_1(c53_466_io_out_1),
    .io_out_2(c53_466_io_out_2)
  );
  C53 c53_467 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_467_io_in_0),
    .io_in_1(c53_467_io_in_1),
    .io_in_2(c53_467_io_in_2),
    .io_in_3(c53_467_io_in_3),
    .io_in_4(c53_467_io_in_4),
    .io_out_0(c53_467_io_out_0),
    .io_out_1(c53_467_io_out_1),
    .io_out_2(c53_467_io_out_2)
  );
  C53 c53_468 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_468_io_in_0),
    .io_in_1(c53_468_io_in_1),
    .io_in_2(c53_468_io_in_2),
    .io_in_3(c53_468_io_in_3),
    .io_in_4(c53_468_io_in_4),
    .io_out_0(c53_468_io_out_0),
    .io_out_1(c53_468_io_out_1),
    .io_out_2(c53_468_io_out_2)
  );
  C53 c53_469 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_469_io_in_0),
    .io_in_1(c53_469_io_in_1),
    .io_in_2(c53_469_io_in_2),
    .io_in_3(c53_469_io_in_3),
    .io_in_4(c53_469_io_in_4),
    .io_out_0(c53_469_io_out_0),
    .io_out_1(c53_469_io_out_1),
    .io_out_2(c53_469_io_out_2)
  );
  C53 c53_470 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_470_io_in_0),
    .io_in_1(c53_470_io_in_1),
    .io_in_2(c53_470_io_in_2),
    .io_in_3(c53_470_io_in_3),
    .io_in_4(c53_470_io_in_4),
    .io_out_0(c53_470_io_out_0),
    .io_out_1(c53_470_io_out_1),
    .io_out_2(c53_470_io_out_2)
  );
  C53 c53_471 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_471_io_in_0),
    .io_in_1(c53_471_io_in_1),
    .io_in_2(c53_471_io_in_2),
    .io_in_3(c53_471_io_in_3),
    .io_in_4(c53_471_io_in_4),
    .io_out_0(c53_471_io_out_0),
    .io_out_1(c53_471_io_out_1),
    .io_out_2(c53_471_io_out_2)
  );
  C53 c53_472 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_472_io_in_0),
    .io_in_1(c53_472_io_in_1),
    .io_in_2(c53_472_io_in_2),
    .io_in_3(c53_472_io_in_3),
    .io_in_4(c53_472_io_in_4),
    .io_out_0(c53_472_io_out_0),
    .io_out_1(c53_472_io_out_1),
    .io_out_2(c53_472_io_out_2)
  );
  C53 c53_473 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_473_io_in_0),
    .io_in_1(c53_473_io_in_1),
    .io_in_2(c53_473_io_in_2),
    .io_in_3(c53_473_io_in_3),
    .io_in_4(c53_473_io_in_4),
    .io_out_0(c53_473_io_out_0),
    .io_out_1(c53_473_io_out_1),
    .io_out_2(c53_473_io_out_2)
  );
  C53 c53_474 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_474_io_in_0),
    .io_in_1(c53_474_io_in_1),
    .io_in_2(c53_474_io_in_2),
    .io_in_3(c53_474_io_in_3),
    .io_in_4(c53_474_io_in_4),
    .io_out_0(c53_474_io_out_0),
    .io_out_1(c53_474_io_out_1),
    .io_out_2(c53_474_io_out_2)
  );
  C53 c53_475 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_475_io_in_0),
    .io_in_1(c53_475_io_in_1),
    .io_in_2(c53_475_io_in_2),
    .io_in_3(c53_475_io_in_3),
    .io_in_4(c53_475_io_in_4),
    .io_out_0(c53_475_io_out_0),
    .io_out_1(c53_475_io_out_1),
    .io_out_2(c53_475_io_out_2)
  );
  C53 c53_476 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_476_io_in_0),
    .io_in_1(c53_476_io_in_1),
    .io_in_2(c53_476_io_in_2),
    .io_in_3(c53_476_io_in_3),
    .io_in_4(c53_476_io_in_4),
    .io_out_0(c53_476_io_out_0),
    .io_out_1(c53_476_io_out_1),
    .io_out_2(c53_476_io_out_2)
  );
  C53 c53_477 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_477_io_in_0),
    .io_in_1(c53_477_io_in_1),
    .io_in_2(c53_477_io_in_2),
    .io_in_3(c53_477_io_in_3),
    .io_in_4(c53_477_io_in_4),
    .io_out_0(c53_477_io_out_0),
    .io_out_1(c53_477_io_out_1),
    .io_out_2(c53_477_io_out_2)
  );
  C53 c53_478 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_478_io_in_0),
    .io_in_1(c53_478_io_in_1),
    .io_in_2(c53_478_io_in_2),
    .io_in_3(c53_478_io_in_3),
    .io_in_4(c53_478_io_in_4),
    .io_out_0(c53_478_io_out_0),
    .io_out_1(c53_478_io_out_1),
    .io_out_2(c53_478_io_out_2)
  );
  C53 c53_479 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_479_io_in_0),
    .io_in_1(c53_479_io_in_1),
    .io_in_2(c53_479_io_in_2),
    .io_in_3(c53_479_io_in_3),
    .io_in_4(c53_479_io_in_4),
    .io_out_0(c53_479_io_out_0),
    .io_out_1(c53_479_io_out_1),
    .io_out_2(c53_479_io_out_2)
  );
  C53 c53_480 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_480_io_in_0),
    .io_in_1(c53_480_io_in_1),
    .io_in_2(c53_480_io_in_2),
    .io_in_3(c53_480_io_in_3),
    .io_in_4(c53_480_io_in_4),
    .io_out_0(c53_480_io_out_0),
    .io_out_1(c53_480_io_out_1),
    .io_out_2(c53_480_io_out_2)
  );
  C53 c53_481 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_481_io_in_0),
    .io_in_1(c53_481_io_in_1),
    .io_in_2(c53_481_io_in_2),
    .io_in_3(c53_481_io_in_3),
    .io_in_4(c53_481_io_in_4),
    .io_out_0(c53_481_io_out_0),
    .io_out_1(c53_481_io_out_1),
    .io_out_2(c53_481_io_out_2)
  );
  C53 c53_482 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_482_io_in_0),
    .io_in_1(c53_482_io_in_1),
    .io_in_2(c53_482_io_in_2),
    .io_in_3(c53_482_io_in_3),
    .io_in_4(c53_482_io_in_4),
    .io_out_0(c53_482_io_out_0),
    .io_out_1(c53_482_io_out_1),
    .io_out_2(c53_482_io_out_2)
  );
  C32 c32_24 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_24_io_in_0),
    .io_in_1(c32_24_io_in_1),
    .io_in_2(c32_24_io_in_2),
    .io_out_0(c32_24_io_out_0),
    .io_out_1(c32_24_io_out_1)
  );
  C53 c53_483 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_483_io_in_0),
    .io_in_1(c53_483_io_in_1),
    .io_in_2(c53_483_io_in_2),
    .io_in_3(c53_483_io_in_3),
    .io_in_4(c53_483_io_in_4),
    .io_out_0(c53_483_io_out_0),
    .io_out_1(c53_483_io_out_1),
    .io_out_2(c53_483_io_out_2)
  );
  C53 c53_484 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_484_io_in_0),
    .io_in_1(c53_484_io_in_1),
    .io_in_2(c53_484_io_in_2),
    .io_in_3(c53_484_io_in_3),
    .io_in_4(c53_484_io_in_4),
    .io_out_0(c53_484_io_out_0),
    .io_out_1(c53_484_io_out_1),
    .io_out_2(c53_484_io_out_2)
  );
  C53 c53_485 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_485_io_in_0),
    .io_in_1(c53_485_io_in_1),
    .io_in_2(c53_485_io_in_2),
    .io_in_3(c53_485_io_in_3),
    .io_in_4(c53_485_io_in_4),
    .io_out_0(c53_485_io_out_0),
    .io_out_1(c53_485_io_out_1),
    .io_out_2(c53_485_io_out_2)
  );
  C32 c32_25 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_25_io_in_0),
    .io_in_1(c32_25_io_in_1),
    .io_in_2(c32_25_io_in_2),
    .io_out_0(c32_25_io_out_0),
    .io_out_1(c32_25_io_out_1)
  );
  C53 c53_486 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_486_io_in_0),
    .io_in_1(c53_486_io_in_1),
    .io_in_2(c53_486_io_in_2),
    .io_in_3(c53_486_io_in_3),
    .io_in_4(c53_486_io_in_4),
    .io_out_0(c53_486_io_out_0),
    .io_out_1(c53_486_io_out_1),
    .io_out_2(c53_486_io_out_2)
  );
  C53 c53_487 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_487_io_in_0),
    .io_in_1(c53_487_io_in_1),
    .io_in_2(c53_487_io_in_2),
    .io_in_3(c53_487_io_in_3),
    .io_in_4(c53_487_io_in_4),
    .io_out_0(c53_487_io_out_0),
    .io_out_1(c53_487_io_out_1),
    .io_out_2(c53_487_io_out_2)
  );
  C53 c53_488 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_488_io_in_0),
    .io_in_1(c53_488_io_in_1),
    .io_in_2(c53_488_io_in_2),
    .io_in_3(c53_488_io_in_3),
    .io_in_4(c53_488_io_in_4),
    .io_out_0(c53_488_io_out_0),
    .io_out_1(c53_488_io_out_1),
    .io_out_2(c53_488_io_out_2)
  );
  C22 c22_24 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_24_io_in_0),
    .io_in_1(c22_24_io_in_1),
    .io_out_0(c22_24_io_out_0),
    .io_out_1(c22_24_io_out_1)
  );
  C53 c53_489 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_489_io_in_0),
    .io_in_1(c53_489_io_in_1),
    .io_in_2(c53_489_io_in_2),
    .io_in_3(c53_489_io_in_3),
    .io_in_4(c53_489_io_in_4),
    .io_out_0(c53_489_io_out_0),
    .io_out_1(c53_489_io_out_1),
    .io_out_2(c53_489_io_out_2)
  );
  C53 c53_490 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_490_io_in_0),
    .io_in_1(c53_490_io_in_1),
    .io_in_2(c53_490_io_in_2),
    .io_in_3(c53_490_io_in_3),
    .io_in_4(c53_490_io_in_4),
    .io_out_0(c53_490_io_out_0),
    .io_out_1(c53_490_io_out_1),
    .io_out_2(c53_490_io_out_2)
  );
  C53 c53_491 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_491_io_in_0),
    .io_in_1(c53_491_io_in_1),
    .io_in_2(c53_491_io_in_2),
    .io_in_3(c53_491_io_in_3),
    .io_in_4(c53_491_io_in_4),
    .io_out_0(c53_491_io_out_0),
    .io_out_1(c53_491_io_out_1),
    .io_out_2(c53_491_io_out_2)
  );
  C22 c22_25 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_25_io_in_0),
    .io_in_1(c22_25_io_in_1),
    .io_out_0(c22_25_io_out_0),
    .io_out_1(c22_25_io_out_1)
  );
  C53 c53_492 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_492_io_in_0),
    .io_in_1(c53_492_io_in_1),
    .io_in_2(c53_492_io_in_2),
    .io_in_3(c53_492_io_in_3),
    .io_in_4(c53_492_io_in_4),
    .io_out_0(c53_492_io_out_0),
    .io_out_1(c53_492_io_out_1),
    .io_out_2(c53_492_io_out_2)
  );
  C53 c53_493 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_493_io_in_0),
    .io_in_1(c53_493_io_in_1),
    .io_in_2(c53_493_io_in_2),
    .io_in_3(c53_493_io_in_3),
    .io_in_4(c53_493_io_in_4),
    .io_out_0(c53_493_io_out_0),
    .io_out_1(c53_493_io_out_1),
    .io_out_2(c53_493_io_out_2)
  );
  C53 c53_494 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_494_io_in_0),
    .io_in_1(c53_494_io_in_1),
    .io_in_2(c53_494_io_in_2),
    .io_in_3(c53_494_io_in_3),
    .io_in_4(c53_494_io_in_4),
    .io_out_0(c53_494_io_out_0),
    .io_out_1(c53_494_io_out_1),
    .io_out_2(c53_494_io_out_2)
  );
  C53 c53_495 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_495_io_in_0),
    .io_in_1(c53_495_io_in_1),
    .io_in_2(c53_495_io_in_2),
    .io_in_3(c53_495_io_in_3),
    .io_in_4(c53_495_io_in_4),
    .io_out_0(c53_495_io_out_0),
    .io_out_1(c53_495_io_out_1),
    .io_out_2(c53_495_io_out_2)
  );
  C53 c53_496 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_496_io_in_0),
    .io_in_1(c53_496_io_in_1),
    .io_in_2(c53_496_io_in_2),
    .io_in_3(c53_496_io_in_3),
    .io_in_4(c53_496_io_in_4),
    .io_out_0(c53_496_io_out_0),
    .io_out_1(c53_496_io_out_1),
    .io_out_2(c53_496_io_out_2)
  );
  C53 c53_497 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_497_io_in_0),
    .io_in_1(c53_497_io_in_1),
    .io_in_2(c53_497_io_in_2),
    .io_in_3(c53_497_io_in_3),
    .io_in_4(c53_497_io_in_4),
    .io_out_0(c53_497_io_out_0),
    .io_out_1(c53_497_io_out_1),
    .io_out_2(c53_497_io_out_2)
  );
  C53 c53_498 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_498_io_in_0),
    .io_in_1(c53_498_io_in_1),
    .io_in_2(c53_498_io_in_2),
    .io_in_3(c53_498_io_in_3),
    .io_in_4(c53_498_io_in_4),
    .io_out_0(c53_498_io_out_0),
    .io_out_1(c53_498_io_out_1),
    .io_out_2(c53_498_io_out_2)
  );
  C53 c53_499 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_499_io_in_0),
    .io_in_1(c53_499_io_in_1),
    .io_in_2(c53_499_io_in_2),
    .io_in_3(c53_499_io_in_3),
    .io_in_4(c53_499_io_in_4),
    .io_out_0(c53_499_io_out_0),
    .io_out_1(c53_499_io_out_1),
    .io_out_2(c53_499_io_out_2)
  );
  C53 c53_500 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_500_io_in_0),
    .io_in_1(c53_500_io_in_1),
    .io_in_2(c53_500_io_in_2),
    .io_in_3(c53_500_io_in_3),
    .io_in_4(c53_500_io_in_4),
    .io_out_0(c53_500_io_out_0),
    .io_out_1(c53_500_io_out_1),
    .io_out_2(c53_500_io_out_2)
  );
  C53 c53_501 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_501_io_in_0),
    .io_in_1(c53_501_io_in_1),
    .io_in_2(c53_501_io_in_2),
    .io_in_3(c53_501_io_in_3),
    .io_in_4(c53_501_io_in_4),
    .io_out_0(c53_501_io_out_0),
    .io_out_1(c53_501_io_out_1),
    .io_out_2(c53_501_io_out_2)
  );
  C53 c53_502 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_502_io_in_0),
    .io_in_1(c53_502_io_in_1),
    .io_in_2(c53_502_io_in_2),
    .io_in_3(c53_502_io_in_3),
    .io_in_4(c53_502_io_in_4),
    .io_out_0(c53_502_io_out_0),
    .io_out_1(c53_502_io_out_1),
    .io_out_2(c53_502_io_out_2)
  );
  C53 c53_503 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_503_io_in_0),
    .io_in_1(c53_503_io_in_1),
    .io_in_2(c53_503_io_in_2),
    .io_in_3(c53_503_io_in_3),
    .io_in_4(c53_503_io_in_4),
    .io_out_0(c53_503_io_out_0),
    .io_out_1(c53_503_io_out_1),
    .io_out_2(c53_503_io_out_2)
  );
  C53 c53_504 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_504_io_in_0),
    .io_in_1(c53_504_io_in_1),
    .io_in_2(c53_504_io_in_2),
    .io_in_3(c53_504_io_in_3),
    .io_in_4(c53_504_io_in_4),
    .io_out_0(c53_504_io_out_0),
    .io_out_1(c53_504_io_out_1),
    .io_out_2(c53_504_io_out_2)
  );
  C53 c53_505 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_505_io_in_0),
    .io_in_1(c53_505_io_in_1),
    .io_in_2(c53_505_io_in_2),
    .io_in_3(c53_505_io_in_3),
    .io_in_4(c53_505_io_in_4),
    .io_out_0(c53_505_io_out_0),
    .io_out_1(c53_505_io_out_1),
    .io_out_2(c53_505_io_out_2)
  );
  C32 c32_26 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_26_io_in_0),
    .io_in_1(c32_26_io_in_1),
    .io_in_2(c32_26_io_in_2),
    .io_out_0(c32_26_io_out_0),
    .io_out_1(c32_26_io_out_1)
  );
  C53 c53_506 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_506_io_in_0),
    .io_in_1(c53_506_io_in_1),
    .io_in_2(c53_506_io_in_2),
    .io_in_3(c53_506_io_in_3),
    .io_in_4(c53_506_io_in_4),
    .io_out_0(c53_506_io_out_0),
    .io_out_1(c53_506_io_out_1),
    .io_out_2(c53_506_io_out_2)
  );
  C53 c53_507 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_507_io_in_0),
    .io_in_1(c53_507_io_in_1),
    .io_in_2(c53_507_io_in_2),
    .io_in_3(c53_507_io_in_3),
    .io_in_4(c53_507_io_in_4),
    .io_out_0(c53_507_io_out_0),
    .io_out_1(c53_507_io_out_1),
    .io_out_2(c53_507_io_out_2)
  );
  C32 c32_27 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_27_io_in_0),
    .io_in_1(c32_27_io_in_1),
    .io_in_2(c32_27_io_in_2),
    .io_out_0(c32_27_io_out_0),
    .io_out_1(c32_27_io_out_1)
  );
  C53 c53_508 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_508_io_in_0),
    .io_in_1(c53_508_io_in_1),
    .io_in_2(c53_508_io_in_2),
    .io_in_3(c53_508_io_in_3),
    .io_in_4(c53_508_io_in_4),
    .io_out_0(c53_508_io_out_0),
    .io_out_1(c53_508_io_out_1),
    .io_out_2(c53_508_io_out_2)
  );
  C53 c53_509 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_509_io_in_0),
    .io_in_1(c53_509_io_in_1),
    .io_in_2(c53_509_io_in_2),
    .io_in_3(c53_509_io_in_3),
    .io_in_4(c53_509_io_in_4),
    .io_out_0(c53_509_io_out_0),
    .io_out_1(c53_509_io_out_1),
    .io_out_2(c53_509_io_out_2)
  );
  C22 c22_26 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_26_io_in_0),
    .io_in_1(c22_26_io_in_1),
    .io_out_0(c22_26_io_out_0),
    .io_out_1(c22_26_io_out_1)
  );
  C53 c53_510 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_510_io_in_0),
    .io_in_1(c53_510_io_in_1),
    .io_in_2(c53_510_io_in_2),
    .io_in_3(c53_510_io_in_3),
    .io_in_4(c53_510_io_in_4),
    .io_out_0(c53_510_io_out_0),
    .io_out_1(c53_510_io_out_1),
    .io_out_2(c53_510_io_out_2)
  );
  C53 c53_511 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_511_io_in_0),
    .io_in_1(c53_511_io_in_1),
    .io_in_2(c53_511_io_in_2),
    .io_in_3(c53_511_io_in_3),
    .io_in_4(c53_511_io_in_4),
    .io_out_0(c53_511_io_out_0),
    .io_out_1(c53_511_io_out_1),
    .io_out_2(c53_511_io_out_2)
  );
  C22 c22_27 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_27_io_in_0),
    .io_in_1(c22_27_io_in_1),
    .io_out_0(c22_27_io_out_0),
    .io_out_1(c22_27_io_out_1)
  );
  C53 c53_512 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_512_io_in_0),
    .io_in_1(c53_512_io_in_1),
    .io_in_2(c53_512_io_in_2),
    .io_in_3(c53_512_io_in_3),
    .io_in_4(c53_512_io_in_4),
    .io_out_0(c53_512_io_out_0),
    .io_out_1(c53_512_io_out_1),
    .io_out_2(c53_512_io_out_2)
  );
  C53 c53_513 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_513_io_in_0),
    .io_in_1(c53_513_io_in_1),
    .io_in_2(c53_513_io_in_2),
    .io_in_3(c53_513_io_in_3),
    .io_in_4(c53_513_io_in_4),
    .io_out_0(c53_513_io_out_0),
    .io_out_1(c53_513_io_out_1),
    .io_out_2(c53_513_io_out_2)
  );
  C53 c53_514 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_514_io_in_0),
    .io_in_1(c53_514_io_in_1),
    .io_in_2(c53_514_io_in_2),
    .io_in_3(c53_514_io_in_3),
    .io_in_4(c53_514_io_in_4),
    .io_out_0(c53_514_io_out_0),
    .io_out_1(c53_514_io_out_1),
    .io_out_2(c53_514_io_out_2)
  );
  C53 c53_515 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_515_io_in_0),
    .io_in_1(c53_515_io_in_1),
    .io_in_2(c53_515_io_in_2),
    .io_in_3(c53_515_io_in_3),
    .io_in_4(c53_515_io_in_4),
    .io_out_0(c53_515_io_out_0),
    .io_out_1(c53_515_io_out_1),
    .io_out_2(c53_515_io_out_2)
  );
  C53 c53_516 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_516_io_in_0),
    .io_in_1(c53_516_io_in_1),
    .io_in_2(c53_516_io_in_2),
    .io_in_3(c53_516_io_in_3),
    .io_in_4(c53_516_io_in_4),
    .io_out_0(c53_516_io_out_0),
    .io_out_1(c53_516_io_out_1),
    .io_out_2(c53_516_io_out_2)
  );
  C53 c53_517 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_517_io_in_0),
    .io_in_1(c53_517_io_in_1),
    .io_in_2(c53_517_io_in_2),
    .io_in_3(c53_517_io_in_3),
    .io_in_4(c53_517_io_in_4),
    .io_out_0(c53_517_io_out_0),
    .io_out_1(c53_517_io_out_1),
    .io_out_2(c53_517_io_out_2)
  );
  C53 c53_518 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_518_io_in_0),
    .io_in_1(c53_518_io_in_1),
    .io_in_2(c53_518_io_in_2),
    .io_in_3(c53_518_io_in_3),
    .io_in_4(c53_518_io_in_4),
    .io_out_0(c53_518_io_out_0),
    .io_out_1(c53_518_io_out_1),
    .io_out_2(c53_518_io_out_2)
  );
  C53 c53_519 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_519_io_in_0),
    .io_in_1(c53_519_io_in_1),
    .io_in_2(c53_519_io_in_2),
    .io_in_3(c53_519_io_in_3),
    .io_in_4(c53_519_io_in_4),
    .io_out_0(c53_519_io_out_0),
    .io_out_1(c53_519_io_out_1),
    .io_out_2(c53_519_io_out_2)
  );
  C53 c53_520 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_520_io_in_0),
    .io_in_1(c53_520_io_in_1),
    .io_in_2(c53_520_io_in_2),
    .io_in_3(c53_520_io_in_3),
    .io_in_4(c53_520_io_in_4),
    .io_out_0(c53_520_io_out_0),
    .io_out_1(c53_520_io_out_1),
    .io_out_2(c53_520_io_out_2)
  );
  C32 c32_28 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_28_io_in_0),
    .io_in_1(c32_28_io_in_1),
    .io_in_2(c32_28_io_in_2),
    .io_out_0(c32_28_io_out_0),
    .io_out_1(c32_28_io_out_1)
  );
  C53 c53_521 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_521_io_in_0),
    .io_in_1(c53_521_io_in_1),
    .io_in_2(c53_521_io_in_2),
    .io_in_3(c53_521_io_in_3),
    .io_in_4(c53_521_io_in_4),
    .io_out_0(c53_521_io_out_0),
    .io_out_1(c53_521_io_out_1),
    .io_out_2(c53_521_io_out_2)
  );
  C32 c32_29 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_29_io_in_0),
    .io_in_1(c32_29_io_in_1),
    .io_in_2(c32_29_io_in_2),
    .io_out_0(c32_29_io_out_0),
    .io_out_1(c32_29_io_out_1)
  );
  C53 c53_522 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_522_io_in_0),
    .io_in_1(c53_522_io_in_1),
    .io_in_2(c53_522_io_in_2),
    .io_in_3(c53_522_io_in_3),
    .io_in_4(c53_522_io_in_4),
    .io_out_0(c53_522_io_out_0),
    .io_out_1(c53_522_io_out_1),
    .io_out_2(c53_522_io_out_2)
  );
  C22 c22_28 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_28_io_in_0),
    .io_in_1(c22_28_io_in_1),
    .io_out_0(c22_28_io_out_0),
    .io_out_1(c22_28_io_out_1)
  );
  C53 c53_523 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_523_io_in_0),
    .io_in_1(c53_523_io_in_1),
    .io_in_2(c53_523_io_in_2),
    .io_in_3(c53_523_io_in_3),
    .io_in_4(c53_523_io_in_4),
    .io_out_0(c53_523_io_out_0),
    .io_out_1(c53_523_io_out_1),
    .io_out_2(c53_523_io_out_2)
  );
  C22 c22_29 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_29_io_in_0),
    .io_in_1(c22_29_io_in_1),
    .io_out_0(c22_29_io_out_0),
    .io_out_1(c22_29_io_out_1)
  );
  C53 c53_524 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_524_io_in_0),
    .io_in_1(c53_524_io_in_1),
    .io_in_2(c53_524_io_in_2),
    .io_in_3(c53_524_io_in_3),
    .io_in_4(c53_524_io_in_4),
    .io_out_0(c53_524_io_out_0),
    .io_out_1(c53_524_io_out_1),
    .io_out_2(c53_524_io_out_2)
  );
  C53 c53_525 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_525_io_in_0),
    .io_in_1(c53_525_io_in_1),
    .io_in_2(c53_525_io_in_2),
    .io_in_3(c53_525_io_in_3),
    .io_in_4(c53_525_io_in_4),
    .io_out_0(c53_525_io_out_0),
    .io_out_1(c53_525_io_out_1),
    .io_out_2(c53_525_io_out_2)
  );
  C53 c53_526 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_526_io_in_0),
    .io_in_1(c53_526_io_in_1),
    .io_in_2(c53_526_io_in_2),
    .io_in_3(c53_526_io_in_3),
    .io_in_4(c53_526_io_in_4),
    .io_out_0(c53_526_io_out_0),
    .io_out_1(c53_526_io_out_1),
    .io_out_2(c53_526_io_out_2)
  );
  C53 c53_527 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_527_io_in_0),
    .io_in_1(c53_527_io_in_1),
    .io_in_2(c53_527_io_in_2),
    .io_in_3(c53_527_io_in_3),
    .io_in_4(c53_527_io_in_4),
    .io_out_0(c53_527_io_out_0),
    .io_out_1(c53_527_io_out_1),
    .io_out_2(c53_527_io_out_2)
  );
  C32 c32_30 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_30_io_in_0),
    .io_in_1(c32_30_io_in_1),
    .io_in_2(c32_30_io_in_2),
    .io_out_0(c32_30_io_out_0),
    .io_out_1(c32_30_io_out_1)
  );
  C32 c32_31 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_31_io_in_0),
    .io_in_1(c32_31_io_in_1),
    .io_in_2(c32_31_io_in_2),
    .io_out_0(c32_31_io_out_0),
    .io_out_1(c32_31_io_out_1)
  );
  C22 c22_30 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_30_io_in_0),
    .io_in_1(c22_30_io_in_1),
    .io_out_0(c22_30_io_out_0),
    .io_out_1(c22_30_io_out_1)
  );
  C22 c22_31 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_31_io_in_0),
    .io_in_1(c22_31_io_in_1),
    .io_out_0(c22_31_io_out_0),
    .io_out_1(c22_31_io_out_1)
  );
  C22 c22_32 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_32_io_in_0),
    .io_in_1(c22_32_io_in_1),
    .io_out_0(c22_32_io_out_0),
    .io_out_1(c22_32_io_out_1)
  );
  C22 c22_33 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_33_io_in_0),
    .io_in_1(c22_33_io_in_1),
    .io_out_0(c22_33_io_out_0),
    .io_out_1(c22_33_io_out_1)
  );
  C22 c22_34 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_34_io_in_0),
    .io_in_1(c22_34_io_in_1),
    .io_out_0(c22_34_io_out_0),
    .io_out_1(c22_34_io_out_1)
  );
  C22 c22_35 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_35_io_in_0),
    .io_in_1(c22_35_io_in_1),
    .io_out_0(c22_35_io_out_0),
    .io_out_1(c22_35_io_out_1)
  );
  C22 c22_36 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_36_io_in_0),
    .io_in_1(c22_36_io_in_1),
    .io_out_0(c22_36_io_out_0),
    .io_out_1(c22_36_io_out_1)
  );
  C32 c32_32 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_32_io_in_0),
    .io_in_1(c32_32_io_in_1),
    .io_in_2(c32_32_io_in_2),
    .io_out_0(c32_32_io_out_0),
    .io_out_1(c32_32_io_out_1)
  );
  C32 c32_33 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_33_io_in_0),
    .io_in_1(c32_33_io_in_1),
    .io_in_2(c32_33_io_in_2),
    .io_out_0(c32_33_io_out_0),
    .io_out_1(c32_33_io_out_1)
  );
  C32 c32_34 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_34_io_in_0),
    .io_in_1(c32_34_io_in_1),
    .io_in_2(c32_34_io_in_2),
    .io_out_0(c32_34_io_out_0),
    .io_out_1(c32_34_io_out_1)
  );
  C53 c53_528 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_528_io_in_0),
    .io_in_1(c53_528_io_in_1),
    .io_in_2(c53_528_io_in_2),
    .io_in_3(c53_528_io_in_3),
    .io_in_4(c53_528_io_in_4),
    .io_out_0(c53_528_io_out_0),
    .io_out_1(c53_528_io_out_1),
    .io_out_2(c53_528_io_out_2)
  );
  C53 c53_529 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_529_io_in_0),
    .io_in_1(c53_529_io_in_1),
    .io_in_2(c53_529_io_in_2),
    .io_in_3(c53_529_io_in_3),
    .io_in_4(c53_529_io_in_4),
    .io_out_0(c53_529_io_out_0),
    .io_out_1(c53_529_io_out_1),
    .io_out_2(c53_529_io_out_2)
  );
  C53 c53_530 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_530_io_in_0),
    .io_in_1(c53_530_io_in_1),
    .io_in_2(c53_530_io_in_2),
    .io_in_3(c53_530_io_in_3),
    .io_in_4(c53_530_io_in_4),
    .io_out_0(c53_530_io_out_0),
    .io_out_1(c53_530_io_out_1),
    .io_out_2(c53_530_io_out_2)
  );
  C53 c53_531 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_531_io_in_0),
    .io_in_1(c53_531_io_in_1),
    .io_in_2(c53_531_io_in_2),
    .io_in_3(c53_531_io_in_3),
    .io_in_4(c53_531_io_in_4),
    .io_out_0(c53_531_io_out_0),
    .io_out_1(c53_531_io_out_1),
    .io_out_2(c53_531_io_out_2)
  );
  C53 c53_532 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_532_io_in_0),
    .io_in_1(c53_532_io_in_1),
    .io_in_2(c53_532_io_in_2),
    .io_in_3(c53_532_io_in_3),
    .io_in_4(c53_532_io_in_4),
    .io_out_0(c53_532_io_out_0),
    .io_out_1(c53_532_io_out_1),
    .io_out_2(c53_532_io_out_2)
  );
  C53 c53_533 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_533_io_in_0),
    .io_in_1(c53_533_io_in_1),
    .io_in_2(c53_533_io_in_2),
    .io_in_3(c53_533_io_in_3),
    .io_in_4(c53_533_io_in_4),
    .io_out_0(c53_533_io_out_0),
    .io_out_1(c53_533_io_out_1),
    .io_out_2(c53_533_io_out_2)
  );
  C53 c53_534 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_534_io_in_0),
    .io_in_1(c53_534_io_in_1),
    .io_in_2(c53_534_io_in_2),
    .io_in_3(c53_534_io_in_3),
    .io_in_4(c53_534_io_in_4),
    .io_out_0(c53_534_io_out_0),
    .io_out_1(c53_534_io_out_1),
    .io_out_2(c53_534_io_out_2)
  );
  C53 c53_535 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_535_io_in_0),
    .io_in_1(c53_535_io_in_1),
    .io_in_2(c53_535_io_in_2),
    .io_in_3(c53_535_io_in_3),
    .io_in_4(c53_535_io_in_4),
    .io_out_0(c53_535_io_out_0),
    .io_out_1(c53_535_io_out_1),
    .io_out_2(c53_535_io_out_2)
  );
  C53 c53_536 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_536_io_in_0),
    .io_in_1(c53_536_io_in_1),
    .io_in_2(c53_536_io_in_2),
    .io_in_3(c53_536_io_in_3),
    .io_in_4(c53_536_io_in_4),
    .io_out_0(c53_536_io_out_0),
    .io_out_1(c53_536_io_out_1),
    .io_out_2(c53_536_io_out_2)
  );
  C22 c22_37 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_37_io_in_0),
    .io_in_1(c22_37_io_in_1),
    .io_out_0(c22_37_io_out_0),
    .io_out_1(c22_37_io_out_1)
  );
  C53 c53_537 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_537_io_in_0),
    .io_in_1(c53_537_io_in_1),
    .io_in_2(c53_537_io_in_2),
    .io_in_3(c53_537_io_in_3),
    .io_in_4(c53_537_io_in_4),
    .io_out_0(c53_537_io_out_0),
    .io_out_1(c53_537_io_out_1),
    .io_out_2(c53_537_io_out_2)
  );
  C22 c22_38 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_38_io_in_0),
    .io_in_1(c22_38_io_in_1),
    .io_out_0(c22_38_io_out_0),
    .io_out_1(c22_38_io_out_1)
  );
  C53 c53_538 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_538_io_in_0),
    .io_in_1(c53_538_io_in_1),
    .io_in_2(c53_538_io_in_2),
    .io_in_3(c53_538_io_in_3),
    .io_in_4(c53_538_io_in_4),
    .io_out_0(c53_538_io_out_0),
    .io_out_1(c53_538_io_out_1),
    .io_out_2(c53_538_io_out_2)
  );
  C22 c22_39 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_39_io_in_0),
    .io_in_1(c22_39_io_in_1),
    .io_out_0(c22_39_io_out_0),
    .io_out_1(c22_39_io_out_1)
  );
  C53 c53_539 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_539_io_in_0),
    .io_in_1(c53_539_io_in_1),
    .io_in_2(c53_539_io_in_2),
    .io_in_3(c53_539_io_in_3),
    .io_in_4(c53_539_io_in_4),
    .io_out_0(c53_539_io_out_0),
    .io_out_1(c53_539_io_out_1),
    .io_out_2(c53_539_io_out_2)
  );
  C22 c22_40 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_40_io_in_0),
    .io_in_1(c22_40_io_in_1),
    .io_out_0(c22_40_io_out_0),
    .io_out_1(c22_40_io_out_1)
  );
  C53 c53_540 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_540_io_in_0),
    .io_in_1(c53_540_io_in_1),
    .io_in_2(c53_540_io_in_2),
    .io_in_3(c53_540_io_in_3),
    .io_in_4(c53_540_io_in_4),
    .io_out_0(c53_540_io_out_0),
    .io_out_1(c53_540_io_out_1),
    .io_out_2(c53_540_io_out_2)
  );
  C22 c22_41 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_41_io_in_0),
    .io_in_1(c22_41_io_in_1),
    .io_out_0(c22_41_io_out_0),
    .io_out_1(c22_41_io_out_1)
  );
  C53 c53_541 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_541_io_in_0),
    .io_in_1(c53_541_io_in_1),
    .io_in_2(c53_541_io_in_2),
    .io_in_3(c53_541_io_in_3),
    .io_in_4(c53_541_io_in_4),
    .io_out_0(c53_541_io_out_0),
    .io_out_1(c53_541_io_out_1),
    .io_out_2(c53_541_io_out_2)
  );
  C32 c32_35 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_35_io_in_0),
    .io_in_1(c32_35_io_in_1),
    .io_in_2(c32_35_io_in_2),
    .io_out_0(c32_35_io_out_0),
    .io_out_1(c32_35_io_out_1)
  );
  C53 c53_542 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_542_io_in_0),
    .io_in_1(c53_542_io_in_1),
    .io_in_2(c53_542_io_in_2),
    .io_in_3(c53_542_io_in_3),
    .io_in_4(c53_542_io_in_4),
    .io_out_0(c53_542_io_out_0),
    .io_out_1(c53_542_io_out_1),
    .io_out_2(c53_542_io_out_2)
  );
  C32 c32_36 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_36_io_in_0),
    .io_in_1(c32_36_io_in_1),
    .io_in_2(c32_36_io_in_2),
    .io_out_0(c32_36_io_out_0),
    .io_out_1(c32_36_io_out_1)
  );
  C53 c53_543 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_543_io_in_0),
    .io_in_1(c53_543_io_in_1),
    .io_in_2(c53_543_io_in_2),
    .io_in_3(c53_543_io_in_3),
    .io_in_4(c53_543_io_in_4),
    .io_out_0(c53_543_io_out_0),
    .io_out_1(c53_543_io_out_1),
    .io_out_2(c53_543_io_out_2)
  );
  C32 c32_37 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_37_io_in_0),
    .io_in_1(c32_37_io_in_1),
    .io_in_2(c32_37_io_in_2),
    .io_out_0(c32_37_io_out_0),
    .io_out_1(c32_37_io_out_1)
  );
  C53 c53_544 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_544_io_in_0),
    .io_in_1(c53_544_io_in_1),
    .io_in_2(c53_544_io_in_2),
    .io_in_3(c53_544_io_in_3),
    .io_in_4(c53_544_io_in_4),
    .io_out_0(c53_544_io_out_0),
    .io_out_1(c53_544_io_out_1),
    .io_out_2(c53_544_io_out_2)
  );
  C53 c53_545 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_545_io_in_0),
    .io_in_1(c53_545_io_in_1),
    .io_in_2(c53_545_io_in_2),
    .io_in_3(c53_545_io_in_3),
    .io_in_4(c53_545_io_in_4),
    .io_out_0(c53_545_io_out_0),
    .io_out_1(c53_545_io_out_1),
    .io_out_2(c53_545_io_out_2)
  );
  C53 c53_546 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_546_io_in_0),
    .io_in_1(c53_546_io_in_1),
    .io_in_2(c53_546_io_in_2),
    .io_in_3(c53_546_io_in_3),
    .io_in_4(c53_546_io_in_4),
    .io_out_0(c53_546_io_out_0),
    .io_out_1(c53_546_io_out_1),
    .io_out_2(c53_546_io_out_2)
  );
  C53 c53_547 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_547_io_in_0),
    .io_in_1(c53_547_io_in_1),
    .io_in_2(c53_547_io_in_2),
    .io_in_3(c53_547_io_in_3),
    .io_in_4(c53_547_io_in_4),
    .io_out_0(c53_547_io_out_0),
    .io_out_1(c53_547_io_out_1),
    .io_out_2(c53_547_io_out_2)
  );
  C53 c53_548 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_548_io_in_0),
    .io_in_1(c53_548_io_in_1),
    .io_in_2(c53_548_io_in_2),
    .io_in_3(c53_548_io_in_3),
    .io_in_4(c53_548_io_in_4),
    .io_out_0(c53_548_io_out_0),
    .io_out_1(c53_548_io_out_1),
    .io_out_2(c53_548_io_out_2)
  );
  C53 c53_549 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_549_io_in_0),
    .io_in_1(c53_549_io_in_1),
    .io_in_2(c53_549_io_in_2),
    .io_in_3(c53_549_io_in_3),
    .io_in_4(c53_549_io_in_4),
    .io_out_0(c53_549_io_out_0),
    .io_out_1(c53_549_io_out_1),
    .io_out_2(c53_549_io_out_2)
  );
  C53 c53_550 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_550_io_in_0),
    .io_in_1(c53_550_io_in_1),
    .io_in_2(c53_550_io_in_2),
    .io_in_3(c53_550_io_in_3),
    .io_in_4(c53_550_io_in_4),
    .io_out_0(c53_550_io_out_0),
    .io_out_1(c53_550_io_out_1),
    .io_out_2(c53_550_io_out_2)
  );
  C53 c53_551 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_551_io_in_0),
    .io_in_1(c53_551_io_in_1),
    .io_in_2(c53_551_io_in_2),
    .io_in_3(c53_551_io_in_3),
    .io_in_4(c53_551_io_in_4),
    .io_out_0(c53_551_io_out_0),
    .io_out_1(c53_551_io_out_1),
    .io_out_2(c53_551_io_out_2)
  );
  C53 c53_552 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_552_io_in_0),
    .io_in_1(c53_552_io_in_1),
    .io_in_2(c53_552_io_in_2),
    .io_in_3(c53_552_io_in_3),
    .io_in_4(c53_552_io_in_4),
    .io_out_0(c53_552_io_out_0),
    .io_out_1(c53_552_io_out_1),
    .io_out_2(c53_552_io_out_2)
  );
  C53 c53_553 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_553_io_in_0),
    .io_in_1(c53_553_io_in_1),
    .io_in_2(c53_553_io_in_2),
    .io_in_3(c53_553_io_in_3),
    .io_in_4(c53_553_io_in_4),
    .io_out_0(c53_553_io_out_0),
    .io_out_1(c53_553_io_out_1),
    .io_out_2(c53_553_io_out_2)
  );
  C53 c53_554 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_554_io_in_0),
    .io_in_1(c53_554_io_in_1),
    .io_in_2(c53_554_io_in_2),
    .io_in_3(c53_554_io_in_3),
    .io_in_4(c53_554_io_in_4),
    .io_out_0(c53_554_io_out_0),
    .io_out_1(c53_554_io_out_1),
    .io_out_2(c53_554_io_out_2)
  );
  C53 c53_555 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_555_io_in_0),
    .io_in_1(c53_555_io_in_1),
    .io_in_2(c53_555_io_in_2),
    .io_in_3(c53_555_io_in_3),
    .io_in_4(c53_555_io_in_4),
    .io_out_0(c53_555_io_out_0),
    .io_out_1(c53_555_io_out_1),
    .io_out_2(c53_555_io_out_2)
  );
  C53 c53_556 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_556_io_in_0),
    .io_in_1(c53_556_io_in_1),
    .io_in_2(c53_556_io_in_2),
    .io_in_3(c53_556_io_in_3),
    .io_in_4(c53_556_io_in_4),
    .io_out_0(c53_556_io_out_0),
    .io_out_1(c53_556_io_out_1),
    .io_out_2(c53_556_io_out_2)
  );
  C53 c53_557 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_557_io_in_0),
    .io_in_1(c53_557_io_in_1),
    .io_in_2(c53_557_io_in_2),
    .io_in_3(c53_557_io_in_3),
    .io_in_4(c53_557_io_in_4),
    .io_out_0(c53_557_io_out_0),
    .io_out_1(c53_557_io_out_1),
    .io_out_2(c53_557_io_out_2)
  );
  C53 c53_558 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_558_io_in_0),
    .io_in_1(c53_558_io_in_1),
    .io_in_2(c53_558_io_in_2),
    .io_in_3(c53_558_io_in_3),
    .io_in_4(c53_558_io_in_4),
    .io_out_0(c53_558_io_out_0),
    .io_out_1(c53_558_io_out_1),
    .io_out_2(c53_558_io_out_2)
  );
  C53 c53_559 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_559_io_in_0),
    .io_in_1(c53_559_io_in_1),
    .io_in_2(c53_559_io_in_2),
    .io_in_3(c53_559_io_in_3),
    .io_in_4(c53_559_io_in_4),
    .io_out_0(c53_559_io_out_0),
    .io_out_1(c53_559_io_out_1),
    .io_out_2(c53_559_io_out_2)
  );
  C53 c53_560 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_560_io_in_0),
    .io_in_1(c53_560_io_in_1),
    .io_in_2(c53_560_io_in_2),
    .io_in_3(c53_560_io_in_3),
    .io_in_4(c53_560_io_in_4),
    .io_out_0(c53_560_io_out_0),
    .io_out_1(c53_560_io_out_1),
    .io_out_2(c53_560_io_out_2)
  );
  C53 c53_561 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_561_io_in_0),
    .io_in_1(c53_561_io_in_1),
    .io_in_2(c53_561_io_in_2),
    .io_in_3(c53_561_io_in_3),
    .io_in_4(c53_561_io_in_4),
    .io_out_0(c53_561_io_out_0),
    .io_out_1(c53_561_io_out_1),
    .io_out_2(c53_561_io_out_2)
  );
  C22 c22_42 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_42_io_in_0),
    .io_in_1(c22_42_io_in_1),
    .io_out_0(c22_42_io_out_0),
    .io_out_1(c22_42_io_out_1)
  );
  C53 c53_562 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_562_io_in_0),
    .io_in_1(c53_562_io_in_1),
    .io_in_2(c53_562_io_in_2),
    .io_in_3(c53_562_io_in_3),
    .io_in_4(c53_562_io_in_4),
    .io_out_0(c53_562_io_out_0),
    .io_out_1(c53_562_io_out_1),
    .io_out_2(c53_562_io_out_2)
  );
  C53 c53_563 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_563_io_in_0),
    .io_in_1(c53_563_io_in_1),
    .io_in_2(c53_563_io_in_2),
    .io_in_3(c53_563_io_in_3),
    .io_in_4(c53_563_io_in_4),
    .io_out_0(c53_563_io_out_0),
    .io_out_1(c53_563_io_out_1),
    .io_out_2(c53_563_io_out_2)
  );
  C22 c22_43 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_43_io_in_0),
    .io_in_1(c22_43_io_in_1),
    .io_out_0(c22_43_io_out_0),
    .io_out_1(c22_43_io_out_1)
  );
  C53 c53_564 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_564_io_in_0),
    .io_in_1(c53_564_io_in_1),
    .io_in_2(c53_564_io_in_2),
    .io_in_3(c53_564_io_in_3),
    .io_in_4(c53_564_io_in_4),
    .io_out_0(c53_564_io_out_0),
    .io_out_1(c53_564_io_out_1),
    .io_out_2(c53_564_io_out_2)
  );
  C53 c53_565 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_565_io_in_0),
    .io_in_1(c53_565_io_in_1),
    .io_in_2(c53_565_io_in_2),
    .io_in_3(c53_565_io_in_3),
    .io_in_4(c53_565_io_in_4),
    .io_out_0(c53_565_io_out_0),
    .io_out_1(c53_565_io_out_1),
    .io_out_2(c53_565_io_out_2)
  );
  C22 c22_44 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_44_io_in_0),
    .io_in_1(c22_44_io_in_1),
    .io_out_0(c22_44_io_out_0),
    .io_out_1(c22_44_io_out_1)
  );
  C53 c53_566 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_566_io_in_0),
    .io_in_1(c53_566_io_in_1),
    .io_in_2(c53_566_io_in_2),
    .io_in_3(c53_566_io_in_3),
    .io_in_4(c53_566_io_in_4),
    .io_out_0(c53_566_io_out_0),
    .io_out_1(c53_566_io_out_1),
    .io_out_2(c53_566_io_out_2)
  );
  C53 c53_567 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_567_io_in_0),
    .io_in_1(c53_567_io_in_1),
    .io_in_2(c53_567_io_in_2),
    .io_in_3(c53_567_io_in_3),
    .io_in_4(c53_567_io_in_4),
    .io_out_0(c53_567_io_out_0),
    .io_out_1(c53_567_io_out_1),
    .io_out_2(c53_567_io_out_2)
  );
  C22 c22_45 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_45_io_in_0),
    .io_in_1(c22_45_io_in_1),
    .io_out_0(c22_45_io_out_0),
    .io_out_1(c22_45_io_out_1)
  );
  C53 c53_568 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_568_io_in_0),
    .io_in_1(c53_568_io_in_1),
    .io_in_2(c53_568_io_in_2),
    .io_in_3(c53_568_io_in_3),
    .io_in_4(c53_568_io_in_4),
    .io_out_0(c53_568_io_out_0),
    .io_out_1(c53_568_io_out_1),
    .io_out_2(c53_568_io_out_2)
  );
  C53 c53_569 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_569_io_in_0),
    .io_in_1(c53_569_io_in_1),
    .io_in_2(c53_569_io_in_2),
    .io_in_3(c53_569_io_in_3),
    .io_in_4(c53_569_io_in_4),
    .io_out_0(c53_569_io_out_0),
    .io_out_1(c53_569_io_out_1),
    .io_out_2(c53_569_io_out_2)
  );
  C22 c22_46 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_46_io_in_0),
    .io_in_1(c22_46_io_in_1),
    .io_out_0(c22_46_io_out_0),
    .io_out_1(c22_46_io_out_1)
  );
  C53 c53_570 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_570_io_in_0),
    .io_in_1(c53_570_io_in_1),
    .io_in_2(c53_570_io_in_2),
    .io_in_3(c53_570_io_in_3),
    .io_in_4(c53_570_io_in_4),
    .io_out_0(c53_570_io_out_0),
    .io_out_1(c53_570_io_out_1),
    .io_out_2(c53_570_io_out_2)
  );
  C53 c53_571 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_571_io_in_0),
    .io_in_1(c53_571_io_in_1),
    .io_in_2(c53_571_io_in_2),
    .io_in_3(c53_571_io_in_3),
    .io_in_4(c53_571_io_in_4),
    .io_out_0(c53_571_io_out_0),
    .io_out_1(c53_571_io_out_1),
    .io_out_2(c53_571_io_out_2)
  );
  C32 c32_38 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_38_io_in_0),
    .io_in_1(c32_38_io_in_1),
    .io_in_2(c32_38_io_in_2),
    .io_out_0(c32_38_io_out_0),
    .io_out_1(c32_38_io_out_1)
  );
  C53 c53_572 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_572_io_in_0),
    .io_in_1(c53_572_io_in_1),
    .io_in_2(c53_572_io_in_2),
    .io_in_3(c53_572_io_in_3),
    .io_in_4(c53_572_io_in_4),
    .io_out_0(c53_572_io_out_0),
    .io_out_1(c53_572_io_out_1),
    .io_out_2(c53_572_io_out_2)
  );
  C53 c53_573 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_573_io_in_0),
    .io_in_1(c53_573_io_in_1),
    .io_in_2(c53_573_io_in_2),
    .io_in_3(c53_573_io_in_3),
    .io_in_4(c53_573_io_in_4),
    .io_out_0(c53_573_io_out_0),
    .io_out_1(c53_573_io_out_1),
    .io_out_2(c53_573_io_out_2)
  );
  C32 c32_39 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_39_io_in_0),
    .io_in_1(c32_39_io_in_1),
    .io_in_2(c32_39_io_in_2),
    .io_out_0(c32_39_io_out_0),
    .io_out_1(c32_39_io_out_1)
  );
  C53 c53_574 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_574_io_in_0),
    .io_in_1(c53_574_io_in_1),
    .io_in_2(c53_574_io_in_2),
    .io_in_3(c53_574_io_in_3),
    .io_in_4(c53_574_io_in_4),
    .io_out_0(c53_574_io_out_0),
    .io_out_1(c53_574_io_out_1),
    .io_out_2(c53_574_io_out_2)
  );
  C53 c53_575 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_575_io_in_0),
    .io_in_1(c53_575_io_in_1),
    .io_in_2(c53_575_io_in_2),
    .io_in_3(c53_575_io_in_3),
    .io_in_4(c53_575_io_in_4),
    .io_out_0(c53_575_io_out_0),
    .io_out_1(c53_575_io_out_1),
    .io_out_2(c53_575_io_out_2)
  );
  C32 c32_40 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_40_io_in_0),
    .io_in_1(c32_40_io_in_1),
    .io_in_2(c32_40_io_in_2),
    .io_out_0(c32_40_io_out_0),
    .io_out_1(c32_40_io_out_1)
  );
  C53 c53_576 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_576_io_in_0),
    .io_in_1(c53_576_io_in_1),
    .io_in_2(c53_576_io_in_2),
    .io_in_3(c53_576_io_in_3),
    .io_in_4(c53_576_io_in_4),
    .io_out_0(c53_576_io_out_0),
    .io_out_1(c53_576_io_out_1),
    .io_out_2(c53_576_io_out_2)
  );
  C53 c53_577 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_577_io_in_0),
    .io_in_1(c53_577_io_in_1),
    .io_in_2(c53_577_io_in_2),
    .io_in_3(c53_577_io_in_3),
    .io_in_4(c53_577_io_in_4),
    .io_out_0(c53_577_io_out_0),
    .io_out_1(c53_577_io_out_1),
    .io_out_2(c53_577_io_out_2)
  );
  C53 c53_578 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_578_io_in_0),
    .io_in_1(c53_578_io_in_1),
    .io_in_2(c53_578_io_in_2),
    .io_in_3(c53_578_io_in_3),
    .io_in_4(c53_578_io_in_4),
    .io_out_0(c53_578_io_out_0),
    .io_out_1(c53_578_io_out_1),
    .io_out_2(c53_578_io_out_2)
  );
  C53 c53_579 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_579_io_in_0),
    .io_in_1(c53_579_io_in_1),
    .io_in_2(c53_579_io_in_2),
    .io_in_3(c53_579_io_in_3),
    .io_in_4(c53_579_io_in_4),
    .io_out_0(c53_579_io_out_0),
    .io_out_1(c53_579_io_out_1),
    .io_out_2(c53_579_io_out_2)
  );
  C53 c53_580 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_580_io_in_0),
    .io_in_1(c53_580_io_in_1),
    .io_in_2(c53_580_io_in_2),
    .io_in_3(c53_580_io_in_3),
    .io_in_4(c53_580_io_in_4),
    .io_out_0(c53_580_io_out_0),
    .io_out_1(c53_580_io_out_1),
    .io_out_2(c53_580_io_out_2)
  );
  C53 c53_581 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_581_io_in_0),
    .io_in_1(c53_581_io_in_1),
    .io_in_2(c53_581_io_in_2),
    .io_in_3(c53_581_io_in_3),
    .io_in_4(c53_581_io_in_4),
    .io_out_0(c53_581_io_out_0),
    .io_out_1(c53_581_io_out_1),
    .io_out_2(c53_581_io_out_2)
  );
  C53 c53_582 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_582_io_in_0),
    .io_in_1(c53_582_io_in_1),
    .io_in_2(c53_582_io_in_2),
    .io_in_3(c53_582_io_in_3),
    .io_in_4(c53_582_io_in_4),
    .io_out_0(c53_582_io_out_0),
    .io_out_1(c53_582_io_out_1),
    .io_out_2(c53_582_io_out_2)
  );
  C53 c53_583 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_583_io_in_0),
    .io_in_1(c53_583_io_in_1),
    .io_in_2(c53_583_io_in_2),
    .io_in_3(c53_583_io_in_3),
    .io_in_4(c53_583_io_in_4),
    .io_out_0(c53_583_io_out_0),
    .io_out_1(c53_583_io_out_1),
    .io_out_2(c53_583_io_out_2)
  );
  C53 c53_584 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_584_io_in_0),
    .io_in_1(c53_584_io_in_1),
    .io_in_2(c53_584_io_in_2),
    .io_in_3(c53_584_io_in_3),
    .io_in_4(c53_584_io_in_4),
    .io_out_0(c53_584_io_out_0),
    .io_out_1(c53_584_io_out_1),
    .io_out_2(c53_584_io_out_2)
  );
  C53 c53_585 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_585_io_in_0),
    .io_in_1(c53_585_io_in_1),
    .io_in_2(c53_585_io_in_2),
    .io_in_3(c53_585_io_in_3),
    .io_in_4(c53_585_io_in_4),
    .io_out_0(c53_585_io_out_0),
    .io_out_1(c53_585_io_out_1),
    .io_out_2(c53_585_io_out_2)
  );
  C53 c53_586 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_586_io_in_0),
    .io_in_1(c53_586_io_in_1),
    .io_in_2(c53_586_io_in_2),
    .io_in_3(c53_586_io_in_3),
    .io_in_4(c53_586_io_in_4),
    .io_out_0(c53_586_io_out_0),
    .io_out_1(c53_586_io_out_1),
    .io_out_2(c53_586_io_out_2)
  );
  C53 c53_587 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_587_io_in_0),
    .io_in_1(c53_587_io_in_1),
    .io_in_2(c53_587_io_in_2),
    .io_in_3(c53_587_io_in_3),
    .io_in_4(c53_587_io_in_4),
    .io_out_0(c53_587_io_out_0),
    .io_out_1(c53_587_io_out_1),
    .io_out_2(c53_587_io_out_2)
  );
  C53 c53_588 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_588_io_in_0),
    .io_in_1(c53_588_io_in_1),
    .io_in_2(c53_588_io_in_2),
    .io_in_3(c53_588_io_in_3),
    .io_in_4(c53_588_io_in_4),
    .io_out_0(c53_588_io_out_0),
    .io_out_1(c53_588_io_out_1),
    .io_out_2(c53_588_io_out_2)
  );
  C53 c53_589 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_589_io_in_0),
    .io_in_1(c53_589_io_in_1),
    .io_in_2(c53_589_io_in_2),
    .io_in_3(c53_589_io_in_3),
    .io_in_4(c53_589_io_in_4),
    .io_out_0(c53_589_io_out_0),
    .io_out_1(c53_589_io_out_1),
    .io_out_2(c53_589_io_out_2)
  );
  C53 c53_590 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_590_io_in_0),
    .io_in_1(c53_590_io_in_1),
    .io_in_2(c53_590_io_in_2),
    .io_in_3(c53_590_io_in_3),
    .io_in_4(c53_590_io_in_4),
    .io_out_0(c53_590_io_out_0),
    .io_out_1(c53_590_io_out_1),
    .io_out_2(c53_590_io_out_2)
  );
  C53 c53_591 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_591_io_in_0),
    .io_in_1(c53_591_io_in_1),
    .io_in_2(c53_591_io_in_2),
    .io_in_3(c53_591_io_in_3),
    .io_in_4(c53_591_io_in_4),
    .io_out_0(c53_591_io_out_0),
    .io_out_1(c53_591_io_out_1),
    .io_out_2(c53_591_io_out_2)
  );
  C53 c53_592 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_592_io_in_0),
    .io_in_1(c53_592_io_in_1),
    .io_in_2(c53_592_io_in_2),
    .io_in_3(c53_592_io_in_3),
    .io_in_4(c53_592_io_in_4),
    .io_out_0(c53_592_io_out_0),
    .io_out_1(c53_592_io_out_1),
    .io_out_2(c53_592_io_out_2)
  );
  C53 c53_593 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_593_io_in_0),
    .io_in_1(c53_593_io_in_1),
    .io_in_2(c53_593_io_in_2),
    .io_in_3(c53_593_io_in_3),
    .io_in_4(c53_593_io_in_4),
    .io_out_0(c53_593_io_out_0),
    .io_out_1(c53_593_io_out_1),
    .io_out_2(c53_593_io_out_2)
  );
  C53 c53_594 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_594_io_in_0),
    .io_in_1(c53_594_io_in_1),
    .io_in_2(c53_594_io_in_2),
    .io_in_3(c53_594_io_in_3),
    .io_in_4(c53_594_io_in_4),
    .io_out_0(c53_594_io_out_0),
    .io_out_1(c53_594_io_out_1),
    .io_out_2(c53_594_io_out_2)
  );
  C53 c53_595 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_595_io_in_0),
    .io_in_1(c53_595_io_in_1),
    .io_in_2(c53_595_io_in_2),
    .io_in_3(c53_595_io_in_3),
    .io_in_4(c53_595_io_in_4),
    .io_out_0(c53_595_io_out_0),
    .io_out_1(c53_595_io_out_1),
    .io_out_2(c53_595_io_out_2)
  );
  C53 c53_596 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_596_io_in_0),
    .io_in_1(c53_596_io_in_1),
    .io_in_2(c53_596_io_in_2),
    .io_in_3(c53_596_io_in_3),
    .io_in_4(c53_596_io_in_4),
    .io_out_0(c53_596_io_out_0),
    .io_out_1(c53_596_io_out_1),
    .io_out_2(c53_596_io_out_2)
  );
  C53 c53_597 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_597_io_in_0),
    .io_in_1(c53_597_io_in_1),
    .io_in_2(c53_597_io_in_2),
    .io_in_3(c53_597_io_in_3),
    .io_in_4(c53_597_io_in_4),
    .io_out_0(c53_597_io_out_0),
    .io_out_1(c53_597_io_out_1),
    .io_out_2(c53_597_io_out_2)
  );
  C53 c53_598 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_598_io_in_0),
    .io_in_1(c53_598_io_in_1),
    .io_in_2(c53_598_io_in_2),
    .io_in_3(c53_598_io_in_3),
    .io_in_4(c53_598_io_in_4),
    .io_out_0(c53_598_io_out_0),
    .io_out_1(c53_598_io_out_1),
    .io_out_2(c53_598_io_out_2)
  );
  C53 c53_599 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_599_io_in_0),
    .io_in_1(c53_599_io_in_1),
    .io_in_2(c53_599_io_in_2),
    .io_in_3(c53_599_io_in_3),
    .io_in_4(c53_599_io_in_4),
    .io_out_0(c53_599_io_out_0),
    .io_out_1(c53_599_io_out_1),
    .io_out_2(c53_599_io_out_2)
  );
  C53 c53_600 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_600_io_in_0),
    .io_in_1(c53_600_io_in_1),
    .io_in_2(c53_600_io_in_2),
    .io_in_3(c53_600_io_in_3),
    .io_in_4(c53_600_io_in_4),
    .io_out_0(c53_600_io_out_0),
    .io_out_1(c53_600_io_out_1),
    .io_out_2(c53_600_io_out_2)
  );
  C53 c53_601 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_601_io_in_0),
    .io_in_1(c53_601_io_in_1),
    .io_in_2(c53_601_io_in_2),
    .io_in_3(c53_601_io_in_3),
    .io_in_4(c53_601_io_in_4),
    .io_out_0(c53_601_io_out_0),
    .io_out_1(c53_601_io_out_1),
    .io_out_2(c53_601_io_out_2)
  );
  C53 c53_602 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_602_io_in_0),
    .io_in_1(c53_602_io_in_1),
    .io_in_2(c53_602_io_in_2),
    .io_in_3(c53_602_io_in_3),
    .io_in_4(c53_602_io_in_4),
    .io_out_0(c53_602_io_out_0),
    .io_out_1(c53_602_io_out_1),
    .io_out_2(c53_602_io_out_2)
  );
  C22 c22_47 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_47_io_in_0),
    .io_in_1(c22_47_io_in_1),
    .io_out_0(c22_47_io_out_0),
    .io_out_1(c22_47_io_out_1)
  );
  C53 c53_603 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_603_io_in_0),
    .io_in_1(c53_603_io_in_1),
    .io_in_2(c53_603_io_in_2),
    .io_in_3(c53_603_io_in_3),
    .io_in_4(c53_603_io_in_4),
    .io_out_0(c53_603_io_out_0),
    .io_out_1(c53_603_io_out_1),
    .io_out_2(c53_603_io_out_2)
  );
  C53 c53_604 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_604_io_in_0),
    .io_in_1(c53_604_io_in_1),
    .io_in_2(c53_604_io_in_2),
    .io_in_3(c53_604_io_in_3),
    .io_in_4(c53_604_io_in_4),
    .io_out_0(c53_604_io_out_0),
    .io_out_1(c53_604_io_out_1),
    .io_out_2(c53_604_io_out_2)
  );
  C53 c53_605 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_605_io_in_0),
    .io_in_1(c53_605_io_in_1),
    .io_in_2(c53_605_io_in_2),
    .io_in_3(c53_605_io_in_3),
    .io_in_4(c53_605_io_in_4),
    .io_out_0(c53_605_io_out_0),
    .io_out_1(c53_605_io_out_1),
    .io_out_2(c53_605_io_out_2)
  );
  C22 c22_48 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_48_io_in_0),
    .io_in_1(c22_48_io_in_1),
    .io_out_0(c22_48_io_out_0),
    .io_out_1(c22_48_io_out_1)
  );
  C53 c53_606 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_606_io_in_0),
    .io_in_1(c53_606_io_in_1),
    .io_in_2(c53_606_io_in_2),
    .io_in_3(c53_606_io_in_3),
    .io_in_4(c53_606_io_in_4),
    .io_out_0(c53_606_io_out_0),
    .io_out_1(c53_606_io_out_1),
    .io_out_2(c53_606_io_out_2)
  );
  C53 c53_607 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_607_io_in_0),
    .io_in_1(c53_607_io_in_1),
    .io_in_2(c53_607_io_in_2),
    .io_in_3(c53_607_io_in_3),
    .io_in_4(c53_607_io_in_4),
    .io_out_0(c53_607_io_out_0),
    .io_out_1(c53_607_io_out_1),
    .io_out_2(c53_607_io_out_2)
  );
  C53 c53_608 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_608_io_in_0),
    .io_in_1(c53_608_io_in_1),
    .io_in_2(c53_608_io_in_2),
    .io_in_3(c53_608_io_in_3),
    .io_in_4(c53_608_io_in_4),
    .io_out_0(c53_608_io_out_0),
    .io_out_1(c53_608_io_out_1),
    .io_out_2(c53_608_io_out_2)
  );
  C22 c22_49 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_49_io_in_0),
    .io_in_1(c22_49_io_in_1),
    .io_out_0(c22_49_io_out_0),
    .io_out_1(c22_49_io_out_1)
  );
  C53 c53_609 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_609_io_in_0),
    .io_in_1(c53_609_io_in_1),
    .io_in_2(c53_609_io_in_2),
    .io_in_3(c53_609_io_in_3),
    .io_in_4(c53_609_io_in_4),
    .io_out_0(c53_609_io_out_0),
    .io_out_1(c53_609_io_out_1),
    .io_out_2(c53_609_io_out_2)
  );
  C53 c53_610 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_610_io_in_0),
    .io_in_1(c53_610_io_in_1),
    .io_in_2(c53_610_io_in_2),
    .io_in_3(c53_610_io_in_3),
    .io_in_4(c53_610_io_in_4),
    .io_out_0(c53_610_io_out_0),
    .io_out_1(c53_610_io_out_1),
    .io_out_2(c53_610_io_out_2)
  );
  C53 c53_611 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_611_io_in_0),
    .io_in_1(c53_611_io_in_1),
    .io_in_2(c53_611_io_in_2),
    .io_in_3(c53_611_io_in_3),
    .io_in_4(c53_611_io_in_4),
    .io_out_0(c53_611_io_out_0),
    .io_out_1(c53_611_io_out_1),
    .io_out_2(c53_611_io_out_2)
  );
  C22 c22_50 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_50_io_in_0),
    .io_in_1(c22_50_io_in_1),
    .io_out_0(c22_50_io_out_0),
    .io_out_1(c22_50_io_out_1)
  );
  C53 c53_612 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_612_io_in_0),
    .io_in_1(c53_612_io_in_1),
    .io_in_2(c53_612_io_in_2),
    .io_in_3(c53_612_io_in_3),
    .io_in_4(c53_612_io_in_4),
    .io_out_0(c53_612_io_out_0),
    .io_out_1(c53_612_io_out_1),
    .io_out_2(c53_612_io_out_2)
  );
  C53 c53_613 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_613_io_in_0),
    .io_in_1(c53_613_io_in_1),
    .io_in_2(c53_613_io_in_2),
    .io_in_3(c53_613_io_in_3),
    .io_in_4(c53_613_io_in_4),
    .io_out_0(c53_613_io_out_0),
    .io_out_1(c53_613_io_out_1),
    .io_out_2(c53_613_io_out_2)
  );
  C53 c53_614 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_614_io_in_0),
    .io_in_1(c53_614_io_in_1),
    .io_in_2(c53_614_io_in_2),
    .io_in_3(c53_614_io_in_3),
    .io_in_4(c53_614_io_in_4),
    .io_out_0(c53_614_io_out_0),
    .io_out_1(c53_614_io_out_1),
    .io_out_2(c53_614_io_out_2)
  );
  C22 c22_51 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_51_io_in_0),
    .io_in_1(c22_51_io_in_1),
    .io_out_0(c22_51_io_out_0),
    .io_out_1(c22_51_io_out_1)
  );
  C53 c53_615 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_615_io_in_0),
    .io_in_1(c53_615_io_in_1),
    .io_in_2(c53_615_io_in_2),
    .io_in_3(c53_615_io_in_3),
    .io_in_4(c53_615_io_in_4),
    .io_out_0(c53_615_io_out_0),
    .io_out_1(c53_615_io_out_1),
    .io_out_2(c53_615_io_out_2)
  );
  C53 c53_616 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_616_io_in_0),
    .io_in_1(c53_616_io_in_1),
    .io_in_2(c53_616_io_in_2),
    .io_in_3(c53_616_io_in_3),
    .io_in_4(c53_616_io_in_4),
    .io_out_0(c53_616_io_out_0),
    .io_out_1(c53_616_io_out_1),
    .io_out_2(c53_616_io_out_2)
  );
  C53 c53_617 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_617_io_in_0),
    .io_in_1(c53_617_io_in_1),
    .io_in_2(c53_617_io_in_2),
    .io_in_3(c53_617_io_in_3),
    .io_in_4(c53_617_io_in_4),
    .io_out_0(c53_617_io_out_0),
    .io_out_1(c53_617_io_out_1),
    .io_out_2(c53_617_io_out_2)
  );
  C32 c32_41 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_41_io_in_0),
    .io_in_1(c32_41_io_in_1),
    .io_in_2(c32_41_io_in_2),
    .io_out_0(c32_41_io_out_0),
    .io_out_1(c32_41_io_out_1)
  );
  C53 c53_618 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_618_io_in_0),
    .io_in_1(c53_618_io_in_1),
    .io_in_2(c53_618_io_in_2),
    .io_in_3(c53_618_io_in_3),
    .io_in_4(c53_618_io_in_4),
    .io_out_0(c53_618_io_out_0),
    .io_out_1(c53_618_io_out_1),
    .io_out_2(c53_618_io_out_2)
  );
  C53 c53_619 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_619_io_in_0),
    .io_in_1(c53_619_io_in_1),
    .io_in_2(c53_619_io_in_2),
    .io_in_3(c53_619_io_in_3),
    .io_in_4(c53_619_io_in_4),
    .io_out_0(c53_619_io_out_0),
    .io_out_1(c53_619_io_out_1),
    .io_out_2(c53_619_io_out_2)
  );
  C53 c53_620 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_620_io_in_0),
    .io_in_1(c53_620_io_in_1),
    .io_in_2(c53_620_io_in_2),
    .io_in_3(c53_620_io_in_3),
    .io_in_4(c53_620_io_in_4),
    .io_out_0(c53_620_io_out_0),
    .io_out_1(c53_620_io_out_1),
    .io_out_2(c53_620_io_out_2)
  );
  C32 c32_42 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_42_io_in_0),
    .io_in_1(c32_42_io_in_1),
    .io_in_2(c32_42_io_in_2),
    .io_out_0(c32_42_io_out_0),
    .io_out_1(c32_42_io_out_1)
  );
  C53 c53_621 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_621_io_in_0),
    .io_in_1(c53_621_io_in_1),
    .io_in_2(c53_621_io_in_2),
    .io_in_3(c53_621_io_in_3),
    .io_in_4(c53_621_io_in_4),
    .io_out_0(c53_621_io_out_0),
    .io_out_1(c53_621_io_out_1),
    .io_out_2(c53_621_io_out_2)
  );
  C53 c53_622 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_622_io_in_0),
    .io_in_1(c53_622_io_in_1),
    .io_in_2(c53_622_io_in_2),
    .io_in_3(c53_622_io_in_3),
    .io_in_4(c53_622_io_in_4),
    .io_out_0(c53_622_io_out_0),
    .io_out_1(c53_622_io_out_1),
    .io_out_2(c53_622_io_out_2)
  );
  C53 c53_623 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_623_io_in_0),
    .io_in_1(c53_623_io_in_1),
    .io_in_2(c53_623_io_in_2),
    .io_in_3(c53_623_io_in_3),
    .io_in_4(c53_623_io_in_4),
    .io_out_0(c53_623_io_out_0),
    .io_out_1(c53_623_io_out_1),
    .io_out_2(c53_623_io_out_2)
  );
  C32 c32_43 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_43_io_in_0),
    .io_in_1(c32_43_io_in_1),
    .io_in_2(c32_43_io_in_2),
    .io_out_0(c32_43_io_out_0),
    .io_out_1(c32_43_io_out_1)
  );
  C53 c53_624 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_624_io_in_0),
    .io_in_1(c53_624_io_in_1),
    .io_in_2(c53_624_io_in_2),
    .io_in_3(c53_624_io_in_3),
    .io_in_4(c53_624_io_in_4),
    .io_out_0(c53_624_io_out_0),
    .io_out_1(c53_624_io_out_1),
    .io_out_2(c53_624_io_out_2)
  );
  C53 c53_625 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_625_io_in_0),
    .io_in_1(c53_625_io_in_1),
    .io_in_2(c53_625_io_in_2),
    .io_in_3(c53_625_io_in_3),
    .io_in_4(c53_625_io_in_4),
    .io_out_0(c53_625_io_out_0),
    .io_out_1(c53_625_io_out_1),
    .io_out_2(c53_625_io_out_2)
  );
  C53 c53_626 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_626_io_in_0),
    .io_in_1(c53_626_io_in_1),
    .io_in_2(c53_626_io_in_2),
    .io_in_3(c53_626_io_in_3),
    .io_in_4(c53_626_io_in_4),
    .io_out_0(c53_626_io_out_0),
    .io_out_1(c53_626_io_out_1),
    .io_out_2(c53_626_io_out_2)
  );
  C53 c53_627 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_627_io_in_0),
    .io_in_1(c53_627_io_in_1),
    .io_in_2(c53_627_io_in_2),
    .io_in_3(c53_627_io_in_3),
    .io_in_4(c53_627_io_in_4),
    .io_out_0(c53_627_io_out_0),
    .io_out_1(c53_627_io_out_1),
    .io_out_2(c53_627_io_out_2)
  );
  C53 c53_628 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_628_io_in_0),
    .io_in_1(c53_628_io_in_1),
    .io_in_2(c53_628_io_in_2),
    .io_in_3(c53_628_io_in_3),
    .io_in_4(c53_628_io_in_4),
    .io_out_0(c53_628_io_out_0),
    .io_out_1(c53_628_io_out_1),
    .io_out_2(c53_628_io_out_2)
  );
  C53 c53_629 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_629_io_in_0),
    .io_in_1(c53_629_io_in_1),
    .io_in_2(c53_629_io_in_2),
    .io_in_3(c53_629_io_in_3),
    .io_in_4(c53_629_io_in_4),
    .io_out_0(c53_629_io_out_0),
    .io_out_1(c53_629_io_out_1),
    .io_out_2(c53_629_io_out_2)
  );
  C53 c53_630 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_630_io_in_0),
    .io_in_1(c53_630_io_in_1),
    .io_in_2(c53_630_io_in_2),
    .io_in_3(c53_630_io_in_3),
    .io_in_4(c53_630_io_in_4),
    .io_out_0(c53_630_io_out_0),
    .io_out_1(c53_630_io_out_1),
    .io_out_2(c53_630_io_out_2)
  );
  C53 c53_631 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_631_io_in_0),
    .io_in_1(c53_631_io_in_1),
    .io_in_2(c53_631_io_in_2),
    .io_in_3(c53_631_io_in_3),
    .io_in_4(c53_631_io_in_4),
    .io_out_0(c53_631_io_out_0),
    .io_out_1(c53_631_io_out_1),
    .io_out_2(c53_631_io_out_2)
  );
  C53 c53_632 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_632_io_in_0),
    .io_in_1(c53_632_io_in_1),
    .io_in_2(c53_632_io_in_2),
    .io_in_3(c53_632_io_in_3),
    .io_in_4(c53_632_io_in_4),
    .io_out_0(c53_632_io_out_0),
    .io_out_1(c53_632_io_out_1),
    .io_out_2(c53_632_io_out_2)
  );
  C53 c53_633 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_633_io_in_0),
    .io_in_1(c53_633_io_in_1),
    .io_in_2(c53_633_io_in_2),
    .io_in_3(c53_633_io_in_3),
    .io_in_4(c53_633_io_in_4),
    .io_out_0(c53_633_io_out_0),
    .io_out_1(c53_633_io_out_1),
    .io_out_2(c53_633_io_out_2)
  );
  C53 c53_634 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_634_io_in_0),
    .io_in_1(c53_634_io_in_1),
    .io_in_2(c53_634_io_in_2),
    .io_in_3(c53_634_io_in_3),
    .io_in_4(c53_634_io_in_4),
    .io_out_0(c53_634_io_out_0),
    .io_out_1(c53_634_io_out_1),
    .io_out_2(c53_634_io_out_2)
  );
  C53 c53_635 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_635_io_in_0),
    .io_in_1(c53_635_io_in_1),
    .io_in_2(c53_635_io_in_2),
    .io_in_3(c53_635_io_in_3),
    .io_in_4(c53_635_io_in_4),
    .io_out_0(c53_635_io_out_0),
    .io_out_1(c53_635_io_out_1),
    .io_out_2(c53_635_io_out_2)
  );
  C53 c53_636 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_636_io_in_0),
    .io_in_1(c53_636_io_in_1),
    .io_in_2(c53_636_io_in_2),
    .io_in_3(c53_636_io_in_3),
    .io_in_4(c53_636_io_in_4),
    .io_out_0(c53_636_io_out_0),
    .io_out_1(c53_636_io_out_1),
    .io_out_2(c53_636_io_out_2)
  );
  C53 c53_637 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_637_io_in_0),
    .io_in_1(c53_637_io_in_1),
    .io_in_2(c53_637_io_in_2),
    .io_in_3(c53_637_io_in_3),
    .io_in_4(c53_637_io_in_4),
    .io_out_0(c53_637_io_out_0),
    .io_out_1(c53_637_io_out_1),
    .io_out_2(c53_637_io_out_2)
  );
  C53 c53_638 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_638_io_in_0),
    .io_in_1(c53_638_io_in_1),
    .io_in_2(c53_638_io_in_2),
    .io_in_3(c53_638_io_in_3),
    .io_in_4(c53_638_io_in_4),
    .io_out_0(c53_638_io_out_0),
    .io_out_1(c53_638_io_out_1),
    .io_out_2(c53_638_io_out_2)
  );
  C53 c53_639 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_639_io_in_0),
    .io_in_1(c53_639_io_in_1),
    .io_in_2(c53_639_io_in_2),
    .io_in_3(c53_639_io_in_3),
    .io_in_4(c53_639_io_in_4),
    .io_out_0(c53_639_io_out_0),
    .io_out_1(c53_639_io_out_1),
    .io_out_2(c53_639_io_out_2)
  );
  C53 c53_640 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_640_io_in_0),
    .io_in_1(c53_640_io_in_1),
    .io_in_2(c53_640_io_in_2),
    .io_in_3(c53_640_io_in_3),
    .io_in_4(c53_640_io_in_4),
    .io_out_0(c53_640_io_out_0),
    .io_out_1(c53_640_io_out_1),
    .io_out_2(c53_640_io_out_2)
  );
  C53 c53_641 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_641_io_in_0),
    .io_in_1(c53_641_io_in_1),
    .io_in_2(c53_641_io_in_2),
    .io_in_3(c53_641_io_in_3),
    .io_in_4(c53_641_io_in_4),
    .io_out_0(c53_641_io_out_0),
    .io_out_1(c53_641_io_out_1),
    .io_out_2(c53_641_io_out_2)
  );
  C53 c53_642 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_642_io_in_0),
    .io_in_1(c53_642_io_in_1),
    .io_in_2(c53_642_io_in_2),
    .io_in_3(c53_642_io_in_3),
    .io_in_4(c53_642_io_in_4),
    .io_out_0(c53_642_io_out_0),
    .io_out_1(c53_642_io_out_1),
    .io_out_2(c53_642_io_out_2)
  );
  C53 c53_643 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_643_io_in_0),
    .io_in_1(c53_643_io_in_1),
    .io_in_2(c53_643_io_in_2),
    .io_in_3(c53_643_io_in_3),
    .io_in_4(c53_643_io_in_4),
    .io_out_0(c53_643_io_out_0),
    .io_out_1(c53_643_io_out_1),
    .io_out_2(c53_643_io_out_2)
  );
  C53 c53_644 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_644_io_in_0),
    .io_in_1(c53_644_io_in_1),
    .io_in_2(c53_644_io_in_2),
    .io_in_3(c53_644_io_in_3),
    .io_in_4(c53_644_io_in_4),
    .io_out_0(c53_644_io_out_0),
    .io_out_1(c53_644_io_out_1),
    .io_out_2(c53_644_io_out_2)
  );
  C53 c53_645 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_645_io_in_0),
    .io_in_1(c53_645_io_in_1),
    .io_in_2(c53_645_io_in_2),
    .io_in_3(c53_645_io_in_3),
    .io_in_4(c53_645_io_in_4),
    .io_out_0(c53_645_io_out_0),
    .io_out_1(c53_645_io_out_1),
    .io_out_2(c53_645_io_out_2)
  );
  C53 c53_646 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_646_io_in_0),
    .io_in_1(c53_646_io_in_1),
    .io_in_2(c53_646_io_in_2),
    .io_in_3(c53_646_io_in_3),
    .io_in_4(c53_646_io_in_4),
    .io_out_0(c53_646_io_out_0),
    .io_out_1(c53_646_io_out_1),
    .io_out_2(c53_646_io_out_2)
  );
  C53 c53_647 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_647_io_in_0),
    .io_in_1(c53_647_io_in_1),
    .io_in_2(c53_647_io_in_2),
    .io_in_3(c53_647_io_in_3),
    .io_in_4(c53_647_io_in_4),
    .io_out_0(c53_647_io_out_0),
    .io_out_1(c53_647_io_out_1),
    .io_out_2(c53_647_io_out_2)
  );
  C53 c53_648 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_648_io_in_0),
    .io_in_1(c53_648_io_in_1),
    .io_in_2(c53_648_io_in_2),
    .io_in_3(c53_648_io_in_3),
    .io_in_4(c53_648_io_in_4),
    .io_out_0(c53_648_io_out_0),
    .io_out_1(c53_648_io_out_1),
    .io_out_2(c53_648_io_out_2)
  );
  C53 c53_649 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_649_io_in_0),
    .io_in_1(c53_649_io_in_1),
    .io_in_2(c53_649_io_in_2),
    .io_in_3(c53_649_io_in_3),
    .io_in_4(c53_649_io_in_4),
    .io_out_0(c53_649_io_out_0),
    .io_out_1(c53_649_io_out_1),
    .io_out_2(c53_649_io_out_2)
  );
  C53 c53_650 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_650_io_in_0),
    .io_in_1(c53_650_io_in_1),
    .io_in_2(c53_650_io_in_2),
    .io_in_3(c53_650_io_in_3),
    .io_in_4(c53_650_io_in_4),
    .io_out_0(c53_650_io_out_0),
    .io_out_1(c53_650_io_out_1),
    .io_out_2(c53_650_io_out_2)
  );
  C53 c53_651 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_651_io_in_0),
    .io_in_1(c53_651_io_in_1),
    .io_in_2(c53_651_io_in_2),
    .io_in_3(c53_651_io_in_3),
    .io_in_4(c53_651_io_in_4),
    .io_out_0(c53_651_io_out_0),
    .io_out_1(c53_651_io_out_1),
    .io_out_2(c53_651_io_out_2)
  );
  C53 c53_652 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_652_io_in_0),
    .io_in_1(c53_652_io_in_1),
    .io_in_2(c53_652_io_in_2),
    .io_in_3(c53_652_io_in_3),
    .io_in_4(c53_652_io_in_4),
    .io_out_0(c53_652_io_out_0),
    .io_out_1(c53_652_io_out_1),
    .io_out_2(c53_652_io_out_2)
  );
  C53 c53_653 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_653_io_in_0),
    .io_in_1(c53_653_io_in_1),
    .io_in_2(c53_653_io_in_2),
    .io_in_3(c53_653_io_in_3),
    .io_in_4(c53_653_io_in_4),
    .io_out_0(c53_653_io_out_0),
    .io_out_1(c53_653_io_out_1),
    .io_out_2(c53_653_io_out_2)
  );
  C53 c53_654 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_654_io_in_0),
    .io_in_1(c53_654_io_in_1),
    .io_in_2(c53_654_io_in_2),
    .io_in_3(c53_654_io_in_3),
    .io_in_4(c53_654_io_in_4),
    .io_out_0(c53_654_io_out_0),
    .io_out_1(c53_654_io_out_1),
    .io_out_2(c53_654_io_out_2)
  );
  C53 c53_655 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_655_io_in_0),
    .io_in_1(c53_655_io_in_1),
    .io_in_2(c53_655_io_in_2),
    .io_in_3(c53_655_io_in_3),
    .io_in_4(c53_655_io_in_4),
    .io_out_0(c53_655_io_out_0),
    .io_out_1(c53_655_io_out_1),
    .io_out_2(c53_655_io_out_2)
  );
  C53 c53_656 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_656_io_in_0),
    .io_in_1(c53_656_io_in_1),
    .io_in_2(c53_656_io_in_2),
    .io_in_3(c53_656_io_in_3),
    .io_in_4(c53_656_io_in_4),
    .io_out_0(c53_656_io_out_0),
    .io_out_1(c53_656_io_out_1),
    .io_out_2(c53_656_io_out_2)
  );
  C53 c53_657 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_657_io_in_0),
    .io_in_1(c53_657_io_in_1),
    .io_in_2(c53_657_io_in_2),
    .io_in_3(c53_657_io_in_3),
    .io_in_4(c53_657_io_in_4),
    .io_out_0(c53_657_io_out_0),
    .io_out_1(c53_657_io_out_1),
    .io_out_2(c53_657_io_out_2)
  );
  C53 c53_658 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_658_io_in_0),
    .io_in_1(c53_658_io_in_1),
    .io_in_2(c53_658_io_in_2),
    .io_in_3(c53_658_io_in_3),
    .io_in_4(c53_658_io_in_4),
    .io_out_0(c53_658_io_out_0),
    .io_out_1(c53_658_io_out_1),
    .io_out_2(c53_658_io_out_2)
  );
  C53 c53_659 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_659_io_in_0),
    .io_in_1(c53_659_io_in_1),
    .io_in_2(c53_659_io_in_2),
    .io_in_3(c53_659_io_in_3),
    .io_in_4(c53_659_io_in_4),
    .io_out_0(c53_659_io_out_0),
    .io_out_1(c53_659_io_out_1),
    .io_out_2(c53_659_io_out_2)
  );
  C53 c53_660 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_660_io_in_0),
    .io_in_1(c53_660_io_in_1),
    .io_in_2(c53_660_io_in_2),
    .io_in_3(c53_660_io_in_3),
    .io_in_4(c53_660_io_in_4),
    .io_out_0(c53_660_io_out_0),
    .io_out_1(c53_660_io_out_1),
    .io_out_2(c53_660_io_out_2)
  );
  C53 c53_661 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_661_io_in_0),
    .io_in_1(c53_661_io_in_1),
    .io_in_2(c53_661_io_in_2),
    .io_in_3(c53_661_io_in_3),
    .io_in_4(c53_661_io_in_4),
    .io_out_0(c53_661_io_out_0),
    .io_out_1(c53_661_io_out_1),
    .io_out_2(c53_661_io_out_2)
  );
  C53 c53_662 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_662_io_in_0),
    .io_in_1(c53_662_io_in_1),
    .io_in_2(c53_662_io_in_2),
    .io_in_3(c53_662_io_in_3),
    .io_in_4(c53_662_io_in_4),
    .io_out_0(c53_662_io_out_0),
    .io_out_1(c53_662_io_out_1),
    .io_out_2(c53_662_io_out_2)
  );
  C53 c53_663 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_663_io_in_0),
    .io_in_1(c53_663_io_in_1),
    .io_in_2(c53_663_io_in_2),
    .io_in_3(c53_663_io_in_3),
    .io_in_4(c53_663_io_in_4),
    .io_out_0(c53_663_io_out_0),
    .io_out_1(c53_663_io_out_1),
    .io_out_2(c53_663_io_out_2)
  );
  C53 c53_664 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_664_io_in_0),
    .io_in_1(c53_664_io_in_1),
    .io_in_2(c53_664_io_in_2),
    .io_in_3(c53_664_io_in_3),
    .io_in_4(c53_664_io_in_4),
    .io_out_0(c53_664_io_out_0),
    .io_out_1(c53_664_io_out_1),
    .io_out_2(c53_664_io_out_2)
  );
  C53 c53_665 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_665_io_in_0),
    .io_in_1(c53_665_io_in_1),
    .io_in_2(c53_665_io_in_2),
    .io_in_3(c53_665_io_in_3),
    .io_in_4(c53_665_io_in_4),
    .io_out_0(c53_665_io_out_0),
    .io_out_1(c53_665_io_out_1),
    .io_out_2(c53_665_io_out_2)
  );
  C53 c53_666 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_666_io_in_0),
    .io_in_1(c53_666_io_in_1),
    .io_in_2(c53_666_io_in_2),
    .io_in_3(c53_666_io_in_3),
    .io_in_4(c53_666_io_in_4),
    .io_out_0(c53_666_io_out_0),
    .io_out_1(c53_666_io_out_1),
    .io_out_2(c53_666_io_out_2)
  );
  C53 c53_667 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_667_io_in_0),
    .io_in_1(c53_667_io_in_1),
    .io_in_2(c53_667_io_in_2),
    .io_in_3(c53_667_io_in_3),
    .io_in_4(c53_667_io_in_4),
    .io_out_0(c53_667_io_out_0),
    .io_out_1(c53_667_io_out_1),
    .io_out_2(c53_667_io_out_2)
  );
  C53 c53_668 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_668_io_in_0),
    .io_in_1(c53_668_io_in_1),
    .io_in_2(c53_668_io_in_2),
    .io_in_3(c53_668_io_in_3),
    .io_in_4(c53_668_io_in_4),
    .io_out_0(c53_668_io_out_0),
    .io_out_1(c53_668_io_out_1),
    .io_out_2(c53_668_io_out_2)
  );
  C53 c53_669 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_669_io_in_0),
    .io_in_1(c53_669_io_in_1),
    .io_in_2(c53_669_io_in_2),
    .io_in_3(c53_669_io_in_3),
    .io_in_4(c53_669_io_in_4),
    .io_out_0(c53_669_io_out_0),
    .io_out_1(c53_669_io_out_1),
    .io_out_2(c53_669_io_out_2)
  );
  C53 c53_670 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_670_io_in_0),
    .io_in_1(c53_670_io_in_1),
    .io_in_2(c53_670_io_in_2),
    .io_in_3(c53_670_io_in_3),
    .io_in_4(c53_670_io_in_4),
    .io_out_0(c53_670_io_out_0),
    .io_out_1(c53_670_io_out_1),
    .io_out_2(c53_670_io_out_2)
  );
  C53 c53_671 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_671_io_in_0),
    .io_in_1(c53_671_io_in_1),
    .io_in_2(c53_671_io_in_2),
    .io_in_3(c53_671_io_in_3),
    .io_in_4(c53_671_io_in_4),
    .io_out_0(c53_671_io_out_0),
    .io_out_1(c53_671_io_out_1),
    .io_out_2(c53_671_io_out_2)
  );
  C53 c53_672 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_672_io_in_0),
    .io_in_1(c53_672_io_in_1),
    .io_in_2(c53_672_io_in_2),
    .io_in_3(c53_672_io_in_3),
    .io_in_4(c53_672_io_in_4),
    .io_out_0(c53_672_io_out_0),
    .io_out_1(c53_672_io_out_1),
    .io_out_2(c53_672_io_out_2)
  );
  C53 c53_673 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_673_io_in_0),
    .io_in_1(c53_673_io_in_1),
    .io_in_2(c53_673_io_in_2),
    .io_in_3(c53_673_io_in_3),
    .io_in_4(c53_673_io_in_4),
    .io_out_0(c53_673_io_out_0),
    .io_out_1(c53_673_io_out_1),
    .io_out_2(c53_673_io_out_2)
  );
  C53 c53_674 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_674_io_in_0),
    .io_in_1(c53_674_io_in_1),
    .io_in_2(c53_674_io_in_2),
    .io_in_3(c53_674_io_in_3),
    .io_in_4(c53_674_io_in_4),
    .io_out_0(c53_674_io_out_0),
    .io_out_1(c53_674_io_out_1),
    .io_out_2(c53_674_io_out_2)
  );
  C53 c53_675 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_675_io_in_0),
    .io_in_1(c53_675_io_in_1),
    .io_in_2(c53_675_io_in_2),
    .io_in_3(c53_675_io_in_3),
    .io_in_4(c53_675_io_in_4),
    .io_out_0(c53_675_io_out_0),
    .io_out_1(c53_675_io_out_1),
    .io_out_2(c53_675_io_out_2)
  );
  C53 c53_676 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_676_io_in_0),
    .io_in_1(c53_676_io_in_1),
    .io_in_2(c53_676_io_in_2),
    .io_in_3(c53_676_io_in_3),
    .io_in_4(c53_676_io_in_4),
    .io_out_0(c53_676_io_out_0),
    .io_out_1(c53_676_io_out_1),
    .io_out_2(c53_676_io_out_2)
  );
  C53 c53_677 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_677_io_in_0),
    .io_in_1(c53_677_io_in_1),
    .io_in_2(c53_677_io_in_2),
    .io_in_3(c53_677_io_in_3),
    .io_in_4(c53_677_io_in_4),
    .io_out_0(c53_677_io_out_0),
    .io_out_1(c53_677_io_out_1),
    .io_out_2(c53_677_io_out_2)
  );
  C53 c53_678 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_678_io_in_0),
    .io_in_1(c53_678_io_in_1),
    .io_in_2(c53_678_io_in_2),
    .io_in_3(c53_678_io_in_3),
    .io_in_4(c53_678_io_in_4),
    .io_out_0(c53_678_io_out_0),
    .io_out_1(c53_678_io_out_1),
    .io_out_2(c53_678_io_out_2)
  );
  C53 c53_679 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_679_io_in_0),
    .io_in_1(c53_679_io_in_1),
    .io_in_2(c53_679_io_in_2),
    .io_in_3(c53_679_io_in_3),
    .io_in_4(c53_679_io_in_4),
    .io_out_0(c53_679_io_out_0),
    .io_out_1(c53_679_io_out_1),
    .io_out_2(c53_679_io_out_2)
  );
  C53 c53_680 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_680_io_in_0),
    .io_in_1(c53_680_io_in_1),
    .io_in_2(c53_680_io_in_2),
    .io_in_3(c53_680_io_in_3),
    .io_in_4(c53_680_io_in_4),
    .io_out_0(c53_680_io_out_0),
    .io_out_1(c53_680_io_out_1),
    .io_out_2(c53_680_io_out_2)
  );
  C53 c53_681 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_681_io_in_0),
    .io_in_1(c53_681_io_in_1),
    .io_in_2(c53_681_io_in_2),
    .io_in_3(c53_681_io_in_3),
    .io_in_4(c53_681_io_in_4),
    .io_out_0(c53_681_io_out_0),
    .io_out_1(c53_681_io_out_1),
    .io_out_2(c53_681_io_out_2)
  );
  C53 c53_682 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_682_io_in_0),
    .io_in_1(c53_682_io_in_1),
    .io_in_2(c53_682_io_in_2),
    .io_in_3(c53_682_io_in_3),
    .io_in_4(c53_682_io_in_4),
    .io_out_0(c53_682_io_out_0),
    .io_out_1(c53_682_io_out_1),
    .io_out_2(c53_682_io_out_2)
  );
  C53 c53_683 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_683_io_in_0),
    .io_in_1(c53_683_io_in_1),
    .io_in_2(c53_683_io_in_2),
    .io_in_3(c53_683_io_in_3),
    .io_in_4(c53_683_io_in_4),
    .io_out_0(c53_683_io_out_0),
    .io_out_1(c53_683_io_out_1),
    .io_out_2(c53_683_io_out_2)
  );
  C53 c53_684 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_684_io_in_0),
    .io_in_1(c53_684_io_in_1),
    .io_in_2(c53_684_io_in_2),
    .io_in_3(c53_684_io_in_3),
    .io_in_4(c53_684_io_in_4),
    .io_out_0(c53_684_io_out_0),
    .io_out_1(c53_684_io_out_1),
    .io_out_2(c53_684_io_out_2)
  );
  C53 c53_685 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_685_io_in_0),
    .io_in_1(c53_685_io_in_1),
    .io_in_2(c53_685_io_in_2),
    .io_in_3(c53_685_io_in_3),
    .io_in_4(c53_685_io_in_4),
    .io_out_0(c53_685_io_out_0),
    .io_out_1(c53_685_io_out_1),
    .io_out_2(c53_685_io_out_2)
  );
  C53 c53_686 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_686_io_in_0),
    .io_in_1(c53_686_io_in_1),
    .io_in_2(c53_686_io_in_2),
    .io_in_3(c53_686_io_in_3),
    .io_in_4(c53_686_io_in_4),
    .io_out_0(c53_686_io_out_0),
    .io_out_1(c53_686_io_out_1),
    .io_out_2(c53_686_io_out_2)
  );
  C53 c53_687 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_687_io_in_0),
    .io_in_1(c53_687_io_in_1),
    .io_in_2(c53_687_io_in_2),
    .io_in_3(c53_687_io_in_3),
    .io_in_4(c53_687_io_in_4),
    .io_out_0(c53_687_io_out_0),
    .io_out_1(c53_687_io_out_1),
    .io_out_2(c53_687_io_out_2)
  );
  C53 c53_688 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_688_io_in_0),
    .io_in_1(c53_688_io_in_1),
    .io_in_2(c53_688_io_in_2),
    .io_in_3(c53_688_io_in_3),
    .io_in_4(c53_688_io_in_4),
    .io_out_0(c53_688_io_out_0),
    .io_out_1(c53_688_io_out_1),
    .io_out_2(c53_688_io_out_2)
  );
  C53 c53_689 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_689_io_in_0),
    .io_in_1(c53_689_io_in_1),
    .io_in_2(c53_689_io_in_2),
    .io_in_3(c53_689_io_in_3),
    .io_in_4(c53_689_io_in_4),
    .io_out_0(c53_689_io_out_0),
    .io_out_1(c53_689_io_out_1),
    .io_out_2(c53_689_io_out_2)
  );
  C53 c53_690 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_690_io_in_0),
    .io_in_1(c53_690_io_in_1),
    .io_in_2(c53_690_io_in_2),
    .io_in_3(c53_690_io_in_3),
    .io_in_4(c53_690_io_in_4),
    .io_out_0(c53_690_io_out_0),
    .io_out_1(c53_690_io_out_1),
    .io_out_2(c53_690_io_out_2)
  );
  C53 c53_691 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_691_io_in_0),
    .io_in_1(c53_691_io_in_1),
    .io_in_2(c53_691_io_in_2),
    .io_in_3(c53_691_io_in_3),
    .io_in_4(c53_691_io_in_4),
    .io_out_0(c53_691_io_out_0),
    .io_out_1(c53_691_io_out_1),
    .io_out_2(c53_691_io_out_2)
  );
  C53 c53_692 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_692_io_in_0),
    .io_in_1(c53_692_io_in_1),
    .io_in_2(c53_692_io_in_2),
    .io_in_3(c53_692_io_in_3),
    .io_in_4(c53_692_io_in_4),
    .io_out_0(c53_692_io_out_0),
    .io_out_1(c53_692_io_out_1),
    .io_out_2(c53_692_io_out_2)
  );
  C53 c53_693 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_693_io_in_0),
    .io_in_1(c53_693_io_in_1),
    .io_in_2(c53_693_io_in_2),
    .io_in_3(c53_693_io_in_3),
    .io_in_4(c53_693_io_in_4),
    .io_out_0(c53_693_io_out_0),
    .io_out_1(c53_693_io_out_1),
    .io_out_2(c53_693_io_out_2)
  );
  C53 c53_694 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_694_io_in_0),
    .io_in_1(c53_694_io_in_1),
    .io_in_2(c53_694_io_in_2),
    .io_in_3(c53_694_io_in_3),
    .io_in_4(c53_694_io_in_4),
    .io_out_0(c53_694_io_out_0),
    .io_out_1(c53_694_io_out_1),
    .io_out_2(c53_694_io_out_2)
  );
  C53 c53_695 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_695_io_in_0),
    .io_in_1(c53_695_io_in_1),
    .io_in_2(c53_695_io_in_2),
    .io_in_3(c53_695_io_in_3),
    .io_in_4(c53_695_io_in_4),
    .io_out_0(c53_695_io_out_0),
    .io_out_1(c53_695_io_out_1),
    .io_out_2(c53_695_io_out_2)
  );
  C53 c53_696 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_696_io_in_0),
    .io_in_1(c53_696_io_in_1),
    .io_in_2(c53_696_io_in_2),
    .io_in_3(c53_696_io_in_3),
    .io_in_4(c53_696_io_in_4),
    .io_out_0(c53_696_io_out_0),
    .io_out_1(c53_696_io_out_1),
    .io_out_2(c53_696_io_out_2)
  );
  C53 c53_697 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_697_io_in_0),
    .io_in_1(c53_697_io_in_1),
    .io_in_2(c53_697_io_in_2),
    .io_in_3(c53_697_io_in_3),
    .io_in_4(c53_697_io_in_4),
    .io_out_0(c53_697_io_out_0),
    .io_out_1(c53_697_io_out_1),
    .io_out_2(c53_697_io_out_2)
  );
  C53 c53_698 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_698_io_in_0),
    .io_in_1(c53_698_io_in_1),
    .io_in_2(c53_698_io_in_2),
    .io_in_3(c53_698_io_in_3),
    .io_in_4(c53_698_io_in_4),
    .io_out_0(c53_698_io_out_0),
    .io_out_1(c53_698_io_out_1),
    .io_out_2(c53_698_io_out_2)
  );
  C32 c32_44 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_44_io_in_0),
    .io_in_1(c32_44_io_in_1),
    .io_in_2(c32_44_io_in_2),
    .io_out_0(c32_44_io_out_0),
    .io_out_1(c32_44_io_out_1)
  );
  C53 c53_699 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_699_io_in_0),
    .io_in_1(c53_699_io_in_1),
    .io_in_2(c53_699_io_in_2),
    .io_in_3(c53_699_io_in_3),
    .io_in_4(c53_699_io_in_4),
    .io_out_0(c53_699_io_out_0),
    .io_out_1(c53_699_io_out_1),
    .io_out_2(c53_699_io_out_2)
  );
  C53 c53_700 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_700_io_in_0),
    .io_in_1(c53_700_io_in_1),
    .io_in_2(c53_700_io_in_2),
    .io_in_3(c53_700_io_in_3),
    .io_in_4(c53_700_io_in_4),
    .io_out_0(c53_700_io_out_0),
    .io_out_1(c53_700_io_out_1),
    .io_out_2(c53_700_io_out_2)
  );
  C53 c53_701 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_701_io_in_0),
    .io_in_1(c53_701_io_in_1),
    .io_in_2(c53_701_io_in_2),
    .io_in_3(c53_701_io_in_3),
    .io_in_4(c53_701_io_in_4),
    .io_out_0(c53_701_io_out_0),
    .io_out_1(c53_701_io_out_1),
    .io_out_2(c53_701_io_out_2)
  );
  C22 c22_52 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_52_io_in_0),
    .io_in_1(c22_52_io_in_1),
    .io_out_0(c22_52_io_out_0),
    .io_out_1(c22_52_io_out_1)
  );
  C53 c53_702 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_702_io_in_0),
    .io_in_1(c53_702_io_in_1),
    .io_in_2(c53_702_io_in_2),
    .io_in_3(c53_702_io_in_3),
    .io_in_4(c53_702_io_in_4),
    .io_out_0(c53_702_io_out_0),
    .io_out_1(c53_702_io_out_1),
    .io_out_2(c53_702_io_out_2)
  );
  C53 c53_703 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_703_io_in_0),
    .io_in_1(c53_703_io_in_1),
    .io_in_2(c53_703_io_in_2),
    .io_in_3(c53_703_io_in_3),
    .io_in_4(c53_703_io_in_4),
    .io_out_0(c53_703_io_out_0),
    .io_out_1(c53_703_io_out_1),
    .io_out_2(c53_703_io_out_2)
  );
  C53 c53_704 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_704_io_in_0),
    .io_in_1(c53_704_io_in_1),
    .io_in_2(c53_704_io_in_2),
    .io_in_3(c53_704_io_in_3),
    .io_in_4(c53_704_io_in_4),
    .io_out_0(c53_704_io_out_0),
    .io_out_1(c53_704_io_out_1),
    .io_out_2(c53_704_io_out_2)
  );
  C22 c22_53 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_53_io_in_0),
    .io_in_1(c22_53_io_in_1),
    .io_out_0(c22_53_io_out_0),
    .io_out_1(c22_53_io_out_1)
  );
  C53 c53_705 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_705_io_in_0),
    .io_in_1(c53_705_io_in_1),
    .io_in_2(c53_705_io_in_2),
    .io_in_3(c53_705_io_in_3),
    .io_in_4(c53_705_io_in_4),
    .io_out_0(c53_705_io_out_0),
    .io_out_1(c53_705_io_out_1),
    .io_out_2(c53_705_io_out_2)
  );
  C53 c53_706 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_706_io_in_0),
    .io_in_1(c53_706_io_in_1),
    .io_in_2(c53_706_io_in_2),
    .io_in_3(c53_706_io_in_3),
    .io_in_4(c53_706_io_in_4),
    .io_out_0(c53_706_io_out_0),
    .io_out_1(c53_706_io_out_1),
    .io_out_2(c53_706_io_out_2)
  );
  C53 c53_707 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_707_io_in_0),
    .io_in_1(c53_707_io_in_1),
    .io_in_2(c53_707_io_in_2),
    .io_in_3(c53_707_io_in_3),
    .io_in_4(c53_707_io_in_4),
    .io_out_0(c53_707_io_out_0),
    .io_out_1(c53_707_io_out_1),
    .io_out_2(c53_707_io_out_2)
  );
  C32 c32_45 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_45_io_in_0),
    .io_in_1(c32_45_io_in_1),
    .io_in_2(c32_45_io_in_2),
    .io_out_0(c32_45_io_out_0),
    .io_out_1(c32_45_io_out_1)
  );
  C53 c53_708 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_708_io_in_0),
    .io_in_1(c53_708_io_in_1),
    .io_in_2(c53_708_io_in_2),
    .io_in_3(c53_708_io_in_3),
    .io_in_4(c53_708_io_in_4),
    .io_out_0(c53_708_io_out_0),
    .io_out_1(c53_708_io_out_1),
    .io_out_2(c53_708_io_out_2)
  );
  C53 c53_709 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_709_io_in_0),
    .io_in_1(c53_709_io_in_1),
    .io_in_2(c53_709_io_in_2),
    .io_in_3(c53_709_io_in_3),
    .io_in_4(c53_709_io_in_4),
    .io_out_0(c53_709_io_out_0),
    .io_out_1(c53_709_io_out_1),
    .io_out_2(c53_709_io_out_2)
  );
  C53 c53_710 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_710_io_in_0),
    .io_in_1(c53_710_io_in_1),
    .io_in_2(c53_710_io_in_2),
    .io_in_3(c53_710_io_in_3),
    .io_in_4(c53_710_io_in_4),
    .io_out_0(c53_710_io_out_0),
    .io_out_1(c53_710_io_out_1),
    .io_out_2(c53_710_io_out_2)
  );
  C22 c22_54 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_54_io_in_0),
    .io_in_1(c22_54_io_in_1),
    .io_out_0(c22_54_io_out_0),
    .io_out_1(c22_54_io_out_1)
  );
  C53 c53_711 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_711_io_in_0),
    .io_in_1(c53_711_io_in_1),
    .io_in_2(c53_711_io_in_2),
    .io_in_3(c53_711_io_in_3),
    .io_in_4(c53_711_io_in_4),
    .io_out_0(c53_711_io_out_0),
    .io_out_1(c53_711_io_out_1),
    .io_out_2(c53_711_io_out_2)
  );
  C53 c53_712 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_712_io_in_0),
    .io_in_1(c53_712_io_in_1),
    .io_in_2(c53_712_io_in_2),
    .io_in_3(c53_712_io_in_3),
    .io_in_4(c53_712_io_in_4),
    .io_out_0(c53_712_io_out_0),
    .io_out_1(c53_712_io_out_1),
    .io_out_2(c53_712_io_out_2)
  );
  C53 c53_713 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_713_io_in_0),
    .io_in_1(c53_713_io_in_1),
    .io_in_2(c53_713_io_in_2),
    .io_in_3(c53_713_io_in_3),
    .io_in_4(c53_713_io_in_4),
    .io_out_0(c53_713_io_out_0),
    .io_out_1(c53_713_io_out_1),
    .io_out_2(c53_713_io_out_2)
  );
  C22 c22_55 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_55_io_in_0),
    .io_in_1(c22_55_io_in_1),
    .io_out_0(c22_55_io_out_0),
    .io_out_1(c22_55_io_out_1)
  );
  C53 c53_714 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_714_io_in_0),
    .io_in_1(c53_714_io_in_1),
    .io_in_2(c53_714_io_in_2),
    .io_in_3(c53_714_io_in_3),
    .io_in_4(c53_714_io_in_4),
    .io_out_0(c53_714_io_out_0),
    .io_out_1(c53_714_io_out_1),
    .io_out_2(c53_714_io_out_2)
  );
  C53 c53_715 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_715_io_in_0),
    .io_in_1(c53_715_io_in_1),
    .io_in_2(c53_715_io_in_2),
    .io_in_3(c53_715_io_in_3),
    .io_in_4(c53_715_io_in_4),
    .io_out_0(c53_715_io_out_0),
    .io_out_1(c53_715_io_out_1),
    .io_out_2(c53_715_io_out_2)
  );
  C53 c53_716 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_716_io_in_0),
    .io_in_1(c53_716_io_in_1),
    .io_in_2(c53_716_io_in_2),
    .io_in_3(c53_716_io_in_3),
    .io_in_4(c53_716_io_in_4),
    .io_out_0(c53_716_io_out_0),
    .io_out_1(c53_716_io_out_1),
    .io_out_2(c53_716_io_out_2)
  );
  C22 c22_56 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_56_io_in_0),
    .io_in_1(c22_56_io_in_1),
    .io_out_0(c22_56_io_out_0),
    .io_out_1(c22_56_io_out_1)
  );
  C53 c53_717 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_717_io_in_0),
    .io_in_1(c53_717_io_in_1),
    .io_in_2(c53_717_io_in_2),
    .io_in_3(c53_717_io_in_3),
    .io_in_4(c53_717_io_in_4),
    .io_out_0(c53_717_io_out_0),
    .io_out_1(c53_717_io_out_1),
    .io_out_2(c53_717_io_out_2)
  );
  C53 c53_718 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_718_io_in_0),
    .io_in_1(c53_718_io_in_1),
    .io_in_2(c53_718_io_in_2),
    .io_in_3(c53_718_io_in_3),
    .io_in_4(c53_718_io_in_4),
    .io_out_0(c53_718_io_out_0),
    .io_out_1(c53_718_io_out_1),
    .io_out_2(c53_718_io_out_2)
  );
  C53 c53_719 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_719_io_in_0),
    .io_in_1(c53_719_io_in_1),
    .io_in_2(c53_719_io_in_2),
    .io_in_3(c53_719_io_in_3),
    .io_in_4(c53_719_io_in_4),
    .io_out_0(c53_719_io_out_0),
    .io_out_1(c53_719_io_out_1),
    .io_out_2(c53_719_io_out_2)
  );
  C22 c22_57 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_57_io_in_0),
    .io_in_1(c22_57_io_in_1),
    .io_out_0(c22_57_io_out_0),
    .io_out_1(c22_57_io_out_1)
  );
  C53 c53_720 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_720_io_in_0),
    .io_in_1(c53_720_io_in_1),
    .io_in_2(c53_720_io_in_2),
    .io_in_3(c53_720_io_in_3),
    .io_in_4(c53_720_io_in_4),
    .io_out_0(c53_720_io_out_0),
    .io_out_1(c53_720_io_out_1),
    .io_out_2(c53_720_io_out_2)
  );
  C53 c53_721 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_721_io_in_0),
    .io_in_1(c53_721_io_in_1),
    .io_in_2(c53_721_io_in_2),
    .io_in_3(c53_721_io_in_3),
    .io_in_4(c53_721_io_in_4),
    .io_out_0(c53_721_io_out_0),
    .io_out_1(c53_721_io_out_1),
    .io_out_2(c53_721_io_out_2)
  );
  C53 c53_722 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_722_io_in_0),
    .io_in_1(c53_722_io_in_1),
    .io_in_2(c53_722_io_in_2),
    .io_in_3(c53_722_io_in_3),
    .io_in_4(c53_722_io_in_4),
    .io_out_0(c53_722_io_out_0),
    .io_out_1(c53_722_io_out_1),
    .io_out_2(c53_722_io_out_2)
  );
  C53 c53_723 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_723_io_in_0),
    .io_in_1(c53_723_io_in_1),
    .io_in_2(c53_723_io_in_2),
    .io_in_3(c53_723_io_in_3),
    .io_in_4(c53_723_io_in_4),
    .io_out_0(c53_723_io_out_0),
    .io_out_1(c53_723_io_out_1),
    .io_out_2(c53_723_io_out_2)
  );
  C53 c53_724 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_724_io_in_0),
    .io_in_1(c53_724_io_in_1),
    .io_in_2(c53_724_io_in_2),
    .io_in_3(c53_724_io_in_3),
    .io_in_4(c53_724_io_in_4),
    .io_out_0(c53_724_io_out_0),
    .io_out_1(c53_724_io_out_1),
    .io_out_2(c53_724_io_out_2)
  );
  C53 c53_725 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_725_io_in_0),
    .io_in_1(c53_725_io_in_1),
    .io_in_2(c53_725_io_in_2),
    .io_in_3(c53_725_io_in_3),
    .io_in_4(c53_725_io_in_4),
    .io_out_0(c53_725_io_out_0),
    .io_out_1(c53_725_io_out_1),
    .io_out_2(c53_725_io_out_2)
  );
  C53 c53_726 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_726_io_in_0),
    .io_in_1(c53_726_io_in_1),
    .io_in_2(c53_726_io_in_2),
    .io_in_3(c53_726_io_in_3),
    .io_in_4(c53_726_io_in_4),
    .io_out_0(c53_726_io_out_0),
    .io_out_1(c53_726_io_out_1),
    .io_out_2(c53_726_io_out_2)
  );
  C53 c53_727 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_727_io_in_0),
    .io_in_1(c53_727_io_in_1),
    .io_in_2(c53_727_io_in_2),
    .io_in_3(c53_727_io_in_3),
    .io_in_4(c53_727_io_in_4),
    .io_out_0(c53_727_io_out_0),
    .io_out_1(c53_727_io_out_1),
    .io_out_2(c53_727_io_out_2)
  );
  C53 c53_728 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_728_io_in_0),
    .io_in_1(c53_728_io_in_1),
    .io_in_2(c53_728_io_in_2),
    .io_in_3(c53_728_io_in_3),
    .io_in_4(c53_728_io_in_4),
    .io_out_0(c53_728_io_out_0),
    .io_out_1(c53_728_io_out_1),
    .io_out_2(c53_728_io_out_2)
  );
  C53 c53_729 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_729_io_in_0),
    .io_in_1(c53_729_io_in_1),
    .io_in_2(c53_729_io_in_2),
    .io_in_3(c53_729_io_in_3),
    .io_in_4(c53_729_io_in_4),
    .io_out_0(c53_729_io_out_0),
    .io_out_1(c53_729_io_out_1),
    .io_out_2(c53_729_io_out_2)
  );
  C53 c53_730 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_730_io_in_0),
    .io_in_1(c53_730_io_in_1),
    .io_in_2(c53_730_io_in_2),
    .io_in_3(c53_730_io_in_3),
    .io_in_4(c53_730_io_in_4),
    .io_out_0(c53_730_io_out_0),
    .io_out_1(c53_730_io_out_1),
    .io_out_2(c53_730_io_out_2)
  );
  C53 c53_731 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_731_io_in_0),
    .io_in_1(c53_731_io_in_1),
    .io_in_2(c53_731_io_in_2),
    .io_in_3(c53_731_io_in_3),
    .io_in_4(c53_731_io_in_4),
    .io_out_0(c53_731_io_out_0),
    .io_out_1(c53_731_io_out_1),
    .io_out_2(c53_731_io_out_2)
  );
  C53 c53_732 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_732_io_in_0),
    .io_in_1(c53_732_io_in_1),
    .io_in_2(c53_732_io_in_2),
    .io_in_3(c53_732_io_in_3),
    .io_in_4(c53_732_io_in_4),
    .io_out_0(c53_732_io_out_0),
    .io_out_1(c53_732_io_out_1),
    .io_out_2(c53_732_io_out_2)
  );
  C53 c53_733 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_733_io_in_0),
    .io_in_1(c53_733_io_in_1),
    .io_in_2(c53_733_io_in_2),
    .io_in_3(c53_733_io_in_3),
    .io_in_4(c53_733_io_in_4),
    .io_out_0(c53_733_io_out_0),
    .io_out_1(c53_733_io_out_1),
    .io_out_2(c53_733_io_out_2)
  );
  C53 c53_734 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_734_io_in_0),
    .io_in_1(c53_734_io_in_1),
    .io_in_2(c53_734_io_in_2),
    .io_in_3(c53_734_io_in_3),
    .io_in_4(c53_734_io_in_4),
    .io_out_0(c53_734_io_out_0),
    .io_out_1(c53_734_io_out_1),
    .io_out_2(c53_734_io_out_2)
  );
  C53 c53_735 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_735_io_in_0),
    .io_in_1(c53_735_io_in_1),
    .io_in_2(c53_735_io_in_2),
    .io_in_3(c53_735_io_in_3),
    .io_in_4(c53_735_io_in_4),
    .io_out_0(c53_735_io_out_0),
    .io_out_1(c53_735_io_out_1),
    .io_out_2(c53_735_io_out_2)
  );
  C53 c53_736 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_736_io_in_0),
    .io_in_1(c53_736_io_in_1),
    .io_in_2(c53_736_io_in_2),
    .io_in_3(c53_736_io_in_3),
    .io_in_4(c53_736_io_in_4),
    .io_out_0(c53_736_io_out_0),
    .io_out_1(c53_736_io_out_1),
    .io_out_2(c53_736_io_out_2)
  );
  C53 c53_737 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_737_io_in_0),
    .io_in_1(c53_737_io_in_1),
    .io_in_2(c53_737_io_in_2),
    .io_in_3(c53_737_io_in_3),
    .io_in_4(c53_737_io_in_4),
    .io_out_0(c53_737_io_out_0),
    .io_out_1(c53_737_io_out_1),
    .io_out_2(c53_737_io_out_2)
  );
  C53 c53_738 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_738_io_in_0),
    .io_in_1(c53_738_io_in_1),
    .io_in_2(c53_738_io_in_2),
    .io_in_3(c53_738_io_in_3),
    .io_in_4(c53_738_io_in_4),
    .io_out_0(c53_738_io_out_0),
    .io_out_1(c53_738_io_out_1),
    .io_out_2(c53_738_io_out_2)
  );
  C53 c53_739 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_739_io_in_0),
    .io_in_1(c53_739_io_in_1),
    .io_in_2(c53_739_io_in_2),
    .io_in_3(c53_739_io_in_3),
    .io_in_4(c53_739_io_in_4),
    .io_out_0(c53_739_io_out_0),
    .io_out_1(c53_739_io_out_1),
    .io_out_2(c53_739_io_out_2)
  );
  C53 c53_740 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_740_io_in_0),
    .io_in_1(c53_740_io_in_1),
    .io_in_2(c53_740_io_in_2),
    .io_in_3(c53_740_io_in_3),
    .io_in_4(c53_740_io_in_4),
    .io_out_0(c53_740_io_out_0),
    .io_out_1(c53_740_io_out_1),
    .io_out_2(c53_740_io_out_2)
  );
  C53 c53_741 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_741_io_in_0),
    .io_in_1(c53_741_io_in_1),
    .io_in_2(c53_741_io_in_2),
    .io_in_3(c53_741_io_in_3),
    .io_in_4(c53_741_io_in_4),
    .io_out_0(c53_741_io_out_0),
    .io_out_1(c53_741_io_out_1),
    .io_out_2(c53_741_io_out_2)
  );
  C53 c53_742 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_742_io_in_0),
    .io_in_1(c53_742_io_in_1),
    .io_in_2(c53_742_io_in_2),
    .io_in_3(c53_742_io_in_3),
    .io_in_4(c53_742_io_in_4),
    .io_out_0(c53_742_io_out_0),
    .io_out_1(c53_742_io_out_1),
    .io_out_2(c53_742_io_out_2)
  );
  C53 c53_743 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_743_io_in_0),
    .io_in_1(c53_743_io_in_1),
    .io_in_2(c53_743_io_in_2),
    .io_in_3(c53_743_io_in_3),
    .io_in_4(c53_743_io_in_4),
    .io_out_0(c53_743_io_out_0),
    .io_out_1(c53_743_io_out_1),
    .io_out_2(c53_743_io_out_2)
  );
  C53 c53_744 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_744_io_in_0),
    .io_in_1(c53_744_io_in_1),
    .io_in_2(c53_744_io_in_2),
    .io_in_3(c53_744_io_in_3),
    .io_in_4(c53_744_io_in_4),
    .io_out_0(c53_744_io_out_0),
    .io_out_1(c53_744_io_out_1),
    .io_out_2(c53_744_io_out_2)
  );
  C53 c53_745 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_745_io_in_0),
    .io_in_1(c53_745_io_in_1),
    .io_in_2(c53_745_io_in_2),
    .io_in_3(c53_745_io_in_3),
    .io_in_4(c53_745_io_in_4),
    .io_out_0(c53_745_io_out_0),
    .io_out_1(c53_745_io_out_1),
    .io_out_2(c53_745_io_out_2)
  );
  C32 c32_46 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_46_io_in_0),
    .io_in_1(c32_46_io_in_1),
    .io_in_2(c32_46_io_in_2),
    .io_out_0(c32_46_io_out_0),
    .io_out_1(c32_46_io_out_1)
  );
  C53 c53_746 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_746_io_in_0),
    .io_in_1(c53_746_io_in_1),
    .io_in_2(c53_746_io_in_2),
    .io_in_3(c53_746_io_in_3),
    .io_in_4(c53_746_io_in_4),
    .io_out_0(c53_746_io_out_0),
    .io_out_1(c53_746_io_out_1),
    .io_out_2(c53_746_io_out_2)
  );
  C53 c53_747 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_747_io_in_0),
    .io_in_1(c53_747_io_in_1),
    .io_in_2(c53_747_io_in_2),
    .io_in_3(c53_747_io_in_3),
    .io_in_4(c53_747_io_in_4),
    .io_out_0(c53_747_io_out_0),
    .io_out_1(c53_747_io_out_1),
    .io_out_2(c53_747_io_out_2)
  );
  C22 c22_58 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_58_io_in_0),
    .io_in_1(c22_58_io_in_1),
    .io_out_0(c22_58_io_out_0),
    .io_out_1(c22_58_io_out_1)
  );
  C53 c53_748 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_748_io_in_0),
    .io_in_1(c53_748_io_in_1),
    .io_in_2(c53_748_io_in_2),
    .io_in_3(c53_748_io_in_3),
    .io_in_4(c53_748_io_in_4),
    .io_out_0(c53_748_io_out_0),
    .io_out_1(c53_748_io_out_1),
    .io_out_2(c53_748_io_out_2)
  );
  C53 c53_749 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_749_io_in_0),
    .io_in_1(c53_749_io_in_1),
    .io_in_2(c53_749_io_in_2),
    .io_in_3(c53_749_io_in_3),
    .io_in_4(c53_749_io_in_4),
    .io_out_0(c53_749_io_out_0),
    .io_out_1(c53_749_io_out_1),
    .io_out_2(c53_749_io_out_2)
  );
  C22 c22_59 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_59_io_in_0),
    .io_in_1(c22_59_io_in_1),
    .io_out_0(c22_59_io_out_0),
    .io_out_1(c22_59_io_out_1)
  );
  C53 c53_750 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_750_io_in_0),
    .io_in_1(c53_750_io_in_1),
    .io_in_2(c53_750_io_in_2),
    .io_in_3(c53_750_io_in_3),
    .io_in_4(c53_750_io_in_4),
    .io_out_0(c53_750_io_out_0),
    .io_out_1(c53_750_io_out_1),
    .io_out_2(c53_750_io_out_2)
  );
  C53 c53_751 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_751_io_in_0),
    .io_in_1(c53_751_io_in_1),
    .io_in_2(c53_751_io_in_2),
    .io_in_3(c53_751_io_in_3),
    .io_in_4(c53_751_io_in_4),
    .io_out_0(c53_751_io_out_0),
    .io_out_1(c53_751_io_out_1),
    .io_out_2(c53_751_io_out_2)
  );
  C32 c32_47 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_47_io_in_0),
    .io_in_1(c32_47_io_in_1),
    .io_in_2(c32_47_io_in_2),
    .io_out_0(c32_47_io_out_0),
    .io_out_1(c32_47_io_out_1)
  );
  C53 c53_752 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_752_io_in_0),
    .io_in_1(c53_752_io_in_1),
    .io_in_2(c53_752_io_in_2),
    .io_in_3(c53_752_io_in_3),
    .io_in_4(c53_752_io_in_4),
    .io_out_0(c53_752_io_out_0),
    .io_out_1(c53_752_io_out_1),
    .io_out_2(c53_752_io_out_2)
  );
  C53 c53_753 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_753_io_in_0),
    .io_in_1(c53_753_io_in_1),
    .io_in_2(c53_753_io_in_2),
    .io_in_3(c53_753_io_in_3),
    .io_in_4(c53_753_io_in_4),
    .io_out_0(c53_753_io_out_0),
    .io_out_1(c53_753_io_out_1),
    .io_out_2(c53_753_io_out_2)
  );
  C22 c22_60 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_60_io_in_0),
    .io_in_1(c22_60_io_in_1),
    .io_out_0(c22_60_io_out_0),
    .io_out_1(c22_60_io_out_1)
  );
  C53 c53_754 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_754_io_in_0),
    .io_in_1(c53_754_io_in_1),
    .io_in_2(c53_754_io_in_2),
    .io_in_3(c53_754_io_in_3),
    .io_in_4(c53_754_io_in_4),
    .io_out_0(c53_754_io_out_0),
    .io_out_1(c53_754_io_out_1),
    .io_out_2(c53_754_io_out_2)
  );
  C53 c53_755 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_755_io_in_0),
    .io_in_1(c53_755_io_in_1),
    .io_in_2(c53_755_io_in_2),
    .io_in_3(c53_755_io_in_3),
    .io_in_4(c53_755_io_in_4),
    .io_out_0(c53_755_io_out_0),
    .io_out_1(c53_755_io_out_1),
    .io_out_2(c53_755_io_out_2)
  );
  C22 c22_61 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_61_io_in_0),
    .io_in_1(c22_61_io_in_1),
    .io_out_0(c22_61_io_out_0),
    .io_out_1(c22_61_io_out_1)
  );
  C53 c53_756 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_756_io_in_0),
    .io_in_1(c53_756_io_in_1),
    .io_in_2(c53_756_io_in_2),
    .io_in_3(c53_756_io_in_3),
    .io_in_4(c53_756_io_in_4),
    .io_out_0(c53_756_io_out_0),
    .io_out_1(c53_756_io_out_1),
    .io_out_2(c53_756_io_out_2)
  );
  C53 c53_757 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_757_io_in_0),
    .io_in_1(c53_757_io_in_1),
    .io_in_2(c53_757_io_in_2),
    .io_in_3(c53_757_io_in_3),
    .io_in_4(c53_757_io_in_4),
    .io_out_0(c53_757_io_out_0),
    .io_out_1(c53_757_io_out_1),
    .io_out_2(c53_757_io_out_2)
  );
  C22 c22_62 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_62_io_in_0),
    .io_in_1(c22_62_io_in_1),
    .io_out_0(c22_62_io_out_0),
    .io_out_1(c22_62_io_out_1)
  );
  C53 c53_758 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_758_io_in_0),
    .io_in_1(c53_758_io_in_1),
    .io_in_2(c53_758_io_in_2),
    .io_in_3(c53_758_io_in_3),
    .io_in_4(c53_758_io_in_4),
    .io_out_0(c53_758_io_out_0),
    .io_out_1(c53_758_io_out_1),
    .io_out_2(c53_758_io_out_2)
  );
  C53 c53_759 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_759_io_in_0),
    .io_in_1(c53_759_io_in_1),
    .io_in_2(c53_759_io_in_2),
    .io_in_3(c53_759_io_in_3),
    .io_in_4(c53_759_io_in_4),
    .io_out_0(c53_759_io_out_0),
    .io_out_1(c53_759_io_out_1),
    .io_out_2(c53_759_io_out_2)
  );
  C22 c22_63 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_63_io_in_0),
    .io_in_1(c22_63_io_in_1),
    .io_out_0(c22_63_io_out_0),
    .io_out_1(c22_63_io_out_1)
  );
  C53 c53_760 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_760_io_in_0),
    .io_in_1(c53_760_io_in_1),
    .io_in_2(c53_760_io_in_2),
    .io_in_3(c53_760_io_in_3),
    .io_in_4(c53_760_io_in_4),
    .io_out_0(c53_760_io_out_0),
    .io_out_1(c53_760_io_out_1),
    .io_out_2(c53_760_io_out_2)
  );
  C53 c53_761 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_761_io_in_0),
    .io_in_1(c53_761_io_in_1),
    .io_in_2(c53_761_io_in_2),
    .io_in_3(c53_761_io_in_3),
    .io_in_4(c53_761_io_in_4),
    .io_out_0(c53_761_io_out_0),
    .io_out_1(c53_761_io_out_1),
    .io_out_2(c53_761_io_out_2)
  );
  C53 c53_762 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_762_io_in_0),
    .io_in_1(c53_762_io_in_1),
    .io_in_2(c53_762_io_in_2),
    .io_in_3(c53_762_io_in_3),
    .io_in_4(c53_762_io_in_4),
    .io_out_0(c53_762_io_out_0),
    .io_out_1(c53_762_io_out_1),
    .io_out_2(c53_762_io_out_2)
  );
  C53 c53_763 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_763_io_in_0),
    .io_in_1(c53_763_io_in_1),
    .io_in_2(c53_763_io_in_2),
    .io_in_3(c53_763_io_in_3),
    .io_in_4(c53_763_io_in_4),
    .io_out_0(c53_763_io_out_0),
    .io_out_1(c53_763_io_out_1),
    .io_out_2(c53_763_io_out_2)
  );
  C53 c53_764 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_764_io_in_0),
    .io_in_1(c53_764_io_in_1),
    .io_in_2(c53_764_io_in_2),
    .io_in_3(c53_764_io_in_3),
    .io_in_4(c53_764_io_in_4),
    .io_out_0(c53_764_io_out_0),
    .io_out_1(c53_764_io_out_1),
    .io_out_2(c53_764_io_out_2)
  );
  C53 c53_765 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_765_io_in_0),
    .io_in_1(c53_765_io_in_1),
    .io_in_2(c53_765_io_in_2),
    .io_in_3(c53_765_io_in_3),
    .io_in_4(c53_765_io_in_4),
    .io_out_0(c53_765_io_out_0),
    .io_out_1(c53_765_io_out_1),
    .io_out_2(c53_765_io_out_2)
  );
  C53 c53_766 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_766_io_in_0),
    .io_in_1(c53_766_io_in_1),
    .io_in_2(c53_766_io_in_2),
    .io_in_3(c53_766_io_in_3),
    .io_in_4(c53_766_io_in_4),
    .io_out_0(c53_766_io_out_0),
    .io_out_1(c53_766_io_out_1),
    .io_out_2(c53_766_io_out_2)
  );
  C53 c53_767 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_767_io_in_0),
    .io_in_1(c53_767_io_in_1),
    .io_in_2(c53_767_io_in_2),
    .io_in_3(c53_767_io_in_3),
    .io_in_4(c53_767_io_in_4),
    .io_out_0(c53_767_io_out_0),
    .io_out_1(c53_767_io_out_1),
    .io_out_2(c53_767_io_out_2)
  );
  C53 c53_768 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_768_io_in_0),
    .io_in_1(c53_768_io_in_1),
    .io_in_2(c53_768_io_in_2),
    .io_in_3(c53_768_io_in_3),
    .io_in_4(c53_768_io_in_4),
    .io_out_0(c53_768_io_out_0),
    .io_out_1(c53_768_io_out_1),
    .io_out_2(c53_768_io_out_2)
  );
  C53 c53_769 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_769_io_in_0),
    .io_in_1(c53_769_io_in_1),
    .io_in_2(c53_769_io_in_2),
    .io_in_3(c53_769_io_in_3),
    .io_in_4(c53_769_io_in_4),
    .io_out_0(c53_769_io_out_0),
    .io_out_1(c53_769_io_out_1),
    .io_out_2(c53_769_io_out_2)
  );
  C53 c53_770 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_770_io_in_0),
    .io_in_1(c53_770_io_in_1),
    .io_in_2(c53_770_io_in_2),
    .io_in_3(c53_770_io_in_3),
    .io_in_4(c53_770_io_in_4),
    .io_out_0(c53_770_io_out_0),
    .io_out_1(c53_770_io_out_1),
    .io_out_2(c53_770_io_out_2)
  );
  C53 c53_771 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_771_io_in_0),
    .io_in_1(c53_771_io_in_1),
    .io_in_2(c53_771_io_in_2),
    .io_in_3(c53_771_io_in_3),
    .io_in_4(c53_771_io_in_4),
    .io_out_0(c53_771_io_out_0),
    .io_out_1(c53_771_io_out_1),
    .io_out_2(c53_771_io_out_2)
  );
  C53 c53_772 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_772_io_in_0),
    .io_in_1(c53_772_io_in_1),
    .io_in_2(c53_772_io_in_2),
    .io_in_3(c53_772_io_in_3),
    .io_in_4(c53_772_io_in_4),
    .io_out_0(c53_772_io_out_0),
    .io_out_1(c53_772_io_out_1),
    .io_out_2(c53_772_io_out_2)
  );
  C53 c53_773 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_773_io_in_0),
    .io_in_1(c53_773_io_in_1),
    .io_in_2(c53_773_io_in_2),
    .io_in_3(c53_773_io_in_3),
    .io_in_4(c53_773_io_in_4),
    .io_out_0(c53_773_io_out_0),
    .io_out_1(c53_773_io_out_1),
    .io_out_2(c53_773_io_out_2)
  );
  C53 c53_774 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_774_io_in_0),
    .io_in_1(c53_774_io_in_1),
    .io_in_2(c53_774_io_in_2),
    .io_in_3(c53_774_io_in_3),
    .io_in_4(c53_774_io_in_4),
    .io_out_0(c53_774_io_out_0),
    .io_out_1(c53_774_io_out_1),
    .io_out_2(c53_774_io_out_2)
  );
  C53 c53_775 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_775_io_in_0),
    .io_in_1(c53_775_io_in_1),
    .io_in_2(c53_775_io_in_2),
    .io_in_3(c53_775_io_in_3),
    .io_in_4(c53_775_io_in_4),
    .io_out_0(c53_775_io_out_0),
    .io_out_1(c53_775_io_out_1),
    .io_out_2(c53_775_io_out_2)
  );
  C53 c53_776 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_776_io_in_0),
    .io_in_1(c53_776_io_in_1),
    .io_in_2(c53_776_io_in_2),
    .io_in_3(c53_776_io_in_3),
    .io_in_4(c53_776_io_in_4),
    .io_out_0(c53_776_io_out_0),
    .io_out_1(c53_776_io_out_1),
    .io_out_2(c53_776_io_out_2)
  );
  C32 c32_48 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_48_io_in_0),
    .io_in_1(c32_48_io_in_1),
    .io_in_2(c32_48_io_in_2),
    .io_out_0(c32_48_io_out_0),
    .io_out_1(c32_48_io_out_1)
  );
  C53 c53_777 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_777_io_in_0),
    .io_in_1(c53_777_io_in_1),
    .io_in_2(c53_777_io_in_2),
    .io_in_3(c53_777_io_in_3),
    .io_in_4(c53_777_io_in_4),
    .io_out_0(c53_777_io_out_0),
    .io_out_1(c53_777_io_out_1),
    .io_out_2(c53_777_io_out_2)
  );
  C22 c22_64 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_64_io_in_0),
    .io_in_1(c22_64_io_in_1),
    .io_out_0(c22_64_io_out_0),
    .io_out_1(c22_64_io_out_1)
  );
  C53 c53_778 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_778_io_in_0),
    .io_in_1(c53_778_io_in_1),
    .io_in_2(c53_778_io_in_2),
    .io_in_3(c53_778_io_in_3),
    .io_in_4(c53_778_io_in_4),
    .io_out_0(c53_778_io_out_0),
    .io_out_1(c53_778_io_out_1),
    .io_out_2(c53_778_io_out_2)
  );
  C22 c22_65 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_65_io_in_0),
    .io_in_1(c22_65_io_in_1),
    .io_out_0(c22_65_io_out_0),
    .io_out_1(c22_65_io_out_1)
  );
  C53 c53_779 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_779_io_in_0),
    .io_in_1(c53_779_io_in_1),
    .io_in_2(c53_779_io_in_2),
    .io_in_3(c53_779_io_in_3),
    .io_in_4(c53_779_io_in_4),
    .io_out_0(c53_779_io_out_0),
    .io_out_1(c53_779_io_out_1),
    .io_out_2(c53_779_io_out_2)
  );
  C32 c32_49 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_49_io_in_0),
    .io_in_1(c32_49_io_in_1),
    .io_in_2(c32_49_io_in_2),
    .io_out_0(c32_49_io_out_0),
    .io_out_1(c32_49_io_out_1)
  );
  C53 c53_780 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_780_io_in_0),
    .io_in_1(c53_780_io_in_1),
    .io_in_2(c53_780_io_in_2),
    .io_in_3(c53_780_io_in_3),
    .io_in_4(c53_780_io_in_4),
    .io_out_0(c53_780_io_out_0),
    .io_out_1(c53_780_io_out_1),
    .io_out_2(c53_780_io_out_2)
  );
  C22 c22_66 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_66_io_in_0),
    .io_in_1(c22_66_io_in_1),
    .io_out_0(c22_66_io_out_0),
    .io_out_1(c22_66_io_out_1)
  );
  C53 c53_781 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_781_io_in_0),
    .io_in_1(c53_781_io_in_1),
    .io_in_2(c53_781_io_in_2),
    .io_in_3(c53_781_io_in_3),
    .io_in_4(c53_781_io_in_4),
    .io_out_0(c53_781_io_out_0),
    .io_out_1(c53_781_io_out_1),
    .io_out_2(c53_781_io_out_2)
  );
  C22 c22_67 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_67_io_in_0),
    .io_in_1(c22_67_io_in_1),
    .io_out_0(c22_67_io_out_0),
    .io_out_1(c22_67_io_out_1)
  );
  C53 c53_782 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_782_io_in_0),
    .io_in_1(c53_782_io_in_1),
    .io_in_2(c53_782_io_in_2),
    .io_in_3(c53_782_io_in_3),
    .io_in_4(c53_782_io_in_4),
    .io_out_0(c53_782_io_out_0),
    .io_out_1(c53_782_io_out_1),
    .io_out_2(c53_782_io_out_2)
  );
  C22 c22_68 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_68_io_in_0),
    .io_in_1(c22_68_io_in_1),
    .io_out_0(c22_68_io_out_0),
    .io_out_1(c22_68_io_out_1)
  );
  C53 c53_783 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_783_io_in_0),
    .io_in_1(c53_783_io_in_1),
    .io_in_2(c53_783_io_in_2),
    .io_in_3(c53_783_io_in_3),
    .io_in_4(c53_783_io_in_4),
    .io_out_0(c53_783_io_out_0),
    .io_out_1(c53_783_io_out_1),
    .io_out_2(c53_783_io_out_2)
  );
  C22 c22_69 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_69_io_in_0),
    .io_in_1(c22_69_io_in_1),
    .io_out_0(c22_69_io_out_0),
    .io_out_1(c22_69_io_out_1)
  );
  C53 c53_784 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_784_io_in_0),
    .io_in_1(c53_784_io_in_1),
    .io_in_2(c53_784_io_in_2),
    .io_in_3(c53_784_io_in_3),
    .io_in_4(c53_784_io_in_4),
    .io_out_0(c53_784_io_out_0),
    .io_out_1(c53_784_io_out_1),
    .io_out_2(c53_784_io_out_2)
  );
  C53 c53_785 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_785_io_in_0),
    .io_in_1(c53_785_io_in_1),
    .io_in_2(c53_785_io_in_2),
    .io_in_3(c53_785_io_in_3),
    .io_in_4(c53_785_io_in_4),
    .io_out_0(c53_785_io_out_0),
    .io_out_1(c53_785_io_out_1),
    .io_out_2(c53_785_io_out_2)
  );
  C53 c53_786 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_786_io_in_0),
    .io_in_1(c53_786_io_in_1),
    .io_in_2(c53_786_io_in_2),
    .io_in_3(c53_786_io_in_3),
    .io_in_4(c53_786_io_in_4),
    .io_out_0(c53_786_io_out_0),
    .io_out_1(c53_786_io_out_1),
    .io_out_2(c53_786_io_out_2)
  );
  C53 c53_787 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_787_io_in_0),
    .io_in_1(c53_787_io_in_1),
    .io_in_2(c53_787_io_in_2),
    .io_in_3(c53_787_io_in_3),
    .io_in_4(c53_787_io_in_4),
    .io_out_0(c53_787_io_out_0),
    .io_out_1(c53_787_io_out_1),
    .io_out_2(c53_787_io_out_2)
  );
  C53 c53_788 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_788_io_in_0),
    .io_in_1(c53_788_io_in_1),
    .io_in_2(c53_788_io_in_2),
    .io_in_3(c53_788_io_in_3),
    .io_in_4(c53_788_io_in_4),
    .io_out_0(c53_788_io_out_0),
    .io_out_1(c53_788_io_out_1),
    .io_out_2(c53_788_io_out_2)
  );
  C53 c53_789 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_789_io_in_0),
    .io_in_1(c53_789_io_in_1),
    .io_in_2(c53_789_io_in_2),
    .io_in_3(c53_789_io_in_3),
    .io_in_4(c53_789_io_in_4),
    .io_out_0(c53_789_io_out_0),
    .io_out_1(c53_789_io_out_1),
    .io_out_2(c53_789_io_out_2)
  );
  C53 c53_790 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_790_io_in_0),
    .io_in_1(c53_790_io_in_1),
    .io_in_2(c53_790_io_in_2),
    .io_in_3(c53_790_io_in_3),
    .io_in_4(c53_790_io_in_4),
    .io_out_0(c53_790_io_out_0),
    .io_out_1(c53_790_io_out_1),
    .io_out_2(c53_790_io_out_2)
  );
  C53 c53_791 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_791_io_in_0),
    .io_in_1(c53_791_io_in_1),
    .io_in_2(c53_791_io_in_2),
    .io_in_3(c53_791_io_in_3),
    .io_in_4(c53_791_io_in_4),
    .io_out_0(c53_791_io_out_0),
    .io_out_1(c53_791_io_out_1),
    .io_out_2(c53_791_io_out_2)
  );
  C32 c32_50 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_50_io_in_0),
    .io_in_1(c32_50_io_in_1),
    .io_in_2(c32_50_io_in_2),
    .io_out_0(c32_50_io_out_0),
    .io_out_1(c32_50_io_out_1)
  );
  C22 c22_70 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_70_io_in_0),
    .io_in_1(c22_70_io_in_1),
    .io_out_0(c22_70_io_out_0),
    .io_out_1(c22_70_io_out_1)
  );
  C22 c22_71 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_71_io_in_0),
    .io_in_1(c22_71_io_in_1),
    .io_out_0(c22_71_io_out_0),
    .io_out_1(c22_71_io_out_1)
  );
  C32 c32_51 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_51_io_in_0),
    .io_in_1(c32_51_io_in_1),
    .io_in_2(c32_51_io_in_2),
    .io_out_0(c32_51_io_out_0),
    .io_out_1(c32_51_io_out_1)
  );
  C22 c22_72 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_72_io_in_0),
    .io_in_1(c22_72_io_in_1),
    .io_out_0(c22_72_io_out_0),
    .io_out_1(c22_72_io_out_1)
  );
  C22 c22_73 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_73_io_in_0),
    .io_in_1(c22_73_io_in_1),
    .io_out_0(c22_73_io_out_0),
    .io_out_1(c22_73_io_out_1)
  );
  C22 c22_74 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_74_io_in_0),
    .io_in_1(c22_74_io_in_1),
    .io_out_0(c22_74_io_out_0),
    .io_out_1(c22_74_io_out_1)
  );
  C22 c22_75 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_75_io_in_0),
    .io_in_1(c22_75_io_in_1),
    .io_out_0(c22_75_io_out_0),
    .io_out_1(c22_75_io_out_1)
  );
  C22 c22_76 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_76_io_in_0),
    .io_in_1(c22_76_io_in_1),
    .io_out_0(c22_76_io_out_0),
    .io_out_1(c22_76_io_out_1)
  );
  C22 c22_77 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_77_io_in_0),
    .io_in_1(c22_77_io_in_1),
    .io_out_0(c22_77_io_out_0),
    .io_out_1(c22_77_io_out_1)
  );
  C22 c22_78 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_78_io_in_0),
    .io_in_1(c22_78_io_in_1),
    .io_out_0(c22_78_io_out_0),
    .io_out_1(c22_78_io_out_1)
  );
  C22 c22_79 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_79_io_in_0),
    .io_in_1(c22_79_io_in_1),
    .io_out_0(c22_79_io_out_0),
    .io_out_1(c22_79_io_out_1)
  );
  C22 c22_80 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_80_io_in_0),
    .io_in_1(c22_80_io_in_1),
    .io_out_0(c22_80_io_out_0),
    .io_out_1(c22_80_io_out_1)
  );
  C22 c22_81 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_81_io_in_0),
    .io_in_1(c22_81_io_in_1),
    .io_out_0(c22_81_io_out_0),
    .io_out_1(c22_81_io_out_1)
  );
  C22 c22_82 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_82_io_in_0),
    .io_in_1(c22_82_io_in_1),
    .io_out_0(c22_82_io_out_0),
    .io_out_1(c22_82_io_out_1)
  );
  C22 c22_83 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_83_io_in_0),
    .io_in_1(c22_83_io_in_1),
    .io_out_0(c22_83_io_out_0),
    .io_out_1(c22_83_io_out_1)
  );
  C22 c22_84 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_84_io_in_0),
    .io_in_1(c22_84_io_in_1),
    .io_out_0(c22_84_io_out_0),
    .io_out_1(c22_84_io_out_1)
  );
  C22 c22_85 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_85_io_in_0),
    .io_in_1(c22_85_io_in_1),
    .io_out_0(c22_85_io_out_0),
    .io_out_1(c22_85_io_out_1)
  );
  C22 c22_86 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_86_io_in_0),
    .io_in_1(c22_86_io_in_1),
    .io_out_0(c22_86_io_out_0),
    .io_out_1(c22_86_io_out_1)
  );
  C32 c32_52 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_52_io_in_0),
    .io_in_1(c32_52_io_in_1),
    .io_in_2(c32_52_io_in_2),
    .io_out_0(c32_52_io_out_0),
    .io_out_1(c32_52_io_out_1)
  );
  C32 c32_53 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_53_io_in_0),
    .io_in_1(c32_53_io_in_1),
    .io_in_2(c32_53_io_in_2),
    .io_out_0(c32_53_io_out_0),
    .io_out_1(c32_53_io_out_1)
  );
  C32 c32_54 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_54_io_in_0),
    .io_in_1(c32_54_io_in_1),
    .io_in_2(c32_54_io_in_2),
    .io_out_0(c32_54_io_out_0),
    .io_out_1(c32_54_io_out_1)
  );
  C32 c32_55 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_55_io_in_0),
    .io_in_1(c32_55_io_in_1),
    .io_in_2(c32_55_io_in_2),
    .io_out_0(c32_55_io_out_0),
    .io_out_1(c32_55_io_out_1)
  );
  C53 c53_792 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_792_io_in_0),
    .io_in_1(c53_792_io_in_1),
    .io_in_2(c53_792_io_in_2),
    .io_in_3(c53_792_io_in_3),
    .io_in_4(c53_792_io_in_4),
    .io_out_0(c53_792_io_out_0),
    .io_out_1(c53_792_io_out_1),
    .io_out_2(c53_792_io_out_2)
  );
  C53 c53_793 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_793_io_in_0),
    .io_in_1(c53_793_io_in_1),
    .io_in_2(c53_793_io_in_2),
    .io_in_3(c53_793_io_in_3),
    .io_in_4(c53_793_io_in_4),
    .io_out_0(c53_793_io_out_0),
    .io_out_1(c53_793_io_out_1),
    .io_out_2(c53_793_io_out_2)
  );
  C53 c53_794 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_794_io_in_0),
    .io_in_1(c53_794_io_in_1),
    .io_in_2(c53_794_io_in_2),
    .io_in_3(c53_794_io_in_3),
    .io_in_4(c53_794_io_in_4),
    .io_out_0(c53_794_io_out_0),
    .io_out_1(c53_794_io_out_1),
    .io_out_2(c53_794_io_out_2)
  );
  C53 c53_795 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_795_io_in_0),
    .io_in_1(c53_795_io_in_1),
    .io_in_2(c53_795_io_in_2),
    .io_in_3(c53_795_io_in_3),
    .io_in_4(c53_795_io_in_4),
    .io_out_0(c53_795_io_out_0),
    .io_out_1(c53_795_io_out_1),
    .io_out_2(c53_795_io_out_2)
  );
  C53 c53_796 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_796_io_in_0),
    .io_in_1(c53_796_io_in_1),
    .io_in_2(c53_796_io_in_2),
    .io_in_3(c53_796_io_in_3),
    .io_in_4(c53_796_io_in_4),
    .io_out_0(c53_796_io_out_0),
    .io_out_1(c53_796_io_out_1),
    .io_out_2(c53_796_io_out_2)
  );
  C53 c53_797 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_797_io_in_0),
    .io_in_1(c53_797_io_in_1),
    .io_in_2(c53_797_io_in_2),
    .io_in_3(c53_797_io_in_3),
    .io_in_4(c53_797_io_in_4),
    .io_out_0(c53_797_io_out_0),
    .io_out_1(c53_797_io_out_1),
    .io_out_2(c53_797_io_out_2)
  );
  C53 c53_798 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_798_io_in_0),
    .io_in_1(c53_798_io_in_1),
    .io_in_2(c53_798_io_in_2),
    .io_in_3(c53_798_io_in_3),
    .io_in_4(c53_798_io_in_4),
    .io_out_0(c53_798_io_out_0),
    .io_out_1(c53_798_io_out_1),
    .io_out_2(c53_798_io_out_2)
  );
  C53 c53_799 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_799_io_in_0),
    .io_in_1(c53_799_io_in_1),
    .io_in_2(c53_799_io_in_2),
    .io_in_3(c53_799_io_in_3),
    .io_in_4(c53_799_io_in_4),
    .io_out_0(c53_799_io_out_0),
    .io_out_1(c53_799_io_out_1),
    .io_out_2(c53_799_io_out_2)
  );
  C53 c53_800 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_800_io_in_0),
    .io_in_1(c53_800_io_in_1),
    .io_in_2(c53_800_io_in_2),
    .io_in_3(c53_800_io_in_3),
    .io_in_4(c53_800_io_in_4),
    .io_out_0(c53_800_io_out_0),
    .io_out_1(c53_800_io_out_1),
    .io_out_2(c53_800_io_out_2)
  );
  C53 c53_801 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_801_io_in_0),
    .io_in_1(c53_801_io_in_1),
    .io_in_2(c53_801_io_in_2),
    .io_in_3(c53_801_io_in_3),
    .io_in_4(c53_801_io_in_4),
    .io_out_0(c53_801_io_out_0),
    .io_out_1(c53_801_io_out_1),
    .io_out_2(c53_801_io_out_2)
  );
  C53 c53_802 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_802_io_in_0),
    .io_in_1(c53_802_io_in_1),
    .io_in_2(c53_802_io_in_2),
    .io_in_3(c53_802_io_in_3),
    .io_in_4(c53_802_io_in_4),
    .io_out_0(c53_802_io_out_0),
    .io_out_1(c53_802_io_out_1),
    .io_out_2(c53_802_io_out_2)
  );
  C53 c53_803 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_803_io_in_0),
    .io_in_1(c53_803_io_in_1),
    .io_in_2(c53_803_io_in_2),
    .io_in_3(c53_803_io_in_3),
    .io_in_4(c53_803_io_in_4),
    .io_out_0(c53_803_io_out_0),
    .io_out_1(c53_803_io_out_1),
    .io_out_2(c53_803_io_out_2)
  );
  C53 c53_804 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_804_io_in_0),
    .io_in_1(c53_804_io_in_1),
    .io_in_2(c53_804_io_in_2),
    .io_in_3(c53_804_io_in_3),
    .io_in_4(c53_804_io_in_4),
    .io_out_0(c53_804_io_out_0),
    .io_out_1(c53_804_io_out_1),
    .io_out_2(c53_804_io_out_2)
  );
  C53 c53_805 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_805_io_in_0),
    .io_in_1(c53_805_io_in_1),
    .io_in_2(c53_805_io_in_2),
    .io_in_3(c53_805_io_in_3),
    .io_in_4(c53_805_io_in_4),
    .io_out_0(c53_805_io_out_0),
    .io_out_1(c53_805_io_out_1),
    .io_out_2(c53_805_io_out_2)
  );
  C53 c53_806 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_806_io_in_0),
    .io_in_1(c53_806_io_in_1),
    .io_in_2(c53_806_io_in_2),
    .io_in_3(c53_806_io_in_3),
    .io_in_4(c53_806_io_in_4),
    .io_out_0(c53_806_io_out_0),
    .io_out_1(c53_806_io_out_1),
    .io_out_2(c53_806_io_out_2)
  );
  C53 c53_807 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_807_io_in_0),
    .io_in_1(c53_807_io_in_1),
    .io_in_2(c53_807_io_in_2),
    .io_in_3(c53_807_io_in_3),
    .io_in_4(c53_807_io_in_4),
    .io_out_0(c53_807_io_out_0),
    .io_out_1(c53_807_io_out_1),
    .io_out_2(c53_807_io_out_2)
  );
  C53 c53_808 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_808_io_in_0),
    .io_in_1(c53_808_io_in_1),
    .io_in_2(c53_808_io_in_2),
    .io_in_3(c53_808_io_in_3),
    .io_in_4(c53_808_io_in_4),
    .io_out_0(c53_808_io_out_0),
    .io_out_1(c53_808_io_out_1),
    .io_out_2(c53_808_io_out_2)
  );
  C22 c22_87 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_87_io_in_0),
    .io_in_1(c22_87_io_in_1),
    .io_out_0(c22_87_io_out_0),
    .io_out_1(c22_87_io_out_1)
  );
  C53 c53_809 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_809_io_in_0),
    .io_in_1(c53_809_io_in_1),
    .io_in_2(c53_809_io_in_2),
    .io_in_3(c53_809_io_in_3),
    .io_in_4(c53_809_io_in_4),
    .io_out_0(c53_809_io_out_0),
    .io_out_1(c53_809_io_out_1),
    .io_out_2(c53_809_io_out_2)
  );
  C22 c22_88 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_88_io_in_0),
    .io_in_1(c22_88_io_in_1),
    .io_out_0(c22_88_io_out_0),
    .io_out_1(c22_88_io_out_1)
  );
  C53 c53_810 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_810_io_in_0),
    .io_in_1(c53_810_io_in_1),
    .io_in_2(c53_810_io_in_2),
    .io_in_3(c53_810_io_in_3),
    .io_in_4(c53_810_io_in_4),
    .io_out_0(c53_810_io_out_0),
    .io_out_1(c53_810_io_out_1),
    .io_out_2(c53_810_io_out_2)
  );
  C22 c22_89 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_89_io_in_0),
    .io_in_1(c22_89_io_in_1),
    .io_out_0(c22_89_io_out_0),
    .io_out_1(c22_89_io_out_1)
  );
  C53 c53_811 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_811_io_in_0),
    .io_in_1(c53_811_io_in_1),
    .io_in_2(c53_811_io_in_2),
    .io_in_3(c53_811_io_in_3),
    .io_in_4(c53_811_io_in_4),
    .io_out_0(c53_811_io_out_0),
    .io_out_1(c53_811_io_out_1),
    .io_out_2(c53_811_io_out_2)
  );
  C22 c22_90 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_90_io_in_0),
    .io_in_1(c22_90_io_in_1),
    .io_out_0(c22_90_io_out_0),
    .io_out_1(c22_90_io_out_1)
  );
  C53 c53_812 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_812_io_in_0),
    .io_in_1(c53_812_io_in_1),
    .io_in_2(c53_812_io_in_2),
    .io_in_3(c53_812_io_in_3),
    .io_in_4(c53_812_io_in_4),
    .io_out_0(c53_812_io_out_0),
    .io_out_1(c53_812_io_out_1),
    .io_out_2(c53_812_io_out_2)
  );
  C22 c22_91 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_91_io_in_0),
    .io_in_1(c22_91_io_in_1),
    .io_out_0(c22_91_io_out_0),
    .io_out_1(c22_91_io_out_1)
  );
  C53 c53_813 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_813_io_in_0),
    .io_in_1(c53_813_io_in_1),
    .io_in_2(c53_813_io_in_2),
    .io_in_3(c53_813_io_in_3),
    .io_in_4(c53_813_io_in_4),
    .io_out_0(c53_813_io_out_0),
    .io_out_1(c53_813_io_out_1),
    .io_out_2(c53_813_io_out_2)
  );
  C22 c22_92 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_92_io_in_0),
    .io_in_1(c22_92_io_in_1),
    .io_out_0(c22_92_io_out_0),
    .io_out_1(c22_92_io_out_1)
  );
  C53 c53_814 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_814_io_in_0),
    .io_in_1(c53_814_io_in_1),
    .io_in_2(c53_814_io_in_2),
    .io_in_3(c53_814_io_in_3),
    .io_in_4(c53_814_io_in_4),
    .io_out_0(c53_814_io_out_0),
    .io_out_1(c53_814_io_out_1),
    .io_out_2(c53_814_io_out_2)
  );
  C22 c22_93 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_93_io_in_0),
    .io_in_1(c22_93_io_in_1),
    .io_out_0(c22_93_io_out_0),
    .io_out_1(c22_93_io_out_1)
  );
  C53 c53_815 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_815_io_in_0),
    .io_in_1(c53_815_io_in_1),
    .io_in_2(c53_815_io_in_2),
    .io_in_3(c53_815_io_in_3),
    .io_in_4(c53_815_io_in_4),
    .io_out_0(c53_815_io_out_0),
    .io_out_1(c53_815_io_out_1),
    .io_out_2(c53_815_io_out_2)
  );
  C22 c22_94 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_94_io_in_0),
    .io_in_1(c22_94_io_in_1),
    .io_out_0(c22_94_io_out_0),
    .io_out_1(c22_94_io_out_1)
  );
  C53 c53_816 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_816_io_in_0),
    .io_in_1(c53_816_io_in_1),
    .io_in_2(c53_816_io_in_2),
    .io_in_3(c53_816_io_in_3),
    .io_in_4(c53_816_io_in_4),
    .io_out_0(c53_816_io_out_0),
    .io_out_1(c53_816_io_out_1),
    .io_out_2(c53_816_io_out_2)
  );
  C22 c22_95 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_95_io_in_0),
    .io_in_1(c22_95_io_in_1),
    .io_out_0(c22_95_io_out_0),
    .io_out_1(c22_95_io_out_1)
  );
  C53 c53_817 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_817_io_in_0),
    .io_in_1(c53_817_io_in_1),
    .io_in_2(c53_817_io_in_2),
    .io_in_3(c53_817_io_in_3),
    .io_in_4(c53_817_io_in_4),
    .io_out_0(c53_817_io_out_0),
    .io_out_1(c53_817_io_out_1),
    .io_out_2(c53_817_io_out_2)
  );
  C22 c22_96 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_96_io_in_0),
    .io_in_1(c22_96_io_in_1),
    .io_out_0(c22_96_io_out_0),
    .io_out_1(c22_96_io_out_1)
  );
  C53 c53_818 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_818_io_in_0),
    .io_in_1(c53_818_io_in_1),
    .io_in_2(c53_818_io_in_2),
    .io_in_3(c53_818_io_in_3),
    .io_in_4(c53_818_io_in_4),
    .io_out_0(c53_818_io_out_0),
    .io_out_1(c53_818_io_out_1),
    .io_out_2(c53_818_io_out_2)
  );
  C22 c22_97 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_97_io_in_0),
    .io_in_1(c22_97_io_in_1),
    .io_out_0(c22_97_io_out_0),
    .io_out_1(c22_97_io_out_1)
  );
  C53 c53_819 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_819_io_in_0),
    .io_in_1(c53_819_io_in_1),
    .io_in_2(c53_819_io_in_2),
    .io_in_3(c53_819_io_in_3),
    .io_in_4(c53_819_io_in_4),
    .io_out_0(c53_819_io_out_0),
    .io_out_1(c53_819_io_out_1),
    .io_out_2(c53_819_io_out_2)
  );
  C22 c22_98 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_98_io_in_0),
    .io_in_1(c22_98_io_in_1),
    .io_out_0(c22_98_io_out_0),
    .io_out_1(c22_98_io_out_1)
  );
  C53 c53_820 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_820_io_in_0),
    .io_in_1(c53_820_io_in_1),
    .io_in_2(c53_820_io_in_2),
    .io_in_3(c53_820_io_in_3),
    .io_in_4(c53_820_io_in_4),
    .io_out_0(c53_820_io_out_0),
    .io_out_1(c53_820_io_out_1),
    .io_out_2(c53_820_io_out_2)
  );
  C32 c32_56 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_56_io_in_0),
    .io_in_1(c32_56_io_in_1),
    .io_in_2(c32_56_io_in_2),
    .io_out_0(c32_56_io_out_0),
    .io_out_1(c32_56_io_out_1)
  );
  C53 c53_821 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_821_io_in_0),
    .io_in_1(c53_821_io_in_1),
    .io_in_2(c53_821_io_in_2),
    .io_in_3(c53_821_io_in_3),
    .io_in_4(c53_821_io_in_4),
    .io_out_0(c53_821_io_out_0),
    .io_out_1(c53_821_io_out_1),
    .io_out_2(c53_821_io_out_2)
  );
  C32 c32_57 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_57_io_in_0),
    .io_in_1(c32_57_io_in_1),
    .io_in_2(c32_57_io_in_2),
    .io_out_0(c32_57_io_out_0),
    .io_out_1(c32_57_io_out_1)
  );
  C53 c53_822 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_822_io_in_0),
    .io_in_1(c53_822_io_in_1),
    .io_in_2(c53_822_io_in_2),
    .io_in_3(c53_822_io_in_3),
    .io_in_4(c53_822_io_in_4),
    .io_out_0(c53_822_io_out_0),
    .io_out_1(c53_822_io_out_1),
    .io_out_2(c53_822_io_out_2)
  );
  C32 c32_58 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_58_io_in_0),
    .io_in_1(c32_58_io_in_1),
    .io_in_2(c32_58_io_in_2),
    .io_out_0(c32_58_io_out_0),
    .io_out_1(c32_58_io_out_1)
  );
  C53 c53_823 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_823_io_in_0),
    .io_in_1(c53_823_io_in_1),
    .io_in_2(c53_823_io_in_2),
    .io_in_3(c53_823_io_in_3),
    .io_in_4(c53_823_io_in_4),
    .io_out_0(c53_823_io_out_0),
    .io_out_1(c53_823_io_out_1),
    .io_out_2(c53_823_io_out_2)
  );
  C32 c32_59 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_59_io_in_0),
    .io_in_1(c32_59_io_in_1),
    .io_in_2(c32_59_io_in_2),
    .io_out_0(c32_59_io_out_0),
    .io_out_1(c32_59_io_out_1)
  );
  C53 c53_824 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_824_io_in_0),
    .io_in_1(c53_824_io_in_1),
    .io_in_2(c53_824_io_in_2),
    .io_in_3(c53_824_io_in_3),
    .io_in_4(c53_824_io_in_4),
    .io_out_0(c53_824_io_out_0),
    .io_out_1(c53_824_io_out_1),
    .io_out_2(c53_824_io_out_2)
  );
  C53 c53_825 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_825_io_in_0),
    .io_in_1(c53_825_io_in_1),
    .io_in_2(c53_825_io_in_2),
    .io_in_3(c53_825_io_in_3),
    .io_in_4(c53_825_io_in_4),
    .io_out_0(c53_825_io_out_0),
    .io_out_1(c53_825_io_out_1),
    .io_out_2(c53_825_io_out_2)
  );
  C53 c53_826 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_826_io_in_0),
    .io_in_1(c53_826_io_in_1),
    .io_in_2(c53_826_io_in_2),
    .io_in_3(c53_826_io_in_3),
    .io_in_4(c53_826_io_in_4),
    .io_out_0(c53_826_io_out_0),
    .io_out_1(c53_826_io_out_1),
    .io_out_2(c53_826_io_out_2)
  );
  C53 c53_827 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_827_io_in_0),
    .io_in_1(c53_827_io_in_1),
    .io_in_2(c53_827_io_in_2),
    .io_in_3(c53_827_io_in_3),
    .io_in_4(c53_827_io_in_4),
    .io_out_0(c53_827_io_out_0),
    .io_out_1(c53_827_io_out_1),
    .io_out_2(c53_827_io_out_2)
  );
  C53 c53_828 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_828_io_in_0),
    .io_in_1(c53_828_io_in_1),
    .io_in_2(c53_828_io_in_2),
    .io_in_3(c53_828_io_in_3),
    .io_in_4(c53_828_io_in_4),
    .io_out_0(c53_828_io_out_0),
    .io_out_1(c53_828_io_out_1),
    .io_out_2(c53_828_io_out_2)
  );
  C53 c53_829 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_829_io_in_0),
    .io_in_1(c53_829_io_in_1),
    .io_in_2(c53_829_io_in_2),
    .io_in_3(c53_829_io_in_3),
    .io_in_4(c53_829_io_in_4),
    .io_out_0(c53_829_io_out_0),
    .io_out_1(c53_829_io_out_1),
    .io_out_2(c53_829_io_out_2)
  );
  C53 c53_830 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_830_io_in_0),
    .io_in_1(c53_830_io_in_1),
    .io_in_2(c53_830_io_in_2),
    .io_in_3(c53_830_io_in_3),
    .io_in_4(c53_830_io_in_4),
    .io_out_0(c53_830_io_out_0),
    .io_out_1(c53_830_io_out_1),
    .io_out_2(c53_830_io_out_2)
  );
  C53 c53_831 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_831_io_in_0),
    .io_in_1(c53_831_io_in_1),
    .io_in_2(c53_831_io_in_2),
    .io_in_3(c53_831_io_in_3),
    .io_in_4(c53_831_io_in_4),
    .io_out_0(c53_831_io_out_0),
    .io_out_1(c53_831_io_out_1),
    .io_out_2(c53_831_io_out_2)
  );
  C53 c53_832 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_832_io_in_0),
    .io_in_1(c53_832_io_in_1),
    .io_in_2(c53_832_io_in_2),
    .io_in_3(c53_832_io_in_3),
    .io_in_4(c53_832_io_in_4),
    .io_out_0(c53_832_io_out_0),
    .io_out_1(c53_832_io_out_1),
    .io_out_2(c53_832_io_out_2)
  );
  C53 c53_833 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_833_io_in_0),
    .io_in_1(c53_833_io_in_1),
    .io_in_2(c53_833_io_in_2),
    .io_in_3(c53_833_io_in_3),
    .io_in_4(c53_833_io_in_4),
    .io_out_0(c53_833_io_out_0),
    .io_out_1(c53_833_io_out_1),
    .io_out_2(c53_833_io_out_2)
  );
  C53 c53_834 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_834_io_in_0),
    .io_in_1(c53_834_io_in_1),
    .io_in_2(c53_834_io_in_2),
    .io_in_3(c53_834_io_in_3),
    .io_in_4(c53_834_io_in_4),
    .io_out_0(c53_834_io_out_0),
    .io_out_1(c53_834_io_out_1),
    .io_out_2(c53_834_io_out_2)
  );
  C53 c53_835 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_835_io_in_0),
    .io_in_1(c53_835_io_in_1),
    .io_in_2(c53_835_io_in_2),
    .io_in_3(c53_835_io_in_3),
    .io_in_4(c53_835_io_in_4),
    .io_out_0(c53_835_io_out_0),
    .io_out_1(c53_835_io_out_1),
    .io_out_2(c53_835_io_out_2)
  );
  C53 c53_836 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_836_io_in_0),
    .io_in_1(c53_836_io_in_1),
    .io_in_2(c53_836_io_in_2),
    .io_in_3(c53_836_io_in_3),
    .io_in_4(c53_836_io_in_4),
    .io_out_0(c53_836_io_out_0),
    .io_out_1(c53_836_io_out_1),
    .io_out_2(c53_836_io_out_2)
  );
  C53 c53_837 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_837_io_in_0),
    .io_in_1(c53_837_io_in_1),
    .io_in_2(c53_837_io_in_2),
    .io_in_3(c53_837_io_in_3),
    .io_in_4(c53_837_io_in_4),
    .io_out_0(c53_837_io_out_0),
    .io_out_1(c53_837_io_out_1),
    .io_out_2(c53_837_io_out_2)
  );
  C53 c53_838 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_838_io_in_0),
    .io_in_1(c53_838_io_in_1),
    .io_in_2(c53_838_io_in_2),
    .io_in_3(c53_838_io_in_3),
    .io_in_4(c53_838_io_in_4),
    .io_out_0(c53_838_io_out_0),
    .io_out_1(c53_838_io_out_1),
    .io_out_2(c53_838_io_out_2)
  );
  C53 c53_839 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_839_io_in_0),
    .io_in_1(c53_839_io_in_1),
    .io_in_2(c53_839_io_in_2),
    .io_in_3(c53_839_io_in_3),
    .io_in_4(c53_839_io_in_4),
    .io_out_0(c53_839_io_out_0),
    .io_out_1(c53_839_io_out_1),
    .io_out_2(c53_839_io_out_2)
  );
  C53 c53_840 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_840_io_in_0),
    .io_in_1(c53_840_io_in_1),
    .io_in_2(c53_840_io_in_2),
    .io_in_3(c53_840_io_in_3),
    .io_in_4(c53_840_io_in_4),
    .io_out_0(c53_840_io_out_0),
    .io_out_1(c53_840_io_out_1),
    .io_out_2(c53_840_io_out_2)
  );
  C53 c53_841 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_841_io_in_0),
    .io_in_1(c53_841_io_in_1),
    .io_in_2(c53_841_io_in_2),
    .io_in_3(c53_841_io_in_3),
    .io_in_4(c53_841_io_in_4),
    .io_out_0(c53_841_io_out_0),
    .io_out_1(c53_841_io_out_1),
    .io_out_2(c53_841_io_out_2)
  );
  C53 c53_842 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_842_io_in_0),
    .io_in_1(c53_842_io_in_1),
    .io_in_2(c53_842_io_in_2),
    .io_in_3(c53_842_io_in_3),
    .io_in_4(c53_842_io_in_4),
    .io_out_0(c53_842_io_out_0),
    .io_out_1(c53_842_io_out_1),
    .io_out_2(c53_842_io_out_2)
  );
  C53 c53_843 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_843_io_in_0),
    .io_in_1(c53_843_io_in_1),
    .io_in_2(c53_843_io_in_2),
    .io_in_3(c53_843_io_in_3),
    .io_in_4(c53_843_io_in_4),
    .io_out_0(c53_843_io_out_0),
    .io_out_1(c53_843_io_out_1),
    .io_out_2(c53_843_io_out_2)
  );
  C53 c53_844 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_844_io_in_0),
    .io_in_1(c53_844_io_in_1),
    .io_in_2(c53_844_io_in_2),
    .io_in_3(c53_844_io_in_3),
    .io_in_4(c53_844_io_in_4),
    .io_out_0(c53_844_io_out_0),
    .io_out_1(c53_844_io_out_1),
    .io_out_2(c53_844_io_out_2)
  );
  C53 c53_845 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_845_io_in_0),
    .io_in_1(c53_845_io_in_1),
    .io_in_2(c53_845_io_in_2),
    .io_in_3(c53_845_io_in_3),
    .io_in_4(c53_845_io_in_4),
    .io_out_0(c53_845_io_out_0),
    .io_out_1(c53_845_io_out_1),
    .io_out_2(c53_845_io_out_2)
  );
  C53 c53_846 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_846_io_in_0),
    .io_in_1(c53_846_io_in_1),
    .io_in_2(c53_846_io_in_2),
    .io_in_3(c53_846_io_in_3),
    .io_in_4(c53_846_io_in_4),
    .io_out_0(c53_846_io_out_0),
    .io_out_1(c53_846_io_out_1),
    .io_out_2(c53_846_io_out_2)
  );
  C53 c53_847 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_847_io_in_0),
    .io_in_1(c53_847_io_in_1),
    .io_in_2(c53_847_io_in_2),
    .io_in_3(c53_847_io_in_3),
    .io_in_4(c53_847_io_in_4),
    .io_out_0(c53_847_io_out_0),
    .io_out_1(c53_847_io_out_1),
    .io_out_2(c53_847_io_out_2)
  );
  C53 c53_848 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_848_io_in_0),
    .io_in_1(c53_848_io_in_1),
    .io_in_2(c53_848_io_in_2),
    .io_in_3(c53_848_io_in_3),
    .io_in_4(c53_848_io_in_4),
    .io_out_0(c53_848_io_out_0),
    .io_out_1(c53_848_io_out_1),
    .io_out_2(c53_848_io_out_2)
  );
  C53 c53_849 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_849_io_in_0),
    .io_in_1(c53_849_io_in_1),
    .io_in_2(c53_849_io_in_2),
    .io_in_3(c53_849_io_in_3),
    .io_in_4(c53_849_io_in_4),
    .io_out_0(c53_849_io_out_0),
    .io_out_1(c53_849_io_out_1),
    .io_out_2(c53_849_io_out_2)
  );
  C53 c53_850 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_850_io_in_0),
    .io_in_1(c53_850_io_in_1),
    .io_in_2(c53_850_io_in_2),
    .io_in_3(c53_850_io_in_3),
    .io_in_4(c53_850_io_in_4),
    .io_out_0(c53_850_io_out_0),
    .io_out_1(c53_850_io_out_1),
    .io_out_2(c53_850_io_out_2)
  );
  C53 c53_851 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_851_io_in_0),
    .io_in_1(c53_851_io_in_1),
    .io_in_2(c53_851_io_in_2),
    .io_in_3(c53_851_io_in_3),
    .io_in_4(c53_851_io_in_4),
    .io_out_0(c53_851_io_out_0),
    .io_out_1(c53_851_io_out_1),
    .io_out_2(c53_851_io_out_2)
  );
  C53 c53_852 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_852_io_in_0),
    .io_in_1(c53_852_io_in_1),
    .io_in_2(c53_852_io_in_2),
    .io_in_3(c53_852_io_in_3),
    .io_in_4(c53_852_io_in_4),
    .io_out_0(c53_852_io_out_0),
    .io_out_1(c53_852_io_out_1),
    .io_out_2(c53_852_io_out_2)
  );
  C53 c53_853 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_853_io_in_0),
    .io_in_1(c53_853_io_in_1),
    .io_in_2(c53_853_io_in_2),
    .io_in_3(c53_853_io_in_3),
    .io_in_4(c53_853_io_in_4),
    .io_out_0(c53_853_io_out_0),
    .io_out_1(c53_853_io_out_1),
    .io_out_2(c53_853_io_out_2)
  );
  C53 c53_854 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_854_io_in_0),
    .io_in_1(c53_854_io_in_1),
    .io_in_2(c53_854_io_in_2),
    .io_in_3(c53_854_io_in_3),
    .io_in_4(c53_854_io_in_4),
    .io_out_0(c53_854_io_out_0),
    .io_out_1(c53_854_io_out_1),
    .io_out_2(c53_854_io_out_2)
  );
  C53 c53_855 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_855_io_in_0),
    .io_in_1(c53_855_io_in_1),
    .io_in_2(c53_855_io_in_2),
    .io_in_3(c53_855_io_in_3),
    .io_in_4(c53_855_io_in_4),
    .io_out_0(c53_855_io_out_0),
    .io_out_1(c53_855_io_out_1),
    .io_out_2(c53_855_io_out_2)
  );
  C53 c53_856 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_856_io_in_0),
    .io_in_1(c53_856_io_in_1),
    .io_in_2(c53_856_io_in_2),
    .io_in_3(c53_856_io_in_3),
    .io_in_4(c53_856_io_in_4),
    .io_out_0(c53_856_io_out_0),
    .io_out_1(c53_856_io_out_1),
    .io_out_2(c53_856_io_out_2)
  );
  C53 c53_857 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_857_io_in_0),
    .io_in_1(c53_857_io_in_1),
    .io_in_2(c53_857_io_in_2),
    .io_in_3(c53_857_io_in_3),
    .io_in_4(c53_857_io_in_4),
    .io_out_0(c53_857_io_out_0),
    .io_out_1(c53_857_io_out_1),
    .io_out_2(c53_857_io_out_2)
  );
  C53 c53_858 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_858_io_in_0),
    .io_in_1(c53_858_io_in_1),
    .io_in_2(c53_858_io_in_2),
    .io_in_3(c53_858_io_in_3),
    .io_in_4(c53_858_io_in_4),
    .io_out_0(c53_858_io_out_0),
    .io_out_1(c53_858_io_out_1),
    .io_out_2(c53_858_io_out_2)
  );
  C53 c53_859 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_859_io_in_0),
    .io_in_1(c53_859_io_in_1),
    .io_in_2(c53_859_io_in_2),
    .io_in_3(c53_859_io_in_3),
    .io_in_4(c53_859_io_in_4),
    .io_out_0(c53_859_io_out_0),
    .io_out_1(c53_859_io_out_1),
    .io_out_2(c53_859_io_out_2)
  );
  C53 c53_860 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_860_io_in_0),
    .io_in_1(c53_860_io_in_1),
    .io_in_2(c53_860_io_in_2),
    .io_in_3(c53_860_io_in_3),
    .io_in_4(c53_860_io_in_4),
    .io_out_0(c53_860_io_out_0),
    .io_out_1(c53_860_io_out_1),
    .io_out_2(c53_860_io_out_2)
  );
  C53 c53_861 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_861_io_in_0),
    .io_in_1(c53_861_io_in_1),
    .io_in_2(c53_861_io_in_2),
    .io_in_3(c53_861_io_in_3),
    .io_in_4(c53_861_io_in_4),
    .io_out_0(c53_861_io_out_0),
    .io_out_1(c53_861_io_out_1),
    .io_out_2(c53_861_io_out_2)
  );
  C53 c53_862 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_862_io_in_0),
    .io_in_1(c53_862_io_in_1),
    .io_in_2(c53_862_io_in_2),
    .io_in_3(c53_862_io_in_3),
    .io_in_4(c53_862_io_in_4),
    .io_out_0(c53_862_io_out_0),
    .io_out_1(c53_862_io_out_1),
    .io_out_2(c53_862_io_out_2)
  );
  C53 c53_863 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_863_io_in_0),
    .io_in_1(c53_863_io_in_1),
    .io_in_2(c53_863_io_in_2),
    .io_in_3(c53_863_io_in_3),
    .io_in_4(c53_863_io_in_4),
    .io_out_0(c53_863_io_out_0),
    .io_out_1(c53_863_io_out_1),
    .io_out_2(c53_863_io_out_2)
  );
  C53 c53_864 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_864_io_in_0),
    .io_in_1(c53_864_io_in_1),
    .io_in_2(c53_864_io_in_2),
    .io_in_3(c53_864_io_in_3),
    .io_in_4(c53_864_io_in_4),
    .io_out_0(c53_864_io_out_0),
    .io_out_1(c53_864_io_out_1),
    .io_out_2(c53_864_io_out_2)
  );
  C53 c53_865 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_865_io_in_0),
    .io_in_1(c53_865_io_in_1),
    .io_in_2(c53_865_io_in_2),
    .io_in_3(c53_865_io_in_3),
    .io_in_4(c53_865_io_in_4),
    .io_out_0(c53_865_io_out_0),
    .io_out_1(c53_865_io_out_1),
    .io_out_2(c53_865_io_out_2)
  );
  C53 c53_866 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_866_io_in_0),
    .io_in_1(c53_866_io_in_1),
    .io_in_2(c53_866_io_in_2),
    .io_in_3(c53_866_io_in_3),
    .io_in_4(c53_866_io_in_4),
    .io_out_0(c53_866_io_out_0),
    .io_out_1(c53_866_io_out_1),
    .io_out_2(c53_866_io_out_2)
  );
  C53 c53_867 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_867_io_in_0),
    .io_in_1(c53_867_io_in_1),
    .io_in_2(c53_867_io_in_2),
    .io_in_3(c53_867_io_in_3),
    .io_in_4(c53_867_io_in_4),
    .io_out_0(c53_867_io_out_0),
    .io_out_1(c53_867_io_out_1),
    .io_out_2(c53_867_io_out_2)
  );
  C53 c53_868 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_868_io_in_0),
    .io_in_1(c53_868_io_in_1),
    .io_in_2(c53_868_io_in_2),
    .io_in_3(c53_868_io_in_3),
    .io_in_4(c53_868_io_in_4),
    .io_out_0(c53_868_io_out_0),
    .io_out_1(c53_868_io_out_1),
    .io_out_2(c53_868_io_out_2)
  );
  C53 c53_869 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_869_io_in_0),
    .io_in_1(c53_869_io_in_1),
    .io_in_2(c53_869_io_in_2),
    .io_in_3(c53_869_io_in_3),
    .io_in_4(c53_869_io_in_4),
    .io_out_0(c53_869_io_out_0),
    .io_out_1(c53_869_io_out_1),
    .io_out_2(c53_869_io_out_2)
  );
  C53 c53_870 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_870_io_in_0),
    .io_in_1(c53_870_io_in_1),
    .io_in_2(c53_870_io_in_2),
    .io_in_3(c53_870_io_in_3),
    .io_in_4(c53_870_io_in_4),
    .io_out_0(c53_870_io_out_0),
    .io_out_1(c53_870_io_out_1),
    .io_out_2(c53_870_io_out_2)
  );
  C53 c53_871 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_871_io_in_0),
    .io_in_1(c53_871_io_in_1),
    .io_in_2(c53_871_io_in_2),
    .io_in_3(c53_871_io_in_3),
    .io_in_4(c53_871_io_in_4),
    .io_out_0(c53_871_io_out_0),
    .io_out_1(c53_871_io_out_1),
    .io_out_2(c53_871_io_out_2)
  );
  C53 c53_872 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_872_io_in_0),
    .io_in_1(c53_872_io_in_1),
    .io_in_2(c53_872_io_in_2),
    .io_in_3(c53_872_io_in_3),
    .io_in_4(c53_872_io_in_4),
    .io_out_0(c53_872_io_out_0),
    .io_out_1(c53_872_io_out_1),
    .io_out_2(c53_872_io_out_2)
  );
  C53 c53_873 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_873_io_in_0),
    .io_in_1(c53_873_io_in_1),
    .io_in_2(c53_873_io_in_2),
    .io_in_3(c53_873_io_in_3),
    .io_in_4(c53_873_io_in_4),
    .io_out_0(c53_873_io_out_0),
    .io_out_1(c53_873_io_out_1),
    .io_out_2(c53_873_io_out_2)
  );
  C53 c53_874 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_874_io_in_0),
    .io_in_1(c53_874_io_in_1),
    .io_in_2(c53_874_io_in_2),
    .io_in_3(c53_874_io_in_3),
    .io_in_4(c53_874_io_in_4),
    .io_out_0(c53_874_io_out_0),
    .io_out_1(c53_874_io_out_1),
    .io_out_2(c53_874_io_out_2)
  );
  C53 c53_875 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_875_io_in_0),
    .io_in_1(c53_875_io_in_1),
    .io_in_2(c53_875_io_in_2),
    .io_in_3(c53_875_io_in_3),
    .io_in_4(c53_875_io_in_4),
    .io_out_0(c53_875_io_out_0),
    .io_out_1(c53_875_io_out_1),
    .io_out_2(c53_875_io_out_2)
  );
  C53 c53_876 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_876_io_in_0),
    .io_in_1(c53_876_io_in_1),
    .io_in_2(c53_876_io_in_2),
    .io_in_3(c53_876_io_in_3),
    .io_in_4(c53_876_io_in_4),
    .io_out_0(c53_876_io_out_0),
    .io_out_1(c53_876_io_out_1),
    .io_out_2(c53_876_io_out_2)
  );
  C53 c53_877 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_877_io_in_0),
    .io_in_1(c53_877_io_in_1),
    .io_in_2(c53_877_io_in_2),
    .io_in_3(c53_877_io_in_3),
    .io_in_4(c53_877_io_in_4),
    .io_out_0(c53_877_io_out_0),
    .io_out_1(c53_877_io_out_1),
    .io_out_2(c53_877_io_out_2)
  );
  C53 c53_878 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_878_io_in_0),
    .io_in_1(c53_878_io_in_1),
    .io_in_2(c53_878_io_in_2),
    .io_in_3(c53_878_io_in_3),
    .io_in_4(c53_878_io_in_4),
    .io_out_0(c53_878_io_out_0),
    .io_out_1(c53_878_io_out_1),
    .io_out_2(c53_878_io_out_2)
  );
  C53 c53_879 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_879_io_in_0),
    .io_in_1(c53_879_io_in_1),
    .io_in_2(c53_879_io_in_2),
    .io_in_3(c53_879_io_in_3),
    .io_in_4(c53_879_io_in_4),
    .io_out_0(c53_879_io_out_0),
    .io_out_1(c53_879_io_out_1),
    .io_out_2(c53_879_io_out_2)
  );
  C53 c53_880 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_880_io_in_0),
    .io_in_1(c53_880_io_in_1),
    .io_in_2(c53_880_io_in_2),
    .io_in_3(c53_880_io_in_3),
    .io_in_4(c53_880_io_in_4),
    .io_out_0(c53_880_io_out_0),
    .io_out_1(c53_880_io_out_1),
    .io_out_2(c53_880_io_out_2)
  );
  C53 c53_881 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_881_io_in_0),
    .io_in_1(c53_881_io_in_1),
    .io_in_2(c53_881_io_in_2),
    .io_in_3(c53_881_io_in_3),
    .io_in_4(c53_881_io_in_4),
    .io_out_0(c53_881_io_out_0),
    .io_out_1(c53_881_io_out_1),
    .io_out_2(c53_881_io_out_2)
  );
  C53 c53_882 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_882_io_in_0),
    .io_in_1(c53_882_io_in_1),
    .io_in_2(c53_882_io_in_2),
    .io_in_3(c53_882_io_in_3),
    .io_in_4(c53_882_io_in_4),
    .io_out_0(c53_882_io_out_0),
    .io_out_1(c53_882_io_out_1),
    .io_out_2(c53_882_io_out_2)
  );
  C53 c53_883 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_883_io_in_0),
    .io_in_1(c53_883_io_in_1),
    .io_in_2(c53_883_io_in_2),
    .io_in_3(c53_883_io_in_3),
    .io_in_4(c53_883_io_in_4),
    .io_out_0(c53_883_io_out_0),
    .io_out_1(c53_883_io_out_1),
    .io_out_2(c53_883_io_out_2)
  );
  C53 c53_884 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_884_io_in_0),
    .io_in_1(c53_884_io_in_1),
    .io_in_2(c53_884_io_in_2),
    .io_in_3(c53_884_io_in_3),
    .io_in_4(c53_884_io_in_4),
    .io_out_0(c53_884_io_out_0),
    .io_out_1(c53_884_io_out_1),
    .io_out_2(c53_884_io_out_2)
  );
  C53 c53_885 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_885_io_in_0),
    .io_in_1(c53_885_io_in_1),
    .io_in_2(c53_885_io_in_2),
    .io_in_3(c53_885_io_in_3),
    .io_in_4(c53_885_io_in_4),
    .io_out_0(c53_885_io_out_0),
    .io_out_1(c53_885_io_out_1),
    .io_out_2(c53_885_io_out_2)
  );
  C53 c53_886 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_886_io_in_0),
    .io_in_1(c53_886_io_in_1),
    .io_in_2(c53_886_io_in_2),
    .io_in_3(c53_886_io_in_3),
    .io_in_4(c53_886_io_in_4),
    .io_out_0(c53_886_io_out_0),
    .io_out_1(c53_886_io_out_1),
    .io_out_2(c53_886_io_out_2)
  );
  C53 c53_887 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_887_io_in_0),
    .io_in_1(c53_887_io_in_1),
    .io_in_2(c53_887_io_in_2),
    .io_in_3(c53_887_io_in_3),
    .io_in_4(c53_887_io_in_4),
    .io_out_0(c53_887_io_out_0),
    .io_out_1(c53_887_io_out_1),
    .io_out_2(c53_887_io_out_2)
  );
  C53 c53_888 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_888_io_in_0),
    .io_in_1(c53_888_io_in_1),
    .io_in_2(c53_888_io_in_2),
    .io_in_3(c53_888_io_in_3),
    .io_in_4(c53_888_io_in_4),
    .io_out_0(c53_888_io_out_0),
    .io_out_1(c53_888_io_out_1),
    .io_out_2(c53_888_io_out_2)
  );
  C53 c53_889 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_889_io_in_0),
    .io_in_1(c53_889_io_in_1),
    .io_in_2(c53_889_io_in_2),
    .io_in_3(c53_889_io_in_3),
    .io_in_4(c53_889_io_in_4),
    .io_out_0(c53_889_io_out_0),
    .io_out_1(c53_889_io_out_1),
    .io_out_2(c53_889_io_out_2)
  );
  C53 c53_890 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_890_io_in_0),
    .io_in_1(c53_890_io_in_1),
    .io_in_2(c53_890_io_in_2),
    .io_in_3(c53_890_io_in_3),
    .io_in_4(c53_890_io_in_4),
    .io_out_0(c53_890_io_out_0),
    .io_out_1(c53_890_io_out_1),
    .io_out_2(c53_890_io_out_2)
  );
  C53 c53_891 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_891_io_in_0),
    .io_in_1(c53_891_io_in_1),
    .io_in_2(c53_891_io_in_2),
    .io_in_3(c53_891_io_in_3),
    .io_in_4(c53_891_io_in_4),
    .io_out_0(c53_891_io_out_0),
    .io_out_1(c53_891_io_out_1),
    .io_out_2(c53_891_io_out_2)
  );
  C53 c53_892 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_892_io_in_0),
    .io_in_1(c53_892_io_in_1),
    .io_in_2(c53_892_io_in_2),
    .io_in_3(c53_892_io_in_3),
    .io_in_4(c53_892_io_in_4),
    .io_out_0(c53_892_io_out_0),
    .io_out_1(c53_892_io_out_1),
    .io_out_2(c53_892_io_out_2)
  );
  C22 c22_99 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_99_io_in_0),
    .io_in_1(c22_99_io_in_1),
    .io_out_0(c22_99_io_out_0),
    .io_out_1(c22_99_io_out_1)
  );
  C53 c53_893 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_893_io_in_0),
    .io_in_1(c53_893_io_in_1),
    .io_in_2(c53_893_io_in_2),
    .io_in_3(c53_893_io_in_3),
    .io_in_4(c53_893_io_in_4),
    .io_out_0(c53_893_io_out_0),
    .io_out_1(c53_893_io_out_1),
    .io_out_2(c53_893_io_out_2)
  );
  C22 c22_100 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_100_io_in_0),
    .io_in_1(c22_100_io_in_1),
    .io_out_0(c22_100_io_out_0),
    .io_out_1(c22_100_io_out_1)
  );
  C53 c53_894 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_894_io_in_0),
    .io_in_1(c53_894_io_in_1),
    .io_in_2(c53_894_io_in_2),
    .io_in_3(c53_894_io_in_3),
    .io_in_4(c53_894_io_in_4),
    .io_out_0(c53_894_io_out_0),
    .io_out_1(c53_894_io_out_1),
    .io_out_2(c53_894_io_out_2)
  );
  C32 c32_60 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_60_io_in_0),
    .io_in_1(c32_60_io_in_1),
    .io_in_2(c32_60_io_in_2),
    .io_out_0(c32_60_io_out_0),
    .io_out_1(c32_60_io_out_1)
  );
  C53 c53_895 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_895_io_in_0),
    .io_in_1(c53_895_io_in_1),
    .io_in_2(c53_895_io_in_2),
    .io_in_3(c53_895_io_in_3),
    .io_in_4(c53_895_io_in_4),
    .io_out_0(c53_895_io_out_0),
    .io_out_1(c53_895_io_out_1),
    .io_out_2(c53_895_io_out_2)
  );
  C22 c22_101 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_101_io_in_0),
    .io_in_1(c22_101_io_in_1),
    .io_out_0(c22_101_io_out_0),
    .io_out_1(c22_101_io_out_1)
  );
  C53 c53_896 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_896_io_in_0),
    .io_in_1(c53_896_io_in_1),
    .io_in_2(c53_896_io_in_2),
    .io_in_3(c53_896_io_in_3),
    .io_in_4(c53_896_io_in_4),
    .io_out_0(c53_896_io_out_0),
    .io_out_1(c53_896_io_out_1),
    .io_out_2(c53_896_io_out_2)
  );
  C22 c22_102 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_102_io_in_0),
    .io_in_1(c22_102_io_in_1),
    .io_out_0(c22_102_io_out_0),
    .io_out_1(c22_102_io_out_1)
  );
  C53 c53_897 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_897_io_in_0),
    .io_in_1(c53_897_io_in_1),
    .io_in_2(c53_897_io_in_2),
    .io_in_3(c53_897_io_in_3),
    .io_in_4(c53_897_io_in_4),
    .io_out_0(c53_897_io_out_0),
    .io_out_1(c53_897_io_out_1),
    .io_out_2(c53_897_io_out_2)
  );
  C22 c22_103 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_103_io_in_0),
    .io_in_1(c22_103_io_in_1),
    .io_out_0(c22_103_io_out_0),
    .io_out_1(c22_103_io_out_1)
  );
  C53 c53_898 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_898_io_in_0),
    .io_in_1(c53_898_io_in_1),
    .io_in_2(c53_898_io_in_2),
    .io_in_3(c53_898_io_in_3),
    .io_in_4(c53_898_io_in_4),
    .io_out_0(c53_898_io_out_0),
    .io_out_1(c53_898_io_out_1),
    .io_out_2(c53_898_io_out_2)
  );
  C22 c22_104 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_104_io_in_0),
    .io_in_1(c22_104_io_in_1),
    .io_out_0(c22_104_io_out_0),
    .io_out_1(c22_104_io_out_1)
  );
  C53 c53_899 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_899_io_in_0),
    .io_in_1(c53_899_io_in_1),
    .io_in_2(c53_899_io_in_2),
    .io_in_3(c53_899_io_in_3),
    .io_in_4(c53_899_io_in_4),
    .io_out_0(c53_899_io_out_0),
    .io_out_1(c53_899_io_out_1),
    .io_out_2(c53_899_io_out_2)
  );
  C32 c32_61 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_61_io_in_0),
    .io_in_1(c32_61_io_in_1),
    .io_in_2(c32_61_io_in_2),
    .io_out_0(c32_61_io_out_0),
    .io_out_1(c32_61_io_out_1)
  );
  C53 c53_900 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_900_io_in_0),
    .io_in_1(c53_900_io_in_1),
    .io_in_2(c53_900_io_in_2),
    .io_in_3(c53_900_io_in_3),
    .io_in_4(c53_900_io_in_4),
    .io_out_0(c53_900_io_out_0),
    .io_out_1(c53_900_io_out_1),
    .io_out_2(c53_900_io_out_2)
  );
  C22 c22_105 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_105_io_in_0),
    .io_in_1(c22_105_io_in_1),
    .io_out_0(c22_105_io_out_0),
    .io_out_1(c22_105_io_out_1)
  );
  C53 c53_901 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_901_io_in_0),
    .io_in_1(c53_901_io_in_1),
    .io_in_2(c53_901_io_in_2),
    .io_in_3(c53_901_io_in_3),
    .io_in_4(c53_901_io_in_4),
    .io_out_0(c53_901_io_out_0),
    .io_out_1(c53_901_io_out_1),
    .io_out_2(c53_901_io_out_2)
  );
  C22 c22_106 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_106_io_in_0),
    .io_in_1(c22_106_io_in_1),
    .io_out_0(c22_106_io_out_0),
    .io_out_1(c22_106_io_out_1)
  );
  C53 c53_902 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_902_io_in_0),
    .io_in_1(c53_902_io_in_1),
    .io_in_2(c53_902_io_in_2),
    .io_in_3(c53_902_io_in_3),
    .io_in_4(c53_902_io_in_4),
    .io_out_0(c53_902_io_out_0),
    .io_out_1(c53_902_io_out_1),
    .io_out_2(c53_902_io_out_2)
  );
  C22 c22_107 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_107_io_in_0),
    .io_in_1(c22_107_io_in_1),
    .io_out_0(c22_107_io_out_0),
    .io_out_1(c22_107_io_out_1)
  );
  C53 c53_903 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_903_io_in_0),
    .io_in_1(c53_903_io_in_1),
    .io_in_2(c53_903_io_in_2),
    .io_in_3(c53_903_io_in_3),
    .io_in_4(c53_903_io_in_4),
    .io_out_0(c53_903_io_out_0),
    .io_out_1(c53_903_io_out_1),
    .io_out_2(c53_903_io_out_2)
  );
  C22 c22_108 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_108_io_in_0),
    .io_in_1(c22_108_io_in_1),
    .io_out_0(c22_108_io_out_0),
    .io_out_1(c22_108_io_out_1)
  );
  C53 c53_904 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_904_io_in_0),
    .io_in_1(c53_904_io_in_1),
    .io_in_2(c53_904_io_in_2),
    .io_in_3(c53_904_io_in_3),
    .io_in_4(c53_904_io_in_4),
    .io_out_0(c53_904_io_out_0),
    .io_out_1(c53_904_io_out_1),
    .io_out_2(c53_904_io_out_2)
  );
  C22 c22_109 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_109_io_in_0),
    .io_in_1(c22_109_io_in_1),
    .io_out_0(c22_109_io_out_0),
    .io_out_1(c22_109_io_out_1)
  );
  C53 c53_905 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_905_io_in_0),
    .io_in_1(c53_905_io_in_1),
    .io_in_2(c53_905_io_in_2),
    .io_in_3(c53_905_io_in_3),
    .io_in_4(c53_905_io_in_4),
    .io_out_0(c53_905_io_out_0),
    .io_out_1(c53_905_io_out_1),
    .io_out_2(c53_905_io_out_2)
  );
  C22 c22_110 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_110_io_in_0),
    .io_in_1(c22_110_io_in_1),
    .io_out_0(c22_110_io_out_0),
    .io_out_1(c22_110_io_out_1)
  );
  C53 c53_906 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_906_io_in_0),
    .io_in_1(c53_906_io_in_1),
    .io_in_2(c53_906_io_in_2),
    .io_in_3(c53_906_io_in_3),
    .io_in_4(c53_906_io_in_4),
    .io_out_0(c53_906_io_out_0),
    .io_out_1(c53_906_io_out_1),
    .io_out_2(c53_906_io_out_2)
  );
  C22 c22_111 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_111_io_in_0),
    .io_in_1(c22_111_io_in_1),
    .io_out_0(c22_111_io_out_0),
    .io_out_1(c22_111_io_out_1)
  );
  C53 c53_907 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_907_io_in_0),
    .io_in_1(c53_907_io_in_1),
    .io_in_2(c53_907_io_in_2),
    .io_in_3(c53_907_io_in_3),
    .io_in_4(c53_907_io_in_4),
    .io_out_0(c53_907_io_out_0),
    .io_out_1(c53_907_io_out_1),
    .io_out_2(c53_907_io_out_2)
  );
  C22 c22_112 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_112_io_in_0),
    .io_in_1(c22_112_io_in_1),
    .io_out_0(c22_112_io_out_0),
    .io_out_1(c22_112_io_out_1)
  );
  C53 c53_908 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_908_io_in_0),
    .io_in_1(c53_908_io_in_1),
    .io_in_2(c53_908_io_in_2),
    .io_in_3(c53_908_io_in_3),
    .io_in_4(c53_908_io_in_4),
    .io_out_0(c53_908_io_out_0),
    .io_out_1(c53_908_io_out_1),
    .io_out_2(c53_908_io_out_2)
  );
  C53 c53_909 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_909_io_in_0),
    .io_in_1(c53_909_io_in_1),
    .io_in_2(c53_909_io_in_2),
    .io_in_3(c53_909_io_in_3),
    .io_in_4(c53_909_io_in_4),
    .io_out_0(c53_909_io_out_0),
    .io_out_1(c53_909_io_out_1),
    .io_out_2(c53_909_io_out_2)
  );
  C53 c53_910 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_910_io_in_0),
    .io_in_1(c53_910_io_in_1),
    .io_in_2(c53_910_io_in_2),
    .io_in_3(c53_910_io_in_3),
    .io_in_4(c53_910_io_in_4),
    .io_out_0(c53_910_io_out_0),
    .io_out_1(c53_910_io_out_1),
    .io_out_2(c53_910_io_out_2)
  );
  C53 c53_911 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_911_io_in_0),
    .io_in_1(c53_911_io_in_1),
    .io_in_2(c53_911_io_in_2),
    .io_in_3(c53_911_io_in_3),
    .io_in_4(c53_911_io_in_4),
    .io_out_0(c53_911_io_out_0),
    .io_out_1(c53_911_io_out_1),
    .io_out_2(c53_911_io_out_2)
  );
  C53 c53_912 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_912_io_in_0),
    .io_in_1(c53_912_io_in_1),
    .io_in_2(c53_912_io_in_2),
    .io_in_3(c53_912_io_in_3),
    .io_in_4(c53_912_io_in_4),
    .io_out_0(c53_912_io_out_0),
    .io_out_1(c53_912_io_out_1),
    .io_out_2(c53_912_io_out_2)
  );
  C53 c53_913 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_913_io_in_0),
    .io_in_1(c53_913_io_in_1),
    .io_in_2(c53_913_io_in_2),
    .io_in_3(c53_913_io_in_3),
    .io_in_4(c53_913_io_in_4),
    .io_out_0(c53_913_io_out_0),
    .io_out_1(c53_913_io_out_1),
    .io_out_2(c53_913_io_out_2)
  );
  C53 c53_914 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_914_io_in_0),
    .io_in_1(c53_914_io_in_1),
    .io_in_2(c53_914_io_in_2),
    .io_in_3(c53_914_io_in_3),
    .io_in_4(c53_914_io_in_4),
    .io_out_0(c53_914_io_out_0),
    .io_out_1(c53_914_io_out_1),
    .io_out_2(c53_914_io_out_2)
  );
  C53 c53_915 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_915_io_in_0),
    .io_in_1(c53_915_io_in_1),
    .io_in_2(c53_915_io_in_2),
    .io_in_3(c53_915_io_in_3),
    .io_in_4(c53_915_io_in_4),
    .io_out_0(c53_915_io_out_0),
    .io_out_1(c53_915_io_out_1),
    .io_out_2(c53_915_io_out_2)
  );
  C53 c53_916 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_916_io_in_0),
    .io_in_1(c53_916_io_in_1),
    .io_in_2(c53_916_io_in_2),
    .io_in_3(c53_916_io_in_3),
    .io_in_4(c53_916_io_in_4),
    .io_out_0(c53_916_io_out_0),
    .io_out_1(c53_916_io_out_1),
    .io_out_2(c53_916_io_out_2)
  );
  C53 c53_917 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_917_io_in_0),
    .io_in_1(c53_917_io_in_1),
    .io_in_2(c53_917_io_in_2),
    .io_in_3(c53_917_io_in_3),
    .io_in_4(c53_917_io_in_4),
    .io_out_0(c53_917_io_out_0),
    .io_out_1(c53_917_io_out_1),
    .io_out_2(c53_917_io_out_2)
  );
  C53 c53_918 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_918_io_in_0),
    .io_in_1(c53_918_io_in_1),
    .io_in_2(c53_918_io_in_2),
    .io_in_3(c53_918_io_in_3),
    .io_in_4(c53_918_io_in_4),
    .io_out_0(c53_918_io_out_0),
    .io_out_1(c53_918_io_out_1),
    .io_out_2(c53_918_io_out_2)
  );
  C53 c53_919 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_919_io_in_0),
    .io_in_1(c53_919_io_in_1),
    .io_in_2(c53_919_io_in_2),
    .io_in_3(c53_919_io_in_3),
    .io_in_4(c53_919_io_in_4),
    .io_out_0(c53_919_io_out_0),
    .io_out_1(c53_919_io_out_1),
    .io_out_2(c53_919_io_out_2)
  );
  C53 c53_920 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_920_io_in_0),
    .io_in_1(c53_920_io_in_1),
    .io_in_2(c53_920_io_in_2),
    .io_in_3(c53_920_io_in_3),
    .io_in_4(c53_920_io_in_4),
    .io_out_0(c53_920_io_out_0),
    .io_out_1(c53_920_io_out_1),
    .io_out_2(c53_920_io_out_2)
  );
  C53 c53_921 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_921_io_in_0),
    .io_in_1(c53_921_io_in_1),
    .io_in_2(c53_921_io_in_2),
    .io_in_3(c53_921_io_in_3),
    .io_in_4(c53_921_io_in_4),
    .io_out_0(c53_921_io_out_0),
    .io_out_1(c53_921_io_out_1),
    .io_out_2(c53_921_io_out_2)
  );
  C53 c53_922 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_922_io_in_0),
    .io_in_1(c53_922_io_in_1),
    .io_in_2(c53_922_io_in_2),
    .io_in_3(c53_922_io_in_3),
    .io_in_4(c53_922_io_in_4),
    .io_out_0(c53_922_io_out_0),
    .io_out_1(c53_922_io_out_1),
    .io_out_2(c53_922_io_out_2)
  );
  C53 c53_923 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_923_io_in_0),
    .io_in_1(c53_923_io_in_1),
    .io_in_2(c53_923_io_in_2),
    .io_in_3(c53_923_io_in_3),
    .io_in_4(c53_923_io_in_4),
    .io_out_0(c53_923_io_out_0),
    .io_out_1(c53_923_io_out_1),
    .io_out_2(c53_923_io_out_2)
  );
  C22 c22_113 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_113_io_in_0),
    .io_in_1(c22_113_io_in_1),
    .io_out_0(c22_113_io_out_0),
    .io_out_1(c22_113_io_out_1)
  );
  C22 c22_114 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_114_io_in_0),
    .io_in_1(c22_114_io_in_1),
    .io_out_0(c22_114_io_out_0),
    .io_out_1(c22_114_io_out_1)
  );
  C32 c32_62 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_62_io_in_0),
    .io_in_1(c32_62_io_in_1),
    .io_in_2(c32_62_io_in_2),
    .io_out_0(c32_62_io_out_0),
    .io_out_1(c32_62_io_out_1)
  );
  C22 c22_115 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_115_io_in_0),
    .io_in_1(c22_115_io_in_1),
    .io_out_0(c22_115_io_out_0),
    .io_out_1(c22_115_io_out_1)
  );
  C22 c22_116 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_116_io_in_0),
    .io_in_1(c22_116_io_in_1),
    .io_out_0(c22_116_io_out_0),
    .io_out_1(c22_116_io_out_1)
  );
  C22 c22_117 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_117_io_in_0),
    .io_in_1(c22_117_io_in_1),
    .io_out_0(c22_117_io_out_0),
    .io_out_1(c22_117_io_out_1)
  );
  C22 c22_118 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_118_io_in_0),
    .io_in_1(c22_118_io_in_1),
    .io_out_0(c22_118_io_out_0),
    .io_out_1(c22_118_io_out_1)
  );
  C32 c32_63 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_63_io_in_0),
    .io_in_1(c32_63_io_in_1),
    .io_in_2(c32_63_io_in_2),
    .io_out_0(c32_63_io_out_0),
    .io_out_1(c32_63_io_out_1)
  );
  C22 c22_119 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_119_io_in_0),
    .io_in_1(c22_119_io_in_1),
    .io_out_0(c22_119_io_out_0),
    .io_out_1(c22_119_io_out_1)
  );
  C22 c22_120 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_120_io_in_0),
    .io_in_1(c22_120_io_in_1),
    .io_out_0(c22_120_io_out_0),
    .io_out_1(c22_120_io_out_1)
  );
  C22 c22_121 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_121_io_in_0),
    .io_in_1(c22_121_io_in_1),
    .io_out_0(c22_121_io_out_0),
    .io_out_1(c22_121_io_out_1)
  );
  C22 c22_122 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_122_io_in_0),
    .io_in_1(c22_122_io_in_1),
    .io_out_0(c22_122_io_out_0),
    .io_out_1(c22_122_io_out_1)
  );
  C22 c22_123 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_123_io_in_0),
    .io_in_1(c22_123_io_in_1),
    .io_out_0(c22_123_io_out_0),
    .io_out_1(c22_123_io_out_1)
  );
  C22 c22_124 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_124_io_in_0),
    .io_in_1(c22_124_io_in_1),
    .io_out_0(c22_124_io_out_0),
    .io_out_1(c22_124_io_out_1)
  );
  C22 c22_125 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_125_io_in_0),
    .io_in_1(c22_125_io_in_1),
    .io_out_0(c22_125_io_out_0),
    .io_out_1(c22_125_io_out_1)
  );
  C22 c22_126 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_126_io_in_0),
    .io_in_1(c22_126_io_in_1),
    .io_out_0(c22_126_io_out_0),
    .io_out_1(c22_126_io_out_1)
  );
  C22 c22_127 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_127_io_in_0),
    .io_in_1(c22_127_io_in_1),
    .io_out_0(c22_127_io_out_0),
    .io_out_1(c22_127_io_out_1)
  );
  C22 c22_128 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_128_io_in_0),
    .io_in_1(c22_128_io_in_1),
    .io_out_0(c22_128_io_out_0),
    .io_out_1(c22_128_io_out_1)
  );
  C22 c22_129 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_129_io_in_0),
    .io_in_1(c22_129_io_in_1),
    .io_out_0(c22_129_io_out_0),
    .io_out_1(c22_129_io_out_1)
  );
  C22 c22_130 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_130_io_in_0),
    .io_in_1(c22_130_io_in_1),
    .io_out_0(c22_130_io_out_0),
    .io_out_1(c22_130_io_out_1)
  );
  C22 c22_131 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_131_io_in_0),
    .io_in_1(c22_131_io_in_1),
    .io_out_0(c22_131_io_out_0),
    .io_out_1(c22_131_io_out_1)
  );
  C22 c22_132 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_132_io_in_0),
    .io_in_1(c22_132_io_in_1),
    .io_out_0(c22_132_io_out_0),
    .io_out_1(c22_132_io_out_1)
  );
  C22 c22_133 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_133_io_in_0),
    .io_in_1(c22_133_io_in_1),
    .io_out_0(c22_133_io_out_0),
    .io_out_1(c22_133_io_out_1)
  );
  C22 c22_134 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_134_io_in_0),
    .io_in_1(c22_134_io_in_1),
    .io_out_0(c22_134_io_out_0),
    .io_out_1(c22_134_io_out_1)
  );
  C22 c22_135 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_135_io_in_0),
    .io_in_1(c22_135_io_in_1),
    .io_out_0(c22_135_io_out_0),
    .io_out_1(c22_135_io_out_1)
  );
  C22 c22_136 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_136_io_in_0),
    .io_in_1(c22_136_io_in_1),
    .io_out_0(c22_136_io_out_0),
    .io_out_1(c22_136_io_out_1)
  );
  C22 c22_137 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_137_io_in_0),
    .io_in_1(c22_137_io_in_1),
    .io_out_0(c22_137_io_out_0),
    .io_out_1(c22_137_io_out_1)
  );
  C22 c22_138 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_138_io_in_0),
    .io_in_1(c22_138_io_in_1),
    .io_out_0(c22_138_io_out_0),
    .io_out_1(c22_138_io_out_1)
  );
  C22 c22_139 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_139_io_in_0),
    .io_in_1(c22_139_io_in_1),
    .io_out_0(c22_139_io_out_0),
    .io_out_1(c22_139_io_out_1)
  );
  C22 c22_140 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_140_io_in_0),
    .io_in_1(c22_140_io_in_1),
    .io_out_0(c22_140_io_out_0),
    .io_out_1(c22_140_io_out_1)
  );
  C22 c22_141 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_141_io_in_0),
    .io_in_1(c22_141_io_in_1),
    .io_out_0(c22_141_io_out_0),
    .io_out_1(c22_141_io_out_1)
  );
  C22 c22_142 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_142_io_in_0),
    .io_in_1(c22_142_io_in_1),
    .io_out_0(c22_142_io_out_0),
    .io_out_1(c22_142_io_out_1)
  );
  C22 c22_143 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_143_io_in_0),
    .io_in_1(c22_143_io_in_1),
    .io_out_0(c22_143_io_out_0),
    .io_out_1(c22_143_io_out_1)
  );
  C22 c22_144 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_144_io_in_0),
    .io_in_1(c22_144_io_in_1),
    .io_out_0(c22_144_io_out_0),
    .io_out_1(c22_144_io_out_1)
  );
  C22 c22_145 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_145_io_in_0),
    .io_in_1(c22_145_io_in_1),
    .io_out_0(c22_145_io_out_0),
    .io_out_1(c22_145_io_out_1)
  );
  C22 c22_146 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_146_io_in_0),
    .io_in_1(c22_146_io_in_1),
    .io_out_0(c22_146_io_out_0),
    .io_out_1(c22_146_io_out_1)
  );
  C22 c22_147 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_147_io_in_0),
    .io_in_1(c22_147_io_in_1),
    .io_out_0(c22_147_io_out_0),
    .io_out_1(c22_147_io_out_1)
  );
  C22 c22_148 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_148_io_in_0),
    .io_in_1(c22_148_io_in_1),
    .io_out_0(c22_148_io_out_0),
    .io_out_1(c22_148_io_out_1)
  );
  C22 c22_149 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_149_io_in_0),
    .io_in_1(c22_149_io_in_1),
    .io_out_0(c22_149_io_out_0),
    .io_out_1(c22_149_io_out_1)
  );
  C22 c22_150 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_150_io_in_0),
    .io_in_1(c22_150_io_in_1),
    .io_out_0(c22_150_io_out_0),
    .io_out_1(c22_150_io_out_1)
  );
  C22 c22_151 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_151_io_in_0),
    .io_in_1(c22_151_io_in_1),
    .io_out_0(c22_151_io_out_0),
    .io_out_1(c22_151_io_out_1)
  );
  C32 c32_64 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_64_io_in_0),
    .io_in_1(c32_64_io_in_1),
    .io_in_2(c32_64_io_in_2),
    .io_out_0(c32_64_io_out_0),
    .io_out_1(c32_64_io_out_1)
  );
  C32 c32_65 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_65_io_in_0),
    .io_in_1(c32_65_io_in_1),
    .io_in_2(c32_65_io_in_2),
    .io_out_0(c32_65_io_out_0),
    .io_out_1(c32_65_io_out_1)
  );
  C32 c32_66 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_66_io_in_0),
    .io_in_1(c32_66_io_in_1),
    .io_in_2(c32_66_io_in_2),
    .io_out_0(c32_66_io_out_0),
    .io_out_1(c32_66_io_out_1)
  );
  C32 c32_67 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_67_io_in_0),
    .io_in_1(c32_67_io_in_1),
    .io_in_2(c32_67_io_in_2),
    .io_out_0(c32_67_io_out_0),
    .io_out_1(c32_67_io_out_1)
  );
  C32 c32_68 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_68_io_in_0),
    .io_in_1(c32_68_io_in_1),
    .io_in_2(c32_68_io_in_2),
    .io_out_0(c32_68_io_out_0),
    .io_out_1(c32_68_io_out_1)
  );
  C53 c53_924 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_924_io_in_0),
    .io_in_1(c53_924_io_in_1),
    .io_in_2(c53_924_io_in_2),
    .io_in_3(c53_924_io_in_3),
    .io_in_4(c53_924_io_in_4),
    .io_out_0(c53_924_io_out_0),
    .io_out_1(c53_924_io_out_1),
    .io_out_2(c53_924_io_out_2)
  );
  C53 c53_925 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_925_io_in_0),
    .io_in_1(c53_925_io_in_1),
    .io_in_2(c53_925_io_in_2),
    .io_in_3(c53_925_io_in_3),
    .io_in_4(c53_925_io_in_4),
    .io_out_0(c53_925_io_out_0),
    .io_out_1(c53_925_io_out_1),
    .io_out_2(c53_925_io_out_2)
  );
  C53 c53_926 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_926_io_in_0),
    .io_in_1(c53_926_io_in_1),
    .io_in_2(c53_926_io_in_2),
    .io_in_3(c53_926_io_in_3),
    .io_in_4(c53_926_io_in_4),
    .io_out_0(c53_926_io_out_0),
    .io_out_1(c53_926_io_out_1),
    .io_out_2(c53_926_io_out_2)
  );
  C53 c53_927 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_927_io_in_0),
    .io_in_1(c53_927_io_in_1),
    .io_in_2(c53_927_io_in_2),
    .io_in_3(c53_927_io_in_3),
    .io_in_4(c53_927_io_in_4),
    .io_out_0(c53_927_io_out_0),
    .io_out_1(c53_927_io_out_1),
    .io_out_2(c53_927_io_out_2)
  );
  C53 c53_928 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_928_io_in_0),
    .io_in_1(c53_928_io_in_1),
    .io_in_2(c53_928_io_in_2),
    .io_in_3(c53_928_io_in_3),
    .io_in_4(c53_928_io_in_4),
    .io_out_0(c53_928_io_out_0),
    .io_out_1(c53_928_io_out_1),
    .io_out_2(c53_928_io_out_2)
  );
  C53 c53_929 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_929_io_in_0),
    .io_in_1(c53_929_io_in_1),
    .io_in_2(c53_929_io_in_2),
    .io_in_3(c53_929_io_in_3),
    .io_in_4(c53_929_io_in_4),
    .io_out_0(c53_929_io_out_0),
    .io_out_1(c53_929_io_out_1),
    .io_out_2(c53_929_io_out_2)
  );
  C53 c53_930 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_930_io_in_0),
    .io_in_1(c53_930_io_in_1),
    .io_in_2(c53_930_io_in_2),
    .io_in_3(c53_930_io_in_3),
    .io_in_4(c53_930_io_in_4),
    .io_out_0(c53_930_io_out_0),
    .io_out_1(c53_930_io_out_1),
    .io_out_2(c53_930_io_out_2)
  );
  C53 c53_931 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_931_io_in_0),
    .io_in_1(c53_931_io_in_1),
    .io_in_2(c53_931_io_in_2),
    .io_in_3(c53_931_io_in_3),
    .io_in_4(c53_931_io_in_4),
    .io_out_0(c53_931_io_out_0),
    .io_out_1(c53_931_io_out_1),
    .io_out_2(c53_931_io_out_2)
  );
  C53 c53_932 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_932_io_in_0),
    .io_in_1(c53_932_io_in_1),
    .io_in_2(c53_932_io_in_2),
    .io_in_3(c53_932_io_in_3),
    .io_in_4(c53_932_io_in_4),
    .io_out_0(c53_932_io_out_0),
    .io_out_1(c53_932_io_out_1),
    .io_out_2(c53_932_io_out_2)
  );
  C53 c53_933 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_933_io_in_0),
    .io_in_1(c53_933_io_in_1),
    .io_in_2(c53_933_io_in_2),
    .io_in_3(c53_933_io_in_3),
    .io_in_4(c53_933_io_in_4),
    .io_out_0(c53_933_io_out_0),
    .io_out_1(c53_933_io_out_1),
    .io_out_2(c53_933_io_out_2)
  );
  C53 c53_934 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_934_io_in_0),
    .io_in_1(c53_934_io_in_1),
    .io_in_2(c53_934_io_in_2),
    .io_in_3(c53_934_io_in_3),
    .io_in_4(c53_934_io_in_4),
    .io_out_0(c53_934_io_out_0),
    .io_out_1(c53_934_io_out_1),
    .io_out_2(c53_934_io_out_2)
  );
  C53 c53_935 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_935_io_in_0),
    .io_in_1(c53_935_io_in_1),
    .io_in_2(c53_935_io_in_2),
    .io_in_3(c53_935_io_in_3),
    .io_in_4(c53_935_io_in_4),
    .io_out_0(c53_935_io_out_0),
    .io_out_1(c53_935_io_out_1),
    .io_out_2(c53_935_io_out_2)
  );
  C53 c53_936 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_936_io_in_0),
    .io_in_1(c53_936_io_in_1),
    .io_in_2(c53_936_io_in_2),
    .io_in_3(c53_936_io_in_3),
    .io_in_4(c53_936_io_in_4),
    .io_out_0(c53_936_io_out_0),
    .io_out_1(c53_936_io_out_1),
    .io_out_2(c53_936_io_out_2)
  );
  C53 c53_937 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_937_io_in_0),
    .io_in_1(c53_937_io_in_1),
    .io_in_2(c53_937_io_in_2),
    .io_in_3(c53_937_io_in_3),
    .io_in_4(c53_937_io_in_4),
    .io_out_0(c53_937_io_out_0),
    .io_out_1(c53_937_io_out_1),
    .io_out_2(c53_937_io_out_2)
  );
  C53 c53_938 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_938_io_in_0),
    .io_in_1(c53_938_io_in_1),
    .io_in_2(c53_938_io_in_2),
    .io_in_3(c53_938_io_in_3),
    .io_in_4(c53_938_io_in_4),
    .io_out_0(c53_938_io_out_0),
    .io_out_1(c53_938_io_out_1),
    .io_out_2(c53_938_io_out_2)
  );
  C53 c53_939 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_939_io_in_0),
    .io_in_1(c53_939_io_in_1),
    .io_in_2(c53_939_io_in_2),
    .io_in_3(c53_939_io_in_3),
    .io_in_4(c53_939_io_in_4),
    .io_out_0(c53_939_io_out_0),
    .io_out_1(c53_939_io_out_1),
    .io_out_2(c53_939_io_out_2)
  );
  C53 c53_940 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_940_io_in_0),
    .io_in_1(c53_940_io_in_1),
    .io_in_2(c53_940_io_in_2),
    .io_in_3(c53_940_io_in_3),
    .io_in_4(c53_940_io_in_4),
    .io_out_0(c53_940_io_out_0),
    .io_out_1(c53_940_io_out_1),
    .io_out_2(c53_940_io_out_2)
  );
  C53 c53_941 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_941_io_in_0),
    .io_in_1(c53_941_io_in_1),
    .io_in_2(c53_941_io_in_2),
    .io_in_3(c53_941_io_in_3),
    .io_in_4(c53_941_io_in_4),
    .io_out_0(c53_941_io_out_0),
    .io_out_1(c53_941_io_out_1),
    .io_out_2(c53_941_io_out_2)
  );
  C53 c53_942 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_942_io_in_0),
    .io_in_1(c53_942_io_in_1),
    .io_in_2(c53_942_io_in_2),
    .io_in_3(c53_942_io_in_3),
    .io_in_4(c53_942_io_in_4),
    .io_out_0(c53_942_io_out_0),
    .io_out_1(c53_942_io_out_1),
    .io_out_2(c53_942_io_out_2)
  );
  C53 c53_943 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_943_io_in_0),
    .io_in_1(c53_943_io_in_1),
    .io_in_2(c53_943_io_in_2),
    .io_in_3(c53_943_io_in_3),
    .io_in_4(c53_943_io_in_4),
    .io_out_0(c53_943_io_out_0),
    .io_out_1(c53_943_io_out_1),
    .io_out_2(c53_943_io_out_2)
  );
  C53 c53_944 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_944_io_in_0),
    .io_in_1(c53_944_io_in_1),
    .io_in_2(c53_944_io_in_2),
    .io_in_3(c53_944_io_in_3),
    .io_in_4(c53_944_io_in_4),
    .io_out_0(c53_944_io_out_0),
    .io_out_1(c53_944_io_out_1),
    .io_out_2(c53_944_io_out_2)
  );
  C53 c53_945 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_945_io_in_0),
    .io_in_1(c53_945_io_in_1),
    .io_in_2(c53_945_io_in_2),
    .io_in_3(c53_945_io_in_3),
    .io_in_4(c53_945_io_in_4),
    .io_out_0(c53_945_io_out_0),
    .io_out_1(c53_945_io_out_1),
    .io_out_2(c53_945_io_out_2)
  );
  C53 c53_946 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_946_io_in_0),
    .io_in_1(c53_946_io_in_1),
    .io_in_2(c53_946_io_in_2),
    .io_in_3(c53_946_io_in_3),
    .io_in_4(c53_946_io_in_4),
    .io_out_0(c53_946_io_out_0),
    .io_out_1(c53_946_io_out_1),
    .io_out_2(c53_946_io_out_2)
  );
  C53 c53_947 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_947_io_in_0),
    .io_in_1(c53_947_io_in_1),
    .io_in_2(c53_947_io_in_2),
    .io_in_3(c53_947_io_in_3),
    .io_in_4(c53_947_io_in_4),
    .io_out_0(c53_947_io_out_0),
    .io_out_1(c53_947_io_out_1),
    .io_out_2(c53_947_io_out_2)
  );
  C53 c53_948 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_948_io_in_0),
    .io_in_1(c53_948_io_in_1),
    .io_in_2(c53_948_io_in_2),
    .io_in_3(c53_948_io_in_3),
    .io_in_4(c53_948_io_in_4),
    .io_out_0(c53_948_io_out_0),
    .io_out_1(c53_948_io_out_1),
    .io_out_2(c53_948_io_out_2)
  );
  C53 c53_949 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_949_io_in_0),
    .io_in_1(c53_949_io_in_1),
    .io_in_2(c53_949_io_in_2),
    .io_in_3(c53_949_io_in_3),
    .io_in_4(c53_949_io_in_4),
    .io_out_0(c53_949_io_out_0),
    .io_out_1(c53_949_io_out_1),
    .io_out_2(c53_949_io_out_2)
  );
  C53 c53_950 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_950_io_in_0),
    .io_in_1(c53_950_io_in_1),
    .io_in_2(c53_950_io_in_2),
    .io_in_3(c53_950_io_in_3),
    .io_in_4(c53_950_io_in_4),
    .io_out_0(c53_950_io_out_0),
    .io_out_1(c53_950_io_out_1),
    .io_out_2(c53_950_io_out_2)
  );
  C53 c53_951 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_951_io_in_0),
    .io_in_1(c53_951_io_in_1),
    .io_in_2(c53_951_io_in_2),
    .io_in_3(c53_951_io_in_3),
    .io_in_4(c53_951_io_in_4),
    .io_out_0(c53_951_io_out_0),
    .io_out_1(c53_951_io_out_1),
    .io_out_2(c53_951_io_out_2)
  );
  C53 c53_952 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_952_io_in_0),
    .io_in_1(c53_952_io_in_1),
    .io_in_2(c53_952_io_in_2),
    .io_in_3(c53_952_io_in_3),
    .io_in_4(c53_952_io_in_4),
    .io_out_0(c53_952_io_out_0),
    .io_out_1(c53_952_io_out_1),
    .io_out_2(c53_952_io_out_2)
  );
  C53 c53_953 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_953_io_in_0),
    .io_in_1(c53_953_io_in_1),
    .io_in_2(c53_953_io_in_2),
    .io_in_3(c53_953_io_in_3),
    .io_in_4(c53_953_io_in_4),
    .io_out_0(c53_953_io_out_0),
    .io_out_1(c53_953_io_out_1),
    .io_out_2(c53_953_io_out_2)
  );
  C53 c53_954 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_954_io_in_0),
    .io_in_1(c53_954_io_in_1),
    .io_in_2(c53_954_io_in_2),
    .io_in_3(c53_954_io_in_3),
    .io_in_4(c53_954_io_in_4),
    .io_out_0(c53_954_io_out_0),
    .io_out_1(c53_954_io_out_1),
    .io_out_2(c53_954_io_out_2)
  );
  C53 c53_955 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_955_io_in_0),
    .io_in_1(c53_955_io_in_1),
    .io_in_2(c53_955_io_in_2),
    .io_in_3(c53_955_io_in_3),
    .io_in_4(c53_955_io_in_4),
    .io_out_0(c53_955_io_out_0),
    .io_out_1(c53_955_io_out_1),
    .io_out_2(c53_955_io_out_2)
  );
  C53 c53_956 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_956_io_in_0),
    .io_in_1(c53_956_io_in_1),
    .io_in_2(c53_956_io_in_2),
    .io_in_3(c53_956_io_in_3),
    .io_in_4(c53_956_io_in_4),
    .io_out_0(c53_956_io_out_0),
    .io_out_1(c53_956_io_out_1),
    .io_out_2(c53_956_io_out_2)
  );
  C53 c53_957 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_957_io_in_0),
    .io_in_1(c53_957_io_in_1),
    .io_in_2(c53_957_io_in_2),
    .io_in_3(c53_957_io_in_3),
    .io_in_4(c53_957_io_in_4),
    .io_out_0(c53_957_io_out_0),
    .io_out_1(c53_957_io_out_1),
    .io_out_2(c53_957_io_out_2)
  );
  C53 c53_958 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_958_io_in_0),
    .io_in_1(c53_958_io_in_1),
    .io_in_2(c53_958_io_in_2),
    .io_in_3(c53_958_io_in_3),
    .io_in_4(c53_958_io_in_4),
    .io_out_0(c53_958_io_out_0),
    .io_out_1(c53_958_io_out_1),
    .io_out_2(c53_958_io_out_2)
  );
  C53 c53_959 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_959_io_in_0),
    .io_in_1(c53_959_io_in_1),
    .io_in_2(c53_959_io_in_2),
    .io_in_3(c53_959_io_in_3),
    .io_in_4(c53_959_io_in_4),
    .io_out_0(c53_959_io_out_0),
    .io_out_1(c53_959_io_out_1),
    .io_out_2(c53_959_io_out_2)
  );
  C53 c53_960 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_960_io_in_0),
    .io_in_1(c53_960_io_in_1),
    .io_in_2(c53_960_io_in_2),
    .io_in_3(c53_960_io_in_3),
    .io_in_4(c53_960_io_in_4),
    .io_out_0(c53_960_io_out_0),
    .io_out_1(c53_960_io_out_1),
    .io_out_2(c53_960_io_out_2)
  );
  C53 c53_961 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_961_io_in_0),
    .io_in_1(c53_961_io_in_1),
    .io_in_2(c53_961_io_in_2),
    .io_in_3(c53_961_io_in_3),
    .io_in_4(c53_961_io_in_4),
    .io_out_0(c53_961_io_out_0),
    .io_out_1(c53_961_io_out_1),
    .io_out_2(c53_961_io_out_2)
  );
  C53 c53_962 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_962_io_in_0),
    .io_in_1(c53_962_io_in_1),
    .io_in_2(c53_962_io_in_2),
    .io_in_3(c53_962_io_in_3),
    .io_in_4(c53_962_io_in_4),
    .io_out_0(c53_962_io_out_0),
    .io_out_1(c53_962_io_out_1),
    .io_out_2(c53_962_io_out_2)
  );
  C53 c53_963 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_963_io_in_0),
    .io_in_1(c53_963_io_in_1),
    .io_in_2(c53_963_io_in_2),
    .io_in_3(c53_963_io_in_3),
    .io_in_4(c53_963_io_in_4),
    .io_out_0(c53_963_io_out_0),
    .io_out_1(c53_963_io_out_1),
    .io_out_2(c53_963_io_out_2)
  );
  C53 c53_964 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_964_io_in_0),
    .io_in_1(c53_964_io_in_1),
    .io_in_2(c53_964_io_in_2),
    .io_in_3(c53_964_io_in_3),
    .io_in_4(c53_964_io_in_4),
    .io_out_0(c53_964_io_out_0),
    .io_out_1(c53_964_io_out_1),
    .io_out_2(c53_964_io_out_2)
  );
  C53 c53_965 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_965_io_in_0),
    .io_in_1(c53_965_io_in_1),
    .io_in_2(c53_965_io_in_2),
    .io_in_3(c53_965_io_in_3),
    .io_in_4(c53_965_io_in_4),
    .io_out_0(c53_965_io_out_0),
    .io_out_1(c53_965_io_out_1),
    .io_out_2(c53_965_io_out_2)
  );
  C53 c53_966 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_966_io_in_0),
    .io_in_1(c53_966_io_in_1),
    .io_in_2(c53_966_io_in_2),
    .io_in_3(c53_966_io_in_3),
    .io_in_4(c53_966_io_in_4),
    .io_out_0(c53_966_io_out_0),
    .io_out_1(c53_966_io_out_1),
    .io_out_2(c53_966_io_out_2)
  );
  C53 c53_967 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_967_io_in_0),
    .io_in_1(c53_967_io_in_1),
    .io_in_2(c53_967_io_in_2),
    .io_in_3(c53_967_io_in_3),
    .io_in_4(c53_967_io_in_4),
    .io_out_0(c53_967_io_out_0),
    .io_out_1(c53_967_io_out_1),
    .io_out_2(c53_967_io_out_2)
  );
  C53 c53_968 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_968_io_in_0),
    .io_in_1(c53_968_io_in_1),
    .io_in_2(c53_968_io_in_2),
    .io_in_3(c53_968_io_in_3),
    .io_in_4(c53_968_io_in_4),
    .io_out_0(c53_968_io_out_0),
    .io_out_1(c53_968_io_out_1),
    .io_out_2(c53_968_io_out_2)
  );
  C53 c53_969 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_969_io_in_0),
    .io_in_1(c53_969_io_in_1),
    .io_in_2(c53_969_io_in_2),
    .io_in_3(c53_969_io_in_3),
    .io_in_4(c53_969_io_in_4),
    .io_out_0(c53_969_io_out_0),
    .io_out_1(c53_969_io_out_1),
    .io_out_2(c53_969_io_out_2)
  );
  C53 c53_970 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_970_io_in_0),
    .io_in_1(c53_970_io_in_1),
    .io_in_2(c53_970_io_in_2),
    .io_in_3(c53_970_io_in_3),
    .io_in_4(c53_970_io_in_4),
    .io_out_0(c53_970_io_out_0),
    .io_out_1(c53_970_io_out_1),
    .io_out_2(c53_970_io_out_2)
  );
  C53 c53_971 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_971_io_in_0),
    .io_in_1(c53_971_io_in_1),
    .io_in_2(c53_971_io_in_2),
    .io_in_3(c53_971_io_in_3),
    .io_in_4(c53_971_io_in_4),
    .io_out_0(c53_971_io_out_0),
    .io_out_1(c53_971_io_out_1),
    .io_out_2(c53_971_io_out_2)
  );
  C53 c53_972 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_972_io_in_0),
    .io_in_1(c53_972_io_in_1),
    .io_in_2(c53_972_io_in_2),
    .io_in_3(c53_972_io_in_3),
    .io_in_4(c53_972_io_in_4),
    .io_out_0(c53_972_io_out_0),
    .io_out_1(c53_972_io_out_1),
    .io_out_2(c53_972_io_out_2)
  );
  C53 c53_973 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_973_io_in_0),
    .io_in_1(c53_973_io_in_1),
    .io_in_2(c53_973_io_in_2),
    .io_in_3(c53_973_io_in_3),
    .io_in_4(c53_973_io_in_4),
    .io_out_0(c53_973_io_out_0),
    .io_out_1(c53_973_io_out_1),
    .io_out_2(c53_973_io_out_2)
  );
  C53 c53_974 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_974_io_in_0),
    .io_in_1(c53_974_io_in_1),
    .io_in_2(c53_974_io_in_2),
    .io_in_3(c53_974_io_in_3),
    .io_in_4(c53_974_io_in_4),
    .io_out_0(c53_974_io_out_0),
    .io_out_1(c53_974_io_out_1),
    .io_out_2(c53_974_io_out_2)
  );
  C53 c53_975 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_975_io_in_0),
    .io_in_1(c53_975_io_in_1),
    .io_in_2(c53_975_io_in_2),
    .io_in_3(c53_975_io_in_3),
    .io_in_4(c53_975_io_in_4),
    .io_out_0(c53_975_io_out_0),
    .io_out_1(c53_975_io_out_1),
    .io_out_2(c53_975_io_out_2)
  );
  C53 c53_976 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_976_io_in_0),
    .io_in_1(c53_976_io_in_1),
    .io_in_2(c53_976_io_in_2),
    .io_in_3(c53_976_io_in_3),
    .io_in_4(c53_976_io_in_4),
    .io_out_0(c53_976_io_out_0),
    .io_out_1(c53_976_io_out_1),
    .io_out_2(c53_976_io_out_2)
  );
  C53 c53_977 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_977_io_in_0),
    .io_in_1(c53_977_io_in_1),
    .io_in_2(c53_977_io_in_2),
    .io_in_3(c53_977_io_in_3),
    .io_in_4(c53_977_io_in_4),
    .io_out_0(c53_977_io_out_0),
    .io_out_1(c53_977_io_out_1),
    .io_out_2(c53_977_io_out_2)
  );
  C53 c53_978 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_978_io_in_0),
    .io_in_1(c53_978_io_in_1),
    .io_in_2(c53_978_io_in_2),
    .io_in_3(c53_978_io_in_3),
    .io_in_4(c53_978_io_in_4),
    .io_out_0(c53_978_io_out_0),
    .io_out_1(c53_978_io_out_1),
    .io_out_2(c53_978_io_out_2)
  );
  C53 c53_979 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_979_io_in_0),
    .io_in_1(c53_979_io_in_1),
    .io_in_2(c53_979_io_in_2),
    .io_in_3(c53_979_io_in_3),
    .io_in_4(c53_979_io_in_4),
    .io_out_0(c53_979_io_out_0),
    .io_out_1(c53_979_io_out_1),
    .io_out_2(c53_979_io_out_2)
  );
  C53 c53_980 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_980_io_in_0),
    .io_in_1(c53_980_io_in_1),
    .io_in_2(c53_980_io_in_2),
    .io_in_3(c53_980_io_in_3),
    .io_in_4(c53_980_io_in_4),
    .io_out_0(c53_980_io_out_0),
    .io_out_1(c53_980_io_out_1),
    .io_out_2(c53_980_io_out_2)
  );
  C53 c53_981 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_981_io_in_0),
    .io_in_1(c53_981_io_in_1),
    .io_in_2(c53_981_io_in_2),
    .io_in_3(c53_981_io_in_3),
    .io_in_4(c53_981_io_in_4),
    .io_out_0(c53_981_io_out_0),
    .io_out_1(c53_981_io_out_1),
    .io_out_2(c53_981_io_out_2)
  );
  C53 c53_982 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_982_io_in_0),
    .io_in_1(c53_982_io_in_1),
    .io_in_2(c53_982_io_in_2),
    .io_in_3(c53_982_io_in_3),
    .io_in_4(c53_982_io_in_4),
    .io_out_0(c53_982_io_out_0),
    .io_out_1(c53_982_io_out_1),
    .io_out_2(c53_982_io_out_2)
  );
  C53 c53_983 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_983_io_in_0),
    .io_in_1(c53_983_io_in_1),
    .io_in_2(c53_983_io_in_2),
    .io_in_3(c53_983_io_in_3),
    .io_in_4(c53_983_io_in_4),
    .io_out_0(c53_983_io_out_0),
    .io_out_1(c53_983_io_out_1),
    .io_out_2(c53_983_io_out_2)
  );
  C53 c53_984 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_984_io_in_0),
    .io_in_1(c53_984_io_in_1),
    .io_in_2(c53_984_io_in_2),
    .io_in_3(c53_984_io_in_3),
    .io_in_4(c53_984_io_in_4),
    .io_out_0(c53_984_io_out_0),
    .io_out_1(c53_984_io_out_1),
    .io_out_2(c53_984_io_out_2)
  );
  C53 c53_985 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_985_io_in_0),
    .io_in_1(c53_985_io_in_1),
    .io_in_2(c53_985_io_in_2),
    .io_in_3(c53_985_io_in_3),
    .io_in_4(c53_985_io_in_4),
    .io_out_0(c53_985_io_out_0),
    .io_out_1(c53_985_io_out_1),
    .io_out_2(c53_985_io_out_2)
  );
  C53 c53_986 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_986_io_in_0),
    .io_in_1(c53_986_io_in_1),
    .io_in_2(c53_986_io_in_2),
    .io_in_3(c53_986_io_in_3),
    .io_in_4(c53_986_io_in_4),
    .io_out_0(c53_986_io_out_0),
    .io_out_1(c53_986_io_out_1),
    .io_out_2(c53_986_io_out_2)
  );
  C53 c53_987 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_987_io_in_0),
    .io_in_1(c53_987_io_in_1),
    .io_in_2(c53_987_io_in_2),
    .io_in_3(c53_987_io_in_3),
    .io_in_4(c53_987_io_in_4),
    .io_out_0(c53_987_io_out_0),
    .io_out_1(c53_987_io_out_1),
    .io_out_2(c53_987_io_out_2)
  );
  C53 c53_988 ( // @[Multiplier.scala 130:25]
    .io_in_0(c53_988_io_in_0),
    .io_in_1(c53_988_io_in_1),
    .io_in_2(c53_988_io_in_2),
    .io_in_3(c53_988_io_in_3),
    .io_in_4(c53_988_io_in_4),
    .io_out_0(c53_988_io_out_0),
    .io_out_1(c53_988_io_out_1),
    .io_out_2(c53_988_io_out_2)
  );
  C32 c32_69 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_69_io_in_0),
    .io_in_1(c32_69_io_in_1),
    .io_in_2(c32_69_io_in_2),
    .io_out_0(c32_69_io_out_0),
    .io_out_1(c32_69_io_out_1)
  );
  C22 c22_152 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_152_io_in_0),
    .io_in_1(c22_152_io_in_1),
    .io_out_0(c22_152_io_out_0),
    .io_out_1(c22_152_io_out_1)
  );
  C32 c32_70 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_70_io_in_0),
    .io_in_1(c32_70_io_in_1),
    .io_in_2(c32_70_io_in_2),
    .io_out_0(c32_70_io_out_0),
    .io_out_1(c32_70_io_out_1)
  );
  C22 c22_153 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_153_io_in_0),
    .io_in_1(c22_153_io_in_1),
    .io_out_0(c22_153_io_out_0),
    .io_out_1(c22_153_io_out_1)
  );
  C22 c22_154 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_154_io_in_0),
    .io_in_1(c22_154_io_in_1),
    .io_out_0(c22_154_io_out_0),
    .io_out_1(c22_154_io_out_1)
  );
  C22 c22_155 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_155_io_in_0),
    .io_in_1(c22_155_io_in_1),
    .io_out_0(c22_155_io_out_0),
    .io_out_1(c22_155_io_out_1)
  );
  C22 c22_156 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_156_io_in_0),
    .io_in_1(c22_156_io_in_1),
    .io_out_0(c22_156_io_out_0),
    .io_out_1(c22_156_io_out_1)
  );
  C32 c32_71 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_71_io_in_0),
    .io_in_1(c32_71_io_in_1),
    .io_in_2(c32_71_io_in_2),
    .io_out_0(c32_71_io_out_0),
    .io_out_1(c32_71_io_out_1)
  );
  C22 c22_157 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_157_io_in_0),
    .io_in_1(c22_157_io_in_1),
    .io_out_0(c22_157_io_out_0),
    .io_out_1(c22_157_io_out_1)
  );
  C22 c22_158 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_158_io_in_0),
    .io_in_1(c22_158_io_in_1),
    .io_out_0(c22_158_io_out_0),
    .io_out_1(c22_158_io_out_1)
  );
  C22 c22_159 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_159_io_in_0),
    .io_in_1(c22_159_io_in_1),
    .io_out_0(c22_159_io_out_0),
    .io_out_1(c22_159_io_out_1)
  );
  C22 c22_160 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_160_io_in_0),
    .io_in_1(c22_160_io_in_1),
    .io_out_0(c22_160_io_out_0),
    .io_out_1(c22_160_io_out_1)
  );
  C22 c22_161 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_161_io_in_0),
    .io_in_1(c22_161_io_in_1),
    .io_out_0(c22_161_io_out_0),
    .io_out_1(c22_161_io_out_1)
  );
  C22 c22_162 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_162_io_in_0),
    .io_in_1(c22_162_io_in_1),
    .io_out_0(c22_162_io_out_0),
    .io_out_1(c22_162_io_out_1)
  );
  C22 c22_163 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_163_io_in_0),
    .io_in_1(c22_163_io_in_1),
    .io_out_0(c22_163_io_out_0),
    .io_out_1(c22_163_io_out_1)
  );
  C22 c22_164 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_164_io_in_0),
    .io_in_1(c22_164_io_in_1),
    .io_out_0(c22_164_io_out_0),
    .io_out_1(c22_164_io_out_1)
  );
  C32 c32_72 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_72_io_in_0),
    .io_in_1(c32_72_io_in_1),
    .io_in_2(c32_72_io_in_2),
    .io_out_0(c32_72_io_out_0),
    .io_out_1(c32_72_io_out_1)
  );
  C22 c22_165 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_165_io_in_0),
    .io_in_1(c22_165_io_in_1),
    .io_out_0(c22_165_io_out_0),
    .io_out_1(c22_165_io_out_1)
  );
  C22 c22_166 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_166_io_in_0),
    .io_in_1(c22_166_io_in_1),
    .io_out_0(c22_166_io_out_0),
    .io_out_1(c22_166_io_out_1)
  );
  C22 c22_167 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_167_io_in_0),
    .io_in_1(c22_167_io_in_1),
    .io_out_0(c22_167_io_out_0),
    .io_out_1(c22_167_io_out_1)
  );
  C22 c22_168 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_168_io_in_0),
    .io_in_1(c22_168_io_in_1),
    .io_out_0(c22_168_io_out_0),
    .io_out_1(c22_168_io_out_1)
  );
  C22 c22_169 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_169_io_in_0),
    .io_in_1(c22_169_io_in_1),
    .io_out_0(c22_169_io_out_0),
    .io_out_1(c22_169_io_out_1)
  );
  C22 c22_170 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_170_io_in_0),
    .io_in_1(c22_170_io_in_1),
    .io_out_0(c22_170_io_out_0),
    .io_out_1(c22_170_io_out_1)
  );
  C22 c22_171 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_171_io_in_0),
    .io_in_1(c22_171_io_in_1),
    .io_out_0(c22_171_io_out_0),
    .io_out_1(c22_171_io_out_1)
  );
  C22 c22_172 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_172_io_in_0),
    .io_in_1(c22_172_io_in_1),
    .io_out_0(c22_172_io_out_0),
    .io_out_1(c22_172_io_out_1)
  );
  C22 c22_173 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_173_io_in_0),
    .io_in_1(c22_173_io_in_1),
    .io_out_0(c22_173_io_out_0),
    .io_out_1(c22_173_io_out_1)
  );
  C22 c22_174 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_174_io_in_0),
    .io_in_1(c22_174_io_in_1),
    .io_out_0(c22_174_io_out_0),
    .io_out_1(c22_174_io_out_1)
  );
  C22 c22_175 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_175_io_in_0),
    .io_in_1(c22_175_io_in_1),
    .io_out_0(c22_175_io_out_0),
    .io_out_1(c22_175_io_out_1)
  );
  C22 c22_176 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_176_io_in_0),
    .io_in_1(c22_176_io_in_1),
    .io_out_0(c22_176_io_out_0),
    .io_out_1(c22_176_io_out_1)
  );
  C22 c22_177 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_177_io_in_0),
    .io_in_1(c22_177_io_in_1),
    .io_out_0(c22_177_io_out_0),
    .io_out_1(c22_177_io_out_1)
  );
  C22 c22_178 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_178_io_in_0),
    .io_in_1(c22_178_io_in_1),
    .io_out_0(c22_178_io_out_0),
    .io_out_1(c22_178_io_out_1)
  );
  C22 c22_179 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_179_io_in_0),
    .io_in_1(c22_179_io_in_1),
    .io_out_0(c22_179_io_out_0),
    .io_out_1(c22_179_io_out_1)
  );
  C22 c22_180 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_180_io_in_0),
    .io_in_1(c22_180_io_in_1),
    .io_out_0(c22_180_io_out_0),
    .io_out_1(c22_180_io_out_1)
  );
  C22 c22_181 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_181_io_in_0),
    .io_in_1(c22_181_io_in_1),
    .io_out_0(c22_181_io_out_0),
    .io_out_1(c22_181_io_out_1)
  );
  C22 c22_182 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_182_io_in_0),
    .io_in_1(c22_182_io_in_1),
    .io_out_0(c22_182_io_out_0),
    .io_out_1(c22_182_io_out_1)
  );
  C22 c22_183 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_183_io_in_0),
    .io_in_1(c22_183_io_in_1),
    .io_out_0(c22_183_io_out_0),
    .io_out_1(c22_183_io_out_1)
  );
  C22 c22_184 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_184_io_in_0),
    .io_in_1(c22_184_io_in_1),
    .io_out_0(c22_184_io_out_0),
    .io_out_1(c22_184_io_out_1)
  );
  C22 c22_185 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_185_io_in_0),
    .io_in_1(c22_185_io_in_1),
    .io_out_0(c22_185_io_out_0),
    .io_out_1(c22_185_io_out_1)
  );
  C22 c22_186 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_186_io_in_0),
    .io_in_1(c22_186_io_in_1),
    .io_out_0(c22_186_io_out_0),
    .io_out_1(c22_186_io_out_1)
  );
  C22 c22_187 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_187_io_in_0),
    .io_in_1(c22_187_io_in_1),
    .io_out_0(c22_187_io_out_0),
    .io_out_1(c22_187_io_out_1)
  );
  C22 c22_188 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_188_io_in_0),
    .io_in_1(c22_188_io_in_1),
    .io_out_0(c22_188_io_out_0),
    .io_out_1(c22_188_io_out_1)
  );
  C22 c22_189 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_189_io_in_0),
    .io_in_1(c22_189_io_in_1),
    .io_out_0(c22_189_io_out_0),
    .io_out_1(c22_189_io_out_1)
  );
  C22 c22_190 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_190_io_in_0),
    .io_in_1(c22_190_io_in_1),
    .io_out_0(c22_190_io_out_0),
    .io_out_1(c22_190_io_out_1)
  );
  C22 c22_191 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_191_io_in_0),
    .io_in_1(c22_191_io_in_1),
    .io_out_0(c22_191_io_out_0),
    .io_out_1(c22_191_io_out_1)
  );
  C22 c22_192 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_192_io_in_0),
    .io_in_1(c22_192_io_in_1),
    .io_out_0(c22_192_io_out_0),
    .io_out_1(c22_192_io_out_1)
  );
  C22 c22_193 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_193_io_in_0),
    .io_in_1(c22_193_io_in_1),
    .io_out_0(c22_193_io_out_0),
    .io_out_1(c22_193_io_out_1)
  );
  C22 c22_194 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_194_io_in_0),
    .io_in_1(c22_194_io_in_1),
    .io_out_0(c22_194_io_out_0),
    .io_out_1(c22_194_io_out_1)
  );
  C22 c22_195 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_195_io_in_0),
    .io_in_1(c22_195_io_in_1),
    .io_out_0(c22_195_io_out_0),
    .io_out_1(c22_195_io_out_1)
  );
  C22 c22_196 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_196_io_in_0),
    .io_in_1(c22_196_io_in_1),
    .io_out_0(c22_196_io_out_0),
    .io_out_1(c22_196_io_out_1)
  );
  C22 c22_197 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_197_io_in_0),
    .io_in_1(c22_197_io_in_1),
    .io_out_0(c22_197_io_out_0),
    .io_out_1(c22_197_io_out_1)
  );
  C22 c22_198 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_198_io_in_0),
    .io_in_1(c22_198_io_in_1),
    .io_out_0(c22_198_io_out_0),
    .io_out_1(c22_198_io_out_1)
  );
  C22 c22_199 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_199_io_in_0),
    .io_in_1(c22_199_io_in_1),
    .io_out_0(c22_199_io_out_0),
    .io_out_1(c22_199_io_out_1)
  );
  C22 c22_200 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_200_io_in_0),
    .io_in_1(c22_200_io_in_1),
    .io_out_0(c22_200_io_out_0),
    .io_out_1(c22_200_io_out_1)
  );
  C22 c22_201 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_201_io_in_0),
    .io_in_1(c22_201_io_in_1),
    .io_out_0(c22_201_io_out_0),
    .io_out_1(c22_201_io_out_1)
  );
  C22 c22_202 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_202_io_in_0),
    .io_in_1(c22_202_io_in_1),
    .io_out_0(c22_202_io_out_0),
    .io_out_1(c22_202_io_out_1)
  );
  C22 c22_203 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_203_io_in_0),
    .io_in_1(c22_203_io_in_1),
    .io_out_0(c22_203_io_out_0),
    .io_out_1(c22_203_io_out_1)
  );
  C22 c22_204 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_204_io_in_0),
    .io_in_1(c22_204_io_in_1),
    .io_out_0(c22_204_io_out_0),
    .io_out_1(c22_204_io_out_1)
  );
  C22 c22_205 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_205_io_in_0),
    .io_in_1(c22_205_io_in_1),
    .io_out_0(c22_205_io_out_0),
    .io_out_1(c22_205_io_out_1)
  );
  C22 c22_206 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_206_io_in_0),
    .io_in_1(c22_206_io_in_1),
    .io_out_0(c22_206_io_out_0),
    .io_out_1(c22_206_io_out_1)
  );
  C22 c22_207 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_207_io_in_0),
    .io_in_1(c22_207_io_in_1),
    .io_out_0(c22_207_io_out_0),
    .io_out_1(c22_207_io_out_1)
  );
  C22 c22_208 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_208_io_in_0),
    .io_in_1(c22_208_io_in_1),
    .io_out_0(c22_208_io_out_0),
    .io_out_1(c22_208_io_out_1)
  );
  C22 c22_209 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_209_io_in_0),
    .io_in_1(c22_209_io_in_1),
    .io_out_0(c22_209_io_out_0),
    .io_out_1(c22_209_io_out_1)
  );
  C22 c22_210 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_210_io_in_0),
    .io_in_1(c22_210_io_in_1),
    .io_out_0(c22_210_io_out_0),
    .io_out_1(c22_210_io_out_1)
  );
  C22 c22_211 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_211_io_in_0),
    .io_in_1(c22_211_io_in_1),
    .io_out_0(c22_211_io_out_0),
    .io_out_1(c22_211_io_out_1)
  );
  C22 c22_212 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_212_io_in_0),
    .io_in_1(c22_212_io_in_1),
    .io_out_0(c22_212_io_out_0),
    .io_out_1(c22_212_io_out_1)
  );
  C22 c22_213 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_213_io_in_0),
    .io_in_1(c22_213_io_in_1),
    .io_out_0(c22_213_io_out_0),
    .io_out_1(c22_213_io_out_1)
  );
  C22 c22_214 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_214_io_in_0),
    .io_in_1(c22_214_io_in_1),
    .io_out_0(c22_214_io_out_0),
    .io_out_1(c22_214_io_out_1)
  );
  C22 c22_215 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_215_io_in_0),
    .io_in_1(c22_215_io_in_1),
    .io_out_0(c22_215_io_out_0),
    .io_out_1(c22_215_io_out_1)
  );
  C22 c22_216 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_216_io_in_0),
    .io_in_1(c22_216_io_in_1),
    .io_out_0(c22_216_io_out_0),
    .io_out_1(c22_216_io_out_1)
  );
  C22 c22_217 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_217_io_in_0),
    .io_in_1(c22_217_io_in_1),
    .io_out_0(c22_217_io_out_0),
    .io_out_1(c22_217_io_out_1)
  );
  C22 c22_218 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_218_io_in_0),
    .io_in_1(c22_218_io_in_1),
    .io_out_0(c22_218_io_out_0),
    .io_out_1(c22_218_io_out_1)
  );
  C22 c22_219 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_219_io_in_0),
    .io_in_1(c22_219_io_in_1),
    .io_out_0(c22_219_io_out_0),
    .io_out_1(c22_219_io_out_1)
  );
  C22 c22_220 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_220_io_in_0),
    .io_in_1(c22_220_io_in_1),
    .io_out_0(c22_220_io_out_0),
    .io_out_1(c22_220_io_out_1)
  );
  C22 c22_221 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_221_io_in_0),
    .io_in_1(c22_221_io_in_1),
    .io_out_0(c22_221_io_out_0),
    .io_out_1(c22_221_io_out_1)
  );
  C22 c22_222 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_222_io_in_0),
    .io_in_1(c22_222_io_in_1),
    .io_out_0(c22_222_io_out_0),
    .io_out_1(c22_222_io_out_1)
  );
  C22 c22_223 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_223_io_in_0),
    .io_in_1(c22_223_io_in_1),
    .io_out_0(c22_223_io_out_0),
    .io_out_1(c22_223_io_out_1)
  );
  C22 c22_224 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_224_io_in_0),
    .io_in_1(c22_224_io_in_1),
    .io_out_0(c22_224_io_out_0),
    .io_out_1(c22_224_io_out_1)
  );
  C22 c22_225 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_225_io_in_0),
    .io_in_1(c22_225_io_in_1),
    .io_out_0(c22_225_io_out_0),
    .io_out_1(c22_225_io_out_1)
  );
  C22 c22_226 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_226_io_in_0),
    .io_in_1(c22_226_io_in_1),
    .io_out_0(c22_226_io_out_0),
    .io_out_1(c22_226_io_out_1)
  );
  C22 c22_227 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_227_io_in_0),
    .io_in_1(c22_227_io_in_1),
    .io_out_0(c22_227_io_out_0),
    .io_out_1(c22_227_io_out_1)
  );
  C22 c22_228 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_228_io_in_0),
    .io_in_1(c22_228_io_in_1),
    .io_out_0(c22_228_io_out_0),
    .io_out_1(c22_228_io_out_1)
  );
  C22 c22_229 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_229_io_in_0),
    .io_in_1(c22_229_io_in_1),
    .io_out_0(c22_229_io_out_0),
    .io_out_1(c22_229_io_out_1)
  );
  C22 c22_230 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_230_io_in_0),
    .io_in_1(c22_230_io_in_1),
    .io_out_0(c22_230_io_out_0),
    .io_out_1(c22_230_io_out_1)
  );
  C22 c22_231 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_231_io_in_0),
    .io_in_1(c22_231_io_in_1),
    .io_out_0(c22_231_io_out_0),
    .io_out_1(c22_231_io_out_1)
  );
  C22 c22_232 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_232_io_in_0),
    .io_in_1(c22_232_io_in_1),
    .io_out_0(c22_232_io_out_0),
    .io_out_1(c22_232_io_out_1)
  );
  C22 c22_233 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_233_io_in_0),
    .io_in_1(c22_233_io_in_1),
    .io_out_0(c22_233_io_out_0),
    .io_out_1(c22_233_io_out_1)
  );
  C22 c22_234 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_234_io_in_0),
    .io_in_1(c22_234_io_in_1),
    .io_out_0(c22_234_io_out_0),
    .io_out_1(c22_234_io_out_1)
  );
  C22 c22_235 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_235_io_in_0),
    .io_in_1(c22_235_io_in_1),
    .io_out_0(c22_235_io_out_0),
    .io_out_1(c22_235_io_out_1)
  );
  C32 c32_73 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_73_io_in_0),
    .io_in_1(c32_73_io_in_1),
    .io_in_2(c32_73_io_in_2),
    .io_out_0(c32_73_io_out_0),
    .io_out_1(c32_73_io_out_1)
  );
  C32 c32_74 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_74_io_in_0),
    .io_in_1(c32_74_io_in_1),
    .io_in_2(c32_74_io_in_2),
    .io_out_0(c32_74_io_out_0),
    .io_out_1(c32_74_io_out_1)
  );
  C32 c32_75 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_75_io_in_0),
    .io_in_1(c32_75_io_in_1),
    .io_in_2(c32_75_io_in_2),
    .io_out_0(c32_75_io_out_0),
    .io_out_1(c32_75_io_out_1)
  );
  C32 c32_76 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_76_io_in_0),
    .io_in_1(c32_76_io_in_1),
    .io_in_2(c32_76_io_in_2),
    .io_out_0(c32_76_io_out_0),
    .io_out_1(c32_76_io_out_1)
  );
  C32 c32_77 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_77_io_in_0),
    .io_in_1(c32_77_io_in_1),
    .io_in_2(c32_77_io_in_2),
    .io_out_0(c32_77_io_out_0),
    .io_out_1(c32_77_io_out_1)
  );
  C32 c32_78 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_78_io_in_0),
    .io_in_1(c32_78_io_in_1),
    .io_in_2(c32_78_io_in_2),
    .io_out_0(c32_78_io_out_0),
    .io_out_1(c32_78_io_out_1)
  );
  C32 c32_79 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_79_io_in_0),
    .io_in_1(c32_79_io_in_1),
    .io_in_2(c32_79_io_in_2),
    .io_out_0(c32_79_io_out_0),
    .io_out_1(c32_79_io_out_1)
  );
  C22 c22_236 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_236_io_in_0),
    .io_in_1(c22_236_io_in_1),
    .io_out_0(c22_236_io_out_0),
    .io_out_1(c22_236_io_out_1)
  );
  C32 c32_80 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_80_io_in_0),
    .io_in_1(c32_80_io_in_1),
    .io_in_2(c32_80_io_in_2),
    .io_out_0(c32_80_io_out_0),
    .io_out_1(c32_80_io_out_1)
  );
  C22 c22_237 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_237_io_in_0),
    .io_in_1(c22_237_io_in_1),
    .io_out_0(c22_237_io_out_0),
    .io_out_1(c22_237_io_out_1)
  );
  C22 c22_238 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_238_io_in_0),
    .io_in_1(c22_238_io_in_1),
    .io_out_0(c22_238_io_out_0),
    .io_out_1(c22_238_io_out_1)
  );
  C22 c22_239 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_239_io_in_0),
    .io_in_1(c22_239_io_in_1),
    .io_out_0(c22_239_io_out_0),
    .io_out_1(c22_239_io_out_1)
  );
  C22 c22_240 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_240_io_in_0),
    .io_in_1(c22_240_io_in_1),
    .io_out_0(c22_240_io_out_0),
    .io_out_1(c22_240_io_out_1)
  );
  C32 c32_81 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_81_io_in_0),
    .io_in_1(c32_81_io_in_1),
    .io_in_2(c32_81_io_in_2),
    .io_out_0(c32_81_io_out_0),
    .io_out_1(c32_81_io_out_1)
  );
  C22 c22_241 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_241_io_in_0),
    .io_in_1(c22_241_io_in_1),
    .io_out_0(c22_241_io_out_0),
    .io_out_1(c22_241_io_out_1)
  );
  C22 c22_242 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_242_io_in_0),
    .io_in_1(c22_242_io_in_1),
    .io_out_0(c22_242_io_out_0),
    .io_out_1(c22_242_io_out_1)
  );
  C22 c22_243 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_243_io_in_0),
    .io_in_1(c22_243_io_in_1),
    .io_out_0(c22_243_io_out_0),
    .io_out_1(c22_243_io_out_1)
  );
  C22 c22_244 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_244_io_in_0),
    .io_in_1(c22_244_io_in_1),
    .io_out_0(c22_244_io_out_0),
    .io_out_1(c22_244_io_out_1)
  );
  C22 c22_245 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_245_io_in_0),
    .io_in_1(c22_245_io_in_1),
    .io_out_0(c22_245_io_out_0),
    .io_out_1(c22_245_io_out_1)
  );
  C22 c22_246 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_246_io_in_0),
    .io_in_1(c22_246_io_in_1),
    .io_out_0(c22_246_io_out_0),
    .io_out_1(c22_246_io_out_1)
  );
  C22 c22_247 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_247_io_in_0),
    .io_in_1(c22_247_io_in_1),
    .io_out_0(c22_247_io_out_0),
    .io_out_1(c22_247_io_out_1)
  );
  C22 c22_248 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_248_io_in_0),
    .io_in_1(c22_248_io_in_1),
    .io_out_0(c22_248_io_out_0),
    .io_out_1(c22_248_io_out_1)
  );
  C32 c32_82 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_82_io_in_0),
    .io_in_1(c32_82_io_in_1),
    .io_in_2(c32_82_io_in_2),
    .io_out_0(c32_82_io_out_0),
    .io_out_1(c32_82_io_out_1)
  );
  C22 c22_249 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_249_io_in_0),
    .io_in_1(c22_249_io_in_1),
    .io_out_0(c22_249_io_out_0),
    .io_out_1(c22_249_io_out_1)
  );
  C22 c22_250 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_250_io_in_0),
    .io_in_1(c22_250_io_in_1),
    .io_out_0(c22_250_io_out_0),
    .io_out_1(c22_250_io_out_1)
  );
  C22 c22_251 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_251_io_in_0),
    .io_in_1(c22_251_io_in_1),
    .io_out_0(c22_251_io_out_0),
    .io_out_1(c22_251_io_out_1)
  );
  C22 c22_252 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_252_io_in_0),
    .io_in_1(c22_252_io_in_1),
    .io_out_0(c22_252_io_out_0),
    .io_out_1(c22_252_io_out_1)
  );
  C22 c22_253 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_253_io_in_0),
    .io_in_1(c22_253_io_in_1),
    .io_out_0(c22_253_io_out_0),
    .io_out_1(c22_253_io_out_1)
  );
  C22 c22_254 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_254_io_in_0),
    .io_in_1(c22_254_io_in_1),
    .io_out_0(c22_254_io_out_0),
    .io_out_1(c22_254_io_out_1)
  );
  C22 c22_255 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_255_io_in_0),
    .io_in_1(c22_255_io_in_1),
    .io_out_0(c22_255_io_out_0),
    .io_out_1(c22_255_io_out_1)
  );
  C22 c22_256 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_256_io_in_0),
    .io_in_1(c22_256_io_in_1),
    .io_out_0(c22_256_io_out_0),
    .io_out_1(c22_256_io_out_1)
  );
  C22 c22_257 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_257_io_in_0),
    .io_in_1(c22_257_io_in_1),
    .io_out_0(c22_257_io_out_0),
    .io_out_1(c22_257_io_out_1)
  );
  C22 c22_258 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_258_io_in_0),
    .io_in_1(c22_258_io_in_1),
    .io_out_0(c22_258_io_out_0),
    .io_out_1(c22_258_io_out_1)
  );
  C22 c22_259 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_259_io_in_0),
    .io_in_1(c22_259_io_in_1),
    .io_out_0(c22_259_io_out_0),
    .io_out_1(c22_259_io_out_1)
  );
  C22 c22_260 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_260_io_in_0),
    .io_in_1(c22_260_io_in_1),
    .io_out_0(c22_260_io_out_0),
    .io_out_1(c22_260_io_out_1)
  );
  C22 c22_261 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_261_io_in_0),
    .io_in_1(c22_261_io_in_1),
    .io_out_0(c22_261_io_out_0),
    .io_out_1(c22_261_io_out_1)
  );
  C22 c22_262 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_262_io_in_0),
    .io_in_1(c22_262_io_in_1),
    .io_out_0(c22_262_io_out_0),
    .io_out_1(c22_262_io_out_1)
  );
  C22 c22_263 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_263_io_in_0),
    .io_in_1(c22_263_io_in_1),
    .io_out_0(c22_263_io_out_0),
    .io_out_1(c22_263_io_out_1)
  );
  C32 c32_83 ( // @[Multiplier.scala 125:25]
    .io_in_0(c32_83_io_in_0),
    .io_in_1(c32_83_io_in_1),
    .io_in_2(c32_83_io_in_2),
    .io_out_0(c32_83_io_out_0),
    .io_out_1(c32_83_io_out_1)
  );
  C22 c22_264 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_264_io_in_0),
    .io_in_1(c22_264_io_in_1),
    .io_out_0(c22_264_io_out_0),
    .io_out_1(c22_264_io_out_1)
  );
  C22 c22_265 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_265_io_in_0),
    .io_in_1(c22_265_io_in_1),
    .io_out_0(c22_265_io_out_0),
    .io_out_1(c22_265_io_out_1)
  );
  C22 c22_266 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_266_io_in_0),
    .io_in_1(c22_266_io_in_1),
    .io_out_0(c22_266_io_out_0),
    .io_out_1(c22_266_io_out_1)
  );
  C22 c22_267 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_267_io_in_0),
    .io_in_1(c22_267_io_in_1),
    .io_out_0(c22_267_io_out_0),
    .io_out_1(c22_267_io_out_1)
  );
  C22 c22_268 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_268_io_in_0),
    .io_in_1(c22_268_io_in_1),
    .io_out_0(c22_268_io_out_0),
    .io_out_1(c22_268_io_out_1)
  );
  C22 c22_269 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_269_io_in_0),
    .io_in_1(c22_269_io_in_1),
    .io_out_0(c22_269_io_out_0),
    .io_out_1(c22_269_io_out_1)
  );
  C22 c22_270 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_270_io_in_0),
    .io_in_1(c22_270_io_in_1),
    .io_out_0(c22_270_io_out_0),
    .io_out_1(c22_270_io_out_1)
  );
  C22 c22_271 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_271_io_in_0),
    .io_in_1(c22_271_io_in_1),
    .io_out_0(c22_271_io_out_0),
    .io_out_1(c22_271_io_out_1)
  );
  C22 c22_272 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_272_io_in_0),
    .io_in_1(c22_272_io_in_1),
    .io_out_0(c22_272_io_out_0),
    .io_out_1(c22_272_io_out_1)
  );
  C22 c22_273 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_273_io_in_0),
    .io_in_1(c22_273_io_in_1),
    .io_out_0(c22_273_io_out_0),
    .io_out_1(c22_273_io_out_1)
  );
  C22 c22_274 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_274_io_in_0),
    .io_in_1(c22_274_io_in_1),
    .io_out_0(c22_274_io_out_0),
    .io_out_1(c22_274_io_out_1)
  );
  C22 c22_275 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_275_io_in_0),
    .io_in_1(c22_275_io_in_1),
    .io_out_0(c22_275_io_out_0),
    .io_out_1(c22_275_io_out_1)
  );
  C22 c22_276 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_276_io_in_0),
    .io_in_1(c22_276_io_in_1),
    .io_out_0(c22_276_io_out_0),
    .io_out_1(c22_276_io_out_1)
  );
  C22 c22_277 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_277_io_in_0),
    .io_in_1(c22_277_io_in_1),
    .io_out_0(c22_277_io_out_0),
    .io_out_1(c22_277_io_out_1)
  );
  C22 c22_278 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_278_io_in_0),
    .io_in_1(c22_278_io_in_1),
    .io_out_0(c22_278_io_out_0),
    .io_out_1(c22_278_io_out_1)
  );
  C22 c22_279 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_279_io_in_0),
    .io_in_1(c22_279_io_in_1),
    .io_out_0(c22_279_io_out_0),
    .io_out_1(c22_279_io_out_1)
  );
  C22 c22_280 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_280_io_in_0),
    .io_in_1(c22_280_io_in_1),
    .io_out_0(c22_280_io_out_0),
    .io_out_1(c22_280_io_out_1)
  );
  C22 c22_281 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_281_io_in_0),
    .io_in_1(c22_281_io_in_1),
    .io_out_0(c22_281_io_out_0),
    .io_out_1(c22_281_io_out_1)
  );
  C22 c22_282 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_282_io_in_0),
    .io_in_1(c22_282_io_in_1),
    .io_out_0(c22_282_io_out_0),
    .io_out_1(c22_282_io_out_1)
  );
  C22 c22_283 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_283_io_in_0),
    .io_in_1(c22_283_io_in_1),
    .io_out_0(c22_283_io_out_0),
    .io_out_1(c22_283_io_out_1)
  );
  C22 c22_284 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_284_io_in_0),
    .io_in_1(c22_284_io_in_1),
    .io_out_0(c22_284_io_out_0),
    .io_out_1(c22_284_io_out_1)
  );
  C22 c22_285 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_285_io_in_0),
    .io_in_1(c22_285_io_in_1),
    .io_out_0(c22_285_io_out_0),
    .io_out_1(c22_285_io_out_1)
  );
  C22 c22_286 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_286_io_in_0),
    .io_in_1(c22_286_io_in_1),
    .io_out_0(c22_286_io_out_0),
    .io_out_1(c22_286_io_out_1)
  );
  C22 c22_287 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_287_io_in_0),
    .io_in_1(c22_287_io_in_1),
    .io_out_0(c22_287_io_out_0),
    .io_out_1(c22_287_io_out_1)
  );
  C22 c22_288 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_288_io_in_0),
    .io_in_1(c22_288_io_in_1),
    .io_out_0(c22_288_io_out_0),
    .io_out_1(c22_288_io_out_1)
  );
  C22 c22_289 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_289_io_in_0),
    .io_in_1(c22_289_io_in_1),
    .io_out_0(c22_289_io_out_0),
    .io_out_1(c22_289_io_out_1)
  );
  C22 c22_290 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_290_io_in_0),
    .io_in_1(c22_290_io_in_1),
    .io_out_0(c22_290_io_out_0),
    .io_out_1(c22_290_io_out_1)
  );
  C22 c22_291 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_291_io_in_0),
    .io_in_1(c22_291_io_in_1),
    .io_out_0(c22_291_io_out_0),
    .io_out_1(c22_291_io_out_1)
  );
  C22 c22_292 ( // @[Multiplier.scala 120:25]
    .io_in_0(c22_292_io_in_0),
    .io_in_1(c22_292_io_in_1),
    .io_out_0(c22_292_io_out_0),
    .io_out_1(c22_292_io_out_1)
  );
  assign io_result = sum + carry_1; // @[Multiplier.scala 181:20]
  assign c22_io_in_0 = r; // @[Multiplier.scala 121:19]
  assign c22_io_in_1 = r_1; // @[Multiplier.scala 121:19]
  assign c22_1_io_in_0 = r_2; // @[Multiplier.scala 121:19]
  assign c22_1_io_in_1 = r_3; // @[Multiplier.scala 121:19]
  assign c32_io_in_0 = r_4; // @[Multiplier.scala 126:19]
  assign c32_io_in_1 = r_5; // @[Multiplier.scala 126:19]
  assign c32_io_in_2 = r_6; // @[Multiplier.scala 126:19]
  assign c32_1_io_in_0 = r_7; // @[Multiplier.scala 126:19]
  assign c32_1_io_in_1 = r_8; // @[Multiplier.scala 126:19]
  assign c32_1_io_in_2 = r_9; // @[Multiplier.scala 126:19]
  assign c53_io_in_0 = r_10; // @[Multiplier.scala 132:13]
  assign c53_io_in_1 = r_11; // @[Multiplier.scala 132:13]
  assign c53_io_in_2 = r_12; // @[Multiplier.scala 132:13]
  assign c53_io_in_3 = r_13; // @[Multiplier.scala 132:13]
  assign c53_io_in_4 = 1'h0; // @[Multiplier.scala 134:24]
  assign c53_1_io_in_0 = r_14; // @[Multiplier.scala 132:13]
  assign c53_1_io_in_1 = r_15; // @[Multiplier.scala 132:13]
  assign c53_1_io_in_2 = r_16; // @[Multiplier.scala 132:13]
  assign c53_1_io_in_3 = r_17; // @[Multiplier.scala 132:13]
  assign c53_1_io_in_4 = c53_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_2_io_in_0 = r_18; // @[Multiplier.scala 132:13]
  assign c53_2_io_in_1 = r_19; // @[Multiplier.scala 132:13]
  assign c53_2_io_in_2 = r_20; // @[Multiplier.scala 132:13]
  assign c53_2_io_in_3 = r_21; // @[Multiplier.scala 132:13]
  assign c53_2_io_in_4 = c53_1_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_3_io_in_0 = r_23; // @[Multiplier.scala 132:13]
  assign c53_3_io_in_1 = r_24; // @[Multiplier.scala 132:13]
  assign c53_3_io_in_2 = r_25; // @[Multiplier.scala 132:13]
  assign c53_3_io_in_3 = r_26; // @[Multiplier.scala 132:13]
  assign c53_3_io_in_4 = c53_2_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_4_io_in_0 = r_28; // @[Multiplier.scala 132:13]
  assign c53_4_io_in_1 = r_29; // @[Multiplier.scala 132:13]
  assign c53_4_io_in_2 = r_30; // @[Multiplier.scala 132:13]
  assign c53_4_io_in_3 = r_31; // @[Multiplier.scala 132:13]
  assign c53_4_io_in_4 = c53_3_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_2_io_in_0 = r_32; // @[Multiplier.scala 121:19]
  assign c22_2_io_in_1 = r_33; // @[Multiplier.scala 121:19]
  assign c53_5_io_in_0 = r_34; // @[Multiplier.scala 132:13]
  assign c53_5_io_in_1 = r_35; // @[Multiplier.scala 132:13]
  assign c53_5_io_in_2 = r_36; // @[Multiplier.scala 132:13]
  assign c53_5_io_in_3 = r_37; // @[Multiplier.scala 132:13]
  assign c53_5_io_in_4 = c53_4_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_3_io_in_0 = r_38; // @[Multiplier.scala 121:19]
  assign c22_3_io_in_1 = r_39; // @[Multiplier.scala 121:19]
  assign c53_6_io_in_0 = r_40; // @[Multiplier.scala 132:13]
  assign c53_6_io_in_1 = r_41; // @[Multiplier.scala 132:13]
  assign c53_6_io_in_2 = r_42; // @[Multiplier.scala 132:13]
  assign c53_6_io_in_3 = r_43; // @[Multiplier.scala 132:13]
  assign c53_6_io_in_4 = c53_5_io_out_1; // @[Multiplier.scala 136:41]
  assign c32_2_io_in_0 = r_44; // @[Multiplier.scala 126:19]
  assign c32_2_io_in_1 = r_45; // @[Multiplier.scala 126:19]
  assign c32_2_io_in_2 = r_46; // @[Multiplier.scala 126:19]
  assign c53_7_io_in_0 = r_47; // @[Multiplier.scala 132:13]
  assign c53_7_io_in_1 = r_48; // @[Multiplier.scala 132:13]
  assign c53_7_io_in_2 = r_49; // @[Multiplier.scala 132:13]
  assign c53_7_io_in_3 = r_50; // @[Multiplier.scala 132:13]
  assign c53_7_io_in_4 = c53_6_io_out_1; // @[Multiplier.scala 136:41]
  assign c32_3_io_in_0 = r_51; // @[Multiplier.scala 126:19]
  assign c32_3_io_in_1 = r_52; // @[Multiplier.scala 126:19]
  assign c32_3_io_in_2 = r_53; // @[Multiplier.scala 126:19]
  assign c53_8_io_in_0 = r_54; // @[Multiplier.scala 132:13]
  assign c53_8_io_in_1 = r_55; // @[Multiplier.scala 132:13]
  assign c53_8_io_in_2 = r_56; // @[Multiplier.scala 132:13]
  assign c53_8_io_in_3 = r_57; // @[Multiplier.scala 132:13]
  assign c53_8_io_in_4 = c53_7_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_9_io_in_0 = r_58; // @[Multiplier.scala 132:13]
  assign c53_9_io_in_1 = r_59; // @[Multiplier.scala 132:13]
  assign c53_9_io_in_2 = r_60; // @[Multiplier.scala 132:13]
  assign c53_9_io_in_3 = r_61; // @[Multiplier.scala 132:13]
  assign c53_9_io_in_4 = 1'h0; // @[Multiplier.scala 134:24]
  assign c53_10_io_in_0 = r_62; // @[Multiplier.scala 132:13]
  assign c53_10_io_in_1 = r_63; // @[Multiplier.scala 132:13]
  assign c53_10_io_in_2 = r_64; // @[Multiplier.scala 132:13]
  assign c53_10_io_in_3 = r_65; // @[Multiplier.scala 132:13]
  assign c53_10_io_in_4 = c53_8_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_11_io_in_0 = r_66; // @[Multiplier.scala 132:13]
  assign c53_11_io_in_1 = r_67; // @[Multiplier.scala 132:13]
  assign c53_11_io_in_2 = r_68; // @[Multiplier.scala 132:13]
  assign c53_11_io_in_3 = r_69; // @[Multiplier.scala 132:13]
  assign c53_11_io_in_4 = c53_9_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_12_io_in_0 = r_70; // @[Multiplier.scala 132:13]
  assign c53_12_io_in_1 = r_71; // @[Multiplier.scala 132:13]
  assign c53_12_io_in_2 = r_72; // @[Multiplier.scala 132:13]
  assign c53_12_io_in_3 = r_73; // @[Multiplier.scala 132:13]
  assign c53_12_io_in_4 = c53_10_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_13_io_in_0 = r_74; // @[Multiplier.scala 132:13]
  assign c53_13_io_in_1 = r_75; // @[Multiplier.scala 132:13]
  assign c53_13_io_in_2 = r_76; // @[Multiplier.scala 132:13]
  assign c53_13_io_in_3 = r_77; // @[Multiplier.scala 132:13]
  assign c53_13_io_in_4 = c53_11_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_14_io_in_0 = r_79; // @[Multiplier.scala 132:13]
  assign c53_14_io_in_1 = r_80; // @[Multiplier.scala 132:13]
  assign c53_14_io_in_2 = r_81; // @[Multiplier.scala 132:13]
  assign c53_14_io_in_3 = r_82; // @[Multiplier.scala 132:13]
  assign c53_14_io_in_4 = c53_12_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_15_io_in_0 = r_83; // @[Multiplier.scala 132:13]
  assign c53_15_io_in_1 = r_84; // @[Multiplier.scala 132:13]
  assign c53_15_io_in_2 = r_85; // @[Multiplier.scala 132:13]
  assign c53_15_io_in_3 = r_86; // @[Multiplier.scala 132:13]
  assign c53_15_io_in_4 = c53_13_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_16_io_in_0 = r_88; // @[Multiplier.scala 132:13]
  assign c53_16_io_in_1 = r_89; // @[Multiplier.scala 132:13]
  assign c53_16_io_in_2 = r_90; // @[Multiplier.scala 132:13]
  assign c53_16_io_in_3 = r_91; // @[Multiplier.scala 132:13]
  assign c53_16_io_in_4 = c53_14_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_17_io_in_0 = r_92; // @[Multiplier.scala 132:13]
  assign c53_17_io_in_1 = r_93; // @[Multiplier.scala 132:13]
  assign c53_17_io_in_2 = r_94; // @[Multiplier.scala 132:13]
  assign c53_17_io_in_3 = r_95; // @[Multiplier.scala 132:13]
  assign c53_17_io_in_4 = c53_15_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_4_io_in_0 = r_96; // @[Multiplier.scala 121:19]
  assign c22_4_io_in_1 = r_97; // @[Multiplier.scala 121:19]
  assign c53_18_io_in_0 = r_98; // @[Multiplier.scala 132:13]
  assign c53_18_io_in_1 = r_99; // @[Multiplier.scala 132:13]
  assign c53_18_io_in_2 = r_100; // @[Multiplier.scala 132:13]
  assign c53_18_io_in_3 = r_101; // @[Multiplier.scala 132:13]
  assign c53_18_io_in_4 = c53_16_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_19_io_in_0 = r_102; // @[Multiplier.scala 132:13]
  assign c53_19_io_in_1 = r_103; // @[Multiplier.scala 132:13]
  assign c53_19_io_in_2 = r_104; // @[Multiplier.scala 132:13]
  assign c53_19_io_in_3 = r_105; // @[Multiplier.scala 132:13]
  assign c53_19_io_in_4 = c53_17_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_5_io_in_0 = r_106; // @[Multiplier.scala 121:19]
  assign c22_5_io_in_1 = r_107; // @[Multiplier.scala 121:19]
  assign c53_20_io_in_0 = r_108; // @[Multiplier.scala 132:13]
  assign c53_20_io_in_1 = r_109; // @[Multiplier.scala 132:13]
  assign c53_20_io_in_2 = r_110; // @[Multiplier.scala 132:13]
  assign c53_20_io_in_3 = r_111; // @[Multiplier.scala 132:13]
  assign c53_20_io_in_4 = c53_18_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_21_io_in_0 = r_112; // @[Multiplier.scala 132:13]
  assign c53_21_io_in_1 = r_113; // @[Multiplier.scala 132:13]
  assign c53_21_io_in_2 = r_114; // @[Multiplier.scala 132:13]
  assign c53_21_io_in_3 = r_115; // @[Multiplier.scala 132:13]
  assign c53_21_io_in_4 = c53_19_io_out_1; // @[Multiplier.scala 136:41]
  assign c32_4_io_in_0 = r_116; // @[Multiplier.scala 126:19]
  assign c32_4_io_in_1 = r_117; // @[Multiplier.scala 126:19]
  assign c32_4_io_in_2 = r_118; // @[Multiplier.scala 126:19]
  assign c53_22_io_in_0 = r_119; // @[Multiplier.scala 132:13]
  assign c53_22_io_in_1 = r_120; // @[Multiplier.scala 132:13]
  assign c53_22_io_in_2 = r_121; // @[Multiplier.scala 132:13]
  assign c53_22_io_in_3 = r_122; // @[Multiplier.scala 132:13]
  assign c53_22_io_in_4 = c53_20_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_23_io_in_0 = r_123; // @[Multiplier.scala 132:13]
  assign c53_23_io_in_1 = r_124; // @[Multiplier.scala 132:13]
  assign c53_23_io_in_2 = r_125; // @[Multiplier.scala 132:13]
  assign c53_23_io_in_3 = r_126; // @[Multiplier.scala 132:13]
  assign c53_23_io_in_4 = c53_21_io_out_1; // @[Multiplier.scala 136:41]
  assign c32_5_io_in_0 = r_127; // @[Multiplier.scala 126:19]
  assign c32_5_io_in_1 = r_128; // @[Multiplier.scala 126:19]
  assign c32_5_io_in_2 = r_129; // @[Multiplier.scala 126:19]
  assign c53_24_io_in_0 = r_130; // @[Multiplier.scala 132:13]
  assign c53_24_io_in_1 = r_131; // @[Multiplier.scala 132:13]
  assign c53_24_io_in_2 = r_132; // @[Multiplier.scala 132:13]
  assign c53_24_io_in_3 = r_133; // @[Multiplier.scala 132:13]
  assign c53_24_io_in_4 = c53_22_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_25_io_in_0 = r_134; // @[Multiplier.scala 132:13]
  assign c53_25_io_in_1 = r_135; // @[Multiplier.scala 132:13]
  assign c53_25_io_in_2 = r_136; // @[Multiplier.scala 132:13]
  assign c53_25_io_in_3 = r_137; // @[Multiplier.scala 132:13]
  assign c53_25_io_in_4 = c53_23_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_26_io_in_0 = r_138; // @[Multiplier.scala 132:13]
  assign c53_26_io_in_1 = r_139; // @[Multiplier.scala 132:13]
  assign c53_26_io_in_2 = r_140; // @[Multiplier.scala 132:13]
  assign c53_26_io_in_3 = r_141; // @[Multiplier.scala 132:13]
  assign c53_26_io_in_4 = 1'h0; // @[Multiplier.scala 134:24]
  assign c53_27_io_in_0 = r_142; // @[Multiplier.scala 132:13]
  assign c53_27_io_in_1 = r_143; // @[Multiplier.scala 132:13]
  assign c53_27_io_in_2 = r_144; // @[Multiplier.scala 132:13]
  assign c53_27_io_in_3 = r_145; // @[Multiplier.scala 132:13]
  assign c53_27_io_in_4 = c53_24_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_28_io_in_0 = r_146; // @[Multiplier.scala 132:13]
  assign c53_28_io_in_1 = r_147; // @[Multiplier.scala 132:13]
  assign c53_28_io_in_2 = r_148; // @[Multiplier.scala 132:13]
  assign c53_28_io_in_3 = r_149; // @[Multiplier.scala 132:13]
  assign c53_28_io_in_4 = c53_25_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_29_io_in_0 = r_150; // @[Multiplier.scala 132:13]
  assign c53_29_io_in_1 = r_151; // @[Multiplier.scala 132:13]
  assign c53_29_io_in_2 = r_152; // @[Multiplier.scala 132:13]
  assign c53_29_io_in_3 = r_153; // @[Multiplier.scala 132:13]
  assign c53_29_io_in_4 = c53_26_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_30_io_in_0 = r_154; // @[Multiplier.scala 132:13]
  assign c53_30_io_in_1 = r_155; // @[Multiplier.scala 132:13]
  assign c53_30_io_in_2 = r_156; // @[Multiplier.scala 132:13]
  assign c53_30_io_in_3 = r_157; // @[Multiplier.scala 132:13]
  assign c53_30_io_in_4 = c53_27_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_31_io_in_0 = r_158; // @[Multiplier.scala 132:13]
  assign c53_31_io_in_1 = r_159; // @[Multiplier.scala 132:13]
  assign c53_31_io_in_2 = r_160; // @[Multiplier.scala 132:13]
  assign c53_31_io_in_3 = r_161; // @[Multiplier.scala 132:13]
  assign c53_31_io_in_4 = c53_28_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_32_io_in_0 = r_162; // @[Multiplier.scala 132:13]
  assign c53_32_io_in_1 = r_163; // @[Multiplier.scala 132:13]
  assign c53_32_io_in_2 = r_164; // @[Multiplier.scala 132:13]
  assign c53_32_io_in_3 = r_165; // @[Multiplier.scala 132:13]
  assign c53_32_io_in_4 = c53_29_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_33_io_in_0 = r_167; // @[Multiplier.scala 132:13]
  assign c53_33_io_in_1 = r_168; // @[Multiplier.scala 132:13]
  assign c53_33_io_in_2 = r_169; // @[Multiplier.scala 132:13]
  assign c53_33_io_in_3 = r_170; // @[Multiplier.scala 132:13]
  assign c53_33_io_in_4 = c53_30_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_34_io_in_0 = r_171; // @[Multiplier.scala 132:13]
  assign c53_34_io_in_1 = r_172; // @[Multiplier.scala 132:13]
  assign c53_34_io_in_2 = r_173; // @[Multiplier.scala 132:13]
  assign c53_34_io_in_3 = r_174; // @[Multiplier.scala 132:13]
  assign c53_34_io_in_4 = c53_31_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_35_io_in_0 = r_175; // @[Multiplier.scala 132:13]
  assign c53_35_io_in_1 = r_176; // @[Multiplier.scala 132:13]
  assign c53_35_io_in_2 = r_177; // @[Multiplier.scala 132:13]
  assign c53_35_io_in_3 = r_178; // @[Multiplier.scala 132:13]
  assign c53_35_io_in_4 = c53_32_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_36_io_in_0 = r_180; // @[Multiplier.scala 132:13]
  assign c53_36_io_in_1 = r_181; // @[Multiplier.scala 132:13]
  assign c53_36_io_in_2 = r_182; // @[Multiplier.scala 132:13]
  assign c53_36_io_in_3 = r_183; // @[Multiplier.scala 132:13]
  assign c53_36_io_in_4 = c53_33_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_37_io_in_0 = r_184; // @[Multiplier.scala 132:13]
  assign c53_37_io_in_1 = r_185; // @[Multiplier.scala 132:13]
  assign c53_37_io_in_2 = r_186; // @[Multiplier.scala 132:13]
  assign c53_37_io_in_3 = r_187; // @[Multiplier.scala 132:13]
  assign c53_37_io_in_4 = c53_34_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_38_io_in_0 = r_188; // @[Multiplier.scala 132:13]
  assign c53_38_io_in_1 = r_189; // @[Multiplier.scala 132:13]
  assign c53_38_io_in_2 = r_190; // @[Multiplier.scala 132:13]
  assign c53_38_io_in_3 = r_191; // @[Multiplier.scala 132:13]
  assign c53_38_io_in_4 = c53_35_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_6_io_in_0 = r_192; // @[Multiplier.scala 121:19]
  assign c22_6_io_in_1 = r_193; // @[Multiplier.scala 121:19]
  assign c53_39_io_in_0 = r_194; // @[Multiplier.scala 132:13]
  assign c53_39_io_in_1 = r_195; // @[Multiplier.scala 132:13]
  assign c53_39_io_in_2 = r_196; // @[Multiplier.scala 132:13]
  assign c53_39_io_in_3 = r_197; // @[Multiplier.scala 132:13]
  assign c53_39_io_in_4 = c53_36_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_40_io_in_0 = r_198; // @[Multiplier.scala 132:13]
  assign c53_40_io_in_1 = r_199; // @[Multiplier.scala 132:13]
  assign c53_40_io_in_2 = r_200; // @[Multiplier.scala 132:13]
  assign c53_40_io_in_3 = r_201; // @[Multiplier.scala 132:13]
  assign c53_40_io_in_4 = c53_37_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_41_io_in_0 = r_202; // @[Multiplier.scala 132:13]
  assign c53_41_io_in_1 = r_203; // @[Multiplier.scala 132:13]
  assign c53_41_io_in_2 = r_204; // @[Multiplier.scala 132:13]
  assign c53_41_io_in_3 = r_205; // @[Multiplier.scala 132:13]
  assign c53_41_io_in_4 = c53_38_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_7_io_in_0 = r_206; // @[Multiplier.scala 121:19]
  assign c22_7_io_in_1 = r_207; // @[Multiplier.scala 121:19]
  assign c53_42_io_in_0 = r_208; // @[Multiplier.scala 132:13]
  assign c53_42_io_in_1 = r_209; // @[Multiplier.scala 132:13]
  assign c53_42_io_in_2 = r_210; // @[Multiplier.scala 132:13]
  assign c53_42_io_in_3 = r_211; // @[Multiplier.scala 132:13]
  assign c53_42_io_in_4 = c53_39_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_43_io_in_0 = r_212; // @[Multiplier.scala 132:13]
  assign c53_43_io_in_1 = r_213; // @[Multiplier.scala 132:13]
  assign c53_43_io_in_2 = r_214; // @[Multiplier.scala 132:13]
  assign c53_43_io_in_3 = r_215; // @[Multiplier.scala 132:13]
  assign c53_43_io_in_4 = c53_40_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_44_io_in_0 = r_216; // @[Multiplier.scala 132:13]
  assign c53_44_io_in_1 = r_217; // @[Multiplier.scala 132:13]
  assign c53_44_io_in_2 = r_218; // @[Multiplier.scala 132:13]
  assign c53_44_io_in_3 = r_219; // @[Multiplier.scala 132:13]
  assign c53_44_io_in_4 = c53_41_io_out_1; // @[Multiplier.scala 136:41]
  assign c32_6_io_in_0 = r_220; // @[Multiplier.scala 126:19]
  assign c32_6_io_in_1 = r_221; // @[Multiplier.scala 126:19]
  assign c32_6_io_in_2 = r_222; // @[Multiplier.scala 126:19]
  assign c53_45_io_in_0 = r_223; // @[Multiplier.scala 132:13]
  assign c53_45_io_in_1 = r_224; // @[Multiplier.scala 132:13]
  assign c53_45_io_in_2 = r_225; // @[Multiplier.scala 132:13]
  assign c53_45_io_in_3 = r_226; // @[Multiplier.scala 132:13]
  assign c53_45_io_in_4 = c53_42_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_46_io_in_0 = r_227; // @[Multiplier.scala 132:13]
  assign c53_46_io_in_1 = r_228; // @[Multiplier.scala 132:13]
  assign c53_46_io_in_2 = r_229; // @[Multiplier.scala 132:13]
  assign c53_46_io_in_3 = r_230; // @[Multiplier.scala 132:13]
  assign c53_46_io_in_4 = c53_43_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_47_io_in_0 = r_231; // @[Multiplier.scala 132:13]
  assign c53_47_io_in_1 = r_232; // @[Multiplier.scala 132:13]
  assign c53_47_io_in_2 = r_233; // @[Multiplier.scala 132:13]
  assign c53_47_io_in_3 = r_234; // @[Multiplier.scala 132:13]
  assign c53_47_io_in_4 = c53_44_io_out_1; // @[Multiplier.scala 136:41]
  assign c32_7_io_in_0 = r_235; // @[Multiplier.scala 126:19]
  assign c32_7_io_in_1 = r_236; // @[Multiplier.scala 126:19]
  assign c32_7_io_in_2 = r_237; // @[Multiplier.scala 126:19]
  assign c53_48_io_in_0 = r_238; // @[Multiplier.scala 132:13]
  assign c53_48_io_in_1 = r_239; // @[Multiplier.scala 132:13]
  assign c53_48_io_in_2 = r_240; // @[Multiplier.scala 132:13]
  assign c53_48_io_in_3 = r_241; // @[Multiplier.scala 132:13]
  assign c53_48_io_in_4 = c53_45_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_49_io_in_0 = r_242; // @[Multiplier.scala 132:13]
  assign c53_49_io_in_1 = r_243; // @[Multiplier.scala 132:13]
  assign c53_49_io_in_2 = r_244; // @[Multiplier.scala 132:13]
  assign c53_49_io_in_3 = r_245; // @[Multiplier.scala 132:13]
  assign c53_49_io_in_4 = c53_46_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_50_io_in_0 = r_246; // @[Multiplier.scala 132:13]
  assign c53_50_io_in_1 = r_247; // @[Multiplier.scala 132:13]
  assign c53_50_io_in_2 = r_248; // @[Multiplier.scala 132:13]
  assign c53_50_io_in_3 = r_249; // @[Multiplier.scala 132:13]
  assign c53_50_io_in_4 = c53_47_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_51_io_in_0 = r_250; // @[Multiplier.scala 132:13]
  assign c53_51_io_in_1 = r_251; // @[Multiplier.scala 132:13]
  assign c53_51_io_in_2 = r_252; // @[Multiplier.scala 132:13]
  assign c53_51_io_in_3 = r_253; // @[Multiplier.scala 132:13]
  assign c53_51_io_in_4 = 1'h0; // @[Multiplier.scala 134:24]
  assign c53_52_io_in_0 = r_254; // @[Multiplier.scala 132:13]
  assign c53_52_io_in_1 = r_255; // @[Multiplier.scala 132:13]
  assign c53_52_io_in_2 = r_256; // @[Multiplier.scala 132:13]
  assign c53_52_io_in_3 = r_257; // @[Multiplier.scala 132:13]
  assign c53_52_io_in_4 = c53_48_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_53_io_in_0 = r_258; // @[Multiplier.scala 132:13]
  assign c53_53_io_in_1 = r_259; // @[Multiplier.scala 132:13]
  assign c53_53_io_in_2 = r_260; // @[Multiplier.scala 132:13]
  assign c53_53_io_in_3 = r_261; // @[Multiplier.scala 132:13]
  assign c53_53_io_in_4 = c53_49_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_54_io_in_0 = r_262; // @[Multiplier.scala 132:13]
  assign c53_54_io_in_1 = r_263; // @[Multiplier.scala 132:13]
  assign c53_54_io_in_2 = r_264; // @[Multiplier.scala 132:13]
  assign c53_54_io_in_3 = r_265; // @[Multiplier.scala 132:13]
  assign c53_54_io_in_4 = c53_50_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_55_io_in_0 = r_266; // @[Multiplier.scala 132:13]
  assign c53_55_io_in_1 = r_267; // @[Multiplier.scala 132:13]
  assign c53_55_io_in_2 = r_268; // @[Multiplier.scala 132:13]
  assign c53_55_io_in_3 = r_269; // @[Multiplier.scala 132:13]
  assign c53_55_io_in_4 = c53_51_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_56_io_in_0 = r_270; // @[Multiplier.scala 132:13]
  assign c53_56_io_in_1 = r_271; // @[Multiplier.scala 132:13]
  assign c53_56_io_in_2 = r_272; // @[Multiplier.scala 132:13]
  assign c53_56_io_in_3 = r_273; // @[Multiplier.scala 132:13]
  assign c53_56_io_in_4 = c53_52_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_57_io_in_0 = r_274; // @[Multiplier.scala 132:13]
  assign c53_57_io_in_1 = r_275; // @[Multiplier.scala 132:13]
  assign c53_57_io_in_2 = r_276; // @[Multiplier.scala 132:13]
  assign c53_57_io_in_3 = r_277; // @[Multiplier.scala 132:13]
  assign c53_57_io_in_4 = c53_53_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_58_io_in_0 = r_278; // @[Multiplier.scala 132:13]
  assign c53_58_io_in_1 = r_279; // @[Multiplier.scala 132:13]
  assign c53_58_io_in_2 = r_280; // @[Multiplier.scala 132:13]
  assign c53_58_io_in_3 = r_281; // @[Multiplier.scala 132:13]
  assign c53_58_io_in_4 = c53_54_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_59_io_in_0 = r_282; // @[Multiplier.scala 132:13]
  assign c53_59_io_in_1 = r_283; // @[Multiplier.scala 132:13]
  assign c53_59_io_in_2 = r_284; // @[Multiplier.scala 132:13]
  assign c53_59_io_in_3 = r_285; // @[Multiplier.scala 132:13]
  assign c53_59_io_in_4 = c53_55_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_60_io_in_0 = r_287; // @[Multiplier.scala 132:13]
  assign c53_60_io_in_1 = r_288; // @[Multiplier.scala 132:13]
  assign c53_60_io_in_2 = r_289; // @[Multiplier.scala 132:13]
  assign c53_60_io_in_3 = r_290; // @[Multiplier.scala 132:13]
  assign c53_60_io_in_4 = c53_56_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_61_io_in_0 = r_291; // @[Multiplier.scala 132:13]
  assign c53_61_io_in_1 = r_292; // @[Multiplier.scala 132:13]
  assign c53_61_io_in_2 = r_293; // @[Multiplier.scala 132:13]
  assign c53_61_io_in_3 = r_294; // @[Multiplier.scala 132:13]
  assign c53_61_io_in_4 = c53_57_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_62_io_in_0 = r_295; // @[Multiplier.scala 132:13]
  assign c53_62_io_in_1 = r_296; // @[Multiplier.scala 132:13]
  assign c53_62_io_in_2 = r_297; // @[Multiplier.scala 132:13]
  assign c53_62_io_in_3 = r_298; // @[Multiplier.scala 132:13]
  assign c53_62_io_in_4 = c53_58_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_63_io_in_0 = r_299; // @[Multiplier.scala 132:13]
  assign c53_63_io_in_1 = r_300; // @[Multiplier.scala 132:13]
  assign c53_63_io_in_2 = r_301; // @[Multiplier.scala 132:13]
  assign c53_63_io_in_3 = r_302; // @[Multiplier.scala 132:13]
  assign c53_63_io_in_4 = c53_59_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_64_io_in_0 = r_304; // @[Multiplier.scala 132:13]
  assign c53_64_io_in_1 = r_305; // @[Multiplier.scala 132:13]
  assign c53_64_io_in_2 = r_306; // @[Multiplier.scala 132:13]
  assign c53_64_io_in_3 = r_307; // @[Multiplier.scala 132:13]
  assign c53_64_io_in_4 = c53_60_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_65_io_in_0 = r_308; // @[Multiplier.scala 132:13]
  assign c53_65_io_in_1 = r_309; // @[Multiplier.scala 132:13]
  assign c53_65_io_in_2 = r_310; // @[Multiplier.scala 132:13]
  assign c53_65_io_in_3 = r_311; // @[Multiplier.scala 132:13]
  assign c53_65_io_in_4 = c53_61_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_66_io_in_0 = r_312; // @[Multiplier.scala 132:13]
  assign c53_66_io_in_1 = r_313; // @[Multiplier.scala 132:13]
  assign c53_66_io_in_2 = r_314; // @[Multiplier.scala 132:13]
  assign c53_66_io_in_3 = r_315; // @[Multiplier.scala 132:13]
  assign c53_66_io_in_4 = c53_62_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_67_io_in_0 = r_316; // @[Multiplier.scala 132:13]
  assign c53_67_io_in_1 = r_317; // @[Multiplier.scala 132:13]
  assign c53_67_io_in_2 = r_318; // @[Multiplier.scala 132:13]
  assign c53_67_io_in_3 = r_319; // @[Multiplier.scala 132:13]
  assign c53_67_io_in_4 = c53_63_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_8_io_in_0 = r_320; // @[Multiplier.scala 121:19]
  assign c22_8_io_in_1 = r_321; // @[Multiplier.scala 121:19]
  assign c53_68_io_in_0 = r_322; // @[Multiplier.scala 132:13]
  assign c53_68_io_in_1 = r_323; // @[Multiplier.scala 132:13]
  assign c53_68_io_in_2 = r_324; // @[Multiplier.scala 132:13]
  assign c53_68_io_in_3 = r_325; // @[Multiplier.scala 132:13]
  assign c53_68_io_in_4 = c53_64_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_69_io_in_0 = r_326; // @[Multiplier.scala 132:13]
  assign c53_69_io_in_1 = r_327; // @[Multiplier.scala 132:13]
  assign c53_69_io_in_2 = r_328; // @[Multiplier.scala 132:13]
  assign c53_69_io_in_3 = r_329; // @[Multiplier.scala 132:13]
  assign c53_69_io_in_4 = c53_65_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_70_io_in_0 = r_330; // @[Multiplier.scala 132:13]
  assign c53_70_io_in_1 = r_331; // @[Multiplier.scala 132:13]
  assign c53_70_io_in_2 = r_332; // @[Multiplier.scala 132:13]
  assign c53_70_io_in_3 = r_333; // @[Multiplier.scala 132:13]
  assign c53_70_io_in_4 = c53_66_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_71_io_in_0 = r_334; // @[Multiplier.scala 132:13]
  assign c53_71_io_in_1 = r_335; // @[Multiplier.scala 132:13]
  assign c53_71_io_in_2 = r_336; // @[Multiplier.scala 132:13]
  assign c53_71_io_in_3 = r_337; // @[Multiplier.scala 132:13]
  assign c53_71_io_in_4 = c53_67_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_9_io_in_0 = r_338; // @[Multiplier.scala 121:19]
  assign c22_9_io_in_1 = r_339; // @[Multiplier.scala 121:19]
  assign c53_72_io_in_0 = r_340; // @[Multiplier.scala 132:13]
  assign c53_72_io_in_1 = r_341; // @[Multiplier.scala 132:13]
  assign c53_72_io_in_2 = r_342; // @[Multiplier.scala 132:13]
  assign c53_72_io_in_3 = r_343; // @[Multiplier.scala 132:13]
  assign c53_72_io_in_4 = c53_68_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_73_io_in_0 = r_344; // @[Multiplier.scala 132:13]
  assign c53_73_io_in_1 = r_345; // @[Multiplier.scala 132:13]
  assign c53_73_io_in_2 = r_346; // @[Multiplier.scala 132:13]
  assign c53_73_io_in_3 = r_347; // @[Multiplier.scala 132:13]
  assign c53_73_io_in_4 = c53_69_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_74_io_in_0 = r_348; // @[Multiplier.scala 132:13]
  assign c53_74_io_in_1 = r_349; // @[Multiplier.scala 132:13]
  assign c53_74_io_in_2 = r_350; // @[Multiplier.scala 132:13]
  assign c53_74_io_in_3 = r_351; // @[Multiplier.scala 132:13]
  assign c53_74_io_in_4 = c53_70_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_75_io_in_0 = r_352; // @[Multiplier.scala 132:13]
  assign c53_75_io_in_1 = r_353; // @[Multiplier.scala 132:13]
  assign c53_75_io_in_2 = r_354; // @[Multiplier.scala 132:13]
  assign c53_75_io_in_3 = r_355; // @[Multiplier.scala 132:13]
  assign c53_75_io_in_4 = c53_71_io_out_1; // @[Multiplier.scala 136:41]
  assign c32_8_io_in_0 = r_356; // @[Multiplier.scala 126:19]
  assign c32_8_io_in_1 = r_357; // @[Multiplier.scala 126:19]
  assign c32_8_io_in_2 = r_358; // @[Multiplier.scala 126:19]
  assign c53_76_io_in_0 = r_359; // @[Multiplier.scala 132:13]
  assign c53_76_io_in_1 = r_360; // @[Multiplier.scala 132:13]
  assign c53_76_io_in_2 = r_361; // @[Multiplier.scala 132:13]
  assign c53_76_io_in_3 = r_362; // @[Multiplier.scala 132:13]
  assign c53_76_io_in_4 = c53_72_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_77_io_in_0 = r_363; // @[Multiplier.scala 132:13]
  assign c53_77_io_in_1 = r_364; // @[Multiplier.scala 132:13]
  assign c53_77_io_in_2 = r_365; // @[Multiplier.scala 132:13]
  assign c53_77_io_in_3 = r_366; // @[Multiplier.scala 132:13]
  assign c53_77_io_in_4 = c53_73_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_78_io_in_0 = r_367; // @[Multiplier.scala 132:13]
  assign c53_78_io_in_1 = r_368; // @[Multiplier.scala 132:13]
  assign c53_78_io_in_2 = r_369; // @[Multiplier.scala 132:13]
  assign c53_78_io_in_3 = r_370; // @[Multiplier.scala 132:13]
  assign c53_78_io_in_4 = c53_74_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_79_io_in_0 = r_371; // @[Multiplier.scala 132:13]
  assign c53_79_io_in_1 = r_372; // @[Multiplier.scala 132:13]
  assign c53_79_io_in_2 = r_373; // @[Multiplier.scala 132:13]
  assign c53_79_io_in_3 = r_374; // @[Multiplier.scala 132:13]
  assign c53_79_io_in_4 = c53_75_io_out_1; // @[Multiplier.scala 136:41]
  assign c32_9_io_in_0 = r_375; // @[Multiplier.scala 126:19]
  assign c32_9_io_in_1 = r_376; // @[Multiplier.scala 126:19]
  assign c32_9_io_in_2 = r_377; // @[Multiplier.scala 126:19]
  assign c53_80_io_in_0 = r_378; // @[Multiplier.scala 132:13]
  assign c53_80_io_in_1 = r_379; // @[Multiplier.scala 132:13]
  assign c53_80_io_in_2 = r_380; // @[Multiplier.scala 132:13]
  assign c53_80_io_in_3 = r_381; // @[Multiplier.scala 132:13]
  assign c53_80_io_in_4 = c53_76_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_81_io_in_0 = r_382; // @[Multiplier.scala 132:13]
  assign c53_81_io_in_1 = r_383; // @[Multiplier.scala 132:13]
  assign c53_81_io_in_2 = r_384; // @[Multiplier.scala 132:13]
  assign c53_81_io_in_3 = r_385; // @[Multiplier.scala 132:13]
  assign c53_81_io_in_4 = c53_77_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_82_io_in_0 = r_386; // @[Multiplier.scala 132:13]
  assign c53_82_io_in_1 = r_387; // @[Multiplier.scala 132:13]
  assign c53_82_io_in_2 = r_388; // @[Multiplier.scala 132:13]
  assign c53_82_io_in_3 = r_389; // @[Multiplier.scala 132:13]
  assign c53_82_io_in_4 = c53_78_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_83_io_in_0 = r_390; // @[Multiplier.scala 132:13]
  assign c53_83_io_in_1 = r_391; // @[Multiplier.scala 132:13]
  assign c53_83_io_in_2 = r_392; // @[Multiplier.scala 132:13]
  assign c53_83_io_in_3 = r_393; // @[Multiplier.scala 132:13]
  assign c53_83_io_in_4 = c53_79_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_84_io_in_0 = r_394; // @[Multiplier.scala 132:13]
  assign c53_84_io_in_1 = r_395; // @[Multiplier.scala 132:13]
  assign c53_84_io_in_2 = r_396; // @[Multiplier.scala 132:13]
  assign c53_84_io_in_3 = r_397; // @[Multiplier.scala 132:13]
  assign c53_84_io_in_4 = 1'h0; // @[Multiplier.scala 134:24]
  assign c53_85_io_in_0 = r_398; // @[Multiplier.scala 132:13]
  assign c53_85_io_in_1 = r_399; // @[Multiplier.scala 132:13]
  assign c53_85_io_in_2 = r_400; // @[Multiplier.scala 132:13]
  assign c53_85_io_in_3 = r_401; // @[Multiplier.scala 132:13]
  assign c53_85_io_in_4 = c53_80_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_86_io_in_0 = r_402; // @[Multiplier.scala 132:13]
  assign c53_86_io_in_1 = r_403; // @[Multiplier.scala 132:13]
  assign c53_86_io_in_2 = r_404; // @[Multiplier.scala 132:13]
  assign c53_86_io_in_3 = r_405; // @[Multiplier.scala 132:13]
  assign c53_86_io_in_4 = c53_81_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_87_io_in_0 = r_406; // @[Multiplier.scala 132:13]
  assign c53_87_io_in_1 = r_407; // @[Multiplier.scala 132:13]
  assign c53_87_io_in_2 = r_408; // @[Multiplier.scala 132:13]
  assign c53_87_io_in_3 = r_409; // @[Multiplier.scala 132:13]
  assign c53_87_io_in_4 = c53_82_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_88_io_in_0 = r_410; // @[Multiplier.scala 132:13]
  assign c53_88_io_in_1 = r_411; // @[Multiplier.scala 132:13]
  assign c53_88_io_in_2 = r_412; // @[Multiplier.scala 132:13]
  assign c53_88_io_in_3 = r_413; // @[Multiplier.scala 132:13]
  assign c53_88_io_in_4 = c53_83_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_89_io_in_0 = r_414; // @[Multiplier.scala 132:13]
  assign c53_89_io_in_1 = r_415; // @[Multiplier.scala 132:13]
  assign c53_89_io_in_2 = r_416; // @[Multiplier.scala 132:13]
  assign c53_89_io_in_3 = r_417; // @[Multiplier.scala 132:13]
  assign c53_89_io_in_4 = c53_84_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_90_io_in_0 = r_418; // @[Multiplier.scala 132:13]
  assign c53_90_io_in_1 = r_419; // @[Multiplier.scala 132:13]
  assign c53_90_io_in_2 = r_420; // @[Multiplier.scala 132:13]
  assign c53_90_io_in_3 = r_421; // @[Multiplier.scala 132:13]
  assign c53_90_io_in_4 = c53_85_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_91_io_in_0 = r_422; // @[Multiplier.scala 132:13]
  assign c53_91_io_in_1 = r_423; // @[Multiplier.scala 132:13]
  assign c53_91_io_in_2 = r_424; // @[Multiplier.scala 132:13]
  assign c53_91_io_in_3 = r_425; // @[Multiplier.scala 132:13]
  assign c53_91_io_in_4 = c53_86_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_92_io_in_0 = r_426; // @[Multiplier.scala 132:13]
  assign c53_92_io_in_1 = r_427; // @[Multiplier.scala 132:13]
  assign c53_92_io_in_2 = r_428; // @[Multiplier.scala 132:13]
  assign c53_92_io_in_3 = r_429; // @[Multiplier.scala 132:13]
  assign c53_92_io_in_4 = c53_87_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_93_io_in_0 = r_430; // @[Multiplier.scala 132:13]
  assign c53_93_io_in_1 = r_431; // @[Multiplier.scala 132:13]
  assign c53_93_io_in_2 = r_432; // @[Multiplier.scala 132:13]
  assign c53_93_io_in_3 = r_433; // @[Multiplier.scala 132:13]
  assign c53_93_io_in_4 = c53_88_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_94_io_in_0 = r_434; // @[Multiplier.scala 132:13]
  assign c53_94_io_in_1 = r_435; // @[Multiplier.scala 132:13]
  assign c53_94_io_in_2 = r_436; // @[Multiplier.scala 132:13]
  assign c53_94_io_in_3 = r_437; // @[Multiplier.scala 132:13]
  assign c53_94_io_in_4 = c53_89_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_95_io_in_0 = r_439; // @[Multiplier.scala 132:13]
  assign c53_95_io_in_1 = r_440; // @[Multiplier.scala 132:13]
  assign c53_95_io_in_2 = r_441; // @[Multiplier.scala 132:13]
  assign c53_95_io_in_3 = r_442; // @[Multiplier.scala 132:13]
  assign c53_95_io_in_4 = c53_90_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_96_io_in_0 = r_443; // @[Multiplier.scala 132:13]
  assign c53_96_io_in_1 = r_444; // @[Multiplier.scala 132:13]
  assign c53_96_io_in_2 = r_445; // @[Multiplier.scala 132:13]
  assign c53_96_io_in_3 = r_446; // @[Multiplier.scala 132:13]
  assign c53_96_io_in_4 = c53_91_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_97_io_in_0 = r_447; // @[Multiplier.scala 132:13]
  assign c53_97_io_in_1 = r_448; // @[Multiplier.scala 132:13]
  assign c53_97_io_in_2 = r_449; // @[Multiplier.scala 132:13]
  assign c53_97_io_in_3 = r_450; // @[Multiplier.scala 132:13]
  assign c53_97_io_in_4 = c53_92_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_98_io_in_0 = r_451; // @[Multiplier.scala 132:13]
  assign c53_98_io_in_1 = r_452; // @[Multiplier.scala 132:13]
  assign c53_98_io_in_2 = r_453; // @[Multiplier.scala 132:13]
  assign c53_98_io_in_3 = r_454; // @[Multiplier.scala 132:13]
  assign c53_98_io_in_4 = c53_93_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_99_io_in_0 = r_455; // @[Multiplier.scala 132:13]
  assign c53_99_io_in_1 = r_456; // @[Multiplier.scala 132:13]
  assign c53_99_io_in_2 = r_457; // @[Multiplier.scala 132:13]
  assign c53_99_io_in_3 = r_458; // @[Multiplier.scala 132:13]
  assign c53_99_io_in_4 = c53_94_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_100_io_in_0 = r_460; // @[Multiplier.scala 132:13]
  assign c53_100_io_in_1 = r_461; // @[Multiplier.scala 132:13]
  assign c53_100_io_in_2 = r_462; // @[Multiplier.scala 132:13]
  assign c53_100_io_in_3 = r_463; // @[Multiplier.scala 132:13]
  assign c53_100_io_in_4 = c53_95_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_101_io_in_0 = r_464; // @[Multiplier.scala 132:13]
  assign c53_101_io_in_1 = r_465; // @[Multiplier.scala 132:13]
  assign c53_101_io_in_2 = r_466; // @[Multiplier.scala 132:13]
  assign c53_101_io_in_3 = r_467; // @[Multiplier.scala 132:13]
  assign c53_101_io_in_4 = c53_96_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_102_io_in_0 = r_468; // @[Multiplier.scala 132:13]
  assign c53_102_io_in_1 = r_469; // @[Multiplier.scala 132:13]
  assign c53_102_io_in_2 = r_470; // @[Multiplier.scala 132:13]
  assign c53_102_io_in_3 = r_471; // @[Multiplier.scala 132:13]
  assign c53_102_io_in_4 = c53_97_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_103_io_in_0 = r_472; // @[Multiplier.scala 132:13]
  assign c53_103_io_in_1 = r_473; // @[Multiplier.scala 132:13]
  assign c53_103_io_in_2 = r_474; // @[Multiplier.scala 132:13]
  assign c53_103_io_in_3 = r_475; // @[Multiplier.scala 132:13]
  assign c53_103_io_in_4 = c53_98_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_104_io_in_0 = r_476; // @[Multiplier.scala 132:13]
  assign c53_104_io_in_1 = r_477; // @[Multiplier.scala 132:13]
  assign c53_104_io_in_2 = r_478; // @[Multiplier.scala 132:13]
  assign c53_104_io_in_3 = r_479; // @[Multiplier.scala 132:13]
  assign c53_104_io_in_4 = c53_99_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_10_io_in_0 = r_480; // @[Multiplier.scala 121:19]
  assign c22_10_io_in_1 = r_481; // @[Multiplier.scala 121:19]
  assign c53_105_io_in_0 = r_482; // @[Multiplier.scala 132:13]
  assign c53_105_io_in_1 = r_483; // @[Multiplier.scala 132:13]
  assign c53_105_io_in_2 = r_484; // @[Multiplier.scala 132:13]
  assign c53_105_io_in_3 = r_485; // @[Multiplier.scala 132:13]
  assign c53_105_io_in_4 = c53_100_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_106_io_in_0 = r_486; // @[Multiplier.scala 132:13]
  assign c53_106_io_in_1 = r_487; // @[Multiplier.scala 132:13]
  assign c53_106_io_in_2 = r_488; // @[Multiplier.scala 132:13]
  assign c53_106_io_in_3 = r_489; // @[Multiplier.scala 132:13]
  assign c53_106_io_in_4 = c53_101_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_107_io_in_0 = r_490; // @[Multiplier.scala 132:13]
  assign c53_107_io_in_1 = r_491; // @[Multiplier.scala 132:13]
  assign c53_107_io_in_2 = r_492; // @[Multiplier.scala 132:13]
  assign c53_107_io_in_3 = r_493; // @[Multiplier.scala 132:13]
  assign c53_107_io_in_4 = c53_102_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_108_io_in_0 = r_494; // @[Multiplier.scala 132:13]
  assign c53_108_io_in_1 = r_495; // @[Multiplier.scala 132:13]
  assign c53_108_io_in_2 = r_496; // @[Multiplier.scala 132:13]
  assign c53_108_io_in_3 = r_497; // @[Multiplier.scala 132:13]
  assign c53_108_io_in_4 = c53_103_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_109_io_in_0 = r_498; // @[Multiplier.scala 132:13]
  assign c53_109_io_in_1 = r_499; // @[Multiplier.scala 132:13]
  assign c53_109_io_in_2 = r_500; // @[Multiplier.scala 132:13]
  assign c53_109_io_in_3 = r_501; // @[Multiplier.scala 132:13]
  assign c53_109_io_in_4 = c53_104_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_11_io_in_0 = r_502; // @[Multiplier.scala 121:19]
  assign c22_11_io_in_1 = r_503; // @[Multiplier.scala 121:19]
  assign c53_110_io_in_0 = r_504; // @[Multiplier.scala 132:13]
  assign c53_110_io_in_1 = r_505; // @[Multiplier.scala 132:13]
  assign c53_110_io_in_2 = r_506; // @[Multiplier.scala 132:13]
  assign c53_110_io_in_3 = r_507; // @[Multiplier.scala 132:13]
  assign c53_110_io_in_4 = c53_105_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_111_io_in_0 = r_508; // @[Multiplier.scala 132:13]
  assign c53_111_io_in_1 = r_509; // @[Multiplier.scala 132:13]
  assign c53_111_io_in_2 = r_510; // @[Multiplier.scala 132:13]
  assign c53_111_io_in_3 = r_511; // @[Multiplier.scala 132:13]
  assign c53_111_io_in_4 = c53_106_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_112_io_in_0 = r_512; // @[Multiplier.scala 132:13]
  assign c53_112_io_in_1 = r_513; // @[Multiplier.scala 132:13]
  assign c53_112_io_in_2 = r_514; // @[Multiplier.scala 132:13]
  assign c53_112_io_in_3 = r_515; // @[Multiplier.scala 132:13]
  assign c53_112_io_in_4 = c53_107_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_113_io_in_0 = r_516; // @[Multiplier.scala 132:13]
  assign c53_113_io_in_1 = r_517; // @[Multiplier.scala 132:13]
  assign c53_113_io_in_2 = r_518; // @[Multiplier.scala 132:13]
  assign c53_113_io_in_3 = r_519; // @[Multiplier.scala 132:13]
  assign c53_113_io_in_4 = c53_108_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_114_io_in_0 = r_520; // @[Multiplier.scala 132:13]
  assign c53_114_io_in_1 = r_521; // @[Multiplier.scala 132:13]
  assign c53_114_io_in_2 = r_522; // @[Multiplier.scala 132:13]
  assign c53_114_io_in_3 = r_523; // @[Multiplier.scala 132:13]
  assign c53_114_io_in_4 = c53_109_io_out_1; // @[Multiplier.scala 136:41]
  assign c32_10_io_in_0 = r_524; // @[Multiplier.scala 126:19]
  assign c32_10_io_in_1 = r_525; // @[Multiplier.scala 126:19]
  assign c32_10_io_in_2 = r_526; // @[Multiplier.scala 126:19]
  assign c53_115_io_in_0 = r_527; // @[Multiplier.scala 132:13]
  assign c53_115_io_in_1 = r_528; // @[Multiplier.scala 132:13]
  assign c53_115_io_in_2 = r_529; // @[Multiplier.scala 132:13]
  assign c53_115_io_in_3 = r_530; // @[Multiplier.scala 132:13]
  assign c53_115_io_in_4 = c53_110_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_116_io_in_0 = r_531; // @[Multiplier.scala 132:13]
  assign c53_116_io_in_1 = r_532; // @[Multiplier.scala 132:13]
  assign c53_116_io_in_2 = r_533; // @[Multiplier.scala 132:13]
  assign c53_116_io_in_3 = r_534; // @[Multiplier.scala 132:13]
  assign c53_116_io_in_4 = c53_111_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_117_io_in_0 = r_535; // @[Multiplier.scala 132:13]
  assign c53_117_io_in_1 = r_536; // @[Multiplier.scala 132:13]
  assign c53_117_io_in_2 = r_537; // @[Multiplier.scala 132:13]
  assign c53_117_io_in_3 = r_538; // @[Multiplier.scala 132:13]
  assign c53_117_io_in_4 = c53_112_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_118_io_in_0 = r_539; // @[Multiplier.scala 132:13]
  assign c53_118_io_in_1 = r_540; // @[Multiplier.scala 132:13]
  assign c53_118_io_in_2 = r_541; // @[Multiplier.scala 132:13]
  assign c53_118_io_in_3 = r_542; // @[Multiplier.scala 132:13]
  assign c53_118_io_in_4 = c53_113_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_119_io_in_0 = r_543; // @[Multiplier.scala 132:13]
  assign c53_119_io_in_1 = r_544; // @[Multiplier.scala 132:13]
  assign c53_119_io_in_2 = r_545; // @[Multiplier.scala 132:13]
  assign c53_119_io_in_3 = r_546; // @[Multiplier.scala 132:13]
  assign c53_119_io_in_4 = c53_114_io_out_1; // @[Multiplier.scala 136:41]
  assign c32_11_io_in_0 = r_547; // @[Multiplier.scala 126:19]
  assign c32_11_io_in_1 = r_548; // @[Multiplier.scala 126:19]
  assign c32_11_io_in_2 = r_549; // @[Multiplier.scala 126:19]
  assign c53_120_io_in_0 = r_550; // @[Multiplier.scala 132:13]
  assign c53_120_io_in_1 = r_551; // @[Multiplier.scala 132:13]
  assign c53_120_io_in_2 = r_552; // @[Multiplier.scala 132:13]
  assign c53_120_io_in_3 = r_553; // @[Multiplier.scala 132:13]
  assign c53_120_io_in_4 = c53_115_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_121_io_in_0 = r_554; // @[Multiplier.scala 132:13]
  assign c53_121_io_in_1 = r_555; // @[Multiplier.scala 132:13]
  assign c53_121_io_in_2 = r_556; // @[Multiplier.scala 132:13]
  assign c53_121_io_in_3 = r_557; // @[Multiplier.scala 132:13]
  assign c53_121_io_in_4 = c53_116_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_122_io_in_0 = r_558; // @[Multiplier.scala 132:13]
  assign c53_122_io_in_1 = r_559; // @[Multiplier.scala 132:13]
  assign c53_122_io_in_2 = r_560; // @[Multiplier.scala 132:13]
  assign c53_122_io_in_3 = r_561; // @[Multiplier.scala 132:13]
  assign c53_122_io_in_4 = c53_117_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_123_io_in_0 = r_562; // @[Multiplier.scala 132:13]
  assign c53_123_io_in_1 = r_563; // @[Multiplier.scala 132:13]
  assign c53_123_io_in_2 = r_564; // @[Multiplier.scala 132:13]
  assign c53_123_io_in_3 = r_565; // @[Multiplier.scala 132:13]
  assign c53_123_io_in_4 = c53_118_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_124_io_in_0 = r_566; // @[Multiplier.scala 132:13]
  assign c53_124_io_in_1 = r_567; // @[Multiplier.scala 132:13]
  assign c53_124_io_in_2 = r_568; // @[Multiplier.scala 132:13]
  assign c53_124_io_in_3 = r_569; // @[Multiplier.scala 132:13]
  assign c53_124_io_in_4 = c53_119_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_125_io_in_0 = r_570; // @[Multiplier.scala 132:13]
  assign c53_125_io_in_1 = r_571; // @[Multiplier.scala 132:13]
  assign c53_125_io_in_2 = r_572; // @[Multiplier.scala 132:13]
  assign c53_125_io_in_3 = r_573; // @[Multiplier.scala 132:13]
  assign c53_125_io_in_4 = 1'h0; // @[Multiplier.scala 134:24]
  assign c53_126_io_in_0 = r_574; // @[Multiplier.scala 132:13]
  assign c53_126_io_in_1 = r_575; // @[Multiplier.scala 132:13]
  assign c53_126_io_in_2 = r_576; // @[Multiplier.scala 132:13]
  assign c53_126_io_in_3 = r_577; // @[Multiplier.scala 132:13]
  assign c53_126_io_in_4 = c53_120_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_127_io_in_0 = r_578; // @[Multiplier.scala 132:13]
  assign c53_127_io_in_1 = r_579; // @[Multiplier.scala 132:13]
  assign c53_127_io_in_2 = r_580; // @[Multiplier.scala 132:13]
  assign c53_127_io_in_3 = r_581; // @[Multiplier.scala 132:13]
  assign c53_127_io_in_4 = c53_121_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_128_io_in_0 = r_582; // @[Multiplier.scala 132:13]
  assign c53_128_io_in_1 = r_583; // @[Multiplier.scala 132:13]
  assign c53_128_io_in_2 = r_584; // @[Multiplier.scala 132:13]
  assign c53_128_io_in_3 = r_585; // @[Multiplier.scala 132:13]
  assign c53_128_io_in_4 = c53_122_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_129_io_in_0 = r_586; // @[Multiplier.scala 132:13]
  assign c53_129_io_in_1 = r_587; // @[Multiplier.scala 132:13]
  assign c53_129_io_in_2 = r_588; // @[Multiplier.scala 132:13]
  assign c53_129_io_in_3 = r_589; // @[Multiplier.scala 132:13]
  assign c53_129_io_in_4 = c53_123_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_130_io_in_0 = r_590; // @[Multiplier.scala 132:13]
  assign c53_130_io_in_1 = r_591; // @[Multiplier.scala 132:13]
  assign c53_130_io_in_2 = r_592; // @[Multiplier.scala 132:13]
  assign c53_130_io_in_3 = r_593; // @[Multiplier.scala 132:13]
  assign c53_130_io_in_4 = c53_124_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_131_io_in_0 = r_594; // @[Multiplier.scala 132:13]
  assign c53_131_io_in_1 = r_595; // @[Multiplier.scala 132:13]
  assign c53_131_io_in_2 = r_596; // @[Multiplier.scala 132:13]
  assign c53_131_io_in_3 = r_597; // @[Multiplier.scala 132:13]
  assign c53_131_io_in_4 = c53_125_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_132_io_in_0 = r_598; // @[Multiplier.scala 132:13]
  assign c53_132_io_in_1 = r_599; // @[Multiplier.scala 132:13]
  assign c53_132_io_in_2 = r_600; // @[Multiplier.scala 132:13]
  assign c53_132_io_in_3 = r_601; // @[Multiplier.scala 132:13]
  assign c53_132_io_in_4 = c53_126_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_133_io_in_0 = r_602; // @[Multiplier.scala 132:13]
  assign c53_133_io_in_1 = r_603; // @[Multiplier.scala 132:13]
  assign c53_133_io_in_2 = r_604; // @[Multiplier.scala 132:13]
  assign c53_133_io_in_3 = r_605; // @[Multiplier.scala 132:13]
  assign c53_133_io_in_4 = c53_127_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_134_io_in_0 = r_606; // @[Multiplier.scala 132:13]
  assign c53_134_io_in_1 = r_607; // @[Multiplier.scala 132:13]
  assign c53_134_io_in_2 = r_608; // @[Multiplier.scala 132:13]
  assign c53_134_io_in_3 = r_609; // @[Multiplier.scala 132:13]
  assign c53_134_io_in_4 = c53_128_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_135_io_in_0 = r_610; // @[Multiplier.scala 132:13]
  assign c53_135_io_in_1 = r_611; // @[Multiplier.scala 132:13]
  assign c53_135_io_in_2 = r_612; // @[Multiplier.scala 132:13]
  assign c53_135_io_in_3 = r_613; // @[Multiplier.scala 132:13]
  assign c53_135_io_in_4 = c53_129_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_136_io_in_0 = r_614; // @[Multiplier.scala 132:13]
  assign c53_136_io_in_1 = r_615; // @[Multiplier.scala 132:13]
  assign c53_136_io_in_2 = r_616; // @[Multiplier.scala 132:13]
  assign c53_136_io_in_3 = r_617; // @[Multiplier.scala 132:13]
  assign c53_136_io_in_4 = c53_130_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_137_io_in_0 = r_618; // @[Multiplier.scala 132:13]
  assign c53_137_io_in_1 = r_619; // @[Multiplier.scala 132:13]
  assign c53_137_io_in_2 = r_620; // @[Multiplier.scala 132:13]
  assign c53_137_io_in_3 = r_621; // @[Multiplier.scala 132:13]
  assign c53_137_io_in_4 = c53_131_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_138_io_in_0 = r_623; // @[Multiplier.scala 132:13]
  assign c53_138_io_in_1 = r_624; // @[Multiplier.scala 132:13]
  assign c53_138_io_in_2 = r_625; // @[Multiplier.scala 132:13]
  assign c53_138_io_in_3 = r_626; // @[Multiplier.scala 132:13]
  assign c53_138_io_in_4 = c53_132_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_139_io_in_0 = r_627; // @[Multiplier.scala 132:13]
  assign c53_139_io_in_1 = r_628; // @[Multiplier.scala 132:13]
  assign c53_139_io_in_2 = r_629; // @[Multiplier.scala 132:13]
  assign c53_139_io_in_3 = r_630; // @[Multiplier.scala 132:13]
  assign c53_139_io_in_4 = c53_133_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_140_io_in_0 = r_631; // @[Multiplier.scala 132:13]
  assign c53_140_io_in_1 = r_632; // @[Multiplier.scala 132:13]
  assign c53_140_io_in_2 = r_633; // @[Multiplier.scala 132:13]
  assign c53_140_io_in_3 = r_634; // @[Multiplier.scala 132:13]
  assign c53_140_io_in_4 = c53_134_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_141_io_in_0 = r_635; // @[Multiplier.scala 132:13]
  assign c53_141_io_in_1 = r_636; // @[Multiplier.scala 132:13]
  assign c53_141_io_in_2 = r_637; // @[Multiplier.scala 132:13]
  assign c53_141_io_in_3 = r_638; // @[Multiplier.scala 132:13]
  assign c53_141_io_in_4 = c53_135_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_142_io_in_0 = r_639; // @[Multiplier.scala 132:13]
  assign c53_142_io_in_1 = r_640; // @[Multiplier.scala 132:13]
  assign c53_142_io_in_2 = r_641; // @[Multiplier.scala 132:13]
  assign c53_142_io_in_3 = r_642; // @[Multiplier.scala 132:13]
  assign c53_142_io_in_4 = c53_136_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_143_io_in_0 = r_643; // @[Multiplier.scala 132:13]
  assign c53_143_io_in_1 = r_644; // @[Multiplier.scala 132:13]
  assign c53_143_io_in_2 = r_645; // @[Multiplier.scala 132:13]
  assign c53_143_io_in_3 = r_646; // @[Multiplier.scala 132:13]
  assign c53_143_io_in_4 = c53_137_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_144_io_in_0 = r_648; // @[Multiplier.scala 132:13]
  assign c53_144_io_in_1 = r_649; // @[Multiplier.scala 132:13]
  assign c53_144_io_in_2 = r_650; // @[Multiplier.scala 132:13]
  assign c53_144_io_in_3 = r_651; // @[Multiplier.scala 132:13]
  assign c53_144_io_in_4 = c53_138_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_145_io_in_0 = r_652; // @[Multiplier.scala 132:13]
  assign c53_145_io_in_1 = r_653; // @[Multiplier.scala 132:13]
  assign c53_145_io_in_2 = r_654; // @[Multiplier.scala 132:13]
  assign c53_145_io_in_3 = r_655; // @[Multiplier.scala 132:13]
  assign c53_145_io_in_4 = c53_139_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_146_io_in_0 = r_656; // @[Multiplier.scala 132:13]
  assign c53_146_io_in_1 = r_657; // @[Multiplier.scala 132:13]
  assign c53_146_io_in_2 = r_658; // @[Multiplier.scala 132:13]
  assign c53_146_io_in_3 = r_659; // @[Multiplier.scala 132:13]
  assign c53_146_io_in_4 = c53_140_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_147_io_in_0 = r_660; // @[Multiplier.scala 132:13]
  assign c53_147_io_in_1 = r_661; // @[Multiplier.scala 132:13]
  assign c53_147_io_in_2 = r_662; // @[Multiplier.scala 132:13]
  assign c53_147_io_in_3 = r_663; // @[Multiplier.scala 132:13]
  assign c53_147_io_in_4 = c53_141_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_148_io_in_0 = r_664; // @[Multiplier.scala 132:13]
  assign c53_148_io_in_1 = r_665; // @[Multiplier.scala 132:13]
  assign c53_148_io_in_2 = r_666; // @[Multiplier.scala 132:13]
  assign c53_148_io_in_3 = r_667; // @[Multiplier.scala 132:13]
  assign c53_148_io_in_4 = c53_142_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_149_io_in_0 = r_668; // @[Multiplier.scala 132:13]
  assign c53_149_io_in_1 = r_669; // @[Multiplier.scala 132:13]
  assign c53_149_io_in_2 = r_670; // @[Multiplier.scala 132:13]
  assign c53_149_io_in_3 = r_671; // @[Multiplier.scala 132:13]
  assign c53_149_io_in_4 = c53_143_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_12_io_in_0 = r_672; // @[Multiplier.scala 121:19]
  assign c22_12_io_in_1 = r_673; // @[Multiplier.scala 121:19]
  assign c53_150_io_in_0 = r_674; // @[Multiplier.scala 132:13]
  assign c53_150_io_in_1 = r_675; // @[Multiplier.scala 132:13]
  assign c53_150_io_in_2 = r_676; // @[Multiplier.scala 132:13]
  assign c53_150_io_in_3 = r_677; // @[Multiplier.scala 132:13]
  assign c53_150_io_in_4 = c53_144_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_151_io_in_0 = r_678; // @[Multiplier.scala 132:13]
  assign c53_151_io_in_1 = r_679; // @[Multiplier.scala 132:13]
  assign c53_151_io_in_2 = r_680; // @[Multiplier.scala 132:13]
  assign c53_151_io_in_3 = r_681; // @[Multiplier.scala 132:13]
  assign c53_151_io_in_4 = c53_145_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_152_io_in_0 = r_682; // @[Multiplier.scala 132:13]
  assign c53_152_io_in_1 = r_683; // @[Multiplier.scala 132:13]
  assign c53_152_io_in_2 = r_684; // @[Multiplier.scala 132:13]
  assign c53_152_io_in_3 = r_685; // @[Multiplier.scala 132:13]
  assign c53_152_io_in_4 = c53_146_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_153_io_in_0 = r_686; // @[Multiplier.scala 132:13]
  assign c53_153_io_in_1 = r_687; // @[Multiplier.scala 132:13]
  assign c53_153_io_in_2 = r_688; // @[Multiplier.scala 132:13]
  assign c53_153_io_in_3 = r_689; // @[Multiplier.scala 132:13]
  assign c53_153_io_in_4 = c53_147_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_154_io_in_0 = r_690; // @[Multiplier.scala 132:13]
  assign c53_154_io_in_1 = r_691; // @[Multiplier.scala 132:13]
  assign c53_154_io_in_2 = r_692; // @[Multiplier.scala 132:13]
  assign c53_154_io_in_3 = r_693; // @[Multiplier.scala 132:13]
  assign c53_154_io_in_4 = c53_148_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_155_io_in_0 = r_694; // @[Multiplier.scala 132:13]
  assign c53_155_io_in_1 = r_695; // @[Multiplier.scala 132:13]
  assign c53_155_io_in_2 = r_696; // @[Multiplier.scala 132:13]
  assign c53_155_io_in_3 = r_697; // @[Multiplier.scala 132:13]
  assign c53_155_io_in_4 = c53_149_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_13_io_in_0 = r_698; // @[Multiplier.scala 121:19]
  assign c22_13_io_in_1 = r_699; // @[Multiplier.scala 121:19]
  assign c53_156_io_in_0 = r_700; // @[Multiplier.scala 132:13]
  assign c53_156_io_in_1 = r_701; // @[Multiplier.scala 132:13]
  assign c53_156_io_in_2 = r_702; // @[Multiplier.scala 132:13]
  assign c53_156_io_in_3 = r_703; // @[Multiplier.scala 132:13]
  assign c53_156_io_in_4 = c53_150_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_157_io_in_0 = r_704; // @[Multiplier.scala 132:13]
  assign c53_157_io_in_1 = r_705; // @[Multiplier.scala 132:13]
  assign c53_157_io_in_2 = r_706; // @[Multiplier.scala 132:13]
  assign c53_157_io_in_3 = r_707; // @[Multiplier.scala 132:13]
  assign c53_157_io_in_4 = c53_151_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_158_io_in_0 = r_708; // @[Multiplier.scala 132:13]
  assign c53_158_io_in_1 = r_709; // @[Multiplier.scala 132:13]
  assign c53_158_io_in_2 = r_710; // @[Multiplier.scala 132:13]
  assign c53_158_io_in_3 = r_711; // @[Multiplier.scala 132:13]
  assign c53_158_io_in_4 = c53_152_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_159_io_in_0 = r_712; // @[Multiplier.scala 132:13]
  assign c53_159_io_in_1 = r_713; // @[Multiplier.scala 132:13]
  assign c53_159_io_in_2 = r_714; // @[Multiplier.scala 132:13]
  assign c53_159_io_in_3 = r_715; // @[Multiplier.scala 132:13]
  assign c53_159_io_in_4 = c53_153_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_160_io_in_0 = r_716; // @[Multiplier.scala 132:13]
  assign c53_160_io_in_1 = r_717; // @[Multiplier.scala 132:13]
  assign c53_160_io_in_2 = r_718; // @[Multiplier.scala 132:13]
  assign c53_160_io_in_3 = r_719; // @[Multiplier.scala 132:13]
  assign c53_160_io_in_4 = c53_154_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_161_io_in_0 = r_720; // @[Multiplier.scala 132:13]
  assign c53_161_io_in_1 = r_721; // @[Multiplier.scala 132:13]
  assign c53_161_io_in_2 = r_722; // @[Multiplier.scala 132:13]
  assign c53_161_io_in_3 = r_723; // @[Multiplier.scala 132:13]
  assign c53_161_io_in_4 = c53_155_io_out_1; // @[Multiplier.scala 136:41]
  assign c32_12_io_in_0 = r_724; // @[Multiplier.scala 126:19]
  assign c32_12_io_in_1 = r_725; // @[Multiplier.scala 126:19]
  assign c32_12_io_in_2 = r_726; // @[Multiplier.scala 126:19]
  assign c53_162_io_in_0 = r_727; // @[Multiplier.scala 132:13]
  assign c53_162_io_in_1 = r_728; // @[Multiplier.scala 132:13]
  assign c53_162_io_in_2 = r_729; // @[Multiplier.scala 132:13]
  assign c53_162_io_in_3 = r_730; // @[Multiplier.scala 132:13]
  assign c53_162_io_in_4 = c53_156_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_163_io_in_0 = r_731; // @[Multiplier.scala 132:13]
  assign c53_163_io_in_1 = r_732; // @[Multiplier.scala 132:13]
  assign c53_163_io_in_2 = r_733; // @[Multiplier.scala 132:13]
  assign c53_163_io_in_3 = r_734; // @[Multiplier.scala 132:13]
  assign c53_163_io_in_4 = c53_157_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_164_io_in_0 = r_735; // @[Multiplier.scala 132:13]
  assign c53_164_io_in_1 = r_736; // @[Multiplier.scala 132:13]
  assign c53_164_io_in_2 = r_737; // @[Multiplier.scala 132:13]
  assign c53_164_io_in_3 = r_738; // @[Multiplier.scala 132:13]
  assign c53_164_io_in_4 = c53_158_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_165_io_in_0 = r_739; // @[Multiplier.scala 132:13]
  assign c53_165_io_in_1 = r_740; // @[Multiplier.scala 132:13]
  assign c53_165_io_in_2 = r_741; // @[Multiplier.scala 132:13]
  assign c53_165_io_in_3 = r_742; // @[Multiplier.scala 132:13]
  assign c53_165_io_in_4 = c53_159_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_166_io_in_0 = r_743; // @[Multiplier.scala 132:13]
  assign c53_166_io_in_1 = r_744; // @[Multiplier.scala 132:13]
  assign c53_166_io_in_2 = r_745; // @[Multiplier.scala 132:13]
  assign c53_166_io_in_3 = r_746; // @[Multiplier.scala 132:13]
  assign c53_166_io_in_4 = c53_160_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_167_io_in_0 = r_747; // @[Multiplier.scala 132:13]
  assign c53_167_io_in_1 = r_748; // @[Multiplier.scala 132:13]
  assign c53_167_io_in_2 = r_749; // @[Multiplier.scala 132:13]
  assign c53_167_io_in_3 = r_750; // @[Multiplier.scala 132:13]
  assign c53_167_io_in_4 = c53_161_io_out_1; // @[Multiplier.scala 136:41]
  assign c32_13_io_in_0 = r_751; // @[Multiplier.scala 126:19]
  assign c32_13_io_in_1 = r_752; // @[Multiplier.scala 126:19]
  assign c32_13_io_in_2 = r_753; // @[Multiplier.scala 126:19]
  assign c53_168_io_in_0 = r_754; // @[Multiplier.scala 132:13]
  assign c53_168_io_in_1 = r_755; // @[Multiplier.scala 132:13]
  assign c53_168_io_in_2 = r_756; // @[Multiplier.scala 132:13]
  assign c53_168_io_in_3 = r_757; // @[Multiplier.scala 132:13]
  assign c53_168_io_in_4 = c53_162_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_169_io_in_0 = r_758; // @[Multiplier.scala 132:13]
  assign c53_169_io_in_1 = r_759; // @[Multiplier.scala 132:13]
  assign c53_169_io_in_2 = r_760; // @[Multiplier.scala 132:13]
  assign c53_169_io_in_3 = r_761; // @[Multiplier.scala 132:13]
  assign c53_169_io_in_4 = c53_163_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_170_io_in_0 = r_762; // @[Multiplier.scala 132:13]
  assign c53_170_io_in_1 = r_763; // @[Multiplier.scala 132:13]
  assign c53_170_io_in_2 = r_764; // @[Multiplier.scala 132:13]
  assign c53_170_io_in_3 = r_765; // @[Multiplier.scala 132:13]
  assign c53_170_io_in_4 = c53_164_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_171_io_in_0 = r_766; // @[Multiplier.scala 132:13]
  assign c53_171_io_in_1 = r_767; // @[Multiplier.scala 132:13]
  assign c53_171_io_in_2 = r_768; // @[Multiplier.scala 132:13]
  assign c53_171_io_in_3 = r_769; // @[Multiplier.scala 132:13]
  assign c53_171_io_in_4 = c53_165_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_172_io_in_0 = r_770; // @[Multiplier.scala 132:13]
  assign c53_172_io_in_1 = r_771; // @[Multiplier.scala 132:13]
  assign c53_172_io_in_2 = r_772; // @[Multiplier.scala 132:13]
  assign c53_172_io_in_3 = r_773; // @[Multiplier.scala 132:13]
  assign c53_172_io_in_4 = c53_166_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_173_io_in_0 = r_774; // @[Multiplier.scala 132:13]
  assign c53_173_io_in_1 = r_775; // @[Multiplier.scala 132:13]
  assign c53_173_io_in_2 = r_776; // @[Multiplier.scala 132:13]
  assign c53_173_io_in_3 = r_777; // @[Multiplier.scala 132:13]
  assign c53_173_io_in_4 = c53_167_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_174_io_in_0 = r_778; // @[Multiplier.scala 132:13]
  assign c53_174_io_in_1 = r_779; // @[Multiplier.scala 132:13]
  assign c53_174_io_in_2 = r_780; // @[Multiplier.scala 132:13]
  assign c53_174_io_in_3 = r_781; // @[Multiplier.scala 132:13]
  assign c53_174_io_in_4 = 1'h0; // @[Multiplier.scala 134:24]
  assign c53_175_io_in_0 = r_782; // @[Multiplier.scala 132:13]
  assign c53_175_io_in_1 = r_783; // @[Multiplier.scala 132:13]
  assign c53_175_io_in_2 = r_784; // @[Multiplier.scala 132:13]
  assign c53_175_io_in_3 = r_785; // @[Multiplier.scala 132:13]
  assign c53_175_io_in_4 = c53_168_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_176_io_in_0 = r_786; // @[Multiplier.scala 132:13]
  assign c53_176_io_in_1 = r_787; // @[Multiplier.scala 132:13]
  assign c53_176_io_in_2 = r_788; // @[Multiplier.scala 132:13]
  assign c53_176_io_in_3 = r_789; // @[Multiplier.scala 132:13]
  assign c53_176_io_in_4 = c53_169_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_177_io_in_0 = r_790; // @[Multiplier.scala 132:13]
  assign c53_177_io_in_1 = r_791; // @[Multiplier.scala 132:13]
  assign c53_177_io_in_2 = r_792; // @[Multiplier.scala 132:13]
  assign c53_177_io_in_3 = r_793; // @[Multiplier.scala 132:13]
  assign c53_177_io_in_4 = c53_170_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_178_io_in_0 = r_794; // @[Multiplier.scala 132:13]
  assign c53_178_io_in_1 = r_795; // @[Multiplier.scala 132:13]
  assign c53_178_io_in_2 = r_796; // @[Multiplier.scala 132:13]
  assign c53_178_io_in_3 = r_797; // @[Multiplier.scala 132:13]
  assign c53_178_io_in_4 = c53_171_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_179_io_in_0 = r_798; // @[Multiplier.scala 132:13]
  assign c53_179_io_in_1 = r_799; // @[Multiplier.scala 132:13]
  assign c53_179_io_in_2 = r_800; // @[Multiplier.scala 132:13]
  assign c53_179_io_in_3 = r_801; // @[Multiplier.scala 132:13]
  assign c53_179_io_in_4 = c53_172_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_180_io_in_0 = r_802; // @[Multiplier.scala 132:13]
  assign c53_180_io_in_1 = r_803; // @[Multiplier.scala 132:13]
  assign c53_180_io_in_2 = r_804; // @[Multiplier.scala 132:13]
  assign c53_180_io_in_3 = r_805; // @[Multiplier.scala 132:13]
  assign c53_180_io_in_4 = c53_173_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_181_io_in_0 = r_806; // @[Multiplier.scala 132:13]
  assign c53_181_io_in_1 = r_807; // @[Multiplier.scala 132:13]
  assign c53_181_io_in_2 = r_808; // @[Multiplier.scala 132:13]
  assign c53_181_io_in_3 = r_809; // @[Multiplier.scala 132:13]
  assign c53_181_io_in_4 = c53_174_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_182_io_in_0 = r_810; // @[Multiplier.scala 132:13]
  assign c53_182_io_in_1 = r_811; // @[Multiplier.scala 132:13]
  assign c53_182_io_in_2 = r_812; // @[Multiplier.scala 132:13]
  assign c53_182_io_in_3 = r_813; // @[Multiplier.scala 132:13]
  assign c53_182_io_in_4 = c53_175_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_183_io_in_0 = r_814; // @[Multiplier.scala 132:13]
  assign c53_183_io_in_1 = r_815; // @[Multiplier.scala 132:13]
  assign c53_183_io_in_2 = r_816; // @[Multiplier.scala 132:13]
  assign c53_183_io_in_3 = r_817; // @[Multiplier.scala 132:13]
  assign c53_183_io_in_4 = c53_176_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_184_io_in_0 = r_818; // @[Multiplier.scala 132:13]
  assign c53_184_io_in_1 = r_819; // @[Multiplier.scala 132:13]
  assign c53_184_io_in_2 = r_820; // @[Multiplier.scala 132:13]
  assign c53_184_io_in_3 = r_821; // @[Multiplier.scala 132:13]
  assign c53_184_io_in_4 = c53_177_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_185_io_in_0 = r_822; // @[Multiplier.scala 132:13]
  assign c53_185_io_in_1 = r_823; // @[Multiplier.scala 132:13]
  assign c53_185_io_in_2 = r_824; // @[Multiplier.scala 132:13]
  assign c53_185_io_in_3 = r_825; // @[Multiplier.scala 132:13]
  assign c53_185_io_in_4 = c53_178_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_186_io_in_0 = r_826; // @[Multiplier.scala 132:13]
  assign c53_186_io_in_1 = r_827; // @[Multiplier.scala 132:13]
  assign c53_186_io_in_2 = r_828; // @[Multiplier.scala 132:13]
  assign c53_186_io_in_3 = r_829; // @[Multiplier.scala 132:13]
  assign c53_186_io_in_4 = c53_179_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_187_io_in_0 = r_830; // @[Multiplier.scala 132:13]
  assign c53_187_io_in_1 = r_831; // @[Multiplier.scala 132:13]
  assign c53_187_io_in_2 = r_832; // @[Multiplier.scala 132:13]
  assign c53_187_io_in_3 = r_833; // @[Multiplier.scala 132:13]
  assign c53_187_io_in_4 = c53_180_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_188_io_in_0 = r_834; // @[Multiplier.scala 132:13]
  assign c53_188_io_in_1 = r_835; // @[Multiplier.scala 132:13]
  assign c53_188_io_in_2 = r_836; // @[Multiplier.scala 132:13]
  assign c53_188_io_in_3 = r_837; // @[Multiplier.scala 132:13]
  assign c53_188_io_in_4 = c53_181_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_189_io_in_0 = r_839; // @[Multiplier.scala 132:13]
  assign c53_189_io_in_1 = r_840; // @[Multiplier.scala 132:13]
  assign c53_189_io_in_2 = r_841; // @[Multiplier.scala 132:13]
  assign c53_189_io_in_3 = r_842; // @[Multiplier.scala 132:13]
  assign c53_189_io_in_4 = c53_182_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_190_io_in_0 = r_843; // @[Multiplier.scala 132:13]
  assign c53_190_io_in_1 = r_844; // @[Multiplier.scala 132:13]
  assign c53_190_io_in_2 = r_845; // @[Multiplier.scala 132:13]
  assign c53_190_io_in_3 = r_846; // @[Multiplier.scala 132:13]
  assign c53_190_io_in_4 = c53_183_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_191_io_in_0 = r_847; // @[Multiplier.scala 132:13]
  assign c53_191_io_in_1 = r_848; // @[Multiplier.scala 132:13]
  assign c53_191_io_in_2 = r_849; // @[Multiplier.scala 132:13]
  assign c53_191_io_in_3 = r_850; // @[Multiplier.scala 132:13]
  assign c53_191_io_in_4 = c53_184_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_192_io_in_0 = r_851; // @[Multiplier.scala 132:13]
  assign c53_192_io_in_1 = r_852; // @[Multiplier.scala 132:13]
  assign c53_192_io_in_2 = r_853; // @[Multiplier.scala 132:13]
  assign c53_192_io_in_3 = r_854; // @[Multiplier.scala 132:13]
  assign c53_192_io_in_4 = c53_185_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_193_io_in_0 = r_855; // @[Multiplier.scala 132:13]
  assign c53_193_io_in_1 = r_856; // @[Multiplier.scala 132:13]
  assign c53_193_io_in_2 = r_857; // @[Multiplier.scala 132:13]
  assign c53_193_io_in_3 = r_858; // @[Multiplier.scala 132:13]
  assign c53_193_io_in_4 = c53_186_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_194_io_in_0 = r_859; // @[Multiplier.scala 132:13]
  assign c53_194_io_in_1 = r_860; // @[Multiplier.scala 132:13]
  assign c53_194_io_in_2 = r_861; // @[Multiplier.scala 132:13]
  assign c53_194_io_in_3 = r_862; // @[Multiplier.scala 132:13]
  assign c53_194_io_in_4 = c53_187_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_195_io_in_0 = r_863; // @[Multiplier.scala 132:13]
  assign c53_195_io_in_1 = r_864; // @[Multiplier.scala 132:13]
  assign c53_195_io_in_2 = r_865; // @[Multiplier.scala 132:13]
  assign c53_195_io_in_3 = r_866; // @[Multiplier.scala 132:13]
  assign c53_195_io_in_4 = c53_188_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_196_io_in_0 = r_868; // @[Multiplier.scala 132:13]
  assign c53_196_io_in_1 = r_869; // @[Multiplier.scala 132:13]
  assign c53_196_io_in_2 = r_870; // @[Multiplier.scala 132:13]
  assign c53_196_io_in_3 = r_871; // @[Multiplier.scala 132:13]
  assign c53_196_io_in_4 = c53_189_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_197_io_in_0 = r_872; // @[Multiplier.scala 132:13]
  assign c53_197_io_in_1 = r_873; // @[Multiplier.scala 132:13]
  assign c53_197_io_in_2 = r_874; // @[Multiplier.scala 132:13]
  assign c53_197_io_in_3 = r_875; // @[Multiplier.scala 132:13]
  assign c53_197_io_in_4 = c53_190_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_198_io_in_0 = r_876; // @[Multiplier.scala 132:13]
  assign c53_198_io_in_1 = r_877; // @[Multiplier.scala 132:13]
  assign c53_198_io_in_2 = r_878; // @[Multiplier.scala 132:13]
  assign c53_198_io_in_3 = r_879; // @[Multiplier.scala 132:13]
  assign c53_198_io_in_4 = c53_191_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_199_io_in_0 = r_880; // @[Multiplier.scala 132:13]
  assign c53_199_io_in_1 = r_881; // @[Multiplier.scala 132:13]
  assign c53_199_io_in_2 = r_882; // @[Multiplier.scala 132:13]
  assign c53_199_io_in_3 = r_883; // @[Multiplier.scala 132:13]
  assign c53_199_io_in_4 = c53_192_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_200_io_in_0 = r_884; // @[Multiplier.scala 132:13]
  assign c53_200_io_in_1 = r_885; // @[Multiplier.scala 132:13]
  assign c53_200_io_in_2 = r_886; // @[Multiplier.scala 132:13]
  assign c53_200_io_in_3 = r_887; // @[Multiplier.scala 132:13]
  assign c53_200_io_in_4 = c53_193_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_201_io_in_0 = r_888; // @[Multiplier.scala 132:13]
  assign c53_201_io_in_1 = r_889; // @[Multiplier.scala 132:13]
  assign c53_201_io_in_2 = r_890; // @[Multiplier.scala 132:13]
  assign c53_201_io_in_3 = r_891; // @[Multiplier.scala 132:13]
  assign c53_201_io_in_4 = c53_194_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_202_io_in_0 = r_892; // @[Multiplier.scala 132:13]
  assign c53_202_io_in_1 = r_893; // @[Multiplier.scala 132:13]
  assign c53_202_io_in_2 = r_894; // @[Multiplier.scala 132:13]
  assign c53_202_io_in_3 = r_895; // @[Multiplier.scala 132:13]
  assign c53_202_io_in_4 = c53_195_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_14_io_in_0 = r_896; // @[Multiplier.scala 121:19]
  assign c22_14_io_in_1 = r_897; // @[Multiplier.scala 121:19]
  assign c53_203_io_in_0 = r_898; // @[Multiplier.scala 132:13]
  assign c53_203_io_in_1 = r_899; // @[Multiplier.scala 132:13]
  assign c53_203_io_in_2 = r_900; // @[Multiplier.scala 132:13]
  assign c53_203_io_in_3 = r_901; // @[Multiplier.scala 132:13]
  assign c53_203_io_in_4 = c53_196_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_204_io_in_0 = r_902; // @[Multiplier.scala 132:13]
  assign c53_204_io_in_1 = r_903; // @[Multiplier.scala 132:13]
  assign c53_204_io_in_2 = r_904; // @[Multiplier.scala 132:13]
  assign c53_204_io_in_3 = r_905; // @[Multiplier.scala 132:13]
  assign c53_204_io_in_4 = c53_197_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_205_io_in_0 = r_906; // @[Multiplier.scala 132:13]
  assign c53_205_io_in_1 = r_907; // @[Multiplier.scala 132:13]
  assign c53_205_io_in_2 = r_908; // @[Multiplier.scala 132:13]
  assign c53_205_io_in_3 = r_909; // @[Multiplier.scala 132:13]
  assign c53_205_io_in_4 = c53_198_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_206_io_in_0 = r_910; // @[Multiplier.scala 132:13]
  assign c53_206_io_in_1 = r_911; // @[Multiplier.scala 132:13]
  assign c53_206_io_in_2 = r_912; // @[Multiplier.scala 132:13]
  assign c53_206_io_in_3 = r_913; // @[Multiplier.scala 132:13]
  assign c53_206_io_in_4 = c53_199_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_207_io_in_0 = r_914; // @[Multiplier.scala 132:13]
  assign c53_207_io_in_1 = r_915; // @[Multiplier.scala 132:13]
  assign c53_207_io_in_2 = r_916; // @[Multiplier.scala 132:13]
  assign c53_207_io_in_3 = r_917; // @[Multiplier.scala 132:13]
  assign c53_207_io_in_4 = c53_200_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_208_io_in_0 = r_918; // @[Multiplier.scala 132:13]
  assign c53_208_io_in_1 = r_919; // @[Multiplier.scala 132:13]
  assign c53_208_io_in_2 = r_920; // @[Multiplier.scala 132:13]
  assign c53_208_io_in_3 = r_921; // @[Multiplier.scala 132:13]
  assign c53_208_io_in_4 = c53_201_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_209_io_in_0 = r_922; // @[Multiplier.scala 132:13]
  assign c53_209_io_in_1 = r_923; // @[Multiplier.scala 132:13]
  assign c53_209_io_in_2 = r_924; // @[Multiplier.scala 132:13]
  assign c53_209_io_in_3 = r_925; // @[Multiplier.scala 132:13]
  assign c53_209_io_in_4 = c53_202_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_15_io_in_0 = r_926; // @[Multiplier.scala 121:19]
  assign c22_15_io_in_1 = r_927; // @[Multiplier.scala 121:19]
  assign c53_210_io_in_0 = r_928; // @[Multiplier.scala 132:13]
  assign c53_210_io_in_1 = r_929; // @[Multiplier.scala 132:13]
  assign c53_210_io_in_2 = r_930; // @[Multiplier.scala 132:13]
  assign c53_210_io_in_3 = r_931; // @[Multiplier.scala 132:13]
  assign c53_210_io_in_4 = c53_203_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_211_io_in_0 = r_932; // @[Multiplier.scala 132:13]
  assign c53_211_io_in_1 = r_933; // @[Multiplier.scala 132:13]
  assign c53_211_io_in_2 = r_934; // @[Multiplier.scala 132:13]
  assign c53_211_io_in_3 = r_935; // @[Multiplier.scala 132:13]
  assign c53_211_io_in_4 = c53_204_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_212_io_in_0 = r_936; // @[Multiplier.scala 132:13]
  assign c53_212_io_in_1 = r_937; // @[Multiplier.scala 132:13]
  assign c53_212_io_in_2 = r_938; // @[Multiplier.scala 132:13]
  assign c53_212_io_in_3 = r_939; // @[Multiplier.scala 132:13]
  assign c53_212_io_in_4 = c53_205_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_213_io_in_0 = r_940; // @[Multiplier.scala 132:13]
  assign c53_213_io_in_1 = r_941; // @[Multiplier.scala 132:13]
  assign c53_213_io_in_2 = r_942; // @[Multiplier.scala 132:13]
  assign c53_213_io_in_3 = r_943; // @[Multiplier.scala 132:13]
  assign c53_213_io_in_4 = c53_206_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_214_io_in_0 = r_944; // @[Multiplier.scala 132:13]
  assign c53_214_io_in_1 = r_945; // @[Multiplier.scala 132:13]
  assign c53_214_io_in_2 = r_946; // @[Multiplier.scala 132:13]
  assign c53_214_io_in_3 = r_947; // @[Multiplier.scala 132:13]
  assign c53_214_io_in_4 = c53_207_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_215_io_in_0 = r_948; // @[Multiplier.scala 132:13]
  assign c53_215_io_in_1 = r_949; // @[Multiplier.scala 132:13]
  assign c53_215_io_in_2 = r_950; // @[Multiplier.scala 132:13]
  assign c53_215_io_in_3 = r_951; // @[Multiplier.scala 132:13]
  assign c53_215_io_in_4 = c53_208_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_216_io_in_0 = r_952; // @[Multiplier.scala 132:13]
  assign c53_216_io_in_1 = r_953; // @[Multiplier.scala 132:13]
  assign c53_216_io_in_2 = r_954; // @[Multiplier.scala 132:13]
  assign c53_216_io_in_3 = r_955; // @[Multiplier.scala 132:13]
  assign c53_216_io_in_4 = c53_209_io_out_1; // @[Multiplier.scala 136:41]
  assign c32_14_io_in_0 = r_956; // @[Multiplier.scala 126:19]
  assign c32_14_io_in_1 = r_957; // @[Multiplier.scala 126:19]
  assign c32_14_io_in_2 = r_958; // @[Multiplier.scala 126:19]
  assign c53_217_io_in_0 = r_959; // @[Multiplier.scala 132:13]
  assign c53_217_io_in_1 = r_960; // @[Multiplier.scala 132:13]
  assign c53_217_io_in_2 = r_961; // @[Multiplier.scala 132:13]
  assign c53_217_io_in_3 = r_962; // @[Multiplier.scala 132:13]
  assign c53_217_io_in_4 = c53_210_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_218_io_in_0 = r_963; // @[Multiplier.scala 132:13]
  assign c53_218_io_in_1 = r_964; // @[Multiplier.scala 132:13]
  assign c53_218_io_in_2 = r_965; // @[Multiplier.scala 132:13]
  assign c53_218_io_in_3 = r_966; // @[Multiplier.scala 132:13]
  assign c53_218_io_in_4 = c53_211_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_219_io_in_0 = r_967; // @[Multiplier.scala 132:13]
  assign c53_219_io_in_1 = r_968; // @[Multiplier.scala 132:13]
  assign c53_219_io_in_2 = r_969; // @[Multiplier.scala 132:13]
  assign c53_219_io_in_3 = r_970; // @[Multiplier.scala 132:13]
  assign c53_219_io_in_4 = c53_212_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_220_io_in_0 = r_971; // @[Multiplier.scala 132:13]
  assign c53_220_io_in_1 = r_972; // @[Multiplier.scala 132:13]
  assign c53_220_io_in_2 = r_973; // @[Multiplier.scala 132:13]
  assign c53_220_io_in_3 = r_974; // @[Multiplier.scala 132:13]
  assign c53_220_io_in_4 = c53_213_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_221_io_in_0 = r_975; // @[Multiplier.scala 132:13]
  assign c53_221_io_in_1 = r_976; // @[Multiplier.scala 132:13]
  assign c53_221_io_in_2 = r_977; // @[Multiplier.scala 132:13]
  assign c53_221_io_in_3 = r_978; // @[Multiplier.scala 132:13]
  assign c53_221_io_in_4 = c53_214_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_222_io_in_0 = r_979; // @[Multiplier.scala 132:13]
  assign c53_222_io_in_1 = r_980; // @[Multiplier.scala 132:13]
  assign c53_222_io_in_2 = r_981; // @[Multiplier.scala 132:13]
  assign c53_222_io_in_3 = r_982; // @[Multiplier.scala 132:13]
  assign c53_222_io_in_4 = c53_215_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_223_io_in_0 = r_983; // @[Multiplier.scala 132:13]
  assign c53_223_io_in_1 = r_984; // @[Multiplier.scala 132:13]
  assign c53_223_io_in_2 = r_985; // @[Multiplier.scala 132:13]
  assign c53_223_io_in_3 = r_986; // @[Multiplier.scala 132:13]
  assign c53_223_io_in_4 = c53_216_io_out_1; // @[Multiplier.scala 136:41]
  assign c32_15_io_in_0 = r_987; // @[Multiplier.scala 126:19]
  assign c32_15_io_in_1 = r_988; // @[Multiplier.scala 126:19]
  assign c32_15_io_in_2 = r_989; // @[Multiplier.scala 126:19]
  assign c53_224_io_in_0 = r_990; // @[Multiplier.scala 132:13]
  assign c53_224_io_in_1 = r_991; // @[Multiplier.scala 132:13]
  assign c53_224_io_in_2 = r_992; // @[Multiplier.scala 132:13]
  assign c53_224_io_in_3 = r_993; // @[Multiplier.scala 132:13]
  assign c53_224_io_in_4 = c53_217_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_225_io_in_0 = r_994; // @[Multiplier.scala 132:13]
  assign c53_225_io_in_1 = r_995; // @[Multiplier.scala 132:13]
  assign c53_225_io_in_2 = r_996; // @[Multiplier.scala 132:13]
  assign c53_225_io_in_3 = r_997; // @[Multiplier.scala 132:13]
  assign c53_225_io_in_4 = c53_218_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_226_io_in_0 = r_998; // @[Multiplier.scala 132:13]
  assign c53_226_io_in_1 = r_999; // @[Multiplier.scala 132:13]
  assign c53_226_io_in_2 = r_1000; // @[Multiplier.scala 132:13]
  assign c53_226_io_in_3 = r_1001; // @[Multiplier.scala 132:13]
  assign c53_226_io_in_4 = c53_219_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_227_io_in_0 = r_1002; // @[Multiplier.scala 132:13]
  assign c53_227_io_in_1 = r_1003; // @[Multiplier.scala 132:13]
  assign c53_227_io_in_2 = r_1004; // @[Multiplier.scala 132:13]
  assign c53_227_io_in_3 = r_1005; // @[Multiplier.scala 132:13]
  assign c53_227_io_in_4 = c53_220_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_228_io_in_0 = r_1006; // @[Multiplier.scala 132:13]
  assign c53_228_io_in_1 = r_1007; // @[Multiplier.scala 132:13]
  assign c53_228_io_in_2 = r_1008; // @[Multiplier.scala 132:13]
  assign c53_228_io_in_3 = r_1009; // @[Multiplier.scala 132:13]
  assign c53_228_io_in_4 = c53_221_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_229_io_in_0 = r_1010; // @[Multiplier.scala 132:13]
  assign c53_229_io_in_1 = r_1011; // @[Multiplier.scala 132:13]
  assign c53_229_io_in_2 = r_1012; // @[Multiplier.scala 132:13]
  assign c53_229_io_in_3 = r_1013; // @[Multiplier.scala 132:13]
  assign c53_229_io_in_4 = c53_222_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_230_io_in_0 = r_1014; // @[Multiplier.scala 132:13]
  assign c53_230_io_in_1 = r_1015; // @[Multiplier.scala 132:13]
  assign c53_230_io_in_2 = r_1016; // @[Multiplier.scala 132:13]
  assign c53_230_io_in_3 = r_1017; // @[Multiplier.scala 132:13]
  assign c53_230_io_in_4 = c53_223_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_231_io_in_0 = r_1018; // @[Multiplier.scala 132:13]
  assign c53_231_io_in_1 = r_1019; // @[Multiplier.scala 132:13]
  assign c53_231_io_in_2 = r_1020; // @[Multiplier.scala 132:13]
  assign c53_231_io_in_3 = r_1021; // @[Multiplier.scala 132:13]
  assign c53_231_io_in_4 = 1'h0; // @[Multiplier.scala 134:24]
  assign c53_232_io_in_0 = r_1022; // @[Multiplier.scala 132:13]
  assign c53_232_io_in_1 = r_1023; // @[Multiplier.scala 132:13]
  assign c53_232_io_in_2 = r_1024; // @[Multiplier.scala 132:13]
  assign c53_232_io_in_3 = r_1025; // @[Multiplier.scala 132:13]
  assign c53_232_io_in_4 = c53_224_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_233_io_in_0 = r_1026; // @[Multiplier.scala 132:13]
  assign c53_233_io_in_1 = r_1027; // @[Multiplier.scala 132:13]
  assign c53_233_io_in_2 = r_1028; // @[Multiplier.scala 132:13]
  assign c53_233_io_in_3 = r_1029; // @[Multiplier.scala 132:13]
  assign c53_233_io_in_4 = c53_225_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_234_io_in_0 = r_1030; // @[Multiplier.scala 132:13]
  assign c53_234_io_in_1 = r_1031; // @[Multiplier.scala 132:13]
  assign c53_234_io_in_2 = r_1032; // @[Multiplier.scala 132:13]
  assign c53_234_io_in_3 = r_1033; // @[Multiplier.scala 132:13]
  assign c53_234_io_in_4 = c53_226_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_235_io_in_0 = r_1034; // @[Multiplier.scala 132:13]
  assign c53_235_io_in_1 = r_1035; // @[Multiplier.scala 132:13]
  assign c53_235_io_in_2 = r_1036; // @[Multiplier.scala 132:13]
  assign c53_235_io_in_3 = r_1037; // @[Multiplier.scala 132:13]
  assign c53_235_io_in_4 = c53_227_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_236_io_in_0 = r_1038; // @[Multiplier.scala 132:13]
  assign c53_236_io_in_1 = r_1039; // @[Multiplier.scala 132:13]
  assign c53_236_io_in_2 = r_1040; // @[Multiplier.scala 132:13]
  assign c53_236_io_in_3 = r_1041; // @[Multiplier.scala 132:13]
  assign c53_236_io_in_4 = c53_228_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_237_io_in_0 = r_1042; // @[Multiplier.scala 132:13]
  assign c53_237_io_in_1 = r_1043; // @[Multiplier.scala 132:13]
  assign c53_237_io_in_2 = r_1044; // @[Multiplier.scala 132:13]
  assign c53_237_io_in_3 = r_1045; // @[Multiplier.scala 132:13]
  assign c53_237_io_in_4 = c53_229_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_238_io_in_0 = r_1046; // @[Multiplier.scala 132:13]
  assign c53_238_io_in_1 = r_1047; // @[Multiplier.scala 132:13]
  assign c53_238_io_in_2 = r_1048; // @[Multiplier.scala 132:13]
  assign c53_238_io_in_3 = r_1049; // @[Multiplier.scala 132:13]
  assign c53_238_io_in_4 = c53_230_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_239_io_in_0 = r_1050; // @[Multiplier.scala 132:13]
  assign c53_239_io_in_1 = r_1051; // @[Multiplier.scala 132:13]
  assign c53_239_io_in_2 = r_1052; // @[Multiplier.scala 132:13]
  assign c53_239_io_in_3 = r_1053; // @[Multiplier.scala 132:13]
  assign c53_239_io_in_4 = c53_231_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_240_io_in_0 = r_1054; // @[Multiplier.scala 132:13]
  assign c53_240_io_in_1 = r_1055; // @[Multiplier.scala 132:13]
  assign c53_240_io_in_2 = r_1056; // @[Multiplier.scala 132:13]
  assign c53_240_io_in_3 = r_1057; // @[Multiplier.scala 132:13]
  assign c53_240_io_in_4 = c53_232_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_241_io_in_0 = r_1058; // @[Multiplier.scala 132:13]
  assign c53_241_io_in_1 = r_1059; // @[Multiplier.scala 132:13]
  assign c53_241_io_in_2 = r_1060; // @[Multiplier.scala 132:13]
  assign c53_241_io_in_3 = r_1061; // @[Multiplier.scala 132:13]
  assign c53_241_io_in_4 = c53_233_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_242_io_in_0 = r_1062; // @[Multiplier.scala 132:13]
  assign c53_242_io_in_1 = r_1063; // @[Multiplier.scala 132:13]
  assign c53_242_io_in_2 = r_1064; // @[Multiplier.scala 132:13]
  assign c53_242_io_in_3 = r_1065; // @[Multiplier.scala 132:13]
  assign c53_242_io_in_4 = c53_234_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_243_io_in_0 = r_1066; // @[Multiplier.scala 132:13]
  assign c53_243_io_in_1 = r_1067; // @[Multiplier.scala 132:13]
  assign c53_243_io_in_2 = r_1068; // @[Multiplier.scala 132:13]
  assign c53_243_io_in_3 = r_1069; // @[Multiplier.scala 132:13]
  assign c53_243_io_in_4 = c53_235_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_244_io_in_0 = r_1070; // @[Multiplier.scala 132:13]
  assign c53_244_io_in_1 = r_1071; // @[Multiplier.scala 132:13]
  assign c53_244_io_in_2 = r_1072; // @[Multiplier.scala 132:13]
  assign c53_244_io_in_3 = r_1073; // @[Multiplier.scala 132:13]
  assign c53_244_io_in_4 = c53_236_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_245_io_in_0 = r_1074; // @[Multiplier.scala 132:13]
  assign c53_245_io_in_1 = r_1075; // @[Multiplier.scala 132:13]
  assign c53_245_io_in_2 = r_1076; // @[Multiplier.scala 132:13]
  assign c53_245_io_in_3 = r_1077; // @[Multiplier.scala 132:13]
  assign c53_245_io_in_4 = c53_237_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_246_io_in_0 = r_1078; // @[Multiplier.scala 132:13]
  assign c53_246_io_in_1 = r_1079; // @[Multiplier.scala 132:13]
  assign c53_246_io_in_2 = r_1080; // @[Multiplier.scala 132:13]
  assign c53_246_io_in_3 = r_1081; // @[Multiplier.scala 132:13]
  assign c53_246_io_in_4 = c53_238_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_247_io_in_0 = r_1082; // @[Multiplier.scala 132:13]
  assign c53_247_io_in_1 = r_1083; // @[Multiplier.scala 132:13]
  assign c53_247_io_in_2 = r_1084; // @[Multiplier.scala 132:13]
  assign c53_247_io_in_3 = r_1085; // @[Multiplier.scala 132:13]
  assign c53_247_io_in_4 = c53_239_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_248_io_in_0 = r_1087; // @[Multiplier.scala 132:13]
  assign c53_248_io_in_1 = r_1088; // @[Multiplier.scala 132:13]
  assign c53_248_io_in_2 = r_1089; // @[Multiplier.scala 132:13]
  assign c53_248_io_in_3 = r_1090; // @[Multiplier.scala 132:13]
  assign c53_248_io_in_4 = c53_240_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_249_io_in_0 = r_1091; // @[Multiplier.scala 132:13]
  assign c53_249_io_in_1 = r_1092; // @[Multiplier.scala 132:13]
  assign c53_249_io_in_2 = r_1093; // @[Multiplier.scala 132:13]
  assign c53_249_io_in_3 = r_1094; // @[Multiplier.scala 132:13]
  assign c53_249_io_in_4 = c53_241_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_250_io_in_0 = r_1095; // @[Multiplier.scala 132:13]
  assign c53_250_io_in_1 = r_1096; // @[Multiplier.scala 132:13]
  assign c53_250_io_in_2 = r_1097; // @[Multiplier.scala 132:13]
  assign c53_250_io_in_3 = r_1098; // @[Multiplier.scala 132:13]
  assign c53_250_io_in_4 = c53_242_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_251_io_in_0 = r_1099; // @[Multiplier.scala 132:13]
  assign c53_251_io_in_1 = r_1100; // @[Multiplier.scala 132:13]
  assign c53_251_io_in_2 = r_1101; // @[Multiplier.scala 132:13]
  assign c53_251_io_in_3 = r_1102; // @[Multiplier.scala 132:13]
  assign c53_251_io_in_4 = c53_243_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_252_io_in_0 = r_1103; // @[Multiplier.scala 132:13]
  assign c53_252_io_in_1 = r_1104; // @[Multiplier.scala 132:13]
  assign c53_252_io_in_2 = r_1105; // @[Multiplier.scala 132:13]
  assign c53_252_io_in_3 = r_1106; // @[Multiplier.scala 132:13]
  assign c53_252_io_in_4 = c53_244_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_253_io_in_0 = r_1107; // @[Multiplier.scala 132:13]
  assign c53_253_io_in_1 = r_1108; // @[Multiplier.scala 132:13]
  assign c53_253_io_in_2 = r_1109; // @[Multiplier.scala 132:13]
  assign c53_253_io_in_3 = r_1110; // @[Multiplier.scala 132:13]
  assign c53_253_io_in_4 = c53_245_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_254_io_in_0 = r_1111; // @[Multiplier.scala 132:13]
  assign c53_254_io_in_1 = r_1112; // @[Multiplier.scala 132:13]
  assign c53_254_io_in_2 = r_1113; // @[Multiplier.scala 132:13]
  assign c53_254_io_in_3 = r_1114; // @[Multiplier.scala 132:13]
  assign c53_254_io_in_4 = c53_246_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_255_io_in_0 = r_1115; // @[Multiplier.scala 132:13]
  assign c53_255_io_in_1 = r_1116; // @[Multiplier.scala 132:13]
  assign c53_255_io_in_2 = r_1117; // @[Multiplier.scala 132:13]
  assign c53_255_io_in_3 = r_1118; // @[Multiplier.scala 132:13]
  assign c53_255_io_in_4 = c53_247_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_256_io_in_0 = r_1120; // @[Multiplier.scala 132:13]
  assign c53_256_io_in_1 = r_1121; // @[Multiplier.scala 132:13]
  assign c53_256_io_in_2 = r_1122; // @[Multiplier.scala 132:13]
  assign c53_256_io_in_3 = r_1123; // @[Multiplier.scala 132:13]
  assign c53_256_io_in_4 = c53_248_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_257_io_in_0 = r_1124; // @[Multiplier.scala 132:13]
  assign c53_257_io_in_1 = r_1125; // @[Multiplier.scala 132:13]
  assign c53_257_io_in_2 = r_1126; // @[Multiplier.scala 132:13]
  assign c53_257_io_in_3 = r_1127; // @[Multiplier.scala 132:13]
  assign c53_257_io_in_4 = c53_249_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_258_io_in_0 = r_1128; // @[Multiplier.scala 132:13]
  assign c53_258_io_in_1 = r_1129; // @[Multiplier.scala 132:13]
  assign c53_258_io_in_2 = r_1130; // @[Multiplier.scala 132:13]
  assign c53_258_io_in_3 = r_1131; // @[Multiplier.scala 132:13]
  assign c53_258_io_in_4 = c53_250_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_259_io_in_0 = r_1132; // @[Multiplier.scala 132:13]
  assign c53_259_io_in_1 = r_1133; // @[Multiplier.scala 132:13]
  assign c53_259_io_in_2 = r_1134; // @[Multiplier.scala 132:13]
  assign c53_259_io_in_3 = r_1135; // @[Multiplier.scala 132:13]
  assign c53_259_io_in_4 = c53_251_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_260_io_in_0 = r_1136; // @[Multiplier.scala 132:13]
  assign c53_260_io_in_1 = r_1137; // @[Multiplier.scala 132:13]
  assign c53_260_io_in_2 = r_1138; // @[Multiplier.scala 132:13]
  assign c53_260_io_in_3 = r_1139; // @[Multiplier.scala 132:13]
  assign c53_260_io_in_4 = c53_252_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_261_io_in_0 = r_1140; // @[Multiplier.scala 132:13]
  assign c53_261_io_in_1 = r_1141; // @[Multiplier.scala 132:13]
  assign c53_261_io_in_2 = r_1142; // @[Multiplier.scala 132:13]
  assign c53_261_io_in_3 = r_1143; // @[Multiplier.scala 132:13]
  assign c53_261_io_in_4 = c53_253_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_262_io_in_0 = r_1144; // @[Multiplier.scala 132:13]
  assign c53_262_io_in_1 = r_1145; // @[Multiplier.scala 132:13]
  assign c53_262_io_in_2 = r_1146; // @[Multiplier.scala 132:13]
  assign c53_262_io_in_3 = r_1147; // @[Multiplier.scala 132:13]
  assign c53_262_io_in_4 = c53_254_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_263_io_in_0 = r_1148; // @[Multiplier.scala 132:13]
  assign c53_263_io_in_1 = r_1149; // @[Multiplier.scala 132:13]
  assign c53_263_io_in_2 = r_1150; // @[Multiplier.scala 132:13]
  assign c53_263_io_in_3 = r_1151; // @[Multiplier.scala 132:13]
  assign c53_263_io_in_4 = c53_255_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_264_io_in_0 = r_1153; // @[Multiplier.scala 132:13]
  assign c53_264_io_in_1 = r_1154; // @[Multiplier.scala 132:13]
  assign c53_264_io_in_2 = r_1155; // @[Multiplier.scala 132:13]
  assign c53_264_io_in_3 = r_1156; // @[Multiplier.scala 132:13]
  assign c53_264_io_in_4 = c53_256_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_265_io_in_0 = r_1157; // @[Multiplier.scala 132:13]
  assign c53_265_io_in_1 = r_1158; // @[Multiplier.scala 132:13]
  assign c53_265_io_in_2 = r_1159; // @[Multiplier.scala 132:13]
  assign c53_265_io_in_3 = r_1160; // @[Multiplier.scala 132:13]
  assign c53_265_io_in_4 = c53_257_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_266_io_in_0 = r_1161; // @[Multiplier.scala 132:13]
  assign c53_266_io_in_1 = r_1162; // @[Multiplier.scala 132:13]
  assign c53_266_io_in_2 = r_1163; // @[Multiplier.scala 132:13]
  assign c53_266_io_in_3 = r_1164; // @[Multiplier.scala 132:13]
  assign c53_266_io_in_4 = c53_258_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_267_io_in_0 = r_1165; // @[Multiplier.scala 132:13]
  assign c53_267_io_in_1 = r_1166; // @[Multiplier.scala 132:13]
  assign c53_267_io_in_2 = r_1167; // @[Multiplier.scala 132:13]
  assign c53_267_io_in_3 = r_1168; // @[Multiplier.scala 132:13]
  assign c53_267_io_in_4 = c53_259_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_268_io_in_0 = r_1169; // @[Multiplier.scala 132:13]
  assign c53_268_io_in_1 = r_1170; // @[Multiplier.scala 132:13]
  assign c53_268_io_in_2 = r_1171; // @[Multiplier.scala 132:13]
  assign c53_268_io_in_3 = r_1172; // @[Multiplier.scala 132:13]
  assign c53_268_io_in_4 = c53_260_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_269_io_in_0 = r_1173; // @[Multiplier.scala 132:13]
  assign c53_269_io_in_1 = r_1174; // @[Multiplier.scala 132:13]
  assign c53_269_io_in_2 = r_1175; // @[Multiplier.scala 132:13]
  assign c53_269_io_in_3 = r_1176; // @[Multiplier.scala 132:13]
  assign c53_269_io_in_4 = c53_261_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_270_io_in_0 = r_1177; // @[Multiplier.scala 132:13]
  assign c53_270_io_in_1 = r_1178; // @[Multiplier.scala 132:13]
  assign c53_270_io_in_2 = r_1179; // @[Multiplier.scala 132:13]
  assign c53_270_io_in_3 = r_1180; // @[Multiplier.scala 132:13]
  assign c53_270_io_in_4 = c53_262_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_271_io_in_0 = r_1181; // @[Multiplier.scala 132:13]
  assign c53_271_io_in_1 = r_1182; // @[Multiplier.scala 132:13]
  assign c53_271_io_in_2 = r_1183; // @[Multiplier.scala 132:13]
  assign c53_271_io_in_3 = r_1184; // @[Multiplier.scala 132:13]
  assign c53_271_io_in_4 = c53_263_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_272_io_in_0 = r_1186; // @[Multiplier.scala 132:13]
  assign c53_272_io_in_1 = r_1187; // @[Multiplier.scala 132:13]
  assign c53_272_io_in_2 = r_1188; // @[Multiplier.scala 132:13]
  assign c53_272_io_in_3 = r_1189; // @[Multiplier.scala 132:13]
  assign c53_272_io_in_4 = c53_264_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_273_io_in_0 = r_1190; // @[Multiplier.scala 132:13]
  assign c53_273_io_in_1 = r_1191; // @[Multiplier.scala 132:13]
  assign c53_273_io_in_2 = r_1192; // @[Multiplier.scala 132:13]
  assign c53_273_io_in_3 = r_1193; // @[Multiplier.scala 132:13]
  assign c53_273_io_in_4 = c53_265_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_274_io_in_0 = r_1194; // @[Multiplier.scala 132:13]
  assign c53_274_io_in_1 = r_1195; // @[Multiplier.scala 132:13]
  assign c53_274_io_in_2 = r_1196; // @[Multiplier.scala 132:13]
  assign c53_274_io_in_3 = r_1197; // @[Multiplier.scala 132:13]
  assign c53_274_io_in_4 = c53_266_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_275_io_in_0 = r_1198; // @[Multiplier.scala 132:13]
  assign c53_275_io_in_1 = r_1199; // @[Multiplier.scala 132:13]
  assign c53_275_io_in_2 = r_1200; // @[Multiplier.scala 132:13]
  assign c53_275_io_in_3 = r_1201; // @[Multiplier.scala 132:13]
  assign c53_275_io_in_4 = c53_267_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_276_io_in_0 = r_1202; // @[Multiplier.scala 132:13]
  assign c53_276_io_in_1 = r_1203; // @[Multiplier.scala 132:13]
  assign c53_276_io_in_2 = r_1204; // @[Multiplier.scala 132:13]
  assign c53_276_io_in_3 = r_1205; // @[Multiplier.scala 132:13]
  assign c53_276_io_in_4 = c53_268_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_277_io_in_0 = r_1206; // @[Multiplier.scala 132:13]
  assign c53_277_io_in_1 = r_1207; // @[Multiplier.scala 132:13]
  assign c53_277_io_in_2 = r_1208; // @[Multiplier.scala 132:13]
  assign c53_277_io_in_3 = r_1209; // @[Multiplier.scala 132:13]
  assign c53_277_io_in_4 = c53_269_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_278_io_in_0 = r_1210; // @[Multiplier.scala 132:13]
  assign c53_278_io_in_1 = r_1211; // @[Multiplier.scala 132:13]
  assign c53_278_io_in_2 = r_1212; // @[Multiplier.scala 132:13]
  assign c53_278_io_in_3 = r_1213; // @[Multiplier.scala 132:13]
  assign c53_278_io_in_4 = c53_270_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_279_io_in_0 = r_1214; // @[Multiplier.scala 132:13]
  assign c53_279_io_in_1 = r_1215; // @[Multiplier.scala 132:13]
  assign c53_279_io_in_2 = r_1216; // @[Multiplier.scala 132:13]
  assign c53_279_io_in_3 = r_1217; // @[Multiplier.scala 132:13]
  assign c53_279_io_in_4 = c53_271_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_280_io_in_0 = r_1219; // @[Multiplier.scala 132:13]
  assign c53_280_io_in_1 = r_1220; // @[Multiplier.scala 132:13]
  assign c53_280_io_in_2 = r_1221; // @[Multiplier.scala 132:13]
  assign c53_280_io_in_3 = r_1222; // @[Multiplier.scala 132:13]
  assign c53_280_io_in_4 = c53_272_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_281_io_in_0 = r_1223; // @[Multiplier.scala 132:13]
  assign c53_281_io_in_1 = r_1224; // @[Multiplier.scala 132:13]
  assign c53_281_io_in_2 = r_1225; // @[Multiplier.scala 132:13]
  assign c53_281_io_in_3 = r_1226; // @[Multiplier.scala 132:13]
  assign c53_281_io_in_4 = c53_273_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_282_io_in_0 = r_1227; // @[Multiplier.scala 132:13]
  assign c53_282_io_in_1 = r_1228; // @[Multiplier.scala 132:13]
  assign c53_282_io_in_2 = r_1229; // @[Multiplier.scala 132:13]
  assign c53_282_io_in_3 = r_1230; // @[Multiplier.scala 132:13]
  assign c53_282_io_in_4 = c53_274_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_283_io_in_0 = r_1231; // @[Multiplier.scala 132:13]
  assign c53_283_io_in_1 = r_1232; // @[Multiplier.scala 132:13]
  assign c53_283_io_in_2 = r_1233; // @[Multiplier.scala 132:13]
  assign c53_283_io_in_3 = r_1234; // @[Multiplier.scala 132:13]
  assign c53_283_io_in_4 = c53_275_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_284_io_in_0 = r_1235; // @[Multiplier.scala 132:13]
  assign c53_284_io_in_1 = r_1236; // @[Multiplier.scala 132:13]
  assign c53_284_io_in_2 = r_1237; // @[Multiplier.scala 132:13]
  assign c53_284_io_in_3 = r_1238; // @[Multiplier.scala 132:13]
  assign c53_284_io_in_4 = c53_276_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_285_io_in_0 = r_1239; // @[Multiplier.scala 132:13]
  assign c53_285_io_in_1 = r_1240; // @[Multiplier.scala 132:13]
  assign c53_285_io_in_2 = r_1241; // @[Multiplier.scala 132:13]
  assign c53_285_io_in_3 = r_1242; // @[Multiplier.scala 132:13]
  assign c53_285_io_in_4 = c53_277_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_286_io_in_0 = r_1243; // @[Multiplier.scala 132:13]
  assign c53_286_io_in_1 = r_1244; // @[Multiplier.scala 132:13]
  assign c53_286_io_in_2 = r_1245; // @[Multiplier.scala 132:13]
  assign c53_286_io_in_3 = r_1246; // @[Multiplier.scala 132:13]
  assign c53_286_io_in_4 = c53_278_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_287_io_in_0 = r_1247; // @[Multiplier.scala 132:13]
  assign c53_287_io_in_1 = r_1248; // @[Multiplier.scala 132:13]
  assign c53_287_io_in_2 = r_1249; // @[Multiplier.scala 132:13]
  assign c53_287_io_in_3 = r_1250; // @[Multiplier.scala 132:13]
  assign c53_287_io_in_4 = c53_279_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_288_io_in_0 = r_1252; // @[Multiplier.scala 132:13]
  assign c53_288_io_in_1 = r_1253; // @[Multiplier.scala 132:13]
  assign c53_288_io_in_2 = r_1254; // @[Multiplier.scala 132:13]
  assign c53_288_io_in_3 = r_1255; // @[Multiplier.scala 132:13]
  assign c53_288_io_in_4 = c53_280_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_289_io_in_0 = r_1256; // @[Multiplier.scala 132:13]
  assign c53_289_io_in_1 = r_1257; // @[Multiplier.scala 132:13]
  assign c53_289_io_in_2 = r_1258; // @[Multiplier.scala 132:13]
  assign c53_289_io_in_3 = r_1259; // @[Multiplier.scala 132:13]
  assign c53_289_io_in_4 = c53_281_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_290_io_in_0 = r_1260; // @[Multiplier.scala 132:13]
  assign c53_290_io_in_1 = r_1261; // @[Multiplier.scala 132:13]
  assign c53_290_io_in_2 = r_1262; // @[Multiplier.scala 132:13]
  assign c53_290_io_in_3 = r_1263; // @[Multiplier.scala 132:13]
  assign c53_290_io_in_4 = c53_282_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_291_io_in_0 = r_1264; // @[Multiplier.scala 132:13]
  assign c53_291_io_in_1 = r_1265; // @[Multiplier.scala 132:13]
  assign c53_291_io_in_2 = r_1266; // @[Multiplier.scala 132:13]
  assign c53_291_io_in_3 = r_1267; // @[Multiplier.scala 132:13]
  assign c53_291_io_in_4 = c53_283_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_292_io_in_0 = r_1268; // @[Multiplier.scala 132:13]
  assign c53_292_io_in_1 = r_1269; // @[Multiplier.scala 132:13]
  assign c53_292_io_in_2 = r_1270; // @[Multiplier.scala 132:13]
  assign c53_292_io_in_3 = r_1271; // @[Multiplier.scala 132:13]
  assign c53_292_io_in_4 = c53_284_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_293_io_in_0 = r_1272; // @[Multiplier.scala 132:13]
  assign c53_293_io_in_1 = r_1273; // @[Multiplier.scala 132:13]
  assign c53_293_io_in_2 = r_1274; // @[Multiplier.scala 132:13]
  assign c53_293_io_in_3 = r_1275; // @[Multiplier.scala 132:13]
  assign c53_293_io_in_4 = c53_285_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_294_io_in_0 = r_1276; // @[Multiplier.scala 132:13]
  assign c53_294_io_in_1 = r_1277; // @[Multiplier.scala 132:13]
  assign c53_294_io_in_2 = r_1278; // @[Multiplier.scala 132:13]
  assign c53_294_io_in_3 = r_1279; // @[Multiplier.scala 132:13]
  assign c53_294_io_in_4 = c53_286_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_295_io_in_0 = r_1280; // @[Multiplier.scala 132:13]
  assign c53_295_io_in_1 = r_1281; // @[Multiplier.scala 132:13]
  assign c53_295_io_in_2 = r_1282; // @[Multiplier.scala 132:13]
  assign c53_295_io_in_3 = r_1283; // @[Multiplier.scala 132:13]
  assign c53_295_io_in_4 = c53_287_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_296_io_in_0 = r_1285; // @[Multiplier.scala 132:13]
  assign c53_296_io_in_1 = r_1286; // @[Multiplier.scala 132:13]
  assign c53_296_io_in_2 = r_1287; // @[Multiplier.scala 132:13]
  assign c53_296_io_in_3 = r_1288; // @[Multiplier.scala 132:13]
  assign c53_296_io_in_4 = c53_288_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_297_io_in_0 = r_1289; // @[Multiplier.scala 132:13]
  assign c53_297_io_in_1 = r_1290; // @[Multiplier.scala 132:13]
  assign c53_297_io_in_2 = r_1291; // @[Multiplier.scala 132:13]
  assign c53_297_io_in_3 = r_1292; // @[Multiplier.scala 132:13]
  assign c53_297_io_in_4 = c53_289_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_298_io_in_0 = r_1293; // @[Multiplier.scala 132:13]
  assign c53_298_io_in_1 = r_1294; // @[Multiplier.scala 132:13]
  assign c53_298_io_in_2 = r_1295; // @[Multiplier.scala 132:13]
  assign c53_298_io_in_3 = r_1296; // @[Multiplier.scala 132:13]
  assign c53_298_io_in_4 = c53_290_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_299_io_in_0 = r_1297; // @[Multiplier.scala 132:13]
  assign c53_299_io_in_1 = r_1298; // @[Multiplier.scala 132:13]
  assign c53_299_io_in_2 = r_1299; // @[Multiplier.scala 132:13]
  assign c53_299_io_in_3 = r_1300; // @[Multiplier.scala 132:13]
  assign c53_299_io_in_4 = c53_291_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_300_io_in_0 = r_1301; // @[Multiplier.scala 132:13]
  assign c53_300_io_in_1 = r_1302; // @[Multiplier.scala 132:13]
  assign c53_300_io_in_2 = r_1303; // @[Multiplier.scala 132:13]
  assign c53_300_io_in_3 = r_1304; // @[Multiplier.scala 132:13]
  assign c53_300_io_in_4 = c53_292_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_301_io_in_0 = r_1305; // @[Multiplier.scala 132:13]
  assign c53_301_io_in_1 = r_1306; // @[Multiplier.scala 132:13]
  assign c53_301_io_in_2 = r_1307; // @[Multiplier.scala 132:13]
  assign c53_301_io_in_3 = r_1308; // @[Multiplier.scala 132:13]
  assign c53_301_io_in_4 = c53_293_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_302_io_in_0 = r_1309; // @[Multiplier.scala 132:13]
  assign c53_302_io_in_1 = r_1310; // @[Multiplier.scala 132:13]
  assign c53_302_io_in_2 = r_1311; // @[Multiplier.scala 132:13]
  assign c53_302_io_in_3 = r_1312; // @[Multiplier.scala 132:13]
  assign c53_302_io_in_4 = c53_294_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_303_io_in_0 = r_1313; // @[Multiplier.scala 132:13]
  assign c53_303_io_in_1 = r_1314; // @[Multiplier.scala 132:13]
  assign c53_303_io_in_2 = r_1315; // @[Multiplier.scala 132:13]
  assign c53_303_io_in_3 = r_1316; // @[Multiplier.scala 132:13]
  assign c53_303_io_in_4 = c53_295_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_304_io_in_0 = r_1317; // @[Multiplier.scala 132:13]
  assign c53_304_io_in_1 = r_1318; // @[Multiplier.scala 132:13]
  assign c53_304_io_in_2 = r_1319; // @[Multiplier.scala 132:13]
  assign c53_304_io_in_3 = r_1320; // @[Multiplier.scala 132:13]
  assign c53_304_io_in_4 = c53_296_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_305_io_in_0 = r_1321; // @[Multiplier.scala 132:13]
  assign c53_305_io_in_1 = r_1322; // @[Multiplier.scala 132:13]
  assign c53_305_io_in_2 = r_1323; // @[Multiplier.scala 132:13]
  assign c53_305_io_in_3 = r_1324; // @[Multiplier.scala 132:13]
  assign c53_305_io_in_4 = c53_297_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_306_io_in_0 = r_1325; // @[Multiplier.scala 132:13]
  assign c53_306_io_in_1 = r_1326; // @[Multiplier.scala 132:13]
  assign c53_306_io_in_2 = r_1327; // @[Multiplier.scala 132:13]
  assign c53_306_io_in_3 = r_1328; // @[Multiplier.scala 132:13]
  assign c53_306_io_in_4 = c53_298_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_307_io_in_0 = r_1329; // @[Multiplier.scala 132:13]
  assign c53_307_io_in_1 = r_1330; // @[Multiplier.scala 132:13]
  assign c53_307_io_in_2 = r_1331; // @[Multiplier.scala 132:13]
  assign c53_307_io_in_3 = r_1332; // @[Multiplier.scala 132:13]
  assign c53_307_io_in_4 = c53_299_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_308_io_in_0 = r_1333; // @[Multiplier.scala 132:13]
  assign c53_308_io_in_1 = r_1334; // @[Multiplier.scala 132:13]
  assign c53_308_io_in_2 = r_1335; // @[Multiplier.scala 132:13]
  assign c53_308_io_in_3 = r_1336; // @[Multiplier.scala 132:13]
  assign c53_308_io_in_4 = c53_300_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_309_io_in_0 = r_1337; // @[Multiplier.scala 132:13]
  assign c53_309_io_in_1 = r_1338; // @[Multiplier.scala 132:13]
  assign c53_309_io_in_2 = r_1339; // @[Multiplier.scala 132:13]
  assign c53_309_io_in_3 = r_1340; // @[Multiplier.scala 132:13]
  assign c53_309_io_in_4 = c53_301_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_310_io_in_0 = r_1341; // @[Multiplier.scala 132:13]
  assign c53_310_io_in_1 = r_1342; // @[Multiplier.scala 132:13]
  assign c53_310_io_in_2 = r_1343; // @[Multiplier.scala 132:13]
  assign c53_310_io_in_3 = r_1344; // @[Multiplier.scala 132:13]
  assign c53_310_io_in_4 = c53_302_io_out_1; // @[Multiplier.scala 136:41]
  assign c32_16_io_in_0 = r_1345; // @[Multiplier.scala 126:19]
  assign c32_16_io_in_1 = r_1346; // @[Multiplier.scala 126:19]
  assign c32_16_io_in_2 = r_1347; // @[Multiplier.scala 126:19]
  assign c53_311_io_in_0 = r_1348; // @[Multiplier.scala 132:13]
  assign c53_311_io_in_1 = r_1349; // @[Multiplier.scala 132:13]
  assign c53_311_io_in_2 = r_1350; // @[Multiplier.scala 132:13]
  assign c53_311_io_in_3 = r_1351; // @[Multiplier.scala 132:13]
  assign c53_311_io_in_4 = c53_304_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_312_io_in_0 = r_1352; // @[Multiplier.scala 132:13]
  assign c53_312_io_in_1 = r_1353; // @[Multiplier.scala 132:13]
  assign c53_312_io_in_2 = r_1354; // @[Multiplier.scala 132:13]
  assign c53_312_io_in_3 = r_1355; // @[Multiplier.scala 132:13]
  assign c53_312_io_in_4 = c53_305_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_313_io_in_0 = r_1356; // @[Multiplier.scala 132:13]
  assign c53_313_io_in_1 = r_1357; // @[Multiplier.scala 132:13]
  assign c53_313_io_in_2 = r_1358; // @[Multiplier.scala 132:13]
  assign c53_313_io_in_3 = r_1359; // @[Multiplier.scala 132:13]
  assign c53_313_io_in_4 = c53_306_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_314_io_in_0 = r_1360; // @[Multiplier.scala 132:13]
  assign c53_314_io_in_1 = r_1361; // @[Multiplier.scala 132:13]
  assign c53_314_io_in_2 = r_1362; // @[Multiplier.scala 132:13]
  assign c53_314_io_in_3 = r_1363; // @[Multiplier.scala 132:13]
  assign c53_314_io_in_4 = c53_307_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_315_io_in_0 = r_1364; // @[Multiplier.scala 132:13]
  assign c53_315_io_in_1 = r_1365; // @[Multiplier.scala 132:13]
  assign c53_315_io_in_2 = r_1366; // @[Multiplier.scala 132:13]
  assign c53_315_io_in_3 = r_1367; // @[Multiplier.scala 132:13]
  assign c53_315_io_in_4 = c53_308_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_316_io_in_0 = r_1368; // @[Multiplier.scala 132:13]
  assign c53_316_io_in_1 = r_1369; // @[Multiplier.scala 132:13]
  assign c53_316_io_in_2 = r_1370; // @[Multiplier.scala 132:13]
  assign c53_316_io_in_3 = r_1371; // @[Multiplier.scala 132:13]
  assign c53_316_io_in_4 = c53_309_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_317_io_in_0 = r_1372; // @[Multiplier.scala 132:13]
  assign c53_317_io_in_1 = r_1373; // @[Multiplier.scala 132:13]
  assign c53_317_io_in_2 = r_1374; // @[Multiplier.scala 132:13]
  assign c53_317_io_in_3 = r_1375; // @[Multiplier.scala 132:13]
  assign c53_317_io_in_4 = c53_310_io_out_1; // @[Multiplier.scala 136:41]
  assign c32_17_io_in_0 = r_1376; // @[Multiplier.scala 126:19]
  assign c32_17_io_in_1 = r_1377; // @[Multiplier.scala 126:19]
  assign c32_17_io_in_2 = r_1378; // @[Multiplier.scala 126:19]
  assign c53_318_io_in_0 = r_1379; // @[Multiplier.scala 132:13]
  assign c53_318_io_in_1 = r_1380; // @[Multiplier.scala 132:13]
  assign c53_318_io_in_2 = r_1381; // @[Multiplier.scala 132:13]
  assign c53_318_io_in_3 = r_1382; // @[Multiplier.scala 132:13]
  assign c53_318_io_in_4 = c53_311_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_319_io_in_0 = r_1383; // @[Multiplier.scala 132:13]
  assign c53_319_io_in_1 = r_1384; // @[Multiplier.scala 132:13]
  assign c53_319_io_in_2 = r_1385; // @[Multiplier.scala 132:13]
  assign c53_319_io_in_3 = r_1386; // @[Multiplier.scala 132:13]
  assign c53_319_io_in_4 = c53_312_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_320_io_in_0 = r_1387; // @[Multiplier.scala 132:13]
  assign c53_320_io_in_1 = r_1388; // @[Multiplier.scala 132:13]
  assign c53_320_io_in_2 = r_1389; // @[Multiplier.scala 132:13]
  assign c53_320_io_in_3 = r_1390; // @[Multiplier.scala 132:13]
  assign c53_320_io_in_4 = c53_313_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_321_io_in_0 = r_1391; // @[Multiplier.scala 132:13]
  assign c53_321_io_in_1 = r_1392; // @[Multiplier.scala 132:13]
  assign c53_321_io_in_2 = r_1393; // @[Multiplier.scala 132:13]
  assign c53_321_io_in_3 = r_1394; // @[Multiplier.scala 132:13]
  assign c53_321_io_in_4 = c53_314_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_322_io_in_0 = r_1395; // @[Multiplier.scala 132:13]
  assign c53_322_io_in_1 = r_1396; // @[Multiplier.scala 132:13]
  assign c53_322_io_in_2 = r_1397; // @[Multiplier.scala 132:13]
  assign c53_322_io_in_3 = r_1398; // @[Multiplier.scala 132:13]
  assign c53_322_io_in_4 = c53_315_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_323_io_in_0 = r_1399; // @[Multiplier.scala 132:13]
  assign c53_323_io_in_1 = r_1400; // @[Multiplier.scala 132:13]
  assign c53_323_io_in_2 = r_1401; // @[Multiplier.scala 132:13]
  assign c53_323_io_in_3 = r_1402; // @[Multiplier.scala 132:13]
  assign c53_323_io_in_4 = c53_316_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_324_io_in_0 = r_1403; // @[Multiplier.scala 132:13]
  assign c53_324_io_in_1 = r_1404; // @[Multiplier.scala 132:13]
  assign c53_324_io_in_2 = r_1405; // @[Multiplier.scala 132:13]
  assign c53_324_io_in_3 = r_1406; // @[Multiplier.scala 132:13]
  assign c53_324_io_in_4 = c53_317_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_16_io_in_0 = r_1407; // @[Multiplier.scala 121:19]
  assign c22_16_io_in_1 = r_1408; // @[Multiplier.scala 121:19]
  assign c53_325_io_in_0 = r_1409; // @[Multiplier.scala 132:13]
  assign c53_325_io_in_1 = r_1410; // @[Multiplier.scala 132:13]
  assign c53_325_io_in_2 = r_1411; // @[Multiplier.scala 132:13]
  assign c53_325_io_in_3 = r_1412; // @[Multiplier.scala 132:13]
  assign c53_325_io_in_4 = c53_318_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_326_io_in_0 = r_1413; // @[Multiplier.scala 132:13]
  assign c53_326_io_in_1 = r_1414; // @[Multiplier.scala 132:13]
  assign c53_326_io_in_2 = r_1415; // @[Multiplier.scala 132:13]
  assign c53_326_io_in_3 = r_1416; // @[Multiplier.scala 132:13]
  assign c53_326_io_in_4 = c53_319_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_327_io_in_0 = r_1417; // @[Multiplier.scala 132:13]
  assign c53_327_io_in_1 = r_1418; // @[Multiplier.scala 132:13]
  assign c53_327_io_in_2 = r_1419; // @[Multiplier.scala 132:13]
  assign c53_327_io_in_3 = r_1420; // @[Multiplier.scala 132:13]
  assign c53_327_io_in_4 = c53_320_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_328_io_in_0 = r_1421; // @[Multiplier.scala 132:13]
  assign c53_328_io_in_1 = r_1422; // @[Multiplier.scala 132:13]
  assign c53_328_io_in_2 = r_1423; // @[Multiplier.scala 132:13]
  assign c53_328_io_in_3 = r_1424; // @[Multiplier.scala 132:13]
  assign c53_328_io_in_4 = c53_321_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_329_io_in_0 = r_1425; // @[Multiplier.scala 132:13]
  assign c53_329_io_in_1 = r_1426; // @[Multiplier.scala 132:13]
  assign c53_329_io_in_2 = r_1427; // @[Multiplier.scala 132:13]
  assign c53_329_io_in_3 = r_1428; // @[Multiplier.scala 132:13]
  assign c53_329_io_in_4 = c53_322_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_330_io_in_0 = r_1429; // @[Multiplier.scala 132:13]
  assign c53_330_io_in_1 = r_1430; // @[Multiplier.scala 132:13]
  assign c53_330_io_in_2 = r_1431; // @[Multiplier.scala 132:13]
  assign c53_330_io_in_3 = r_1432; // @[Multiplier.scala 132:13]
  assign c53_330_io_in_4 = c53_323_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_331_io_in_0 = r_1433; // @[Multiplier.scala 132:13]
  assign c53_331_io_in_1 = r_1434; // @[Multiplier.scala 132:13]
  assign c53_331_io_in_2 = r_1435; // @[Multiplier.scala 132:13]
  assign c53_331_io_in_3 = r_1436; // @[Multiplier.scala 132:13]
  assign c53_331_io_in_4 = c53_324_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_17_io_in_0 = r_1437; // @[Multiplier.scala 121:19]
  assign c22_17_io_in_1 = r_1438; // @[Multiplier.scala 121:19]
  assign c53_332_io_in_0 = r_1439; // @[Multiplier.scala 132:13]
  assign c53_332_io_in_1 = r_1440; // @[Multiplier.scala 132:13]
  assign c53_332_io_in_2 = r_1441; // @[Multiplier.scala 132:13]
  assign c53_332_io_in_3 = r_1442; // @[Multiplier.scala 132:13]
  assign c53_332_io_in_4 = c53_325_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_333_io_in_0 = r_1443; // @[Multiplier.scala 132:13]
  assign c53_333_io_in_1 = r_1444; // @[Multiplier.scala 132:13]
  assign c53_333_io_in_2 = r_1445; // @[Multiplier.scala 132:13]
  assign c53_333_io_in_3 = r_1446; // @[Multiplier.scala 132:13]
  assign c53_333_io_in_4 = c53_326_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_334_io_in_0 = r_1447; // @[Multiplier.scala 132:13]
  assign c53_334_io_in_1 = r_1448; // @[Multiplier.scala 132:13]
  assign c53_334_io_in_2 = r_1449; // @[Multiplier.scala 132:13]
  assign c53_334_io_in_3 = r_1450; // @[Multiplier.scala 132:13]
  assign c53_334_io_in_4 = c53_327_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_335_io_in_0 = r_1451; // @[Multiplier.scala 132:13]
  assign c53_335_io_in_1 = r_1452; // @[Multiplier.scala 132:13]
  assign c53_335_io_in_2 = r_1453; // @[Multiplier.scala 132:13]
  assign c53_335_io_in_3 = r_1454; // @[Multiplier.scala 132:13]
  assign c53_335_io_in_4 = c53_328_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_336_io_in_0 = r_1455; // @[Multiplier.scala 132:13]
  assign c53_336_io_in_1 = r_1456; // @[Multiplier.scala 132:13]
  assign c53_336_io_in_2 = r_1457; // @[Multiplier.scala 132:13]
  assign c53_336_io_in_3 = r_1458; // @[Multiplier.scala 132:13]
  assign c53_336_io_in_4 = c53_329_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_337_io_in_0 = r_1459; // @[Multiplier.scala 132:13]
  assign c53_337_io_in_1 = r_1460; // @[Multiplier.scala 132:13]
  assign c53_337_io_in_2 = r_1461; // @[Multiplier.scala 132:13]
  assign c53_337_io_in_3 = r_1462; // @[Multiplier.scala 132:13]
  assign c53_337_io_in_4 = c53_330_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_338_io_in_0 = r_1463; // @[Multiplier.scala 132:13]
  assign c53_338_io_in_1 = r_1464; // @[Multiplier.scala 132:13]
  assign c53_338_io_in_2 = r_1465; // @[Multiplier.scala 132:13]
  assign c53_338_io_in_3 = r_1466; // @[Multiplier.scala 132:13]
  assign c53_338_io_in_4 = c53_331_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_339_io_in_0 = r_1468; // @[Multiplier.scala 132:13]
  assign c53_339_io_in_1 = r_1469; // @[Multiplier.scala 132:13]
  assign c53_339_io_in_2 = r_1470; // @[Multiplier.scala 132:13]
  assign c53_339_io_in_3 = r_1471; // @[Multiplier.scala 132:13]
  assign c53_339_io_in_4 = c53_332_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_340_io_in_0 = r_1472; // @[Multiplier.scala 132:13]
  assign c53_340_io_in_1 = r_1473; // @[Multiplier.scala 132:13]
  assign c53_340_io_in_2 = r_1474; // @[Multiplier.scala 132:13]
  assign c53_340_io_in_3 = r_1475; // @[Multiplier.scala 132:13]
  assign c53_340_io_in_4 = c53_333_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_341_io_in_0 = r_1476; // @[Multiplier.scala 132:13]
  assign c53_341_io_in_1 = r_1477; // @[Multiplier.scala 132:13]
  assign c53_341_io_in_2 = r_1478; // @[Multiplier.scala 132:13]
  assign c53_341_io_in_3 = r_1479; // @[Multiplier.scala 132:13]
  assign c53_341_io_in_4 = c53_334_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_342_io_in_0 = r_1480; // @[Multiplier.scala 132:13]
  assign c53_342_io_in_1 = r_1481; // @[Multiplier.scala 132:13]
  assign c53_342_io_in_2 = r_1482; // @[Multiplier.scala 132:13]
  assign c53_342_io_in_3 = r_1483; // @[Multiplier.scala 132:13]
  assign c53_342_io_in_4 = c53_335_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_343_io_in_0 = r_1484; // @[Multiplier.scala 132:13]
  assign c53_343_io_in_1 = r_1485; // @[Multiplier.scala 132:13]
  assign c53_343_io_in_2 = r_1486; // @[Multiplier.scala 132:13]
  assign c53_343_io_in_3 = r_1487; // @[Multiplier.scala 132:13]
  assign c53_343_io_in_4 = c53_336_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_344_io_in_0 = r_1488; // @[Multiplier.scala 132:13]
  assign c53_344_io_in_1 = r_1489; // @[Multiplier.scala 132:13]
  assign c53_344_io_in_2 = r_1490; // @[Multiplier.scala 132:13]
  assign c53_344_io_in_3 = r_1491; // @[Multiplier.scala 132:13]
  assign c53_344_io_in_4 = c53_337_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_345_io_in_0 = r_1492; // @[Multiplier.scala 132:13]
  assign c53_345_io_in_1 = r_1493; // @[Multiplier.scala 132:13]
  assign c53_345_io_in_2 = r_1494; // @[Multiplier.scala 132:13]
  assign c53_345_io_in_3 = r_1495; // @[Multiplier.scala 132:13]
  assign c53_345_io_in_4 = c53_338_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_346_io_in_0 = r_1497; // @[Multiplier.scala 132:13]
  assign c53_346_io_in_1 = r_1498; // @[Multiplier.scala 132:13]
  assign c53_346_io_in_2 = r_1499; // @[Multiplier.scala 132:13]
  assign c53_346_io_in_3 = r_1500; // @[Multiplier.scala 132:13]
  assign c53_346_io_in_4 = c53_339_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_347_io_in_0 = r_1501; // @[Multiplier.scala 132:13]
  assign c53_347_io_in_1 = r_1502; // @[Multiplier.scala 132:13]
  assign c53_347_io_in_2 = r_1503; // @[Multiplier.scala 132:13]
  assign c53_347_io_in_3 = r_1504; // @[Multiplier.scala 132:13]
  assign c53_347_io_in_4 = c53_340_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_348_io_in_0 = r_1505; // @[Multiplier.scala 132:13]
  assign c53_348_io_in_1 = r_1506; // @[Multiplier.scala 132:13]
  assign c53_348_io_in_2 = r_1507; // @[Multiplier.scala 132:13]
  assign c53_348_io_in_3 = r_1508; // @[Multiplier.scala 132:13]
  assign c53_348_io_in_4 = c53_341_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_349_io_in_0 = r_1509; // @[Multiplier.scala 132:13]
  assign c53_349_io_in_1 = r_1510; // @[Multiplier.scala 132:13]
  assign c53_349_io_in_2 = r_1511; // @[Multiplier.scala 132:13]
  assign c53_349_io_in_3 = r_1512; // @[Multiplier.scala 132:13]
  assign c53_349_io_in_4 = c53_342_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_350_io_in_0 = r_1513; // @[Multiplier.scala 132:13]
  assign c53_350_io_in_1 = r_1514; // @[Multiplier.scala 132:13]
  assign c53_350_io_in_2 = r_1515; // @[Multiplier.scala 132:13]
  assign c53_350_io_in_3 = r_1516; // @[Multiplier.scala 132:13]
  assign c53_350_io_in_4 = c53_343_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_351_io_in_0 = r_1517; // @[Multiplier.scala 132:13]
  assign c53_351_io_in_1 = r_1518; // @[Multiplier.scala 132:13]
  assign c53_351_io_in_2 = r_1519; // @[Multiplier.scala 132:13]
  assign c53_351_io_in_3 = r_1520; // @[Multiplier.scala 132:13]
  assign c53_351_io_in_4 = c53_344_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_352_io_in_0 = r_1521; // @[Multiplier.scala 132:13]
  assign c53_352_io_in_1 = r_1522; // @[Multiplier.scala 132:13]
  assign c53_352_io_in_2 = r_1523; // @[Multiplier.scala 132:13]
  assign c53_352_io_in_3 = r_1524; // @[Multiplier.scala 132:13]
  assign c53_352_io_in_4 = c53_345_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_353_io_in_0 = r_1525; // @[Multiplier.scala 132:13]
  assign c53_353_io_in_1 = r_1526; // @[Multiplier.scala 132:13]
  assign c53_353_io_in_2 = r_1527; // @[Multiplier.scala 132:13]
  assign c53_353_io_in_3 = r_1528; // @[Multiplier.scala 132:13]
  assign c53_353_io_in_4 = c53_346_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_354_io_in_0 = r_1529; // @[Multiplier.scala 132:13]
  assign c53_354_io_in_1 = r_1530; // @[Multiplier.scala 132:13]
  assign c53_354_io_in_2 = r_1531; // @[Multiplier.scala 132:13]
  assign c53_354_io_in_3 = r_1532; // @[Multiplier.scala 132:13]
  assign c53_354_io_in_4 = c53_347_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_355_io_in_0 = r_1533; // @[Multiplier.scala 132:13]
  assign c53_355_io_in_1 = r_1534; // @[Multiplier.scala 132:13]
  assign c53_355_io_in_2 = r_1535; // @[Multiplier.scala 132:13]
  assign c53_355_io_in_3 = r_1536; // @[Multiplier.scala 132:13]
  assign c53_355_io_in_4 = c53_348_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_356_io_in_0 = r_1537; // @[Multiplier.scala 132:13]
  assign c53_356_io_in_1 = r_1538; // @[Multiplier.scala 132:13]
  assign c53_356_io_in_2 = r_1539; // @[Multiplier.scala 132:13]
  assign c53_356_io_in_3 = r_1540; // @[Multiplier.scala 132:13]
  assign c53_356_io_in_4 = c53_349_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_357_io_in_0 = r_1541; // @[Multiplier.scala 132:13]
  assign c53_357_io_in_1 = r_1542; // @[Multiplier.scala 132:13]
  assign c53_357_io_in_2 = r_1543; // @[Multiplier.scala 132:13]
  assign c53_357_io_in_3 = r_1544; // @[Multiplier.scala 132:13]
  assign c53_357_io_in_4 = c53_350_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_358_io_in_0 = r_1545; // @[Multiplier.scala 132:13]
  assign c53_358_io_in_1 = r_1546; // @[Multiplier.scala 132:13]
  assign c53_358_io_in_2 = r_1547; // @[Multiplier.scala 132:13]
  assign c53_358_io_in_3 = r_1548; // @[Multiplier.scala 132:13]
  assign c53_358_io_in_4 = c53_351_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_359_io_in_0 = r_1549; // @[Multiplier.scala 132:13]
  assign c53_359_io_in_1 = r_1550; // @[Multiplier.scala 132:13]
  assign c53_359_io_in_2 = r_1551; // @[Multiplier.scala 132:13]
  assign c53_359_io_in_3 = r_1552; // @[Multiplier.scala 132:13]
  assign c53_359_io_in_4 = c53_352_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_360_io_in_0 = r_1553; // @[Multiplier.scala 132:13]
  assign c53_360_io_in_1 = r_1554; // @[Multiplier.scala 132:13]
  assign c53_360_io_in_2 = r_1555; // @[Multiplier.scala 132:13]
  assign c53_360_io_in_3 = r_1556; // @[Multiplier.scala 132:13]
  assign c53_360_io_in_4 = c53_353_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_361_io_in_0 = r_1557; // @[Multiplier.scala 132:13]
  assign c53_361_io_in_1 = r_1558; // @[Multiplier.scala 132:13]
  assign c53_361_io_in_2 = r_1559; // @[Multiplier.scala 132:13]
  assign c53_361_io_in_3 = r_1560; // @[Multiplier.scala 132:13]
  assign c53_361_io_in_4 = c53_354_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_362_io_in_0 = r_1561; // @[Multiplier.scala 132:13]
  assign c53_362_io_in_1 = r_1562; // @[Multiplier.scala 132:13]
  assign c53_362_io_in_2 = r_1563; // @[Multiplier.scala 132:13]
  assign c53_362_io_in_3 = r_1564; // @[Multiplier.scala 132:13]
  assign c53_362_io_in_4 = c53_355_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_363_io_in_0 = r_1565; // @[Multiplier.scala 132:13]
  assign c53_363_io_in_1 = r_1566; // @[Multiplier.scala 132:13]
  assign c53_363_io_in_2 = r_1567; // @[Multiplier.scala 132:13]
  assign c53_363_io_in_3 = r_1568; // @[Multiplier.scala 132:13]
  assign c53_363_io_in_4 = c53_356_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_364_io_in_0 = r_1569; // @[Multiplier.scala 132:13]
  assign c53_364_io_in_1 = r_1570; // @[Multiplier.scala 132:13]
  assign c53_364_io_in_2 = r_1571; // @[Multiplier.scala 132:13]
  assign c53_364_io_in_3 = r_1572; // @[Multiplier.scala 132:13]
  assign c53_364_io_in_4 = c53_357_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_365_io_in_0 = r_1573; // @[Multiplier.scala 132:13]
  assign c53_365_io_in_1 = r_1574; // @[Multiplier.scala 132:13]
  assign c53_365_io_in_2 = r_1575; // @[Multiplier.scala 132:13]
  assign c53_365_io_in_3 = r_1576; // @[Multiplier.scala 132:13]
  assign c53_365_io_in_4 = c53_358_io_out_1; // @[Multiplier.scala 136:41]
  assign c32_18_io_in_0 = r_1577; // @[Multiplier.scala 126:19]
  assign c32_18_io_in_1 = r_1578; // @[Multiplier.scala 126:19]
  assign c32_18_io_in_2 = r_1579; // @[Multiplier.scala 126:19]
  assign c53_366_io_in_0 = r_1580; // @[Multiplier.scala 132:13]
  assign c53_366_io_in_1 = r_1581; // @[Multiplier.scala 132:13]
  assign c53_366_io_in_2 = r_1582; // @[Multiplier.scala 132:13]
  assign c53_366_io_in_3 = r_1583; // @[Multiplier.scala 132:13]
  assign c53_366_io_in_4 = c53_360_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_367_io_in_0 = r_1584; // @[Multiplier.scala 132:13]
  assign c53_367_io_in_1 = r_1585; // @[Multiplier.scala 132:13]
  assign c53_367_io_in_2 = r_1586; // @[Multiplier.scala 132:13]
  assign c53_367_io_in_3 = r_1587; // @[Multiplier.scala 132:13]
  assign c53_367_io_in_4 = c53_361_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_368_io_in_0 = r_1588; // @[Multiplier.scala 132:13]
  assign c53_368_io_in_1 = r_1589; // @[Multiplier.scala 132:13]
  assign c53_368_io_in_2 = r_1590; // @[Multiplier.scala 132:13]
  assign c53_368_io_in_3 = r_1591; // @[Multiplier.scala 132:13]
  assign c53_368_io_in_4 = c53_362_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_369_io_in_0 = r_1592; // @[Multiplier.scala 132:13]
  assign c53_369_io_in_1 = r_1593; // @[Multiplier.scala 132:13]
  assign c53_369_io_in_2 = r_1594; // @[Multiplier.scala 132:13]
  assign c53_369_io_in_3 = r_1595; // @[Multiplier.scala 132:13]
  assign c53_369_io_in_4 = c53_363_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_370_io_in_0 = r_1596; // @[Multiplier.scala 132:13]
  assign c53_370_io_in_1 = r_1597; // @[Multiplier.scala 132:13]
  assign c53_370_io_in_2 = r_1598; // @[Multiplier.scala 132:13]
  assign c53_370_io_in_3 = r_1599; // @[Multiplier.scala 132:13]
  assign c53_370_io_in_4 = c53_364_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_371_io_in_0 = r_1600; // @[Multiplier.scala 132:13]
  assign c53_371_io_in_1 = r_1601; // @[Multiplier.scala 132:13]
  assign c53_371_io_in_2 = r_1602; // @[Multiplier.scala 132:13]
  assign c53_371_io_in_3 = r_1603; // @[Multiplier.scala 132:13]
  assign c53_371_io_in_4 = c53_365_io_out_1; // @[Multiplier.scala 136:41]
  assign c32_19_io_in_0 = r_1604; // @[Multiplier.scala 126:19]
  assign c32_19_io_in_1 = r_1605; // @[Multiplier.scala 126:19]
  assign c32_19_io_in_2 = r_1606; // @[Multiplier.scala 126:19]
  assign c53_372_io_in_0 = r_1607; // @[Multiplier.scala 132:13]
  assign c53_372_io_in_1 = r_1608; // @[Multiplier.scala 132:13]
  assign c53_372_io_in_2 = r_1609; // @[Multiplier.scala 132:13]
  assign c53_372_io_in_3 = r_1610; // @[Multiplier.scala 132:13]
  assign c53_372_io_in_4 = c53_366_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_373_io_in_0 = r_1611; // @[Multiplier.scala 132:13]
  assign c53_373_io_in_1 = r_1612; // @[Multiplier.scala 132:13]
  assign c53_373_io_in_2 = r_1613; // @[Multiplier.scala 132:13]
  assign c53_373_io_in_3 = r_1614; // @[Multiplier.scala 132:13]
  assign c53_373_io_in_4 = c53_367_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_374_io_in_0 = r_1615; // @[Multiplier.scala 132:13]
  assign c53_374_io_in_1 = r_1616; // @[Multiplier.scala 132:13]
  assign c53_374_io_in_2 = r_1617; // @[Multiplier.scala 132:13]
  assign c53_374_io_in_3 = r_1618; // @[Multiplier.scala 132:13]
  assign c53_374_io_in_4 = c53_368_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_375_io_in_0 = r_1619; // @[Multiplier.scala 132:13]
  assign c53_375_io_in_1 = r_1620; // @[Multiplier.scala 132:13]
  assign c53_375_io_in_2 = r_1621; // @[Multiplier.scala 132:13]
  assign c53_375_io_in_3 = r_1622; // @[Multiplier.scala 132:13]
  assign c53_375_io_in_4 = c53_369_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_376_io_in_0 = r_1623; // @[Multiplier.scala 132:13]
  assign c53_376_io_in_1 = r_1624; // @[Multiplier.scala 132:13]
  assign c53_376_io_in_2 = r_1625; // @[Multiplier.scala 132:13]
  assign c53_376_io_in_3 = r_1626; // @[Multiplier.scala 132:13]
  assign c53_376_io_in_4 = c53_370_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_377_io_in_0 = r_1627; // @[Multiplier.scala 132:13]
  assign c53_377_io_in_1 = r_1628; // @[Multiplier.scala 132:13]
  assign c53_377_io_in_2 = r_1629; // @[Multiplier.scala 132:13]
  assign c53_377_io_in_3 = r_1630; // @[Multiplier.scala 132:13]
  assign c53_377_io_in_4 = c53_371_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_18_io_in_0 = r_1631; // @[Multiplier.scala 121:19]
  assign c22_18_io_in_1 = r_1632; // @[Multiplier.scala 121:19]
  assign c53_378_io_in_0 = r_1633; // @[Multiplier.scala 132:13]
  assign c53_378_io_in_1 = r_1634; // @[Multiplier.scala 132:13]
  assign c53_378_io_in_2 = r_1635; // @[Multiplier.scala 132:13]
  assign c53_378_io_in_3 = r_1636; // @[Multiplier.scala 132:13]
  assign c53_378_io_in_4 = c53_372_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_379_io_in_0 = r_1637; // @[Multiplier.scala 132:13]
  assign c53_379_io_in_1 = r_1638; // @[Multiplier.scala 132:13]
  assign c53_379_io_in_2 = r_1639; // @[Multiplier.scala 132:13]
  assign c53_379_io_in_3 = r_1640; // @[Multiplier.scala 132:13]
  assign c53_379_io_in_4 = c53_373_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_380_io_in_0 = r_1641; // @[Multiplier.scala 132:13]
  assign c53_380_io_in_1 = r_1642; // @[Multiplier.scala 132:13]
  assign c53_380_io_in_2 = r_1643; // @[Multiplier.scala 132:13]
  assign c53_380_io_in_3 = r_1644; // @[Multiplier.scala 132:13]
  assign c53_380_io_in_4 = c53_374_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_381_io_in_0 = r_1645; // @[Multiplier.scala 132:13]
  assign c53_381_io_in_1 = r_1646; // @[Multiplier.scala 132:13]
  assign c53_381_io_in_2 = r_1647; // @[Multiplier.scala 132:13]
  assign c53_381_io_in_3 = r_1648; // @[Multiplier.scala 132:13]
  assign c53_381_io_in_4 = c53_375_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_382_io_in_0 = r_1649; // @[Multiplier.scala 132:13]
  assign c53_382_io_in_1 = r_1650; // @[Multiplier.scala 132:13]
  assign c53_382_io_in_2 = r_1651; // @[Multiplier.scala 132:13]
  assign c53_382_io_in_3 = r_1652; // @[Multiplier.scala 132:13]
  assign c53_382_io_in_4 = c53_376_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_383_io_in_0 = r_1653; // @[Multiplier.scala 132:13]
  assign c53_383_io_in_1 = r_1654; // @[Multiplier.scala 132:13]
  assign c53_383_io_in_2 = r_1655; // @[Multiplier.scala 132:13]
  assign c53_383_io_in_3 = r_1656; // @[Multiplier.scala 132:13]
  assign c53_383_io_in_4 = c53_377_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_19_io_in_0 = r_1657; // @[Multiplier.scala 121:19]
  assign c22_19_io_in_1 = r_1658; // @[Multiplier.scala 121:19]
  assign c53_384_io_in_0 = r_1659; // @[Multiplier.scala 132:13]
  assign c53_384_io_in_1 = r_1660; // @[Multiplier.scala 132:13]
  assign c53_384_io_in_2 = r_1661; // @[Multiplier.scala 132:13]
  assign c53_384_io_in_3 = r_1662; // @[Multiplier.scala 132:13]
  assign c53_384_io_in_4 = c53_378_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_385_io_in_0 = r_1663; // @[Multiplier.scala 132:13]
  assign c53_385_io_in_1 = r_1664; // @[Multiplier.scala 132:13]
  assign c53_385_io_in_2 = r_1665; // @[Multiplier.scala 132:13]
  assign c53_385_io_in_3 = r_1666; // @[Multiplier.scala 132:13]
  assign c53_385_io_in_4 = c53_379_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_386_io_in_0 = r_1667; // @[Multiplier.scala 132:13]
  assign c53_386_io_in_1 = r_1668; // @[Multiplier.scala 132:13]
  assign c53_386_io_in_2 = r_1669; // @[Multiplier.scala 132:13]
  assign c53_386_io_in_3 = r_1670; // @[Multiplier.scala 132:13]
  assign c53_386_io_in_4 = c53_380_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_387_io_in_0 = r_1671; // @[Multiplier.scala 132:13]
  assign c53_387_io_in_1 = r_1672; // @[Multiplier.scala 132:13]
  assign c53_387_io_in_2 = r_1673; // @[Multiplier.scala 132:13]
  assign c53_387_io_in_3 = r_1674; // @[Multiplier.scala 132:13]
  assign c53_387_io_in_4 = c53_381_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_388_io_in_0 = r_1675; // @[Multiplier.scala 132:13]
  assign c53_388_io_in_1 = r_1676; // @[Multiplier.scala 132:13]
  assign c53_388_io_in_2 = r_1677; // @[Multiplier.scala 132:13]
  assign c53_388_io_in_3 = r_1678; // @[Multiplier.scala 132:13]
  assign c53_388_io_in_4 = c53_382_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_389_io_in_0 = r_1679; // @[Multiplier.scala 132:13]
  assign c53_389_io_in_1 = r_1680; // @[Multiplier.scala 132:13]
  assign c53_389_io_in_2 = r_1681; // @[Multiplier.scala 132:13]
  assign c53_389_io_in_3 = r_1682; // @[Multiplier.scala 132:13]
  assign c53_389_io_in_4 = c53_383_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_390_io_in_0 = r_1684; // @[Multiplier.scala 132:13]
  assign c53_390_io_in_1 = r_1685; // @[Multiplier.scala 132:13]
  assign c53_390_io_in_2 = r_1686; // @[Multiplier.scala 132:13]
  assign c53_390_io_in_3 = r_1687; // @[Multiplier.scala 132:13]
  assign c53_390_io_in_4 = c53_384_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_391_io_in_0 = r_1688; // @[Multiplier.scala 132:13]
  assign c53_391_io_in_1 = r_1689; // @[Multiplier.scala 132:13]
  assign c53_391_io_in_2 = r_1690; // @[Multiplier.scala 132:13]
  assign c53_391_io_in_3 = r_1691; // @[Multiplier.scala 132:13]
  assign c53_391_io_in_4 = c53_385_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_392_io_in_0 = r_1692; // @[Multiplier.scala 132:13]
  assign c53_392_io_in_1 = r_1693; // @[Multiplier.scala 132:13]
  assign c53_392_io_in_2 = r_1694; // @[Multiplier.scala 132:13]
  assign c53_392_io_in_3 = r_1695; // @[Multiplier.scala 132:13]
  assign c53_392_io_in_4 = c53_386_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_393_io_in_0 = r_1696; // @[Multiplier.scala 132:13]
  assign c53_393_io_in_1 = r_1697; // @[Multiplier.scala 132:13]
  assign c53_393_io_in_2 = r_1698; // @[Multiplier.scala 132:13]
  assign c53_393_io_in_3 = r_1699; // @[Multiplier.scala 132:13]
  assign c53_393_io_in_4 = c53_387_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_394_io_in_0 = r_1700; // @[Multiplier.scala 132:13]
  assign c53_394_io_in_1 = r_1701; // @[Multiplier.scala 132:13]
  assign c53_394_io_in_2 = r_1702; // @[Multiplier.scala 132:13]
  assign c53_394_io_in_3 = r_1703; // @[Multiplier.scala 132:13]
  assign c53_394_io_in_4 = c53_388_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_395_io_in_0 = r_1704; // @[Multiplier.scala 132:13]
  assign c53_395_io_in_1 = r_1705; // @[Multiplier.scala 132:13]
  assign c53_395_io_in_2 = r_1706; // @[Multiplier.scala 132:13]
  assign c53_395_io_in_3 = r_1707; // @[Multiplier.scala 132:13]
  assign c53_395_io_in_4 = c53_389_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_396_io_in_0 = r_1709; // @[Multiplier.scala 132:13]
  assign c53_396_io_in_1 = r_1710; // @[Multiplier.scala 132:13]
  assign c53_396_io_in_2 = r_1711; // @[Multiplier.scala 132:13]
  assign c53_396_io_in_3 = r_1712; // @[Multiplier.scala 132:13]
  assign c53_396_io_in_4 = c53_390_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_397_io_in_0 = r_1713; // @[Multiplier.scala 132:13]
  assign c53_397_io_in_1 = r_1714; // @[Multiplier.scala 132:13]
  assign c53_397_io_in_2 = r_1715; // @[Multiplier.scala 132:13]
  assign c53_397_io_in_3 = r_1716; // @[Multiplier.scala 132:13]
  assign c53_397_io_in_4 = c53_391_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_398_io_in_0 = r_1717; // @[Multiplier.scala 132:13]
  assign c53_398_io_in_1 = r_1718; // @[Multiplier.scala 132:13]
  assign c53_398_io_in_2 = r_1719; // @[Multiplier.scala 132:13]
  assign c53_398_io_in_3 = r_1720; // @[Multiplier.scala 132:13]
  assign c53_398_io_in_4 = c53_392_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_399_io_in_0 = r_1721; // @[Multiplier.scala 132:13]
  assign c53_399_io_in_1 = r_1722; // @[Multiplier.scala 132:13]
  assign c53_399_io_in_2 = r_1723; // @[Multiplier.scala 132:13]
  assign c53_399_io_in_3 = r_1724; // @[Multiplier.scala 132:13]
  assign c53_399_io_in_4 = c53_393_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_400_io_in_0 = r_1725; // @[Multiplier.scala 132:13]
  assign c53_400_io_in_1 = r_1726; // @[Multiplier.scala 132:13]
  assign c53_400_io_in_2 = r_1727; // @[Multiplier.scala 132:13]
  assign c53_400_io_in_3 = r_1728; // @[Multiplier.scala 132:13]
  assign c53_400_io_in_4 = c53_394_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_401_io_in_0 = r_1729; // @[Multiplier.scala 132:13]
  assign c53_401_io_in_1 = r_1730; // @[Multiplier.scala 132:13]
  assign c53_401_io_in_2 = r_1731; // @[Multiplier.scala 132:13]
  assign c53_401_io_in_3 = r_1732; // @[Multiplier.scala 132:13]
  assign c53_401_io_in_4 = c53_395_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_402_io_in_0 = r_1733; // @[Multiplier.scala 132:13]
  assign c53_402_io_in_1 = r_1734; // @[Multiplier.scala 132:13]
  assign c53_402_io_in_2 = r_1735; // @[Multiplier.scala 132:13]
  assign c53_402_io_in_3 = r_1736; // @[Multiplier.scala 132:13]
  assign c53_402_io_in_4 = c53_396_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_403_io_in_0 = r_1737; // @[Multiplier.scala 132:13]
  assign c53_403_io_in_1 = r_1738; // @[Multiplier.scala 132:13]
  assign c53_403_io_in_2 = r_1739; // @[Multiplier.scala 132:13]
  assign c53_403_io_in_3 = r_1740; // @[Multiplier.scala 132:13]
  assign c53_403_io_in_4 = c53_397_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_404_io_in_0 = r_1741; // @[Multiplier.scala 132:13]
  assign c53_404_io_in_1 = r_1742; // @[Multiplier.scala 132:13]
  assign c53_404_io_in_2 = r_1743; // @[Multiplier.scala 132:13]
  assign c53_404_io_in_3 = r_1744; // @[Multiplier.scala 132:13]
  assign c53_404_io_in_4 = c53_398_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_405_io_in_0 = r_1745; // @[Multiplier.scala 132:13]
  assign c53_405_io_in_1 = r_1746; // @[Multiplier.scala 132:13]
  assign c53_405_io_in_2 = r_1747; // @[Multiplier.scala 132:13]
  assign c53_405_io_in_3 = r_1748; // @[Multiplier.scala 132:13]
  assign c53_405_io_in_4 = c53_399_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_406_io_in_0 = r_1749; // @[Multiplier.scala 132:13]
  assign c53_406_io_in_1 = r_1750; // @[Multiplier.scala 132:13]
  assign c53_406_io_in_2 = r_1751; // @[Multiplier.scala 132:13]
  assign c53_406_io_in_3 = r_1752; // @[Multiplier.scala 132:13]
  assign c53_406_io_in_4 = c53_400_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_407_io_in_0 = r_1753; // @[Multiplier.scala 132:13]
  assign c53_407_io_in_1 = r_1754; // @[Multiplier.scala 132:13]
  assign c53_407_io_in_2 = r_1755; // @[Multiplier.scala 132:13]
  assign c53_407_io_in_3 = r_1756; // @[Multiplier.scala 132:13]
  assign c53_407_io_in_4 = c53_401_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_408_io_in_0 = r_1757; // @[Multiplier.scala 132:13]
  assign c53_408_io_in_1 = r_1758; // @[Multiplier.scala 132:13]
  assign c53_408_io_in_2 = r_1759; // @[Multiplier.scala 132:13]
  assign c53_408_io_in_3 = r_1760; // @[Multiplier.scala 132:13]
  assign c53_408_io_in_4 = c53_402_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_409_io_in_0 = r_1761; // @[Multiplier.scala 132:13]
  assign c53_409_io_in_1 = r_1762; // @[Multiplier.scala 132:13]
  assign c53_409_io_in_2 = r_1763; // @[Multiplier.scala 132:13]
  assign c53_409_io_in_3 = r_1764; // @[Multiplier.scala 132:13]
  assign c53_409_io_in_4 = c53_403_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_410_io_in_0 = r_1765; // @[Multiplier.scala 132:13]
  assign c53_410_io_in_1 = r_1766; // @[Multiplier.scala 132:13]
  assign c53_410_io_in_2 = r_1767; // @[Multiplier.scala 132:13]
  assign c53_410_io_in_3 = r_1768; // @[Multiplier.scala 132:13]
  assign c53_410_io_in_4 = c53_404_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_411_io_in_0 = r_1769; // @[Multiplier.scala 132:13]
  assign c53_411_io_in_1 = r_1770; // @[Multiplier.scala 132:13]
  assign c53_411_io_in_2 = r_1771; // @[Multiplier.scala 132:13]
  assign c53_411_io_in_3 = r_1772; // @[Multiplier.scala 132:13]
  assign c53_411_io_in_4 = c53_405_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_412_io_in_0 = r_1773; // @[Multiplier.scala 132:13]
  assign c53_412_io_in_1 = r_1774; // @[Multiplier.scala 132:13]
  assign c53_412_io_in_2 = r_1775; // @[Multiplier.scala 132:13]
  assign c53_412_io_in_3 = r_1776; // @[Multiplier.scala 132:13]
  assign c53_412_io_in_4 = c53_406_io_out_1; // @[Multiplier.scala 136:41]
  assign c32_20_io_in_0 = r_1777; // @[Multiplier.scala 126:19]
  assign c32_20_io_in_1 = r_1778; // @[Multiplier.scala 126:19]
  assign c32_20_io_in_2 = r_1779; // @[Multiplier.scala 126:19]
  assign c53_413_io_in_0 = r_1780; // @[Multiplier.scala 132:13]
  assign c53_413_io_in_1 = r_1781; // @[Multiplier.scala 132:13]
  assign c53_413_io_in_2 = r_1782; // @[Multiplier.scala 132:13]
  assign c53_413_io_in_3 = r_1783; // @[Multiplier.scala 132:13]
  assign c53_413_io_in_4 = c53_408_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_414_io_in_0 = r_1784; // @[Multiplier.scala 132:13]
  assign c53_414_io_in_1 = r_1785; // @[Multiplier.scala 132:13]
  assign c53_414_io_in_2 = r_1786; // @[Multiplier.scala 132:13]
  assign c53_414_io_in_3 = r_1787; // @[Multiplier.scala 132:13]
  assign c53_414_io_in_4 = c53_409_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_415_io_in_0 = r_1788; // @[Multiplier.scala 132:13]
  assign c53_415_io_in_1 = r_1789; // @[Multiplier.scala 132:13]
  assign c53_415_io_in_2 = r_1790; // @[Multiplier.scala 132:13]
  assign c53_415_io_in_3 = r_1791; // @[Multiplier.scala 132:13]
  assign c53_415_io_in_4 = c53_410_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_416_io_in_0 = r_1792; // @[Multiplier.scala 132:13]
  assign c53_416_io_in_1 = r_1793; // @[Multiplier.scala 132:13]
  assign c53_416_io_in_2 = r_1794; // @[Multiplier.scala 132:13]
  assign c53_416_io_in_3 = r_1795; // @[Multiplier.scala 132:13]
  assign c53_416_io_in_4 = c53_411_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_417_io_in_0 = r_1796; // @[Multiplier.scala 132:13]
  assign c53_417_io_in_1 = r_1797; // @[Multiplier.scala 132:13]
  assign c53_417_io_in_2 = r_1798; // @[Multiplier.scala 132:13]
  assign c53_417_io_in_3 = r_1799; // @[Multiplier.scala 132:13]
  assign c53_417_io_in_4 = c53_412_io_out_1; // @[Multiplier.scala 136:41]
  assign c32_21_io_in_0 = r_1800; // @[Multiplier.scala 126:19]
  assign c32_21_io_in_1 = r_1801; // @[Multiplier.scala 126:19]
  assign c32_21_io_in_2 = r_1802; // @[Multiplier.scala 126:19]
  assign c53_418_io_in_0 = r_1803; // @[Multiplier.scala 132:13]
  assign c53_418_io_in_1 = r_1804; // @[Multiplier.scala 132:13]
  assign c53_418_io_in_2 = r_1805; // @[Multiplier.scala 132:13]
  assign c53_418_io_in_3 = r_1806; // @[Multiplier.scala 132:13]
  assign c53_418_io_in_4 = c53_413_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_419_io_in_0 = r_1807; // @[Multiplier.scala 132:13]
  assign c53_419_io_in_1 = r_1808; // @[Multiplier.scala 132:13]
  assign c53_419_io_in_2 = r_1809; // @[Multiplier.scala 132:13]
  assign c53_419_io_in_3 = r_1810; // @[Multiplier.scala 132:13]
  assign c53_419_io_in_4 = c53_414_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_420_io_in_0 = r_1811; // @[Multiplier.scala 132:13]
  assign c53_420_io_in_1 = r_1812; // @[Multiplier.scala 132:13]
  assign c53_420_io_in_2 = r_1813; // @[Multiplier.scala 132:13]
  assign c53_420_io_in_3 = r_1814; // @[Multiplier.scala 132:13]
  assign c53_420_io_in_4 = c53_415_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_421_io_in_0 = r_1815; // @[Multiplier.scala 132:13]
  assign c53_421_io_in_1 = r_1816; // @[Multiplier.scala 132:13]
  assign c53_421_io_in_2 = r_1817; // @[Multiplier.scala 132:13]
  assign c53_421_io_in_3 = r_1818; // @[Multiplier.scala 132:13]
  assign c53_421_io_in_4 = c53_416_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_422_io_in_0 = r_1819; // @[Multiplier.scala 132:13]
  assign c53_422_io_in_1 = r_1820; // @[Multiplier.scala 132:13]
  assign c53_422_io_in_2 = r_1821; // @[Multiplier.scala 132:13]
  assign c53_422_io_in_3 = r_1822; // @[Multiplier.scala 132:13]
  assign c53_422_io_in_4 = c53_417_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_20_io_in_0 = r_1823; // @[Multiplier.scala 121:19]
  assign c22_20_io_in_1 = r_1824; // @[Multiplier.scala 121:19]
  assign c53_423_io_in_0 = r_1825; // @[Multiplier.scala 132:13]
  assign c53_423_io_in_1 = r_1826; // @[Multiplier.scala 132:13]
  assign c53_423_io_in_2 = r_1827; // @[Multiplier.scala 132:13]
  assign c53_423_io_in_3 = r_1828; // @[Multiplier.scala 132:13]
  assign c53_423_io_in_4 = c53_418_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_424_io_in_0 = r_1829; // @[Multiplier.scala 132:13]
  assign c53_424_io_in_1 = r_1830; // @[Multiplier.scala 132:13]
  assign c53_424_io_in_2 = r_1831; // @[Multiplier.scala 132:13]
  assign c53_424_io_in_3 = r_1832; // @[Multiplier.scala 132:13]
  assign c53_424_io_in_4 = c53_419_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_425_io_in_0 = r_1833; // @[Multiplier.scala 132:13]
  assign c53_425_io_in_1 = r_1834; // @[Multiplier.scala 132:13]
  assign c53_425_io_in_2 = r_1835; // @[Multiplier.scala 132:13]
  assign c53_425_io_in_3 = r_1836; // @[Multiplier.scala 132:13]
  assign c53_425_io_in_4 = c53_420_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_426_io_in_0 = r_1837; // @[Multiplier.scala 132:13]
  assign c53_426_io_in_1 = r_1838; // @[Multiplier.scala 132:13]
  assign c53_426_io_in_2 = r_1839; // @[Multiplier.scala 132:13]
  assign c53_426_io_in_3 = r_1840; // @[Multiplier.scala 132:13]
  assign c53_426_io_in_4 = c53_421_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_427_io_in_0 = r_1841; // @[Multiplier.scala 132:13]
  assign c53_427_io_in_1 = r_1842; // @[Multiplier.scala 132:13]
  assign c53_427_io_in_2 = r_1843; // @[Multiplier.scala 132:13]
  assign c53_427_io_in_3 = r_1844; // @[Multiplier.scala 132:13]
  assign c53_427_io_in_4 = c53_422_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_21_io_in_0 = r_1845; // @[Multiplier.scala 121:19]
  assign c22_21_io_in_1 = r_1846; // @[Multiplier.scala 121:19]
  assign c53_428_io_in_0 = r_1847; // @[Multiplier.scala 132:13]
  assign c53_428_io_in_1 = r_1848; // @[Multiplier.scala 132:13]
  assign c53_428_io_in_2 = r_1849; // @[Multiplier.scala 132:13]
  assign c53_428_io_in_3 = r_1850; // @[Multiplier.scala 132:13]
  assign c53_428_io_in_4 = c53_423_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_429_io_in_0 = r_1851; // @[Multiplier.scala 132:13]
  assign c53_429_io_in_1 = r_1852; // @[Multiplier.scala 132:13]
  assign c53_429_io_in_2 = r_1853; // @[Multiplier.scala 132:13]
  assign c53_429_io_in_3 = r_1854; // @[Multiplier.scala 132:13]
  assign c53_429_io_in_4 = c53_424_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_430_io_in_0 = r_1855; // @[Multiplier.scala 132:13]
  assign c53_430_io_in_1 = r_1856; // @[Multiplier.scala 132:13]
  assign c53_430_io_in_2 = r_1857; // @[Multiplier.scala 132:13]
  assign c53_430_io_in_3 = r_1858; // @[Multiplier.scala 132:13]
  assign c53_430_io_in_4 = c53_425_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_431_io_in_0 = r_1859; // @[Multiplier.scala 132:13]
  assign c53_431_io_in_1 = r_1860; // @[Multiplier.scala 132:13]
  assign c53_431_io_in_2 = r_1861; // @[Multiplier.scala 132:13]
  assign c53_431_io_in_3 = r_1862; // @[Multiplier.scala 132:13]
  assign c53_431_io_in_4 = c53_426_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_432_io_in_0 = r_1863; // @[Multiplier.scala 132:13]
  assign c53_432_io_in_1 = r_1864; // @[Multiplier.scala 132:13]
  assign c53_432_io_in_2 = r_1865; // @[Multiplier.scala 132:13]
  assign c53_432_io_in_3 = r_1866; // @[Multiplier.scala 132:13]
  assign c53_432_io_in_4 = c53_427_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_433_io_in_0 = r_1868; // @[Multiplier.scala 132:13]
  assign c53_433_io_in_1 = r_1869; // @[Multiplier.scala 132:13]
  assign c53_433_io_in_2 = r_1870; // @[Multiplier.scala 132:13]
  assign c53_433_io_in_3 = r_1871; // @[Multiplier.scala 132:13]
  assign c53_433_io_in_4 = c53_428_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_434_io_in_0 = r_1872; // @[Multiplier.scala 132:13]
  assign c53_434_io_in_1 = r_1873; // @[Multiplier.scala 132:13]
  assign c53_434_io_in_2 = r_1874; // @[Multiplier.scala 132:13]
  assign c53_434_io_in_3 = r_1875; // @[Multiplier.scala 132:13]
  assign c53_434_io_in_4 = c53_429_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_435_io_in_0 = r_1876; // @[Multiplier.scala 132:13]
  assign c53_435_io_in_1 = r_1877; // @[Multiplier.scala 132:13]
  assign c53_435_io_in_2 = r_1878; // @[Multiplier.scala 132:13]
  assign c53_435_io_in_3 = r_1879; // @[Multiplier.scala 132:13]
  assign c53_435_io_in_4 = c53_430_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_436_io_in_0 = r_1880; // @[Multiplier.scala 132:13]
  assign c53_436_io_in_1 = r_1881; // @[Multiplier.scala 132:13]
  assign c53_436_io_in_2 = r_1882; // @[Multiplier.scala 132:13]
  assign c53_436_io_in_3 = r_1883; // @[Multiplier.scala 132:13]
  assign c53_436_io_in_4 = c53_431_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_437_io_in_0 = r_1884; // @[Multiplier.scala 132:13]
  assign c53_437_io_in_1 = r_1885; // @[Multiplier.scala 132:13]
  assign c53_437_io_in_2 = r_1886; // @[Multiplier.scala 132:13]
  assign c53_437_io_in_3 = r_1887; // @[Multiplier.scala 132:13]
  assign c53_437_io_in_4 = c53_432_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_438_io_in_0 = r_1889; // @[Multiplier.scala 132:13]
  assign c53_438_io_in_1 = r_1890; // @[Multiplier.scala 132:13]
  assign c53_438_io_in_2 = r_1891; // @[Multiplier.scala 132:13]
  assign c53_438_io_in_3 = r_1892; // @[Multiplier.scala 132:13]
  assign c53_438_io_in_4 = c53_433_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_439_io_in_0 = r_1893; // @[Multiplier.scala 132:13]
  assign c53_439_io_in_1 = r_1894; // @[Multiplier.scala 132:13]
  assign c53_439_io_in_2 = r_1895; // @[Multiplier.scala 132:13]
  assign c53_439_io_in_3 = r_1896; // @[Multiplier.scala 132:13]
  assign c53_439_io_in_4 = c53_434_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_440_io_in_0 = r_1897; // @[Multiplier.scala 132:13]
  assign c53_440_io_in_1 = r_1898; // @[Multiplier.scala 132:13]
  assign c53_440_io_in_2 = r_1899; // @[Multiplier.scala 132:13]
  assign c53_440_io_in_3 = r_1900; // @[Multiplier.scala 132:13]
  assign c53_440_io_in_4 = c53_435_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_441_io_in_0 = r_1901; // @[Multiplier.scala 132:13]
  assign c53_441_io_in_1 = r_1902; // @[Multiplier.scala 132:13]
  assign c53_441_io_in_2 = r_1903; // @[Multiplier.scala 132:13]
  assign c53_441_io_in_3 = r_1904; // @[Multiplier.scala 132:13]
  assign c53_441_io_in_4 = c53_436_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_442_io_in_0 = r_1905; // @[Multiplier.scala 132:13]
  assign c53_442_io_in_1 = r_1906; // @[Multiplier.scala 132:13]
  assign c53_442_io_in_2 = r_1907; // @[Multiplier.scala 132:13]
  assign c53_442_io_in_3 = r_1908; // @[Multiplier.scala 132:13]
  assign c53_442_io_in_4 = c53_437_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_443_io_in_0 = r_1909; // @[Multiplier.scala 132:13]
  assign c53_443_io_in_1 = r_1910; // @[Multiplier.scala 132:13]
  assign c53_443_io_in_2 = r_1911; // @[Multiplier.scala 132:13]
  assign c53_443_io_in_3 = r_1912; // @[Multiplier.scala 132:13]
  assign c53_443_io_in_4 = c53_438_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_444_io_in_0 = r_1913; // @[Multiplier.scala 132:13]
  assign c53_444_io_in_1 = r_1914; // @[Multiplier.scala 132:13]
  assign c53_444_io_in_2 = r_1915; // @[Multiplier.scala 132:13]
  assign c53_444_io_in_3 = r_1916; // @[Multiplier.scala 132:13]
  assign c53_444_io_in_4 = c53_439_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_445_io_in_0 = r_1917; // @[Multiplier.scala 132:13]
  assign c53_445_io_in_1 = r_1918; // @[Multiplier.scala 132:13]
  assign c53_445_io_in_2 = r_1919; // @[Multiplier.scala 132:13]
  assign c53_445_io_in_3 = r_1920; // @[Multiplier.scala 132:13]
  assign c53_445_io_in_4 = c53_440_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_446_io_in_0 = r_1921; // @[Multiplier.scala 132:13]
  assign c53_446_io_in_1 = r_1922; // @[Multiplier.scala 132:13]
  assign c53_446_io_in_2 = r_1923; // @[Multiplier.scala 132:13]
  assign c53_446_io_in_3 = r_1924; // @[Multiplier.scala 132:13]
  assign c53_446_io_in_4 = c53_441_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_447_io_in_0 = r_1925; // @[Multiplier.scala 132:13]
  assign c53_447_io_in_1 = r_1926; // @[Multiplier.scala 132:13]
  assign c53_447_io_in_2 = r_1927; // @[Multiplier.scala 132:13]
  assign c53_447_io_in_3 = r_1928; // @[Multiplier.scala 132:13]
  assign c53_447_io_in_4 = c53_442_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_448_io_in_0 = r_1929; // @[Multiplier.scala 132:13]
  assign c53_448_io_in_1 = r_1930; // @[Multiplier.scala 132:13]
  assign c53_448_io_in_2 = r_1931; // @[Multiplier.scala 132:13]
  assign c53_448_io_in_3 = r_1932; // @[Multiplier.scala 132:13]
  assign c53_448_io_in_4 = c53_443_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_449_io_in_0 = r_1933; // @[Multiplier.scala 132:13]
  assign c53_449_io_in_1 = r_1934; // @[Multiplier.scala 132:13]
  assign c53_449_io_in_2 = r_1935; // @[Multiplier.scala 132:13]
  assign c53_449_io_in_3 = r_1936; // @[Multiplier.scala 132:13]
  assign c53_449_io_in_4 = c53_444_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_450_io_in_0 = r_1937; // @[Multiplier.scala 132:13]
  assign c53_450_io_in_1 = r_1938; // @[Multiplier.scala 132:13]
  assign c53_450_io_in_2 = r_1939; // @[Multiplier.scala 132:13]
  assign c53_450_io_in_3 = r_1940; // @[Multiplier.scala 132:13]
  assign c53_450_io_in_4 = c53_445_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_451_io_in_0 = r_1941; // @[Multiplier.scala 132:13]
  assign c53_451_io_in_1 = r_1942; // @[Multiplier.scala 132:13]
  assign c53_451_io_in_2 = r_1943; // @[Multiplier.scala 132:13]
  assign c53_451_io_in_3 = r_1944; // @[Multiplier.scala 132:13]
  assign c53_451_io_in_4 = c53_446_io_out_1; // @[Multiplier.scala 136:41]
  assign c32_22_io_in_0 = r_1945; // @[Multiplier.scala 126:19]
  assign c32_22_io_in_1 = r_1946; // @[Multiplier.scala 126:19]
  assign c32_22_io_in_2 = r_1947; // @[Multiplier.scala 126:19]
  assign c53_452_io_in_0 = r_1948; // @[Multiplier.scala 132:13]
  assign c53_452_io_in_1 = r_1949; // @[Multiplier.scala 132:13]
  assign c53_452_io_in_2 = r_1950; // @[Multiplier.scala 132:13]
  assign c53_452_io_in_3 = r_1951; // @[Multiplier.scala 132:13]
  assign c53_452_io_in_4 = c53_448_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_453_io_in_0 = r_1952; // @[Multiplier.scala 132:13]
  assign c53_453_io_in_1 = r_1953; // @[Multiplier.scala 132:13]
  assign c53_453_io_in_2 = r_1954; // @[Multiplier.scala 132:13]
  assign c53_453_io_in_3 = r_1955; // @[Multiplier.scala 132:13]
  assign c53_453_io_in_4 = c53_449_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_454_io_in_0 = r_1956; // @[Multiplier.scala 132:13]
  assign c53_454_io_in_1 = r_1957; // @[Multiplier.scala 132:13]
  assign c53_454_io_in_2 = r_1958; // @[Multiplier.scala 132:13]
  assign c53_454_io_in_3 = r_1959; // @[Multiplier.scala 132:13]
  assign c53_454_io_in_4 = c53_450_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_455_io_in_0 = r_1960; // @[Multiplier.scala 132:13]
  assign c53_455_io_in_1 = r_1961; // @[Multiplier.scala 132:13]
  assign c53_455_io_in_2 = r_1962; // @[Multiplier.scala 132:13]
  assign c53_455_io_in_3 = r_1963; // @[Multiplier.scala 132:13]
  assign c53_455_io_in_4 = c53_451_io_out_1; // @[Multiplier.scala 136:41]
  assign c32_23_io_in_0 = r_1964; // @[Multiplier.scala 126:19]
  assign c32_23_io_in_1 = r_1965; // @[Multiplier.scala 126:19]
  assign c32_23_io_in_2 = r_1966; // @[Multiplier.scala 126:19]
  assign c53_456_io_in_0 = r_1967; // @[Multiplier.scala 132:13]
  assign c53_456_io_in_1 = r_1968; // @[Multiplier.scala 132:13]
  assign c53_456_io_in_2 = r_1969; // @[Multiplier.scala 132:13]
  assign c53_456_io_in_3 = r_1970; // @[Multiplier.scala 132:13]
  assign c53_456_io_in_4 = c53_452_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_457_io_in_0 = r_1971; // @[Multiplier.scala 132:13]
  assign c53_457_io_in_1 = r_1972; // @[Multiplier.scala 132:13]
  assign c53_457_io_in_2 = r_1973; // @[Multiplier.scala 132:13]
  assign c53_457_io_in_3 = r_1974; // @[Multiplier.scala 132:13]
  assign c53_457_io_in_4 = c53_453_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_458_io_in_0 = r_1975; // @[Multiplier.scala 132:13]
  assign c53_458_io_in_1 = r_1976; // @[Multiplier.scala 132:13]
  assign c53_458_io_in_2 = r_1977; // @[Multiplier.scala 132:13]
  assign c53_458_io_in_3 = r_1978; // @[Multiplier.scala 132:13]
  assign c53_458_io_in_4 = c53_454_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_459_io_in_0 = r_1979; // @[Multiplier.scala 132:13]
  assign c53_459_io_in_1 = r_1980; // @[Multiplier.scala 132:13]
  assign c53_459_io_in_2 = r_1981; // @[Multiplier.scala 132:13]
  assign c53_459_io_in_3 = r_1982; // @[Multiplier.scala 132:13]
  assign c53_459_io_in_4 = c53_455_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_22_io_in_0 = r_1983; // @[Multiplier.scala 121:19]
  assign c22_22_io_in_1 = r_1984; // @[Multiplier.scala 121:19]
  assign c53_460_io_in_0 = r_1985; // @[Multiplier.scala 132:13]
  assign c53_460_io_in_1 = r_1986; // @[Multiplier.scala 132:13]
  assign c53_460_io_in_2 = r_1987; // @[Multiplier.scala 132:13]
  assign c53_460_io_in_3 = r_1988; // @[Multiplier.scala 132:13]
  assign c53_460_io_in_4 = c53_456_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_461_io_in_0 = r_1989; // @[Multiplier.scala 132:13]
  assign c53_461_io_in_1 = r_1990; // @[Multiplier.scala 132:13]
  assign c53_461_io_in_2 = r_1991; // @[Multiplier.scala 132:13]
  assign c53_461_io_in_3 = r_1992; // @[Multiplier.scala 132:13]
  assign c53_461_io_in_4 = c53_457_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_462_io_in_0 = r_1993; // @[Multiplier.scala 132:13]
  assign c53_462_io_in_1 = r_1994; // @[Multiplier.scala 132:13]
  assign c53_462_io_in_2 = r_1995; // @[Multiplier.scala 132:13]
  assign c53_462_io_in_3 = r_1996; // @[Multiplier.scala 132:13]
  assign c53_462_io_in_4 = c53_458_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_463_io_in_0 = r_1997; // @[Multiplier.scala 132:13]
  assign c53_463_io_in_1 = r_1998; // @[Multiplier.scala 132:13]
  assign c53_463_io_in_2 = r_1999; // @[Multiplier.scala 132:13]
  assign c53_463_io_in_3 = r_2000; // @[Multiplier.scala 132:13]
  assign c53_463_io_in_4 = c53_459_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_23_io_in_0 = r_2001; // @[Multiplier.scala 121:19]
  assign c22_23_io_in_1 = r_2002; // @[Multiplier.scala 121:19]
  assign c53_464_io_in_0 = r_2003; // @[Multiplier.scala 132:13]
  assign c53_464_io_in_1 = r_2004; // @[Multiplier.scala 132:13]
  assign c53_464_io_in_2 = r_2005; // @[Multiplier.scala 132:13]
  assign c53_464_io_in_3 = r_2006; // @[Multiplier.scala 132:13]
  assign c53_464_io_in_4 = c53_460_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_465_io_in_0 = r_2007; // @[Multiplier.scala 132:13]
  assign c53_465_io_in_1 = r_2008; // @[Multiplier.scala 132:13]
  assign c53_465_io_in_2 = r_2009; // @[Multiplier.scala 132:13]
  assign c53_465_io_in_3 = r_2010; // @[Multiplier.scala 132:13]
  assign c53_465_io_in_4 = c53_461_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_466_io_in_0 = r_2011; // @[Multiplier.scala 132:13]
  assign c53_466_io_in_1 = r_2012; // @[Multiplier.scala 132:13]
  assign c53_466_io_in_2 = r_2013; // @[Multiplier.scala 132:13]
  assign c53_466_io_in_3 = r_2014; // @[Multiplier.scala 132:13]
  assign c53_466_io_in_4 = c53_462_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_467_io_in_0 = r_2015; // @[Multiplier.scala 132:13]
  assign c53_467_io_in_1 = r_2016; // @[Multiplier.scala 132:13]
  assign c53_467_io_in_2 = r_2017; // @[Multiplier.scala 132:13]
  assign c53_467_io_in_3 = r_2018; // @[Multiplier.scala 132:13]
  assign c53_467_io_in_4 = c53_463_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_468_io_in_0 = r_2020; // @[Multiplier.scala 132:13]
  assign c53_468_io_in_1 = r_2021; // @[Multiplier.scala 132:13]
  assign c53_468_io_in_2 = r_2022; // @[Multiplier.scala 132:13]
  assign c53_468_io_in_3 = r_2023; // @[Multiplier.scala 132:13]
  assign c53_468_io_in_4 = c53_464_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_469_io_in_0 = r_2024; // @[Multiplier.scala 132:13]
  assign c53_469_io_in_1 = r_2025; // @[Multiplier.scala 132:13]
  assign c53_469_io_in_2 = r_2026; // @[Multiplier.scala 132:13]
  assign c53_469_io_in_3 = r_2027; // @[Multiplier.scala 132:13]
  assign c53_469_io_in_4 = c53_465_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_470_io_in_0 = r_2028; // @[Multiplier.scala 132:13]
  assign c53_470_io_in_1 = r_2029; // @[Multiplier.scala 132:13]
  assign c53_470_io_in_2 = r_2030; // @[Multiplier.scala 132:13]
  assign c53_470_io_in_3 = r_2031; // @[Multiplier.scala 132:13]
  assign c53_470_io_in_4 = c53_466_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_471_io_in_0 = r_2032; // @[Multiplier.scala 132:13]
  assign c53_471_io_in_1 = r_2033; // @[Multiplier.scala 132:13]
  assign c53_471_io_in_2 = r_2034; // @[Multiplier.scala 132:13]
  assign c53_471_io_in_3 = r_2035; // @[Multiplier.scala 132:13]
  assign c53_471_io_in_4 = c53_467_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_472_io_in_0 = r_2037; // @[Multiplier.scala 132:13]
  assign c53_472_io_in_1 = r_2038; // @[Multiplier.scala 132:13]
  assign c53_472_io_in_2 = r_2039; // @[Multiplier.scala 132:13]
  assign c53_472_io_in_3 = r_2040; // @[Multiplier.scala 132:13]
  assign c53_472_io_in_4 = c53_468_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_473_io_in_0 = r_2041; // @[Multiplier.scala 132:13]
  assign c53_473_io_in_1 = r_2042; // @[Multiplier.scala 132:13]
  assign c53_473_io_in_2 = r_2043; // @[Multiplier.scala 132:13]
  assign c53_473_io_in_3 = r_2044; // @[Multiplier.scala 132:13]
  assign c53_473_io_in_4 = c53_469_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_474_io_in_0 = r_2045; // @[Multiplier.scala 132:13]
  assign c53_474_io_in_1 = r_2046; // @[Multiplier.scala 132:13]
  assign c53_474_io_in_2 = r_2047; // @[Multiplier.scala 132:13]
  assign c53_474_io_in_3 = r_2048; // @[Multiplier.scala 132:13]
  assign c53_474_io_in_4 = c53_470_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_475_io_in_0 = r_2049; // @[Multiplier.scala 132:13]
  assign c53_475_io_in_1 = r_2050; // @[Multiplier.scala 132:13]
  assign c53_475_io_in_2 = r_2051; // @[Multiplier.scala 132:13]
  assign c53_475_io_in_3 = r_2052; // @[Multiplier.scala 132:13]
  assign c53_475_io_in_4 = c53_471_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_476_io_in_0 = r_2053; // @[Multiplier.scala 132:13]
  assign c53_476_io_in_1 = r_2054; // @[Multiplier.scala 132:13]
  assign c53_476_io_in_2 = r_2055; // @[Multiplier.scala 132:13]
  assign c53_476_io_in_3 = r_2056; // @[Multiplier.scala 132:13]
  assign c53_476_io_in_4 = c53_472_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_477_io_in_0 = r_2057; // @[Multiplier.scala 132:13]
  assign c53_477_io_in_1 = r_2058; // @[Multiplier.scala 132:13]
  assign c53_477_io_in_2 = r_2059; // @[Multiplier.scala 132:13]
  assign c53_477_io_in_3 = r_2060; // @[Multiplier.scala 132:13]
  assign c53_477_io_in_4 = c53_473_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_478_io_in_0 = r_2061; // @[Multiplier.scala 132:13]
  assign c53_478_io_in_1 = r_2062; // @[Multiplier.scala 132:13]
  assign c53_478_io_in_2 = r_2063; // @[Multiplier.scala 132:13]
  assign c53_478_io_in_3 = r_2064; // @[Multiplier.scala 132:13]
  assign c53_478_io_in_4 = c53_474_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_479_io_in_0 = r_2065; // @[Multiplier.scala 132:13]
  assign c53_479_io_in_1 = r_2066; // @[Multiplier.scala 132:13]
  assign c53_479_io_in_2 = r_2067; // @[Multiplier.scala 132:13]
  assign c53_479_io_in_3 = r_2068; // @[Multiplier.scala 132:13]
  assign c53_479_io_in_4 = c53_475_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_480_io_in_0 = r_2069; // @[Multiplier.scala 132:13]
  assign c53_480_io_in_1 = r_2070; // @[Multiplier.scala 132:13]
  assign c53_480_io_in_2 = r_2071; // @[Multiplier.scala 132:13]
  assign c53_480_io_in_3 = r_2072; // @[Multiplier.scala 132:13]
  assign c53_480_io_in_4 = c53_476_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_481_io_in_0 = r_2073; // @[Multiplier.scala 132:13]
  assign c53_481_io_in_1 = r_2074; // @[Multiplier.scala 132:13]
  assign c53_481_io_in_2 = r_2075; // @[Multiplier.scala 132:13]
  assign c53_481_io_in_3 = r_2076; // @[Multiplier.scala 132:13]
  assign c53_481_io_in_4 = c53_477_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_482_io_in_0 = r_2077; // @[Multiplier.scala 132:13]
  assign c53_482_io_in_1 = r_2078; // @[Multiplier.scala 132:13]
  assign c53_482_io_in_2 = r_2079; // @[Multiplier.scala 132:13]
  assign c53_482_io_in_3 = r_2080; // @[Multiplier.scala 132:13]
  assign c53_482_io_in_4 = c53_478_io_out_1; // @[Multiplier.scala 136:41]
  assign c32_24_io_in_0 = r_2081; // @[Multiplier.scala 126:19]
  assign c32_24_io_in_1 = r_2082; // @[Multiplier.scala 126:19]
  assign c32_24_io_in_2 = r_2083; // @[Multiplier.scala 126:19]
  assign c53_483_io_in_0 = r_2084; // @[Multiplier.scala 132:13]
  assign c53_483_io_in_1 = r_2085; // @[Multiplier.scala 132:13]
  assign c53_483_io_in_2 = r_2086; // @[Multiplier.scala 132:13]
  assign c53_483_io_in_3 = r_2087; // @[Multiplier.scala 132:13]
  assign c53_483_io_in_4 = c53_480_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_484_io_in_0 = r_2088; // @[Multiplier.scala 132:13]
  assign c53_484_io_in_1 = r_2089; // @[Multiplier.scala 132:13]
  assign c53_484_io_in_2 = r_2090; // @[Multiplier.scala 132:13]
  assign c53_484_io_in_3 = r_2091; // @[Multiplier.scala 132:13]
  assign c53_484_io_in_4 = c53_481_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_485_io_in_0 = r_2092; // @[Multiplier.scala 132:13]
  assign c53_485_io_in_1 = r_2093; // @[Multiplier.scala 132:13]
  assign c53_485_io_in_2 = r_2094; // @[Multiplier.scala 132:13]
  assign c53_485_io_in_3 = r_2095; // @[Multiplier.scala 132:13]
  assign c53_485_io_in_4 = c53_482_io_out_1; // @[Multiplier.scala 136:41]
  assign c32_25_io_in_0 = r_2096; // @[Multiplier.scala 126:19]
  assign c32_25_io_in_1 = r_2097; // @[Multiplier.scala 126:19]
  assign c32_25_io_in_2 = r_2098; // @[Multiplier.scala 126:19]
  assign c53_486_io_in_0 = r_2099; // @[Multiplier.scala 132:13]
  assign c53_486_io_in_1 = r_2100; // @[Multiplier.scala 132:13]
  assign c53_486_io_in_2 = r_2101; // @[Multiplier.scala 132:13]
  assign c53_486_io_in_3 = r_2102; // @[Multiplier.scala 132:13]
  assign c53_486_io_in_4 = c53_483_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_487_io_in_0 = r_2103; // @[Multiplier.scala 132:13]
  assign c53_487_io_in_1 = r_2104; // @[Multiplier.scala 132:13]
  assign c53_487_io_in_2 = r_2105; // @[Multiplier.scala 132:13]
  assign c53_487_io_in_3 = r_2106; // @[Multiplier.scala 132:13]
  assign c53_487_io_in_4 = c53_484_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_488_io_in_0 = r_2107; // @[Multiplier.scala 132:13]
  assign c53_488_io_in_1 = r_2108; // @[Multiplier.scala 132:13]
  assign c53_488_io_in_2 = r_2109; // @[Multiplier.scala 132:13]
  assign c53_488_io_in_3 = r_2110; // @[Multiplier.scala 132:13]
  assign c53_488_io_in_4 = c53_485_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_24_io_in_0 = r_2111; // @[Multiplier.scala 121:19]
  assign c22_24_io_in_1 = r_2112; // @[Multiplier.scala 121:19]
  assign c53_489_io_in_0 = r_2113; // @[Multiplier.scala 132:13]
  assign c53_489_io_in_1 = r_2114; // @[Multiplier.scala 132:13]
  assign c53_489_io_in_2 = r_2115; // @[Multiplier.scala 132:13]
  assign c53_489_io_in_3 = r_2116; // @[Multiplier.scala 132:13]
  assign c53_489_io_in_4 = c53_486_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_490_io_in_0 = r_2117; // @[Multiplier.scala 132:13]
  assign c53_490_io_in_1 = r_2118; // @[Multiplier.scala 132:13]
  assign c53_490_io_in_2 = r_2119; // @[Multiplier.scala 132:13]
  assign c53_490_io_in_3 = r_2120; // @[Multiplier.scala 132:13]
  assign c53_490_io_in_4 = c53_487_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_491_io_in_0 = r_2121; // @[Multiplier.scala 132:13]
  assign c53_491_io_in_1 = r_2122; // @[Multiplier.scala 132:13]
  assign c53_491_io_in_2 = r_2123; // @[Multiplier.scala 132:13]
  assign c53_491_io_in_3 = r_2124; // @[Multiplier.scala 132:13]
  assign c53_491_io_in_4 = c53_488_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_25_io_in_0 = r_2125; // @[Multiplier.scala 121:19]
  assign c22_25_io_in_1 = r_2126; // @[Multiplier.scala 121:19]
  assign c53_492_io_in_0 = r_2127; // @[Multiplier.scala 132:13]
  assign c53_492_io_in_1 = r_2128; // @[Multiplier.scala 132:13]
  assign c53_492_io_in_2 = r_2129; // @[Multiplier.scala 132:13]
  assign c53_492_io_in_3 = r_2130; // @[Multiplier.scala 132:13]
  assign c53_492_io_in_4 = c53_489_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_493_io_in_0 = r_2131; // @[Multiplier.scala 132:13]
  assign c53_493_io_in_1 = r_2132; // @[Multiplier.scala 132:13]
  assign c53_493_io_in_2 = r_2133; // @[Multiplier.scala 132:13]
  assign c53_493_io_in_3 = r_2134; // @[Multiplier.scala 132:13]
  assign c53_493_io_in_4 = c53_490_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_494_io_in_0 = r_2135; // @[Multiplier.scala 132:13]
  assign c53_494_io_in_1 = r_2136; // @[Multiplier.scala 132:13]
  assign c53_494_io_in_2 = r_2137; // @[Multiplier.scala 132:13]
  assign c53_494_io_in_3 = r_2138; // @[Multiplier.scala 132:13]
  assign c53_494_io_in_4 = c53_491_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_495_io_in_0 = r_2140; // @[Multiplier.scala 132:13]
  assign c53_495_io_in_1 = r_2141; // @[Multiplier.scala 132:13]
  assign c53_495_io_in_2 = r_2142; // @[Multiplier.scala 132:13]
  assign c53_495_io_in_3 = r_2143; // @[Multiplier.scala 132:13]
  assign c53_495_io_in_4 = c53_492_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_496_io_in_0 = r_2144; // @[Multiplier.scala 132:13]
  assign c53_496_io_in_1 = r_2145; // @[Multiplier.scala 132:13]
  assign c53_496_io_in_2 = r_2146; // @[Multiplier.scala 132:13]
  assign c53_496_io_in_3 = r_2147; // @[Multiplier.scala 132:13]
  assign c53_496_io_in_4 = c53_493_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_497_io_in_0 = r_2148; // @[Multiplier.scala 132:13]
  assign c53_497_io_in_1 = r_2149; // @[Multiplier.scala 132:13]
  assign c53_497_io_in_2 = r_2150; // @[Multiplier.scala 132:13]
  assign c53_497_io_in_3 = r_2151; // @[Multiplier.scala 132:13]
  assign c53_497_io_in_4 = c53_494_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_498_io_in_0 = r_2153; // @[Multiplier.scala 132:13]
  assign c53_498_io_in_1 = r_2154; // @[Multiplier.scala 132:13]
  assign c53_498_io_in_2 = r_2155; // @[Multiplier.scala 132:13]
  assign c53_498_io_in_3 = r_2156; // @[Multiplier.scala 132:13]
  assign c53_498_io_in_4 = c53_495_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_499_io_in_0 = r_2157; // @[Multiplier.scala 132:13]
  assign c53_499_io_in_1 = r_2158; // @[Multiplier.scala 132:13]
  assign c53_499_io_in_2 = r_2159; // @[Multiplier.scala 132:13]
  assign c53_499_io_in_3 = r_2160; // @[Multiplier.scala 132:13]
  assign c53_499_io_in_4 = c53_496_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_500_io_in_0 = r_2161; // @[Multiplier.scala 132:13]
  assign c53_500_io_in_1 = r_2162; // @[Multiplier.scala 132:13]
  assign c53_500_io_in_2 = r_2163; // @[Multiplier.scala 132:13]
  assign c53_500_io_in_3 = r_2164; // @[Multiplier.scala 132:13]
  assign c53_500_io_in_4 = c53_497_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_501_io_in_0 = r_2165; // @[Multiplier.scala 132:13]
  assign c53_501_io_in_1 = r_2166; // @[Multiplier.scala 132:13]
  assign c53_501_io_in_2 = r_2167; // @[Multiplier.scala 132:13]
  assign c53_501_io_in_3 = r_2168; // @[Multiplier.scala 132:13]
  assign c53_501_io_in_4 = c53_498_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_502_io_in_0 = r_2169; // @[Multiplier.scala 132:13]
  assign c53_502_io_in_1 = r_2170; // @[Multiplier.scala 132:13]
  assign c53_502_io_in_2 = r_2171; // @[Multiplier.scala 132:13]
  assign c53_502_io_in_3 = r_2172; // @[Multiplier.scala 132:13]
  assign c53_502_io_in_4 = c53_499_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_503_io_in_0 = r_2173; // @[Multiplier.scala 132:13]
  assign c53_503_io_in_1 = r_2174; // @[Multiplier.scala 132:13]
  assign c53_503_io_in_2 = r_2175; // @[Multiplier.scala 132:13]
  assign c53_503_io_in_3 = r_2176; // @[Multiplier.scala 132:13]
  assign c53_503_io_in_4 = c53_500_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_504_io_in_0 = r_2177; // @[Multiplier.scala 132:13]
  assign c53_504_io_in_1 = r_2178; // @[Multiplier.scala 132:13]
  assign c53_504_io_in_2 = r_2179; // @[Multiplier.scala 132:13]
  assign c53_504_io_in_3 = r_2180; // @[Multiplier.scala 132:13]
  assign c53_504_io_in_4 = c53_501_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_505_io_in_0 = r_2181; // @[Multiplier.scala 132:13]
  assign c53_505_io_in_1 = r_2182; // @[Multiplier.scala 132:13]
  assign c53_505_io_in_2 = r_2183; // @[Multiplier.scala 132:13]
  assign c53_505_io_in_3 = r_2184; // @[Multiplier.scala 132:13]
  assign c53_505_io_in_4 = c53_502_io_out_1; // @[Multiplier.scala 136:41]
  assign c32_26_io_in_0 = r_2185; // @[Multiplier.scala 126:19]
  assign c32_26_io_in_1 = r_2186; // @[Multiplier.scala 126:19]
  assign c32_26_io_in_2 = r_2187; // @[Multiplier.scala 126:19]
  assign c53_506_io_in_0 = r_2188; // @[Multiplier.scala 132:13]
  assign c53_506_io_in_1 = r_2189; // @[Multiplier.scala 132:13]
  assign c53_506_io_in_2 = r_2190; // @[Multiplier.scala 132:13]
  assign c53_506_io_in_3 = r_2191; // @[Multiplier.scala 132:13]
  assign c53_506_io_in_4 = c53_504_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_507_io_in_0 = r_2192; // @[Multiplier.scala 132:13]
  assign c53_507_io_in_1 = r_2193; // @[Multiplier.scala 132:13]
  assign c53_507_io_in_2 = r_2194; // @[Multiplier.scala 132:13]
  assign c53_507_io_in_3 = r_2195; // @[Multiplier.scala 132:13]
  assign c53_507_io_in_4 = c53_505_io_out_1; // @[Multiplier.scala 136:41]
  assign c32_27_io_in_0 = r_2196; // @[Multiplier.scala 126:19]
  assign c32_27_io_in_1 = r_2197; // @[Multiplier.scala 126:19]
  assign c32_27_io_in_2 = r_2198; // @[Multiplier.scala 126:19]
  assign c53_508_io_in_0 = r_2199; // @[Multiplier.scala 132:13]
  assign c53_508_io_in_1 = r_2200; // @[Multiplier.scala 132:13]
  assign c53_508_io_in_2 = r_2201; // @[Multiplier.scala 132:13]
  assign c53_508_io_in_3 = r_2202; // @[Multiplier.scala 132:13]
  assign c53_508_io_in_4 = c53_506_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_509_io_in_0 = r_2203; // @[Multiplier.scala 132:13]
  assign c53_509_io_in_1 = r_2204; // @[Multiplier.scala 132:13]
  assign c53_509_io_in_2 = r_2205; // @[Multiplier.scala 132:13]
  assign c53_509_io_in_3 = r_2206; // @[Multiplier.scala 132:13]
  assign c53_509_io_in_4 = c53_507_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_26_io_in_0 = r_2207; // @[Multiplier.scala 121:19]
  assign c22_26_io_in_1 = r_2208; // @[Multiplier.scala 121:19]
  assign c53_510_io_in_0 = r_2209; // @[Multiplier.scala 132:13]
  assign c53_510_io_in_1 = r_2210; // @[Multiplier.scala 132:13]
  assign c53_510_io_in_2 = r_2211; // @[Multiplier.scala 132:13]
  assign c53_510_io_in_3 = r_2212; // @[Multiplier.scala 132:13]
  assign c53_510_io_in_4 = c53_508_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_511_io_in_0 = r_2213; // @[Multiplier.scala 132:13]
  assign c53_511_io_in_1 = r_2214; // @[Multiplier.scala 132:13]
  assign c53_511_io_in_2 = r_2215; // @[Multiplier.scala 132:13]
  assign c53_511_io_in_3 = r_2216; // @[Multiplier.scala 132:13]
  assign c53_511_io_in_4 = c53_509_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_27_io_in_0 = r_2217; // @[Multiplier.scala 121:19]
  assign c22_27_io_in_1 = r_2218; // @[Multiplier.scala 121:19]
  assign c53_512_io_in_0 = r_2219; // @[Multiplier.scala 132:13]
  assign c53_512_io_in_1 = r_2220; // @[Multiplier.scala 132:13]
  assign c53_512_io_in_2 = r_2221; // @[Multiplier.scala 132:13]
  assign c53_512_io_in_3 = r_2222; // @[Multiplier.scala 132:13]
  assign c53_512_io_in_4 = c53_510_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_513_io_in_0 = r_2223; // @[Multiplier.scala 132:13]
  assign c53_513_io_in_1 = r_2224; // @[Multiplier.scala 132:13]
  assign c53_513_io_in_2 = r_2225; // @[Multiplier.scala 132:13]
  assign c53_513_io_in_3 = r_2226; // @[Multiplier.scala 132:13]
  assign c53_513_io_in_4 = c53_511_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_514_io_in_0 = r_2228; // @[Multiplier.scala 132:13]
  assign c53_514_io_in_1 = r_2229; // @[Multiplier.scala 132:13]
  assign c53_514_io_in_2 = r_2230; // @[Multiplier.scala 132:13]
  assign c53_514_io_in_3 = r_2231; // @[Multiplier.scala 132:13]
  assign c53_514_io_in_4 = c53_512_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_515_io_in_0 = r_2232; // @[Multiplier.scala 132:13]
  assign c53_515_io_in_1 = r_2233; // @[Multiplier.scala 132:13]
  assign c53_515_io_in_2 = r_2234; // @[Multiplier.scala 132:13]
  assign c53_515_io_in_3 = r_2235; // @[Multiplier.scala 132:13]
  assign c53_515_io_in_4 = c53_513_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_516_io_in_0 = r_2237; // @[Multiplier.scala 132:13]
  assign c53_516_io_in_1 = r_2238; // @[Multiplier.scala 132:13]
  assign c53_516_io_in_2 = r_2239; // @[Multiplier.scala 132:13]
  assign c53_516_io_in_3 = r_2240; // @[Multiplier.scala 132:13]
  assign c53_516_io_in_4 = c53_514_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_517_io_in_0 = r_2241; // @[Multiplier.scala 132:13]
  assign c53_517_io_in_1 = r_2242; // @[Multiplier.scala 132:13]
  assign c53_517_io_in_2 = r_2243; // @[Multiplier.scala 132:13]
  assign c53_517_io_in_3 = r_2244; // @[Multiplier.scala 132:13]
  assign c53_517_io_in_4 = c53_515_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_518_io_in_0 = r_2245; // @[Multiplier.scala 132:13]
  assign c53_518_io_in_1 = r_2246; // @[Multiplier.scala 132:13]
  assign c53_518_io_in_2 = r_2247; // @[Multiplier.scala 132:13]
  assign c53_518_io_in_3 = r_2248; // @[Multiplier.scala 132:13]
  assign c53_518_io_in_4 = c53_516_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_519_io_in_0 = r_2249; // @[Multiplier.scala 132:13]
  assign c53_519_io_in_1 = r_2250; // @[Multiplier.scala 132:13]
  assign c53_519_io_in_2 = r_2251; // @[Multiplier.scala 132:13]
  assign c53_519_io_in_3 = r_2252; // @[Multiplier.scala 132:13]
  assign c53_519_io_in_4 = c53_517_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_520_io_in_0 = r_2253; // @[Multiplier.scala 132:13]
  assign c53_520_io_in_1 = r_2254; // @[Multiplier.scala 132:13]
  assign c53_520_io_in_2 = r_2255; // @[Multiplier.scala 132:13]
  assign c53_520_io_in_3 = r_2256; // @[Multiplier.scala 132:13]
  assign c53_520_io_in_4 = c53_518_io_out_1; // @[Multiplier.scala 136:41]
  assign c32_28_io_in_0 = r_2257; // @[Multiplier.scala 126:19]
  assign c32_28_io_in_1 = r_2258; // @[Multiplier.scala 126:19]
  assign c32_28_io_in_2 = r_2259; // @[Multiplier.scala 126:19]
  assign c53_521_io_in_0 = r_2260; // @[Multiplier.scala 132:13]
  assign c53_521_io_in_1 = r_2261; // @[Multiplier.scala 132:13]
  assign c53_521_io_in_2 = r_2262; // @[Multiplier.scala 132:13]
  assign c53_521_io_in_3 = r_2263; // @[Multiplier.scala 132:13]
  assign c53_521_io_in_4 = c53_520_io_out_1; // @[Multiplier.scala 136:41]
  assign c32_29_io_in_0 = r_2264; // @[Multiplier.scala 126:19]
  assign c32_29_io_in_1 = r_2265; // @[Multiplier.scala 126:19]
  assign c32_29_io_in_2 = r_2266; // @[Multiplier.scala 126:19]
  assign c53_522_io_in_0 = r_2267; // @[Multiplier.scala 132:13]
  assign c53_522_io_in_1 = r_2268; // @[Multiplier.scala 132:13]
  assign c53_522_io_in_2 = r_2269; // @[Multiplier.scala 132:13]
  assign c53_522_io_in_3 = r_2270; // @[Multiplier.scala 132:13]
  assign c53_522_io_in_4 = c53_521_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_28_io_in_0 = r_2271; // @[Multiplier.scala 121:19]
  assign c22_28_io_in_1 = r_2272; // @[Multiplier.scala 121:19]
  assign c53_523_io_in_0 = r_2273; // @[Multiplier.scala 132:13]
  assign c53_523_io_in_1 = r_2274; // @[Multiplier.scala 132:13]
  assign c53_523_io_in_2 = r_2275; // @[Multiplier.scala 132:13]
  assign c53_523_io_in_3 = r_2276; // @[Multiplier.scala 132:13]
  assign c53_523_io_in_4 = c53_522_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_29_io_in_0 = r_2277; // @[Multiplier.scala 121:19]
  assign c22_29_io_in_1 = r_2278; // @[Multiplier.scala 121:19]
  assign c53_524_io_in_0 = r_2279; // @[Multiplier.scala 132:13]
  assign c53_524_io_in_1 = r_2280; // @[Multiplier.scala 132:13]
  assign c53_524_io_in_2 = r_2281; // @[Multiplier.scala 132:13]
  assign c53_524_io_in_3 = r_2282; // @[Multiplier.scala 132:13]
  assign c53_524_io_in_4 = c53_523_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_525_io_in_0 = r_2284; // @[Multiplier.scala 132:13]
  assign c53_525_io_in_1 = r_2285; // @[Multiplier.scala 132:13]
  assign c53_525_io_in_2 = r_2286; // @[Multiplier.scala 132:13]
  assign c53_525_io_in_3 = r_2287; // @[Multiplier.scala 132:13]
  assign c53_525_io_in_4 = c53_524_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_526_io_in_0 = r_2289; // @[Multiplier.scala 132:13]
  assign c53_526_io_in_1 = r_2290; // @[Multiplier.scala 132:13]
  assign c53_526_io_in_2 = r_2291; // @[Multiplier.scala 132:13]
  assign c53_526_io_in_3 = r_2292; // @[Multiplier.scala 132:13]
  assign c53_526_io_in_4 = c53_525_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_527_io_in_0 = r_2293; // @[Multiplier.scala 132:13]
  assign c53_527_io_in_1 = r_2294; // @[Multiplier.scala 132:13]
  assign c53_527_io_in_2 = r_2295; // @[Multiplier.scala 132:13]
  assign c53_527_io_in_3 = r_2296; // @[Multiplier.scala 132:13]
  assign c53_527_io_in_4 = c53_526_io_out_1; // @[Multiplier.scala 136:41]
  assign c32_30_io_in_0 = r_2297; // @[Multiplier.scala 126:19]
  assign c32_30_io_in_1 = r_2298; // @[Multiplier.scala 126:19]
  assign c32_30_io_in_2 = r_2299; // @[Multiplier.scala 126:19]
  assign c32_31_io_in_0 = r_2300; // @[Multiplier.scala 126:19]
  assign c32_31_io_in_1 = r_2301; // @[Multiplier.scala 126:19]
  assign c32_31_io_in_2 = r_2302; // @[Multiplier.scala 126:19]
  assign c22_30_io_in_0 = r_2303; // @[Multiplier.scala 121:19]
  assign c22_30_io_in_1 = r_2304; // @[Multiplier.scala 121:19]
  assign c22_31_io_in_0 = r_2305; // @[Multiplier.scala 121:19]
  assign c22_31_io_in_1 = r_2306; // @[Multiplier.scala 121:19]
  assign c22_32_io_in_0 = c22_1_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_32_io_in_1 = c22_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_33_io_in_0 = c32_io_out_0; // @[Multiplier.scala 127:35]
  assign c22_33_io_in_1 = c22_1_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_34_io_in_0 = c32_1_io_out_0; // @[Multiplier.scala 127:35]
  assign c22_34_io_in_1 = c32_io_out_1; // @[Multiplier.scala 128:41]
  assign c22_35_io_in_0 = c53_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_35_io_in_1 = c32_1_io_out_1; // @[Multiplier.scala 128:41]
  assign c22_36_io_in_0 = c53_1_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_36_io_in_1 = c53_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_32_io_in_0 = c53_2_io_out_0; // @[Multiplier.scala 135:39]
  assign c32_32_io_in_1 = r_22; // @[Multiplier.scala 126:19]
  assign c32_32_io_in_2 = c53_1_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_33_io_in_0 = c53_3_io_out_0; // @[Multiplier.scala 135:39]
  assign c32_33_io_in_1 = r_27; // @[Multiplier.scala 126:19]
  assign c32_33_io_in_2 = c53_2_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_34_io_in_0 = c53_4_io_out_0; // @[Multiplier.scala 135:39]
  assign c32_34_io_in_1 = c22_2_io_out_0; // @[Multiplier.scala 122:35]
  assign c32_34_io_in_2 = c53_3_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_528_io_in_0 = c53_5_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_528_io_in_1 = c22_3_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_528_io_in_2 = c53_4_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_528_io_in_3 = c22_2_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_528_io_in_4 = 1'h0; // @[Multiplier.scala 134:24]
  assign c53_529_io_in_0 = c53_6_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_529_io_in_1 = c32_2_io_out_0; // @[Multiplier.scala 127:35]
  assign c53_529_io_in_2 = c53_5_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_529_io_in_3 = c22_3_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_529_io_in_4 = c53_528_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_530_io_in_0 = c53_7_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_530_io_in_1 = c32_3_io_out_0; // @[Multiplier.scala 127:35]
  assign c53_530_io_in_2 = c53_6_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_530_io_in_3 = c32_2_io_out_1; // @[Multiplier.scala 128:41]
  assign c53_530_io_in_4 = c53_529_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_531_io_in_0 = c53_8_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_531_io_in_1 = c53_9_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_531_io_in_2 = c53_7_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_531_io_in_3 = c32_3_io_out_1; // @[Multiplier.scala 128:41]
  assign c53_531_io_in_4 = c53_530_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_532_io_in_0 = c53_10_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_532_io_in_1 = c53_11_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_532_io_in_2 = c53_8_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_532_io_in_3 = c53_9_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_532_io_in_4 = c53_531_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_533_io_in_0 = c53_12_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_533_io_in_1 = c53_13_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_533_io_in_2 = r_78; // @[Multiplier.scala 132:13]
  assign c53_533_io_in_3 = c53_10_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_533_io_in_4 = c53_532_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_534_io_in_0 = c53_14_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_534_io_in_1 = c53_15_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_534_io_in_2 = r_87; // @[Multiplier.scala 132:13]
  assign c53_534_io_in_3 = c53_12_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_534_io_in_4 = c53_533_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_535_io_in_0 = c53_16_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_535_io_in_1 = c53_17_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_535_io_in_2 = c22_4_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_535_io_in_3 = c53_14_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_535_io_in_4 = c53_534_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_536_io_in_0 = c53_18_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_536_io_in_1 = c53_19_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_536_io_in_2 = c22_5_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_536_io_in_3 = c53_16_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_536_io_in_4 = c53_535_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_37_io_in_0 = c53_17_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_37_io_in_1 = c22_4_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_537_io_in_0 = c53_20_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_537_io_in_1 = c53_21_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_537_io_in_2 = c32_4_io_out_0; // @[Multiplier.scala 127:35]
  assign c53_537_io_in_3 = c53_18_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_537_io_in_4 = c53_536_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_38_io_in_0 = c53_19_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_38_io_in_1 = c22_5_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_538_io_in_0 = c53_22_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_538_io_in_1 = c53_23_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_538_io_in_2 = c32_5_io_out_0; // @[Multiplier.scala 127:35]
  assign c53_538_io_in_3 = c53_20_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_538_io_in_4 = c53_537_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_39_io_in_0 = c53_21_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_39_io_in_1 = c32_4_io_out_1; // @[Multiplier.scala 128:41]
  assign c53_539_io_in_0 = c53_24_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_539_io_in_1 = c53_25_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_539_io_in_2 = c53_26_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_539_io_in_3 = c53_22_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_539_io_in_4 = c53_538_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_40_io_in_0 = c53_23_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_40_io_in_1 = c32_5_io_out_1; // @[Multiplier.scala 128:41]
  assign c53_540_io_in_0 = c53_27_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_540_io_in_1 = c53_28_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_540_io_in_2 = c53_29_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_540_io_in_3 = c53_24_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_540_io_in_4 = c53_539_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_41_io_in_0 = c53_25_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_41_io_in_1 = c53_26_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_541_io_in_0 = c53_30_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_541_io_in_1 = c53_31_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_541_io_in_2 = c53_32_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_541_io_in_3 = r_166; // @[Multiplier.scala 132:13]
  assign c53_541_io_in_4 = c53_540_io_out_1; // @[Multiplier.scala 136:41]
  assign c32_35_io_in_0 = c53_27_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_35_io_in_1 = c53_28_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_35_io_in_2 = c53_29_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_542_io_in_0 = c53_33_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_542_io_in_1 = c53_34_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_542_io_in_2 = c53_35_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_542_io_in_3 = r_179; // @[Multiplier.scala 132:13]
  assign c53_542_io_in_4 = c53_541_io_out_1; // @[Multiplier.scala 136:41]
  assign c32_36_io_in_0 = c53_30_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_36_io_in_1 = c53_31_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_36_io_in_2 = c53_32_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_543_io_in_0 = c53_36_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_543_io_in_1 = c53_37_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_543_io_in_2 = c53_38_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_543_io_in_3 = c22_6_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_543_io_in_4 = c53_542_io_out_1; // @[Multiplier.scala 136:41]
  assign c32_37_io_in_0 = c53_33_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_37_io_in_1 = c53_34_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_37_io_in_2 = c53_35_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_544_io_in_0 = c53_39_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_544_io_in_1 = c53_40_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_544_io_in_2 = c53_41_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_544_io_in_3 = c22_7_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_544_io_in_4 = c53_543_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_545_io_in_0 = c53_36_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_545_io_in_1 = c53_37_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_545_io_in_2 = c53_38_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_545_io_in_3 = c22_6_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_545_io_in_4 = 1'h0; // @[Multiplier.scala 134:24]
  assign c53_546_io_in_0 = c53_42_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_546_io_in_1 = c53_43_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_546_io_in_2 = c53_44_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_546_io_in_3 = c32_6_io_out_0; // @[Multiplier.scala 127:35]
  assign c53_546_io_in_4 = c53_544_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_547_io_in_0 = c53_39_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_547_io_in_1 = c53_40_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_547_io_in_2 = c53_41_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_547_io_in_3 = c22_7_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_547_io_in_4 = c53_545_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_548_io_in_0 = c53_45_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_548_io_in_1 = c53_46_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_548_io_in_2 = c53_47_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_548_io_in_3 = c32_7_io_out_0; // @[Multiplier.scala 127:35]
  assign c53_548_io_in_4 = c53_546_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_549_io_in_0 = c53_42_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_549_io_in_1 = c53_43_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_549_io_in_2 = c53_44_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_549_io_in_3 = c32_6_io_out_1; // @[Multiplier.scala 128:41]
  assign c53_549_io_in_4 = c53_547_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_550_io_in_0 = c53_48_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_550_io_in_1 = c53_49_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_550_io_in_2 = c53_50_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_550_io_in_3 = c53_51_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_550_io_in_4 = c53_548_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_551_io_in_0 = c53_45_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_551_io_in_1 = c53_46_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_551_io_in_2 = c53_47_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_551_io_in_3 = c32_7_io_out_1; // @[Multiplier.scala 128:41]
  assign c53_551_io_in_4 = c53_549_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_552_io_in_0 = c53_52_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_552_io_in_1 = c53_53_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_552_io_in_2 = c53_54_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_552_io_in_3 = c53_55_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_552_io_in_4 = c53_550_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_553_io_in_0 = c53_48_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_553_io_in_1 = c53_49_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_553_io_in_2 = c53_50_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_553_io_in_3 = c53_51_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_553_io_in_4 = c53_551_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_554_io_in_0 = c53_56_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_554_io_in_1 = c53_57_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_554_io_in_2 = c53_58_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_554_io_in_3 = c53_59_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_554_io_in_4 = c53_552_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_555_io_in_0 = r_286; // @[Multiplier.scala 132:13]
  assign c53_555_io_in_1 = c53_52_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_555_io_in_2 = c53_53_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_555_io_in_3 = c53_54_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_555_io_in_4 = c53_553_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_556_io_in_0 = c53_60_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_556_io_in_1 = c53_61_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_556_io_in_2 = c53_62_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_556_io_in_3 = c53_63_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_556_io_in_4 = c53_554_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_557_io_in_0 = r_303; // @[Multiplier.scala 132:13]
  assign c53_557_io_in_1 = c53_56_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_557_io_in_2 = c53_57_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_557_io_in_3 = c53_58_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_557_io_in_4 = c53_555_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_558_io_in_0 = c53_64_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_558_io_in_1 = c53_65_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_558_io_in_2 = c53_66_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_558_io_in_3 = c53_67_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_558_io_in_4 = c53_556_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_559_io_in_0 = c22_8_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_559_io_in_1 = c53_60_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_559_io_in_2 = c53_61_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_559_io_in_3 = c53_62_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_559_io_in_4 = c53_557_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_560_io_in_0 = c53_68_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_560_io_in_1 = c53_69_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_560_io_in_2 = c53_70_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_560_io_in_3 = c53_71_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_560_io_in_4 = c53_558_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_561_io_in_0 = c22_9_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_561_io_in_1 = c53_64_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_561_io_in_2 = c53_65_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_561_io_in_3 = c53_66_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_561_io_in_4 = c53_559_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_42_io_in_0 = c53_67_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_42_io_in_1 = c22_8_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_562_io_in_0 = c53_72_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_562_io_in_1 = c53_73_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_562_io_in_2 = c53_74_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_562_io_in_3 = c53_75_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_562_io_in_4 = c53_560_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_563_io_in_0 = c32_8_io_out_0; // @[Multiplier.scala 127:35]
  assign c53_563_io_in_1 = c53_68_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_563_io_in_2 = c53_69_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_563_io_in_3 = c53_70_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_563_io_in_4 = c53_561_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_43_io_in_0 = c53_71_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_43_io_in_1 = c22_9_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_564_io_in_0 = c53_76_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_564_io_in_1 = c53_77_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_564_io_in_2 = c53_78_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_564_io_in_3 = c53_79_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_564_io_in_4 = c53_562_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_565_io_in_0 = c32_9_io_out_0; // @[Multiplier.scala 127:35]
  assign c53_565_io_in_1 = c53_72_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_565_io_in_2 = c53_73_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_565_io_in_3 = c53_74_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_565_io_in_4 = c53_563_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_44_io_in_0 = c53_75_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_44_io_in_1 = c32_8_io_out_1; // @[Multiplier.scala 128:41]
  assign c53_566_io_in_0 = c53_80_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_566_io_in_1 = c53_81_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_566_io_in_2 = c53_82_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_566_io_in_3 = c53_83_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_566_io_in_4 = c53_564_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_567_io_in_0 = c53_84_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_567_io_in_1 = c53_76_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_567_io_in_2 = c53_77_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_567_io_in_3 = c53_78_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_567_io_in_4 = c53_565_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_45_io_in_0 = c53_79_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_45_io_in_1 = c32_9_io_out_1; // @[Multiplier.scala 128:41]
  assign c53_568_io_in_0 = c53_85_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_568_io_in_1 = c53_86_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_568_io_in_2 = c53_87_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_568_io_in_3 = c53_88_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_568_io_in_4 = c53_566_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_569_io_in_0 = c53_89_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_569_io_in_1 = c53_80_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_569_io_in_2 = c53_81_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_569_io_in_3 = c53_82_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_569_io_in_4 = c53_567_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_46_io_in_0 = c53_83_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_46_io_in_1 = c53_84_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_570_io_in_0 = c53_90_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_570_io_in_1 = c53_91_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_570_io_in_2 = c53_92_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_570_io_in_3 = c53_93_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_570_io_in_4 = c53_568_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_571_io_in_0 = c53_94_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_571_io_in_1 = r_438; // @[Multiplier.scala 132:13]
  assign c53_571_io_in_2 = c53_85_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_571_io_in_3 = c53_86_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_571_io_in_4 = c53_569_io_out_1; // @[Multiplier.scala 136:41]
  assign c32_38_io_in_0 = c53_87_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_38_io_in_1 = c53_88_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_38_io_in_2 = c53_89_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_572_io_in_0 = c53_95_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_572_io_in_1 = c53_96_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_572_io_in_2 = c53_97_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_572_io_in_3 = c53_98_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_572_io_in_4 = c53_570_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_573_io_in_0 = c53_99_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_573_io_in_1 = r_459; // @[Multiplier.scala 132:13]
  assign c53_573_io_in_2 = c53_90_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_573_io_in_3 = c53_91_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_573_io_in_4 = c53_571_io_out_1; // @[Multiplier.scala 136:41]
  assign c32_39_io_in_0 = c53_92_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_39_io_in_1 = c53_93_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_39_io_in_2 = c53_94_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_574_io_in_0 = c53_100_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_574_io_in_1 = c53_101_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_574_io_in_2 = c53_102_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_574_io_in_3 = c53_103_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_574_io_in_4 = c53_572_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_575_io_in_0 = c53_104_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_575_io_in_1 = c22_10_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_575_io_in_2 = c53_95_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_575_io_in_3 = c53_96_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_575_io_in_4 = c53_573_io_out_1; // @[Multiplier.scala 136:41]
  assign c32_40_io_in_0 = c53_97_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_40_io_in_1 = c53_98_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_40_io_in_2 = c53_99_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_576_io_in_0 = c53_105_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_576_io_in_1 = c53_106_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_576_io_in_2 = c53_107_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_576_io_in_3 = c53_108_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_576_io_in_4 = c53_574_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_577_io_in_0 = c53_109_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_577_io_in_1 = c22_11_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_577_io_in_2 = c53_100_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_577_io_in_3 = c53_101_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_577_io_in_4 = c53_575_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_578_io_in_0 = c53_102_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_578_io_in_1 = c53_103_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_578_io_in_2 = c53_104_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_578_io_in_3 = c22_10_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_578_io_in_4 = 1'h0; // @[Multiplier.scala 134:24]
  assign c53_579_io_in_0 = c53_110_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_579_io_in_1 = c53_111_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_579_io_in_2 = c53_112_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_579_io_in_3 = c53_113_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_579_io_in_4 = c53_576_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_580_io_in_0 = c53_114_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_580_io_in_1 = c32_10_io_out_0; // @[Multiplier.scala 127:35]
  assign c53_580_io_in_2 = c53_105_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_580_io_in_3 = c53_106_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_580_io_in_4 = c53_577_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_581_io_in_0 = c53_107_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_581_io_in_1 = c53_108_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_581_io_in_2 = c53_109_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_581_io_in_3 = c22_11_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_581_io_in_4 = c53_578_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_582_io_in_0 = c53_115_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_582_io_in_1 = c53_116_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_582_io_in_2 = c53_117_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_582_io_in_3 = c53_118_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_582_io_in_4 = c53_579_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_583_io_in_0 = c53_119_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_583_io_in_1 = c32_11_io_out_0; // @[Multiplier.scala 127:35]
  assign c53_583_io_in_2 = c53_110_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_583_io_in_3 = c53_111_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_583_io_in_4 = c53_580_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_584_io_in_0 = c53_112_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_584_io_in_1 = c53_113_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_584_io_in_2 = c53_114_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_584_io_in_3 = c32_10_io_out_1; // @[Multiplier.scala 128:41]
  assign c53_584_io_in_4 = c53_581_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_585_io_in_0 = c53_120_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_585_io_in_1 = c53_121_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_585_io_in_2 = c53_122_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_585_io_in_3 = c53_123_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_585_io_in_4 = c53_582_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_586_io_in_0 = c53_124_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_586_io_in_1 = c53_125_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_586_io_in_2 = c53_115_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_586_io_in_3 = c53_116_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_586_io_in_4 = c53_583_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_587_io_in_0 = c53_117_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_587_io_in_1 = c53_118_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_587_io_in_2 = c53_119_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_587_io_in_3 = c32_11_io_out_1; // @[Multiplier.scala 128:41]
  assign c53_587_io_in_4 = c53_584_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_588_io_in_0 = c53_126_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_588_io_in_1 = c53_127_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_588_io_in_2 = c53_128_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_588_io_in_3 = c53_129_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_588_io_in_4 = c53_585_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_589_io_in_0 = c53_130_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_589_io_in_1 = c53_131_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_589_io_in_2 = c53_120_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_589_io_in_3 = c53_121_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_589_io_in_4 = c53_586_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_590_io_in_0 = c53_122_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_590_io_in_1 = c53_123_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_590_io_in_2 = c53_124_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_590_io_in_3 = c53_125_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_590_io_in_4 = c53_587_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_591_io_in_0 = c53_132_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_591_io_in_1 = c53_133_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_591_io_in_2 = c53_134_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_591_io_in_3 = c53_135_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_591_io_in_4 = c53_588_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_592_io_in_0 = c53_136_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_592_io_in_1 = c53_137_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_592_io_in_2 = r_622; // @[Multiplier.scala 132:13]
  assign c53_592_io_in_3 = c53_126_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_592_io_in_4 = c53_589_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_593_io_in_0 = c53_127_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_593_io_in_1 = c53_128_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_593_io_in_2 = c53_129_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_593_io_in_3 = c53_130_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_593_io_in_4 = c53_590_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_594_io_in_0 = c53_138_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_594_io_in_1 = c53_139_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_594_io_in_2 = c53_140_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_594_io_in_3 = c53_141_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_594_io_in_4 = c53_591_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_595_io_in_0 = c53_142_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_595_io_in_1 = c53_143_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_595_io_in_2 = r_647; // @[Multiplier.scala 132:13]
  assign c53_595_io_in_3 = c53_132_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_595_io_in_4 = c53_592_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_596_io_in_0 = c53_133_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_596_io_in_1 = c53_134_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_596_io_in_2 = c53_135_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_596_io_in_3 = c53_136_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_596_io_in_4 = c53_593_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_597_io_in_0 = c53_144_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_597_io_in_1 = c53_145_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_597_io_in_2 = c53_146_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_597_io_in_3 = c53_147_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_597_io_in_4 = c53_594_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_598_io_in_0 = c53_148_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_598_io_in_1 = c53_149_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_598_io_in_2 = c22_12_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_598_io_in_3 = c53_138_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_598_io_in_4 = c53_595_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_599_io_in_0 = c53_139_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_599_io_in_1 = c53_140_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_599_io_in_2 = c53_141_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_599_io_in_3 = c53_142_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_599_io_in_4 = c53_596_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_600_io_in_0 = c53_150_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_600_io_in_1 = c53_151_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_600_io_in_2 = c53_152_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_600_io_in_3 = c53_153_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_600_io_in_4 = c53_597_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_601_io_in_0 = c53_154_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_601_io_in_1 = c53_155_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_601_io_in_2 = c22_13_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_601_io_in_3 = c53_144_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_601_io_in_4 = c53_598_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_602_io_in_0 = c53_145_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_602_io_in_1 = c53_146_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_602_io_in_2 = c53_147_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_602_io_in_3 = c53_148_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_602_io_in_4 = c53_599_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_47_io_in_0 = c53_149_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_47_io_in_1 = c22_12_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_603_io_in_0 = c53_156_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_603_io_in_1 = c53_157_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_603_io_in_2 = c53_158_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_603_io_in_3 = c53_159_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_603_io_in_4 = c53_600_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_604_io_in_0 = c53_160_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_604_io_in_1 = c53_161_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_604_io_in_2 = c32_12_io_out_0; // @[Multiplier.scala 127:35]
  assign c53_604_io_in_3 = c53_150_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_604_io_in_4 = c53_601_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_605_io_in_0 = c53_151_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_605_io_in_1 = c53_152_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_605_io_in_2 = c53_153_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_605_io_in_3 = c53_154_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_605_io_in_4 = c53_602_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_48_io_in_0 = c53_155_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_48_io_in_1 = c22_13_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_606_io_in_0 = c53_162_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_606_io_in_1 = c53_163_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_606_io_in_2 = c53_164_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_606_io_in_3 = c53_165_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_606_io_in_4 = c53_603_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_607_io_in_0 = c53_166_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_607_io_in_1 = c53_167_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_607_io_in_2 = c32_13_io_out_0; // @[Multiplier.scala 127:35]
  assign c53_607_io_in_3 = c53_156_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_607_io_in_4 = c53_604_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_608_io_in_0 = c53_157_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_608_io_in_1 = c53_158_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_608_io_in_2 = c53_159_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_608_io_in_3 = c53_160_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_608_io_in_4 = c53_605_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_49_io_in_0 = c53_161_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_49_io_in_1 = c32_12_io_out_1; // @[Multiplier.scala 128:41]
  assign c53_609_io_in_0 = c53_168_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_609_io_in_1 = c53_169_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_609_io_in_2 = c53_170_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_609_io_in_3 = c53_171_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_609_io_in_4 = c53_606_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_610_io_in_0 = c53_172_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_610_io_in_1 = c53_173_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_610_io_in_2 = c53_174_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_610_io_in_3 = c53_162_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_610_io_in_4 = c53_607_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_611_io_in_0 = c53_163_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_611_io_in_1 = c53_164_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_611_io_in_2 = c53_165_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_611_io_in_3 = c53_166_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_611_io_in_4 = c53_608_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_50_io_in_0 = c53_167_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_50_io_in_1 = c32_13_io_out_1; // @[Multiplier.scala 128:41]
  assign c53_612_io_in_0 = c53_175_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_612_io_in_1 = c53_176_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_612_io_in_2 = c53_177_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_612_io_in_3 = c53_178_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_612_io_in_4 = c53_609_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_613_io_in_0 = c53_179_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_613_io_in_1 = c53_180_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_613_io_in_2 = c53_181_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_613_io_in_3 = c53_168_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_613_io_in_4 = c53_610_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_614_io_in_0 = c53_169_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_614_io_in_1 = c53_170_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_614_io_in_2 = c53_171_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_614_io_in_3 = c53_172_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_614_io_in_4 = c53_611_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_51_io_in_0 = c53_173_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_51_io_in_1 = c53_174_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_615_io_in_0 = c53_182_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_615_io_in_1 = c53_183_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_615_io_in_2 = c53_184_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_615_io_in_3 = c53_185_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_615_io_in_4 = c53_612_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_616_io_in_0 = c53_186_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_616_io_in_1 = c53_187_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_616_io_in_2 = c53_188_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_616_io_in_3 = r_838; // @[Multiplier.scala 132:13]
  assign c53_616_io_in_4 = c53_613_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_617_io_in_0 = c53_175_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_617_io_in_1 = c53_176_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_617_io_in_2 = c53_177_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_617_io_in_3 = c53_178_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_617_io_in_4 = c53_614_io_out_1; // @[Multiplier.scala 136:41]
  assign c32_41_io_in_0 = c53_179_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_41_io_in_1 = c53_180_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_41_io_in_2 = c53_181_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_618_io_in_0 = c53_189_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_618_io_in_1 = c53_190_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_618_io_in_2 = c53_191_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_618_io_in_3 = c53_192_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_618_io_in_4 = c53_615_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_619_io_in_0 = c53_193_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_619_io_in_1 = c53_194_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_619_io_in_2 = c53_195_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_619_io_in_3 = r_867; // @[Multiplier.scala 132:13]
  assign c53_619_io_in_4 = c53_616_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_620_io_in_0 = c53_182_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_620_io_in_1 = c53_183_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_620_io_in_2 = c53_184_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_620_io_in_3 = c53_185_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_620_io_in_4 = c53_617_io_out_1; // @[Multiplier.scala 136:41]
  assign c32_42_io_in_0 = c53_186_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_42_io_in_1 = c53_187_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_42_io_in_2 = c53_188_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_621_io_in_0 = c53_196_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_621_io_in_1 = c53_197_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_621_io_in_2 = c53_198_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_621_io_in_3 = c53_199_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_621_io_in_4 = c53_618_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_622_io_in_0 = c53_200_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_622_io_in_1 = c53_201_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_622_io_in_2 = c53_202_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_622_io_in_3 = c22_14_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_622_io_in_4 = c53_619_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_623_io_in_0 = c53_189_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_623_io_in_1 = c53_190_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_623_io_in_2 = c53_191_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_623_io_in_3 = c53_192_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_623_io_in_4 = c53_620_io_out_1; // @[Multiplier.scala 136:41]
  assign c32_43_io_in_0 = c53_193_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_43_io_in_1 = c53_194_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_43_io_in_2 = c53_195_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_624_io_in_0 = c53_203_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_624_io_in_1 = c53_204_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_624_io_in_2 = c53_205_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_624_io_in_3 = c53_206_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_624_io_in_4 = c53_621_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_625_io_in_0 = c53_207_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_625_io_in_1 = c53_208_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_625_io_in_2 = c53_209_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_625_io_in_3 = c22_15_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_625_io_in_4 = c53_622_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_626_io_in_0 = c53_196_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_626_io_in_1 = c53_197_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_626_io_in_2 = c53_198_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_626_io_in_3 = c53_199_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_626_io_in_4 = c53_623_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_627_io_in_0 = c53_200_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_627_io_in_1 = c53_201_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_627_io_in_2 = c53_202_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_627_io_in_3 = c22_14_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_627_io_in_4 = 1'h0; // @[Multiplier.scala 134:24]
  assign c53_628_io_in_0 = c53_210_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_628_io_in_1 = c53_211_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_628_io_in_2 = c53_212_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_628_io_in_3 = c53_213_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_628_io_in_4 = c53_624_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_629_io_in_0 = c53_214_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_629_io_in_1 = c53_215_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_629_io_in_2 = c53_216_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_629_io_in_3 = c32_14_io_out_0; // @[Multiplier.scala 127:35]
  assign c53_629_io_in_4 = c53_625_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_630_io_in_0 = c53_203_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_630_io_in_1 = c53_204_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_630_io_in_2 = c53_205_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_630_io_in_3 = c53_206_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_630_io_in_4 = c53_626_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_631_io_in_0 = c53_207_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_631_io_in_1 = c53_208_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_631_io_in_2 = c53_209_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_631_io_in_3 = c22_15_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_631_io_in_4 = c53_627_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_632_io_in_0 = c53_217_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_632_io_in_1 = c53_218_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_632_io_in_2 = c53_219_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_632_io_in_3 = c53_220_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_632_io_in_4 = c53_628_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_633_io_in_0 = c53_221_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_633_io_in_1 = c53_222_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_633_io_in_2 = c53_223_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_633_io_in_3 = c32_15_io_out_0; // @[Multiplier.scala 127:35]
  assign c53_633_io_in_4 = c53_629_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_634_io_in_0 = c53_210_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_634_io_in_1 = c53_211_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_634_io_in_2 = c53_212_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_634_io_in_3 = c53_213_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_634_io_in_4 = c53_630_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_635_io_in_0 = c53_214_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_635_io_in_1 = c53_215_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_635_io_in_2 = c53_216_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_635_io_in_3 = c32_14_io_out_1; // @[Multiplier.scala 128:41]
  assign c53_635_io_in_4 = c53_631_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_636_io_in_0 = c53_224_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_636_io_in_1 = c53_225_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_636_io_in_2 = c53_226_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_636_io_in_3 = c53_227_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_636_io_in_4 = c53_632_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_637_io_in_0 = c53_228_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_637_io_in_1 = c53_229_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_637_io_in_2 = c53_230_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_637_io_in_3 = c53_231_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_637_io_in_4 = c53_633_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_638_io_in_0 = c53_217_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_638_io_in_1 = c53_218_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_638_io_in_2 = c53_219_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_638_io_in_3 = c53_220_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_638_io_in_4 = c53_634_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_639_io_in_0 = c53_221_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_639_io_in_1 = c53_222_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_639_io_in_2 = c53_223_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_639_io_in_3 = c32_15_io_out_1; // @[Multiplier.scala 128:41]
  assign c53_639_io_in_4 = c53_635_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_640_io_in_0 = c53_232_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_640_io_in_1 = c53_233_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_640_io_in_2 = c53_234_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_640_io_in_3 = c53_235_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_640_io_in_4 = c53_636_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_641_io_in_0 = c53_236_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_641_io_in_1 = c53_237_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_641_io_in_2 = c53_238_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_641_io_in_3 = c53_239_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_641_io_in_4 = c53_637_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_642_io_in_0 = c53_224_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_642_io_in_1 = c53_225_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_642_io_in_2 = c53_226_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_642_io_in_3 = c53_227_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_642_io_in_4 = c53_638_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_643_io_in_0 = c53_228_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_643_io_in_1 = c53_229_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_643_io_in_2 = c53_230_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_643_io_in_3 = c53_231_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_643_io_in_4 = c53_639_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_644_io_in_0 = c53_240_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_644_io_in_1 = c53_241_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_644_io_in_2 = c53_242_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_644_io_in_3 = c53_243_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_644_io_in_4 = c53_640_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_645_io_in_0 = c53_244_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_645_io_in_1 = c53_245_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_645_io_in_2 = c53_246_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_645_io_in_3 = c53_247_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_645_io_in_4 = c53_641_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_646_io_in_0 = r_1086; // @[Multiplier.scala 132:13]
  assign c53_646_io_in_1 = c53_232_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_646_io_in_2 = c53_233_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_646_io_in_3 = c53_234_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_646_io_in_4 = c53_642_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_647_io_in_0 = c53_235_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_647_io_in_1 = c53_236_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_647_io_in_2 = c53_237_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_647_io_in_3 = c53_238_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_647_io_in_4 = c53_643_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_648_io_in_0 = c53_248_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_648_io_in_1 = c53_249_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_648_io_in_2 = c53_250_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_648_io_in_3 = c53_251_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_648_io_in_4 = c53_644_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_649_io_in_0 = c53_252_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_649_io_in_1 = c53_253_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_649_io_in_2 = c53_254_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_649_io_in_3 = c53_255_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_649_io_in_4 = c53_645_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_650_io_in_0 = r_1119; // @[Multiplier.scala 132:13]
  assign c53_650_io_in_1 = c53_240_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_650_io_in_2 = c53_241_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_650_io_in_3 = c53_242_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_650_io_in_4 = c53_646_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_651_io_in_0 = c53_243_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_651_io_in_1 = c53_244_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_651_io_in_2 = c53_245_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_651_io_in_3 = c53_246_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_651_io_in_4 = c53_647_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_652_io_in_0 = c53_256_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_652_io_in_1 = c53_257_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_652_io_in_2 = c53_258_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_652_io_in_3 = c53_259_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_652_io_in_4 = c53_648_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_653_io_in_0 = c53_260_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_653_io_in_1 = c53_261_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_653_io_in_2 = c53_262_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_653_io_in_3 = c53_263_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_653_io_in_4 = c53_649_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_654_io_in_0 = r_1152; // @[Multiplier.scala 132:13]
  assign c53_654_io_in_1 = c53_248_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_654_io_in_2 = c53_249_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_654_io_in_3 = c53_250_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_654_io_in_4 = c53_650_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_655_io_in_0 = c53_251_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_655_io_in_1 = c53_252_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_655_io_in_2 = c53_253_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_655_io_in_3 = c53_254_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_655_io_in_4 = c53_651_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_656_io_in_0 = c53_264_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_656_io_in_1 = c53_265_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_656_io_in_2 = c53_266_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_656_io_in_3 = c53_267_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_656_io_in_4 = c53_652_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_657_io_in_0 = c53_268_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_657_io_in_1 = c53_269_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_657_io_in_2 = c53_270_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_657_io_in_3 = c53_271_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_657_io_in_4 = c53_653_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_658_io_in_0 = r_1185; // @[Multiplier.scala 132:13]
  assign c53_658_io_in_1 = c53_256_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_658_io_in_2 = c53_257_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_658_io_in_3 = c53_258_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_658_io_in_4 = c53_654_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_659_io_in_0 = c53_259_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_659_io_in_1 = c53_260_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_659_io_in_2 = c53_261_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_659_io_in_3 = c53_262_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_659_io_in_4 = c53_655_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_660_io_in_0 = c53_272_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_660_io_in_1 = c53_273_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_660_io_in_2 = c53_274_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_660_io_in_3 = c53_275_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_660_io_in_4 = c53_656_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_661_io_in_0 = c53_276_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_661_io_in_1 = c53_277_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_661_io_in_2 = c53_278_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_661_io_in_3 = c53_279_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_661_io_in_4 = c53_657_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_662_io_in_0 = r_1218; // @[Multiplier.scala 132:13]
  assign c53_662_io_in_1 = c53_264_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_662_io_in_2 = c53_265_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_662_io_in_3 = c53_266_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_662_io_in_4 = c53_658_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_663_io_in_0 = c53_267_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_663_io_in_1 = c53_268_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_663_io_in_2 = c53_269_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_663_io_in_3 = c53_270_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_663_io_in_4 = c53_659_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_664_io_in_0 = c53_280_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_664_io_in_1 = c53_281_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_664_io_in_2 = c53_282_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_664_io_in_3 = c53_283_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_664_io_in_4 = c53_660_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_665_io_in_0 = c53_284_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_665_io_in_1 = c53_285_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_665_io_in_2 = c53_286_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_665_io_in_3 = c53_287_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_665_io_in_4 = c53_661_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_666_io_in_0 = r_1251; // @[Multiplier.scala 132:13]
  assign c53_666_io_in_1 = c53_272_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_666_io_in_2 = c53_273_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_666_io_in_3 = c53_274_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_666_io_in_4 = c53_662_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_667_io_in_0 = c53_275_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_667_io_in_1 = c53_276_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_667_io_in_2 = c53_277_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_667_io_in_3 = c53_278_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_667_io_in_4 = c53_663_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_668_io_in_0 = c53_288_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_668_io_in_1 = c53_289_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_668_io_in_2 = c53_290_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_668_io_in_3 = c53_291_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_668_io_in_4 = c53_664_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_669_io_in_0 = c53_292_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_669_io_in_1 = c53_293_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_669_io_in_2 = c53_294_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_669_io_in_3 = c53_295_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_669_io_in_4 = c53_665_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_670_io_in_0 = r_1284; // @[Multiplier.scala 132:13]
  assign c53_670_io_in_1 = c53_280_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_670_io_in_2 = c53_281_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_670_io_in_3 = c53_282_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_670_io_in_4 = c53_666_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_671_io_in_0 = c53_283_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_671_io_in_1 = c53_284_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_671_io_in_2 = c53_285_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_671_io_in_3 = c53_286_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_671_io_in_4 = c53_667_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_672_io_in_0 = c53_296_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_672_io_in_1 = c53_297_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_672_io_in_2 = c53_298_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_672_io_in_3 = c53_299_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_672_io_in_4 = c53_668_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_673_io_in_0 = c53_300_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_673_io_in_1 = c53_301_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_673_io_in_2 = c53_302_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_673_io_in_3 = c53_303_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_673_io_in_4 = c53_669_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_674_io_in_0 = c53_288_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_674_io_in_1 = c53_289_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_674_io_in_2 = c53_290_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_674_io_in_3 = c53_291_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_674_io_in_4 = c53_670_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_675_io_in_0 = c53_292_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_675_io_in_1 = c53_293_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_675_io_in_2 = c53_294_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_675_io_in_3 = c53_295_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_675_io_in_4 = c53_671_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_676_io_in_0 = c53_304_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_676_io_in_1 = c53_305_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_676_io_in_2 = c53_306_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_676_io_in_3 = c53_307_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_676_io_in_4 = c53_672_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_677_io_in_0 = c53_308_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_677_io_in_1 = c53_309_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_677_io_in_2 = c53_310_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_677_io_in_3 = c32_16_io_out_0; // @[Multiplier.scala 127:35]
  assign c53_677_io_in_4 = c53_673_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_678_io_in_0 = c53_303_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_678_io_in_1 = c53_296_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_678_io_in_2 = c53_297_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_678_io_in_3 = c53_298_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_678_io_in_4 = c53_674_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_679_io_in_0 = c53_299_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_679_io_in_1 = c53_300_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_679_io_in_2 = c53_301_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_679_io_in_3 = c53_302_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_679_io_in_4 = c53_675_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_680_io_in_0 = c53_311_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_680_io_in_1 = c53_312_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_680_io_in_2 = c53_313_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_680_io_in_3 = c53_314_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_680_io_in_4 = c53_676_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_681_io_in_0 = c53_315_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_681_io_in_1 = c53_316_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_681_io_in_2 = c53_317_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_681_io_in_3 = c32_17_io_out_0; // @[Multiplier.scala 127:35]
  assign c53_681_io_in_4 = c53_677_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_682_io_in_0 = c53_304_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_682_io_in_1 = c53_305_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_682_io_in_2 = c53_306_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_682_io_in_3 = c53_307_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_682_io_in_4 = c53_678_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_683_io_in_0 = c53_308_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_683_io_in_1 = c53_309_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_683_io_in_2 = c53_310_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_683_io_in_3 = c32_16_io_out_1; // @[Multiplier.scala 128:41]
  assign c53_683_io_in_4 = c53_679_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_684_io_in_0 = c53_318_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_684_io_in_1 = c53_319_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_684_io_in_2 = c53_320_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_684_io_in_3 = c53_321_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_684_io_in_4 = c53_680_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_685_io_in_0 = c53_322_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_685_io_in_1 = c53_323_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_685_io_in_2 = c53_324_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_685_io_in_3 = c22_16_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_685_io_in_4 = c53_681_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_686_io_in_0 = c53_311_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_686_io_in_1 = c53_312_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_686_io_in_2 = c53_313_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_686_io_in_3 = c53_314_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_686_io_in_4 = c53_682_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_687_io_in_0 = c53_315_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_687_io_in_1 = c53_316_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_687_io_in_2 = c53_317_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_687_io_in_3 = c32_17_io_out_1; // @[Multiplier.scala 128:41]
  assign c53_687_io_in_4 = c53_683_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_688_io_in_0 = c53_325_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_688_io_in_1 = c53_326_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_688_io_in_2 = c53_327_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_688_io_in_3 = c53_328_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_688_io_in_4 = c53_684_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_689_io_in_0 = c53_329_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_689_io_in_1 = c53_330_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_689_io_in_2 = c53_331_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_689_io_in_3 = c22_17_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_689_io_in_4 = c53_685_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_690_io_in_0 = c53_318_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_690_io_in_1 = c53_319_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_690_io_in_2 = c53_320_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_690_io_in_3 = c53_321_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_690_io_in_4 = c53_686_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_691_io_in_0 = c53_322_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_691_io_in_1 = c53_323_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_691_io_in_2 = c53_324_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_691_io_in_3 = c22_16_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_691_io_in_4 = c53_687_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_692_io_in_0 = c53_332_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_692_io_in_1 = c53_333_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_692_io_in_2 = c53_334_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_692_io_in_3 = c53_335_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_692_io_in_4 = c53_688_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_693_io_in_0 = c53_336_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_693_io_in_1 = c53_337_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_693_io_in_2 = c53_338_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_693_io_in_3 = r_1467; // @[Multiplier.scala 132:13]
  assign c53_693_io_in_4 = c53_689_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_694_io_in_0 = c53_325_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_694_io_in_1 = c53_326_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_694_io_in_2 = c53_327_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_694_io_in_3 = c53_328_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_694_io_in_4 = c53_690_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_695_io_in_0 = c53_329_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_695_io_in_1 = c53_330_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_695_io_in_2 = c53_331_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_695_io_in_3 = c22_17_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_695_io_in_4 = c53_691_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_696_io_in_0 = c53_339_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_696_io_in_1 = c53_340_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_696_io_in_2 = c53_341_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_696_io_in_3 = c53_342_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_696_io_in_4 = c53_692_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_697_io_in_0 = c53_343_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_697_io_in_1 = c53_344_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_697_io_in_2 = c53_345_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_697_io_in_3 = r_1496; // @[Multiplier.scala 132:13]
  assign c53_697_io_in_4 = c53_693_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_698_io_in_0 = c53_332_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_698_io_in_1 = c53_333_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_698_io_in_2 = c53_334_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_698_io_in_3 = c53_335_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_698_io_in_4 = c53_694_io_out_1; // @[Multiplier.scala 136:41]
  assign c32_44_io_in_0 = c53_336_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_44_io_in_1 = c53_337_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_44_io_in_2 = c53_338_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_699_io_in_0 = c53_346_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_699_io_in_1 = c53_347_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_699_io_in_2 = c53_348_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_699_io_in_3 = c53_349_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_699_io_in_4 = c53_696_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_700_io_in_0 = c53_350_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_700_io_in_1 = c53_351_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_700_io_in_2 = c53_352_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_700_io_in_3 = c53_339_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_700_io_in_4 = c53_697_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_701_io_in_0 = c53_340_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_701_io_in_1 = c53_341_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_701_io_in_2 = c53_342_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_701_io_in_3 = c53_343_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_701_io_in_4 = c53_698_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_52_io_in_0 = c53_344_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_52_io_in_1 = c53_345_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_702_io_in_0 = c53_353_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_702_io_in_1 = c53_354_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_702_io_in_2 = c53_355_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_702_io_in_3 = c53_356_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_702_io_in_4 = c53_699_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_703_io_in_0 = c53_357_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_703_io_in_1 = c53_358_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_703_io_in_2 = c53_359_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_703_io_in_3 = c53_346_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_703_io_in_4 = c53_700_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_704_io_in_0 = c53_347_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_704_io_in_1 = c53_348_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_704_io_in_2 = c53_349_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_704_io_in_3 = c53_350_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_704_io_in_4 = c53_701_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_53_io_in_0 = c53_351_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_53_io_in_1 = c53_352_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_705_io_in_0 = c53_360_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_705_io_in_1 = c53_361_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_705_io_in_2 = c53_362_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_705_io_in_3 = c53_363_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_705_io_in_4 = c53_702_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_706_io_in_0 = c53_364_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_706_io_in_1 = c53_365_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_706_io_in_2 = c32_18_io_out_0; // @[Multiplier.scala 127:35]
  assign c53_706_io_in_3 = c53_359_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_706_io_in_4 = c53_703_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_707_io_in_0 = c53_353_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_707_io_in_1 = c53_354_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_707_io_in_2 = c53_355_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_707_io_in_3 = c53_356_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_707_io_in_4 = c53_704_io_out_1; // @[Multiplier.scala 136:41]
  assign c32_45_io_in_0 = c53_357_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_45_io_in_1 = c53_358_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_45_io_in_2 = c53_359_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_708_io_in_0 = c53_366_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_708_io_in_1 = c53_367_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_708_io_in_2 = c53_368_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_708_io_in_3 = c53_369_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_708_io_in_4 = c53_705_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_709_io_in_0 = c53_370_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_709_io_in_1 = c53_371_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_709_io_in_2 = c32_19_io_out_0; // @[Multiplier.scala 127:35]
  assign c53_709_io_in_3 = c53_360_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_709_io_in_4 = c53_706_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_710_io_in_0 = c53_361_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_710_io_in_1 = c53_362_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_710_io_in_2 = c53_363_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_710_io_in_3 = c53_364_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_710_io_in_4 = c53_707_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_54_io_in_0 = c53_365_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_54_io_in_1 = c32_18_io_out_1; // @[Multiplier.scala 128:41]
  assign c53_711_io_in_0 = c53_372_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_711_io_in_1 = c53_373_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_711_io_in_2 = c53_374_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_711_io_in_3 = c53_375_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_711_io_in_4 = c53_708_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_712_io_in_0 = c53_376_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_712_io_in_1 = c53_377_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_712_io_in_2 = c22_18_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_712_io_in_3 = c53_366_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_712_io_in_4 = c53_709_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_713_io_in_0 = c53_367_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_713_io_in_1 = c53_368_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_713_io_in_2 = c53_369_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_713_io_in_3 = c53_370_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_713_io_in_4 = c53_710_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_55_io_in_0 = c53_371_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_55_io_in_1 = c32_19_io_out_1; // @[Multiplier.scala 128:41]
  assign c53_714_io_in_0 = c53_378_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_714_io_in_1 = c53_379_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_714_io_in_2 = c53_380_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_714_io_in_3 = c53_381_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_714_io_in_4 = c53_711_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_715_io_in_0 = c53_382_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_715_io_in_1 = c53_383_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_715_io_in_2 = c22_19_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_715_io_in_3 = c53_372_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_715_io_in_4 = c53_712_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_716_io_in_0 = c53_373_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_716_io_in_1 = c53_374_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_716_io_in_2 = c53_375_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_716_io_in_3 = c53_376_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_716_io_in_4 = c53_713_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_56_io_in_0 = c53_377_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_56_io_in_1 = c22_18_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_717_io_in_0 = c53_384_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_717_io_in_1 = c53_385_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_717_io_in_2 = c53_386_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_717_io_in_3 = c53_387_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_717_io_in_4 = c53_714_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_718_io_in_0 = c53_388_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_718_io_in_1 = c53_389_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_718_io_in_2 = r_1683; // @[Multiplier.scala 132:13]
  assign c53_718_io_in_3 = c53_378_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_718_io_in_4 = c53_715_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_719_io_in_0 = c53_379_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_719_io_in_1 = c53_380_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_719_io_in_2 = c53_381_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_719_io_in_3 = c53_382_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_719_io_in_4 = c53_716_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_57_io_in_0 = c53_383_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_57_io_in_1 = c22_19_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_720_io_in_0 = c53_390_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_720_io_in_1 = c53_391_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_720_io_in_2 = c53_392_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_720_io_in_3 = c53_393_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_720_io_in_4 = c53_717_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_721_io_in_0 = c53_394_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_721_io_in_1 = c53_395_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_721_io_in_2 = r_1708; // @[Multiplier.scala 132:13]
  assign c53_721_io_in_3 = c53_384_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_721_io_in_4 = c53_718_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_722_io_in_0 = c53_385_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_722_io_in_1 = c53_386_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_722_io_in_2 = c53_387_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_722_io_in_3 = c53_388_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_722_io_in_4 = c53_719_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_723_io_in_0 = c53_396_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_723_io_in_1 = c53_397_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_723_io_in_2 = c53_398_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_723_io_in_3 = c53_399_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_723_io_in_4 = c53_720_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_724_io_in_0 = c53_400_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_724_io_in_1 = c53_401_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_724_io_in_2 = c53_390_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_724_io_in_3 = c53_391_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_724_io_in_4 = c53_721_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_725_io_in_0 = c53_392_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_725_io_in_1 = c53_393_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_725_io_in_2 = c53_394_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_725_io_in_3 = c53_395_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_725_io_in_4 = c53_722_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_726_io_in_0 = c53_402_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_726_io_in_1 = c53_403_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_726_io_in_2 = c53_404_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_726_io_in_3 = c53_405_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_726_io_in_4 = c53_723_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_727_io_in_0 = c53_406_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_727_io_in_1 = c53_407_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_727_io_in_2 = c53_396_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_727_io_in_3 = c53_397_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_727_io_in_4 = c53_724_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_728_io_in_0 = c53_398_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_728_io_in_1 = c53_399_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_728_io_in_2 = c53_400_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_728_io_in_3 = c53_401_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_728_io_in_4 = c53_725_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_729_io_in_0 = c53_408_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_729_io_in_1 = c53_409_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_729_io_in_2 = c53_410_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_729_io_in_3 = c53_411_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_729_io_in_4 = c53_726_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_730_io_in_0 = c53_412_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_730_io_in_1 = c32_20_io_out_0; // @[Multiplier.scala 127:35]
  assign c53_730_io_in_2 = c53_407_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_730_io_in_3 = c53_402_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_730_io_in_4 = c53_727_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_731_io_in_0 = c53_403_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_731_io_in_1 = c53_404_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_731_io_in_2 = c53_405_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_731_io_in_3 = c53_406_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_731_io_in_4 = c53_728_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_732_io_in_0 = c53_413_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_732_io_in_1 = c53_414_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_732_io_in_2 = c53_415_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_732_io_in_3 = c53_416_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_732_io_in_4 = c53_729_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_733_io_in_0 = c53_417_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_733_io_in_1 = c32_21_io_out_0; // @[Multiplier.scala 127:35]
  assign c53_733_io_in_2 = c53_408_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_733_io_in_3 = c53_409_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_733_io_in_4 = c53_730_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_734_io_in_0 = c53_410_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_734_io_in_1 = c53_411_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_734_io_in_2 = c53_412_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_734_io_in_3 = c32_20_io_out_1; // @[Multiplier.scala 128:41]
  assign c53_734_io_in_4 = c53_731_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_735_io_in_0 = c53_418_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_735_io_in_1 = c53_419_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_735_io_in_2 = c53_420_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_735_io_in_3 = c53_421_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_735_io_in_4 = c53_732_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_736_io_in_0 = c53_422_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_736_io_in_1 = c22_20_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_736_io_in_2 = c53_413_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_736_io_in_3 = c53_414_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_736_io_in_4 = c53_733_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_737_io_in_0 = c53_415_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_737_io_in_1 = c53_416_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_737_io_in_2 = c53_417_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_737_io_in_3 = c32_21_io_out_1; // @[Multiplier.scala 128:41]
  assign c53_737_io_in_4 = c53_734_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_738_io_in_0 = c53_423_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_738_io_in_1 = c53_424_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_738_io_in_2 = c53_425_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_738_io_in_3 = c53_426_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_738_io_in_4 = c53_735_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_739_io_in_0 = c53_427_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_739_io_in_1 = c22_21_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_739_io_in_2 = c53_418_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_739_io_in_3 = c53_419_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_739_io_in_4 = c53_736_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_740_io_in_0 = c53_420_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_740_io_in_1 = c53_421_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_740_io_in_2 = c53_422_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_740_io_in_3 = c22_20_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_740_io_in_4 = c53_737_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_741_io_in_0 = c53_428_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_741_io_in_1 = c53_429_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_741_io_in_2 = c53_430_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_741_io_in_3 = c53_431_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_741_io_in_4 = c53_738_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_742_io_in_0 = c53_432_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_742_io_in_1 = r_1867; // @[Multiplier.scala 132:13]
  assign c53_742_io_in_2 = c53_423_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_742_io_in_3 = c53_424_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_742_io_in_4 = c53_739_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_743_io_in_0 = c53_425_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_743_io_in_1 = c53_426_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_743_io_in_2 = c53_427_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_743_io_in_3 = c22_21_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_743_io_in_4 = c53_740_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_744_io_in_0 = c53_433_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_744_io_in_1 = c53_434_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_744_io_in_2 = c53_435_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_744_io_in_3 = c53_436_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_744_io_in_4 = c53_741_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_745_io_in_0 = c53_437_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_745_io_in_1 = r_1888; // @[Multiplier.scala 132:13]
  assign c53_745_io_in_2 = c53_428_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_745_io_in_3 = c53_429_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_745_io_in_4 = c53_742_io_out_1; // @[Multiplier.scala 136:41]
  assign c32_46_io_in_0 = c53_430_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_46_io_in_1 = c53_431_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_46_io_in_2 = c53_432_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_746_io_in_0 = c53_438_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_746_io_in_1 = c53_439_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_746_io_in_2 = c53_440_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_746_io_in_3 = c53_441_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_746_io_in_4 = c53_744_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_747_io_in_0 = c53_442_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_747_io_in_1 = c53_433_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_747_io_in_2 = c53_434_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_747_io_in_3 = c53_435_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_747_io_in_4 = c53_745_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_58_io_in_0 = c53_436_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_58_io_in_1 = c53_437_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_748_io_in_0 = c53_443_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_748_io_in_1 = c53_444_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_748_io_in_2 = c53_445_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_748_io_in_3 = c53_446_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_748_io_in_4 = c53_746_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_749_io_in_0 = c53_447_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_749_io_in_1 = c53_438_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_749_io_in_2 = c53_439_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_749_io_in_3 = c53_440_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_749_io_in_4 = c53_747_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_59_io_in_0 = c53_441_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_59_io_in_1 = c53_442_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_750_io_in_0 = c53_448_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_750_io_in_1 = c53_449_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_750_io_in_2 = c53_450_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_750_io_in_3 = c53_451_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_750_io_in_4 = c53_748_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_751_io_in_0 = c32_22_io_out_0; // @[Multiplier.scala 127:35]
  assign c53_751_io_in_1 = c53_447_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_751_io_in_2 = c53_443_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_751_io_in_3 = c53_444_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_751_io_in_4 = c53_749_io_out_1; // @[Multiplier.scala 136:41]
  assign c32_47_io_in_0 = c53_445_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_47_io_in_1 = c53_446_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_47_io_in_2 = c53_447_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_752_io_in_0 = c53_452_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_752_io_in_1 = c53_453_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_752_io_in_2 = c53_454_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_752_io_in_3 = c53_455_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_752_io_in_4 = c53_750_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_753_io_in_0 = c32_23_io_out_0; // @[Multiplier.scala 127:35]
  assign c53_753_io_in_1 = c53_448_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_753_io_in_2 = c53_449_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_753_io_in_3 = c53_450_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_753_io_in_4 = c53_751_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_60_io_in_0 = c53_451_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_60_io_in_1 = c32_22_io_out_1; // @[Multiplier.scala 128:41]
  assign c53_754_io_in_0 = c53_456_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_754_io_in_1 = c53_457_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_754_io_in_2 = c53_458_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_754_io_in_3 = c53_459_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_754_io_in_4 = c53_752_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_755_io_in_0 = c22_22_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_755_io_in_1 = c53_452_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_755_io_in_2 = c53_453_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_755_io_in_3 = c53_454_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_755_io_in_4 = c53_753_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_61_io_in_0 = c53_455_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_61_io_in_1 = c32_23_io_out_1; // @[Multiplier.scala 128:41]
  assign c53_756_io_in_0 = c53_460_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_756_io_in_1 = c53_461_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_756_io_in_2 = c53_462_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_756_io_in_3 = c53_463_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_756_io_in_4 = c53_754_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_757_io_in_0 = c22_23_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_757_io_in_1 = c53_456_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_757_io_in_2 = c53_457_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_757_io_in_3 = c53_458_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_757_io_in_4 = c53_755_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_62_io_in_0 = c53_459_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_62_io_in_1 = c22_22_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_758_io_in_0 = c53_464_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_758_io_in_1 = c53_465_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_758_io_in_2 = c53_466_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_758_io_in_3 = c53_467_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_758_io_in_4 = c53_756_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_759_io_in_0 = r_2019; // @[Multiplier.scala 132:13]
  assign c53_759_io_in_1 = c53_460_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_759_io_in_2 = c53_461_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_759_io_in_3 = c53_462_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_759_io_in_4 = c53_757_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_63_io_in_0 = c53_463_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_63_io_in_1 = c22_23_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_760_io_in_0 = c53_468_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_760_io_in_1 = c53_469_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_760_io_in_2 = c53_470_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_760_io_in_3 = c53_471_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_760_io_in_4 = c53_758_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_761_io_in_0 = r_2036; // @[Multiplier.scala 132:13]
  assign c53_761_io_in_1 = c53_464_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_761_io_in_2 = c53_465_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_761_io_in_3 = c53_466_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_761_io_in_4 = c53_759_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_762_io_in_0 = c53_472_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_762_io_in_1 = c53_473_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_762_io_in_2 = c53_474_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_762_io_in_3 = c53_475_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_762_io_in_4 = c53_760_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_763_io_in_0 = c53_468_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_763_io_in_1 = c53_469_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_763_io_in_2 = c53_470_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_763_io_in_3 = c53_471_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_763_io_in_4 = c53_761_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_764_io_in_0 = c53_476_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_764_io_in_1 = c53_477_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_764_io_in_2 = c53_478_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_764_io_in_3 = c53_479_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_764_io_in_4 = c53_762_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_765_io_in_0 = c53_472_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_765_io_in_1 = c53_473_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_765_io_in_2 = c53_474_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_765_io_in_3 = c53_475_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_765_io_in_4 = c53_763_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_766_io_in_0 = c53_480_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_766_io_in_1 = c53_481_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_766_io_in_2 = c53_482_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_766_io_in_3 = c32_24_io_out_0; // @[Multiplier.scala 127:35]
  assign c53_766_io_in_4 = c53_764_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_767_io_in_0 = c53_479_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_767_io_in_1 = c53_476_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_767_io_in_2 = c53_477_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_767_io_in_3 = c53_478_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_767_io_in_4 = c53_765_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_768_io_in_0 = c53_483_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_768_io_in_1 = c53_484_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_768_io_in_2 = c53_485_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_768_io_in_3 = c32_25_io_out_0; // @[Multiplier.scala 127:35]
  assign c53_768_io_in_4 = c53_766_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_769_io_in_0 = c53_480_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_769_io_in_1 = c53_481_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_769_io_in_2 = c53_482_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_769_io_in_3 = c32_24_io_out_1; // @[Multiplier.scala 128:41]
  assign c53_769_io_in_4 = c53_767_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_770_io_in_0 = c53_486_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_770_io_in_1 = c53_487_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_770_io_in_2 = c53_488_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_770_io_in_3 = c22_24_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_770_io_in_4 = c53_768_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_771_io_in_0 = c53_483_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_771_io_in_1 = c53_484_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_771_io_in_2 = c53_485_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_771_io_in_3 = c32_25_io_out_1; // @[Multiplier.scala 128:41]
  assign c53_771_io_in_4 = c53_769_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_772_io_in_0 = c53_489_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_772_io_in_1 = c53_490_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_772_io_in_2 = c53_491_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_772_io_in_3 = c22_25_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_772_io_in_4 = c53_770_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_773_io_in_0 = c53_486_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_773_io_in_1 = c53_487_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_773_io_in_2 = c53_488_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_773_io_in_3 = c22_24_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_773_io_in_4 = c53_771_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_774_io_in_0 = c53_492_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_774_io_in_1 = c53_493_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_774_io_in_2 = c53_494_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_774_io_in_3 = r_2139; // @[Multiplier.scala 132:13]
  assign c53_774_io_in_4 = c53_772_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_775_io_in_0 = c53_489_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_775_io_in_1 = c53_490_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_775_io_in_2 = c53_491_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_775_io_in_3 = c22_25_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_775_io_in_4 = c53_773_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_776_io_in_0 = c53_495_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_776_io_in_1 = c53_496_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_776_io_in_2 = c53_497_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_776_io_in_3 = r_2152; // @[Multiplier.scala 132:13]
  assign c53_776_io_in_4 = c53_774_io_out_1; // @[Multiplier.scala 136:41]
  assign c32_48_io_in_0 = c53_492_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_48_io_in_1 = c53_493_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_48_io_in_2 = c53_494_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_777_io_in_0 = c53_498_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_777_io_in_1 = c53_499_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_777_io_in_2 = c53_500_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_777_io_in_3 = c53_495_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_777_io_in_4 = c53_776_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_64_io_in_0 = c53_496_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_64_io_in_1 = c53_497_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_778_io_in_0 = c53_501_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_778_io_in_1 = c53_502_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_778_io_in_2 = c53_503_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_778_io_in_3 = c53_498_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_778_io_in_4 = c53_777_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_65_io_in_0 = c53_499_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_65_io_in_1 = c53_500_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_779_io_in_0 = c53_504_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_779_io_in_1 = c53_505_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_779_io_in_2 = c32_26_io_out_0; // @[Multiplier.scala 127:35]
  assign c53_779_io_in_3 = c53_503_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_779_io_in_4 = c53_778_io_out_1; // @[Multiplier.scala 136:41]
  assign c32_49_io_in_0 = c53_501_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_49_io_in_1 = c53_502_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_49_io_in_2 = c53_503_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_780_io_in_0 = c53_506_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_780_io_in_1 = c53_507_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_780_io_in_2 = c32_27_io_out_0; // @[Multiplier.scala 127:35]
  assign c53_780_io_in_3 = c53_504_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_780_io_in_4 = c53_779_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_66_io_in_0 = c53_505_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_66_io_in_1 = c32_26_io_out_1; // @[Multiplier.scala 128:41]
  assign c53_781_io_in_0 = c53_508_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_781_io_in_1 = c53_509_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_781_io_in_2 = c22_26_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_781_io_in_3 = c53_506_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_781_io_in_4 = c53_780_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_67_io_in_0 = c53_507_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_67_io_in_1 = c32_27_io_out_1; // @[Multiplier.scala 128:41]
  assign c53_782_io_in_0 = c53_510_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_782_io_in_1 = c53_511_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_782_io_in_2 = c22_27_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_782_io_in_3 = c53_508_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_782_io_in_4 = c53_781_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_68_io_in_0 = c53_509_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_68_io_in_1 = c22_26_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_783_io_in_0 = c53_512_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_783_io_in_1 = c53_513_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_783_io_in_2 = r_2227; // @[Multiplier.scala 132:13]
  assign c53_783_io_in_3 = c53_510_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_783_io_in_4 = c53_782_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_69_io_in_0 = c53_511_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_69_io_in_1 = c22_27_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_784_io_in_0 = c53_514_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_784_io_in_1 = c53_515_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_784_io_in_2 = r_2236; // @[Multiplier.scala 132:13]
  assign c53_784_io_in_3 = c53_512_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_784_io_in_4 = c53_783_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_785_io_in_0 = c53_516_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_785_io_in_1 = c53_517_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_785_io_in_2 = c53_514_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_785_io_in_3 = c53_515_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_785_io_in_4 = c53_784_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_786_io_in_0 = c53_518_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_786_io_in_1 = c53_519_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_786_io_in_2 = c53_516_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_786_io_in_3 = c53_517_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_786_io_in_4 = c53_785_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_787_io_in_0 = c53_520_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_787_io_in_1 = c32_28_io_out_0; // @[Multiplier.scala 127:35]
  assign c53_787_io_in_2 = c53_519_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_787_io_in_3 = c53_518_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_787_io_in_4 = c53_786_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_788_io_in_0 = c53_521_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_788_io_in_1 = c32_29_io_out_0; // @[Multiplier.scala 127:35]
  assign c53_788_io_in_2 = c53_520_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_788_io_in_3 = c32_28_io_out_1; // @[Multiplier.scala 128:41]
  assign c53_788_io_in_4 = c53_787_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_789_io_in_0 = c53_522_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_789_io_in_1 = c22_28_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_789_io_in_2 = c53_521_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_789_io_in_3 = c32_29_io_out_1; // @[Multiplier.scala 128:41]
  assign c53_789_io_in_4 = c53_788_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_790_io_in_0 = c53_523_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_790_io_in_1 = c22_29_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_790_io_in_2 = c53_522_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_790_io_in_3 = c22_28_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_790_io_in_4 = c53_789_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_791_io_in_0 = c53_524_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_791_io_in_1 = r_2283; // @[Multiplier.scala 132:13]
  assign c53_791_io_in_2 = c53_523_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_791_io_in_3 = c22_29_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_791_io_in_4 = c53_790_io_out_1; // @[Multiplier.scala 136:41]
  assign c32_50_io_in_0 = c53_525_io_out_0; // @[Multiplier.scala 135:39]
  assign c32_50_io_in_1 = r_2288; // @[Multiplier.scala 126:19]
  assign c32_50_io_in_2 = c53_524_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_70_io_in_0 = c53_526_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_70_io_in_1 = c53_525_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_71_io_in_0 = c53_527_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_71_io_in_1 = c53_526_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_51_io_in_0 = c32_30_io_out_0; // @[Multiplier.scala 127:35]
  assign c32_51_io_in_1 = c53_527_io_out_1; // @[Multiplier.scala 136:41]
  assign c32_51_io_in_2 = c53_527_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_72_io_in_0 = c32_31_io_out_0; // @[Multiplier.scala 127:35]
  assign c22_72_io_in_1 = c32_30_io_out_1; // @[Multiplier.scala 128:41]
  assign c22_73_io_in_0 = c22_30_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_73_io_in_1 = c32_31_io_out_1; // @[Multiplier.scala 128:41]
  assign c22_74_io_in_0 = c22_31_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_74_io_in_1 = c22_30_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_75_io_in_0 = c22_33_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_75_io_in_1 = c22_32_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_76_io_in_0 = c22_34_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_76_io_in_1 = c22_33_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_77_io_in_0 = c22_35_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_77_io_in_1 = c22_34_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_78_io_in_0 = c22_36_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_78_io_in_1 = c22_35_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_79_io_in_0 = c32_32_io_out_0; // @[Multiplier.scala 127:35]
  assign c22_79_io_in_1 = c22_36_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_80_io_in_0 = c32_33_io_out_0; // @[Multiplier.scala 127:35]
  assign c22_80_io_in_1 = c32_32_io_out_1; // @[Multiplier.scala 128:41]
  assign c22_81_io_in_0 = c32_34_io_out_0; // @[Multiplier.scala 127:35]
  assign c22_81_io_in_1 = c32_33_io_out_1; // @[Multiplier.scala 128:41]
  assign c22_82_io_in_0 = c53_528_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_82_io_in_1 = c32_34_io_out_1; // @[Multiplier.scala 128:41]
  assign c22_83_io_in_0 = c53_529_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_83_io_in_1 = c53_528_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_84_io_in_0 = c53_530_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_84_io_in_1 = c53_529_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_85_io_in_0 = c53_531_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_85_io_in_1 = c53_530_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_86_io_in_0 = c53_532_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_86_io_in_1 = c53_531_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_52_io_in_0 = c53_533_io_out_0; // @[Multiplier.scala 135:39]
  assign c32_52_io_in_1 = c53_11_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_52_io_in_2 = c53_532_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_53_io_in_0 = c53_534_io_out_0; // @[Multiplier.scala 135:39]
  assign c32_53_io_in_1 = c53_13_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_53_io_in_2 = c53_533_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_54_io_in_0 = c53_535_io_out_0; // @[Multiplier.scala 135:39]
  assign c32_54_io_in_1 = c53_15_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_54_io_in_2 = c53_534_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_55_io_in_0 = c53_536_io_out_0; // @[Multiplier.scala 135:39]
  assign c32_55_io_in_1 = c22_37_io_out_0; // @[Multiplier.scala 122:35]
  assign c32_55_io_in_2 = c53_535_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_792_io_in_0 = c53_537_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_792_io_in_1 = c22_38_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_792_io_in_2 = c53_536_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_792_io_in_3 = c22_37_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_792_io_in_4 = 1'h0; // @[Multiplier.scala 134:24]
  assign c53_793_io_in_0 = c53_538_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_793_io_in_1 = c22_39_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_793_io_in_2 = c53_537_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_793_io_in_3 = c22_38_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_793_io_in_4 = c53_792_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_794_io_in_0 = c53_539_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_794_io_in_1 = c22_40_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_794_io_in_2 = c53_538_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_794_io_in_3 = c22_39_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_794_io_in_4 = c53_793_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_795_io_in_0 = c53_540_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_795_io_in_1 = c22_41_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_795_io_in_2 = c53_539_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_795_io_in_3 = c22_40_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_795_io_in_4 = c53_794_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_796_io_in_0 = c53_541_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_796_io_in_1 = c32_35_io_out_0; // @[Multiplier.scala 127:35]
  assign c53_796_io_in_2 = c53_540_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_796_io_in_3 = c22_41_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_796_io_in_4 = c53_795_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_797_io_in_0 = c53_542_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_797_io_in_1 = c32_36_io_out_0; // @[Multiplier.scala 127:35]
  assign c53_797_io_in_2 = c53_541_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_797_io_in_3 = c32_35_io_out_1; // @[Multiplier.scala 128:41]
  assign c53_797_io_in_4 = c53_796_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_798_io_in_0 = c53_543_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_798_io_in_1 = c32_37_io_out_0; // @[Multiplier.scala 127:35]
  assign c53_798_io_in_2 = c53_542_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_798_io_in_3 = c32_36_io_out_1; // @[Multiplier.scala 128:41]
  assign c53_798_io_in_4 = c53_797_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_799_io_in_0 = c53_544_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_799_io_in_1 = c53_545_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_799_io_in_2 = c53_543_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_799_io_in_3 = c32_37_io_out_1; // @[Multiplier.scala 128:41]
  assign c53_799_io_in_4 = c53_798_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_800_io_in_0 = c53_546_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_800_io_in_1 = c53_547_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_800_io_in_2 = c53_544_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_800_io_in_3 = c53_545_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_800_io_in_4 = c53_799_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_801_io_in_0 = c53_548_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_801_io_in_1 = c53_549_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_801_io_in_2 = c53_546_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_801_io_in_3 = c53_547_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_801_io_in_4 = c53_800_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_802_io_in_0 = c53_550_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_802_io_in_1 = c53_551_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_802_io_in_2 = c53_548_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_802_io_in_3 = c53_549_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_802_io_in_4 = c53_801_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_803_io_in_0 = c53_552_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_803_io_in_1 = c53_553_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_803_io_in_2 = c53_550_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_803_io_in_3 = c53_551_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_803_io_in_4 = c53_802_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_804_io_in_0 = c53_554_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_804_io_in_1 = c53_555_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_804_io_in_2 = c53_55_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_804_io_in_3 = c53_552_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_804_io_in_4 = c53_803_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_805_io_in_0 = c53_556_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_805_io_in_1 = c53_557_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_805_io_in_2 = c53_59_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_805_io_in_3 = c53_554_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_805_io_in_4 = c53_804_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_806_io_in_0 = c53_558_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_806_io_in_1 = c53_559_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_806_io_in_2 = c53_63_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_806_io_in_3 = c53_556_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_806_io_in_4 = c53_805_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_807_io_in_0 = c53_560_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_807_io_in_1 = c53_561_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_807_io_in_2 = c22_42_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_807_io_in_3 = c53_558_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_807_io_in_4 = c53_806_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_808_io_in_0 = c53_562_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_808_io_in_1 = c53_563_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_808_io_in_2 = c22_43_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_808_io_in_3 = c53_560_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_808_io_in_4 = c53_807_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_87_io_in_0 = c53_561_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_87_io_in_1 = c22_42_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_809_io_in_0 = c53_564_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_809_io_in_1 = c53_565_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_809_io_in_2 = c22_44_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_809_io_in_3 = c53_562_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_809_io_in_4 = c53_808_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_88_io_in_0 = c53_563_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_88_io_in_1 = c22_43_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_810_io_in_0 = c53_566_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_810_io_in_1 = c53_567_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_810_io_in_2 = c22_45_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_810_io_in_3 = c53_564_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_810_io_in_4 = c53_809_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_89_io_in_0 = c53_565_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_89_io_in_1 = c22_44_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_811_io_in_0 = c53_568_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_811_io_in_1 = c53_569_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_811_io_in_2 = c22_46_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_811_io_in_3 = c53_566_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_811_io_in_4 = c53_810_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_90_io_in_0 = c53_567_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_90_io_in_1 = c22_45_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_812_io_in_0 = c53_570_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_812_io_in_1 = c53_571_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_812_io_in_2 = c32_38_io_out_0; // @[Multiplier.scala 127:35]
  assign c53_812_io_in_3 = c53_568_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_812_io_in_4 = c53_811_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_91_io_in_0 = c53_569_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_91_io_in_1 = c22_46_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_813_io_in_0 = c53_572_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_813_io_in_1 = c53_573_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_813_io_in_2 = c32_39_io_out_0; // @[Multiplier.scala 127:35]
  assign c53_813_io_in_3 = c53_570_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_813_io_in_4 = c53_812_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_92_io_in_0 = c53_571_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_92_io_in_1 = c32_38_io_out_1; // @[Multiplier.scala 128:41]
  assign c53_814_io_in_0 = c53_574_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_814_io_in_1 = c53_575_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_814_io_in_2 = c32_40_io_out_0; // @[Multiplier.scala 127:35]
  assign c53_814_io_in_3 = c53_572_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_814_io_in_4 = c53_813_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_93_io_in_0 = c53_573_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_93_io_in_1 = c32_39_io_out_1; // @[Multiplier.scala 128:41]
  assign c53_815_io_in_0 = c53_576_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_815_io_in_1 = c53_577_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_815_io_in_2 = c53_578_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_815_io_in_3 = c53_574_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_815_io_in_4 = c53_814_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_94_io_in_0 = c53_575_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_94_io_in_1 = c32_40_io_out_1; // @[Multiplier.scala 128:41]
  assign c53_816_io_in_0 = c53_579_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_816_io_in_1 = c53_580_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_816_io_in_2 = c53_581_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_816_io_in_3 = c53_576_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_816_io_in_4 = c53_815_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_95_io_in_0 = c53_577_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_95_io_in_1 = c53_578_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_817_io_in_0 = c53_582_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_817_io_in_1 = c53_583_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_817_io_in_2 = c53_584_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_817_io_in_3 = c53_579_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_817_io_in_4 = c53_816_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_96_io_in_0 = c53_580_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_96_io_in_1 = c53_581_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_818_io_in_0 = c53_585_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_818_io_in_1 = c53_586_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_818_io_in_2 = c53_587_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_818_io_in_3 = c53_582_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_818_io_in_4 = c53_817_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_97_io_in_0 = c53_583_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_97_io_in_1 = c53_584_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_819_io_in_0 = c53_588_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_819_io_in_1 = c53_589_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_819_io_in_2 = c53_590_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_819_io_in_3 = c53_585_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_819_io_in_4 = c53_818_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_98_io_in_0 = c53_586_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_98_io_in_1 = c53_587_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_820_io_in_0 = c53_591_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_820_io_in_1 = c53_592_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_820_io_in_2 = c53_593_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_820_io_in_3 = c53_131_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_820_io_in_4 = c53_819_io_out_1; // @[Multiplier.scala 136:41]
  assign c32_56_io_in_0 = c53_588_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_56_io_in_1 = c53_589_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_56_io_in_2 = c53_590_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_821_io_in_0 = c53_594_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_821_io_in_1 = c53_595_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_821_io_in_2 = c53_596_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_821_io_in_3 = c53_137_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_821_io_in_4 = c53_820_io_out_1; // @[Multiplier.scala 136:41]
  assign c32_57_io_in_0 = c53_591_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_57_io_in_1 = c53_592_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_57_io_in_2 = c53_593_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_822_io_in_0 = c53_597_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_822_io_in_1 = c53_598_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_822_io_in_2 = c53_599_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_822_io_in_3 = c53_143_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_822_io_in_4 = c53_821_io_out_1; // @[Multiplier.scala 136:41]
  assign c32_58_io_in_0 = c53_594_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_58_io_in_1 = c53_595_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_58_io_in_2 = c53_596_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_823_io_in_0 = c53_600_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_823_io_in_1 = c53_601_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_823_io_in_2 = c53_602_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_823_io_in_3 = c22_47_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_823_io_in_4 = c53_822_io_out_1; // @[Multiplier.scala 136:41]
  assign c32_59_io_in_0 = c53_597_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_59_io_in_1 = c53_598_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_59_io_in_2 = c53_599_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_824_io_in_0 = c53_603_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_824_io_in_1 = c53_604_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_824_io_in_2 = c53_605_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_824_io_in_3 = c22_48_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_824_io_in_4 = c53_823_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_825_io_in_0 = c53_600_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_825_io_in_1 = c53_601_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_825_io_in_2 = c53_602_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_825_io_in_3 = c22_47_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_825_io_in_4 = 1'h0; // @[Multiplier.scala 134:24]
  assign c53_826_io_in_0 = c53_606_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_826_io_in_1 = c53_607_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_826_io_in_2 = c53_608_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_826_io_in_3 = c22_49_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_826_io_in_4 = c53_824_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_827_io_in_0 = c53_603_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_827_io_in_1 = c53_604_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_827_io_in_2 = c53_605_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_827_io_in_3 = c22_48_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_827_io_in_4 = c53_825_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_828_io_in_0 = c53_609_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_828_io_in_1 = c53_610_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_828_io_in_2 = c53_611_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_828_io_in_3 = c22_50_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_828_io_in_4 = c53_826_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_829_io_in_0 = c53_606_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_829_io_in_1 = c53_607_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_829_io_in_2 = c53_608_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_829_io_in_3 = c22_49_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_829_io_in_4 = c53_827_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_830_io_in_0 = c53_612_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_830_io_in_1 = c53_613_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_830_io_in_2 = c53_614_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_830_io_in_3 = c22_51_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_830_io_in_4 = c53_828_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_831_io_in_0 = c53_609_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_831_io_in_1 = c53_610_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_831_io_in_2 = c53_611_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_831_io_in_3 = c22_50_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_831_io_in_4 = c53_829_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_832_io_in_0 = c53_615_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_832_io_in_1 = c53_616_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_832_io_in_2 = c53_617_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_832_io_in_3 = c32_41_io_out_0; // @[Multiplier.scala 127:35]
  assign c53_832_io_in_4 = c53_830_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_833_io_in_0 = c53_612_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_833_io_in_1 = c53_613_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_833_io_in_2 = c53_614_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_833_io_in_3 = c22_51_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_833_io_in_4 = c53_831_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_834_io_in_0 = c53_618_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_834_io_in_1 = c53_619_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_834_io_in_2 = c53_620_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_834_io_in_3 = c32_42_io_out_0; // @[Multiplier.scala 127:35]
  assign c53_834_io_in_4 = c53_832_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_835_io_in_0 = c53_615_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_835_io_in_1 = c53_616_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_835_io_in_2 = c53_617_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_835_io_in_3 = c32_41_io_out_1; // @[Multiplier.scala 128:41]
  assign c53_835_io_in_4 = c53_833_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_836_io_in_0 = c53_621_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_836_io_in_1 = c53_622_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_836_io_in_2 = c53_623_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_836_io_in_3 = c32_43_io_out_0; // @[Multiplier.scala 127:35]
  assign c53_836_io_in_4 = c53_834_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_837_io_in_0 = c53_618_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_837_io_in_1 = c53_619_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_837_io_in_2 = c53_620_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_837_io_in_3 = c32_42_io_out_1; // @[Multiplier.scala 128:41]
  assign c53_837_io_in_4 = c53_835_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_838_io_in_0 = c53_624_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_838_io_in_1 = c53_625_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_838_io_in_2 = c53_626_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_838_io_in_3 = c53_627_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_838_io_in_4 = c53_836_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_839_io_in_0 = c53_621_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_839_io_in_1 = c53_622_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_839_io_in_2 = c53_623_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_839_io_in_3 = c32_43_io_out_1; // @[Multiplier.scala 128:41]
  assign c53_839_io_in_4 = c53_837_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_840_io_in_0 = c53_628_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_840_io_in_1 = c53_629_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_840_io_in_2 = c53_630_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_840_io_in_3 = c53_631_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_840_io_in_4 = c53_838_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_841_io_in_0 = c53_624_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_841_io_in_1 = c53_625_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_841_io_in_2 = c53_626_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_841_io_in_3 = c53_627_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_841_io_in_4 = c53_839_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_842_io_in_0 = c53_632_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_842_io_in_1 = c53_633_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_842_io_in_2 = c53_634_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_842_io_in_3 = c53_635_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_842_io_in_4 = c53_840_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_843_io_in_0 = c53_628_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_843_io_in_1 = c53_629_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_843_io_in_2 = c53_630_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_843_io_in_3 = c53_631_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_843_io_in_4 = c53_841_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_844_io_in_0 = c53_636_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_844_io_in_1 = c53_637_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_844_io_in_2 = c53_638_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_844_io_in_3 = c53_639_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_844_io_in_4 = c53_842_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_845_io_in_0 = c53_632_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_845_io_in_1 = c53_633_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_845_io_in_2 = c53_634_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_845_io_in_3 = c53_635_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_845_io_in_4 = c53_843_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_846_io_in_0 = c53_640_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_846_io_in_1 = c53_641_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_846_io_in_2 = c53_642_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_846_io_in_3 = c53_643_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_846_io_in_4 = c53_844_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_847_io_in_0 = c53_636_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_847_io_in_1 = c53_637_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_847_io_in_2 = c53_638_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_847_io_in_3 = c53_639_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_847_io_in_4 = c53_845_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_848_io_in_0 = c53_644_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_848_io_in_1 = c53_645_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_848_io_in_2 = c53_646_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_848_io_in_3 = c53_647_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_848_io_in_4 = c53_846_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_849_io_in_0 = c53_239_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_849_io_in_1 = c53_640_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_849_io_in_2 = c53_641_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_849_io_in_3 = c53_642_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_849_io_in_4 = c53_847_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_850_io_in_0 = c53_648_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_850_io_in_1 = c53_649_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_850_io_in_2 = c53_650_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_850_io_in_3 = c53_651_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_850_io_in_4 = c53_848_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_851_io_in_0 = c53_247_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_851_io_in_1 = c53_644_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_851_io_in_2 = c53_645_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_851_io_in_3 = c53_646_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_851_io_in_4 = c53_849_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_852_io_in_0 = c53_652_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_852_io_in_1 = c53_653_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_852_io_in_2 = c53_654_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_852_io_in_3 = c53_655_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_852_io_in_4 = c53_850_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_853_io_in_0 = c53_255_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_853_io_in_1 = c53_648_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_853_io_in_2 = c53_649_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_853_io_in_3 = c53_650_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_853_io_in_4 = c53_851_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_854_io_in_0 = c53_656_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_854_io_in_1 = c53_657_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_854_io_in_2 = c53_658_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_854_io_in_3 = c53_659_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_854_io_in_4 = c53_852_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_855_io_in_0 = c53_263_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_855_io_in_1 = c53_652_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_855_io_in_2 = c53_653_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_855_io_in_3 = c53_654_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_855_io_in_4 = c53_853_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_856_io_in_0 = c53_660_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_856_io_in_1 = c53_661_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_856_io_in_2 = c53_662_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_856_io_in_3 = c53_663_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_856_io_in_4 = c53_854_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_857_io_in_0 = c53_271_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_857_io_in_1 = c53_656_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_857_io_in_2 = c53_657_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_857_io_in_3 = c53_658_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_857_io_in_4 = c53_855_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_858_io_in_0 = c53_664_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_858_io_in_1 = c53_665_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_858_io_in_2 = c53_666_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_858_io_in_3 = c53_667_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_858_io_in_4 = c53_856_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_859_io_in_0 = c53_279_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_859_io_in_1 = c53_660_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_859_io_in_2 = c53_661_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_859_io_in_3 = c53_662_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_859_io_in_4 = c53_857_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_860_io_in_0 = c53_668_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_860_io_in_1 = c53_669_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_860_io_in_2 = c53_670_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_860_io_in_3 = c53_671_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_860_io_in_4 = c53_858_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_861_io_in_0 = c53_287_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_861_io_in_1 = c53_664_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_861_io_in_2 = c53_665_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_861_io_in_3 = c53_666_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_861_io_in_4 = c53_859_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_862_io_in_0 = c53_672_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_862_io_in_1 = c53_673_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_862_io_in_2 = c53_674_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_862_io_in_3 = c53_675_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_862_io_in_4 = c53_860_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_863_io_in_0 = c53_668_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_863_io_in_1 = c53_669_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_863_io_in_2 = c53_670_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_863_io_in_3 = c53_671_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_863_io_in_4 = c53_861_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_864_io_in_0 = c53_676_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_864_io_in_1 = c53_677_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_864_io_in_2 = c53_678_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_864_io_in_3 = c53_679_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_864_io_in_4 = c53_862_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_865_io_in_0 = c53_303_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_865_io_in_1 = c53_672_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_865_io_in_2 = c53_673_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_865_io_in_3 = c53_674_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_865_io_in_4 = c53_863_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_866_io_in_0 = c53_680_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_866_io_in_1 = c53_681_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_866_io_in_2 = c53_682_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_866_io_in_3 = c53_683_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_866_io_in_4 = c53_864_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_867_io_in_0 = c53_676_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_867_io_in_1 = c53_677_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_867_io_in_2 = c53_678_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_867_io_in_3 = c53_679_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_867_io_in_4 = c53_865_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_868_io_in_0 = c53_684_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_868_io_in_1 = c53_685_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_868_io_in_2 = c53_686_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_868_io_in_3 = c53_687_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_868_io_in_4 = c53_866_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_869_io_in_0 = c53_680_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_869_io_in_1 = c53_681_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_869_io_in_2 = c53_682_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_869_io_in_3 = c53_683_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_869_io_in_4 = c53_867_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_870_io_in_0 = c53_688_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_870_io_in_1 = c53_689_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_870_io_in_2 = c53_690_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_870_io_in_3 = c53_691_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_870_io_in_4 = c53_868_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_871_io_in_0 = c53_684_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_871_io_in_1 = c53_685_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_871_io_in_2 = c53_686_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_871_io_in_3 = c53_687_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_871_io_in_4 = c53_869_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_872_io_in_0 = c53_692_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_872_io_in_1 = c53_693_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_872_io_in_2 = c53_694_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_872_io_in_3 = c53_695_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_872_io_in_4 = c53_870_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_873_io_in_0 = c53_688_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_873_io_in_1 = c53_689_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_873_io_in_2 = c53_690_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_873_io_in_3 = c53_691_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_873_io_in_4 = c53_871_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_874_io_in_0 = c53_696_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_874_io_in_1 = c53_697_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_874_io_in_2 = c53_698_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_874_io_in_3 = c32_44_io_out_0; // @[Multiplier.scala 127:35]
  assign c53_874_io_in_4 = c53_872_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_875_io_in_0 = c53_695_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_875_io_in_1 = c53_692_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_875_io_in_2 = c53_693_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_875_io_in_3 = c53_694_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_875_io_in_4 = c53_873_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_876_io_in_0 = c53_699_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_876_io_in_1 = c53_700_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_876_io_in_2 = c53_701_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_876_io_in_3 = c22_52_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_876_io_in_4 = c53_874_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_877_io_in_0 = c53_696_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_877_io_in_1 = c53_697_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_877_io_in_2 = c53_698_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_877_io_in_3 = c32_44_io_out_1; // @[Multiplier.scala 128:41]
  assign c53_877_io_in_4 = c53_875_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_878_io_in_0 = c53_702_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_878_io_in_1 = c53_703_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_878_io_in_2 = c53_704_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_878_io_in_3 = c22_53_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_878_io_in_4 = c53_876_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_879_io_in_0 = c53_699_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_879_io_in_1 = c53_700_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_879_io_in_2 = c53_701_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_879_io_in_3 = c22_52_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_879_io_in_4 = c53_877_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_880_io_in_0 = c53_705_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_880_io_in_1 = c53_706_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_880_io_in_2 = c53_707_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_880_io_in_3 = c32_45_io_out_0; // @[Multiplier.scala 127:35]
  assign c53_880_io_in_4 = c53_878_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_881_io_in_0 = c53_702_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_881_io_in_1 = c53_703_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_881_io_in_2 = c53_704_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_881_io_in_3 = c22_53_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_881_io_in_4 = c53_879_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_882_io_in_0 = c53_708_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_882_io_in_1 = c53_709_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_882_io_in_2 = c53_710_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_882_io_in_3 = c22_54_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_882_io_in_4 = c53_880_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_883_io_in_0 = c53_705_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_883_io_in_1 = c53_706_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_883_io_in_2 = c53_707_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_883_io_in_3 = c32_45_io_out_1; // @[Multiplier.scala 128:41]
  assign c53_883_io_in_4 = c53_881_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_884_io_in_0 = c53_711_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_884_io_in_1 = c53_712_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_884_io_in_2 = c53_713_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_884_io_in_3 = c22_55_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_884_io_in_4 = c53_882_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_885_io_in_0 = c53_708_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_885_io_in_1 = c53_709_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_885_io_in_2 = c53_710_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_885_io_in_3 = c22_54_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_885_io_in_4 = c53_883_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_886_io_in_0 = c53_714_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_886_io_in_1 = c53_715_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_886_io_in_2 = c53_716_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_886_io_in_3 = c22_56_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_886_io_in_4 = c53_884_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_887_io_in_0 = c53_711_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_887_io_in_1 = c53_712_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_887_io_in_2 = c53_713_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_887_io_in_3 = c22_55_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_887_io_in_4 = c53_885_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_888_io_in_0 = c53_717_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_888_io_in_1 = c53_718_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_888_io_in_2 = c53_719_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_888_io_in_3 = c22_57_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_888_io_in_4 = c53_886_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_889_io_in_0 = c53_714_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_889_io_in_1 = c53_715_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_889_io_in_2 = c53_716_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_889_io_in_3 = c22_56_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_889_io_in_4 = c53_887_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_890_io_in_0 = c53_720_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_890_io_in_1 = c53_721_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_890_io_in_2 = c53_722_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_890_io_in_3 = c53_389_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_890_io_in_4 = c53_888_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_891_io_in_0 = c53_717_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_891_io_in_1 = c53_718_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_891_io_in_2 = c53_719_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_891_io_in_3 = c22_57_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_891_io_in_4 = c53_889_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_892_io_in_0 = c53_723_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_892_io_in_1 = c53_724_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_892_io_in_2 = c53_725_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_892_io_in_3 = c53_720_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_892_io_in_4 = c53_890_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_99_io_in_0 = c53_721_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_99_io_in_1 = c53_722_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_893_io_in_0 = c53_726_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_893_io_in_1 = c53_727_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_893_io_in_2 = c53_728_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_893_io_in_3 = c53_723_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_893_io_in_4 = c53_892_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_100_io_in_0 = c53_724_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_100_io_in_1 = c53_725_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_894_io_in_0 = c53_729_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_894_io_in_1 = c53_730_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_894_io_in_2 = c53_731_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_894_io_in_3 = c53_407_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_894_io_in_4 = c53_893_io_out_1; // @[Multiplier.scala 136:41]
  assign c32_60_io_in_0 = c53_726_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_60_io_in_1 = c53_727_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_60_io_in_2 = c53_728_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_895_io_in_0 = c53_732_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_895_io_in_1 = c53_733_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_895_io_in_2 = c53_734_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_895_io_in_3 = c53_729_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_895_io_in_4 = c53_894_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_101_io_in_0 = c53_730_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_101_io_in_1 = c53_731_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_896_io_in_0 = c53_735_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_896_io_in_1 = c53_736_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_896_io_in_2 = c53_737_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_896_io_in_3 = c53_732_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_896_io_in_4 = c53_895_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_102_io_in_0 = c53_733_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_102_io_in_1 = c53_734_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_897_io_in_0 = c53_738_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_897_io_in_1 = c53_739_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_897_io_in_2 = c53_740_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_897_io_in_3 = c53_735_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_897_io_in_4 = c53_896_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_103_io_in_0 = c53_736_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_103_io_in_1 = c53_737_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_898_io_in_0 = c53_741_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_898_io_in_1 = c53_742_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_898_io_in_2 = c53_743_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_898_io_in_3 = c53_738_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_898_io_in_4 = c53_897_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_104_io_in_0 = c53_739_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_104_io_in_1 = c53_740_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_899_io_in_0 = c53_744_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_899_io_in_1 = c53_745_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_899_io_in_2 = c32_46_io_out_0; // @[Multiplier.scala 127:35]
  assign c53_899_io_in_3 = c53_743_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_899_io_in_4 = c53_898_io_out_1; // @[Multiplier.scala 136:41]
  assign c32_61_io_in_0 = c53_741_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_61_io_in_1 = c53_742_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_61_io_in_2 = c53_743_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_900_io_in_0 = c53_746_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_900_io_in_1 = c53_747_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_900_io_in_2 = c22_58_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_900_io_in_3 = c53_744_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_900_io_in_4 = c53_899_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_105_io_in_0 = c53_745_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_105_io_in_1 = c32_46_io_out_1; // @[Multiplier.scala 128:41]
  assign c53_901_io_in_0 = c53_748_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_901_io_in_1 = c53_749_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_901_io_in_2 = c22_59_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_901_io_in_3 = c53_746_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_901_io_in_4 = c53_900_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_106_io_in_0 = c53_747_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_106_io_in_1 = c22_58_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_902_io_in_0 = c53_750_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_902_io_in_1 = c53_751_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_902_io_in_2 = c32_47_io_out_0; // @[Multiplier.scala 127:35]
  assign c53_902_io_in_3 = c53_748_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_902_io_in_4 = c53_901_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_107_io_in_0 = c53_749_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_107_io_in_1 = c22_59_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_903_io_in_0 = c53_752_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_903_io_in_1 = c53_753_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_903_io_in_2 = c22_60_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_903_io_in_3 = c53_750_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_903_io_in_4 = c53_902_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_108_io_in_0 = c53_751_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_108_io_in_1 = c32_47_io_out_1; // @[Multiplier.scala 128:41]
  assign c53_904_io_in_0 = c53_754_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_904_io_in_1 = c53_755_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_904_io_in_2 = c22_61_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_904_io_in_3 = c53_752_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_904_io_in_4 = c53_903_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_109_io_in_0 = c53_753_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_109_io_in_1 = c22_60_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_905_io_in_0 = c53_756_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_905_io_in_1 = c53_757_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_905_io_in_2 = c22_62_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_905_io_in_3 = c53_754_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_905_io_in_4 = c53_904_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_110_io_in_0 = c53_755_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_110_io_in_1 = c22_61_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_906_io_in_0 = c53_758_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_906_io_in_1 = c53_759_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_906_io_in_2 = c22_63_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_906_io_in_3 = c53_756_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_906_io_in_4 = c53_905_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_111_io_in_0 = c53_757_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_111_io_in_1 = c22_62_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_907_io_in_0 = c53_760_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_907_io_in_1 = c53_761_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_907_io_in_2 = c53_467_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_907_io_in_3 = c53_758_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_907_io_in_4 = c53_906_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_112_io_in_0 = c53_759_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_112_io_in_1 = c22_63_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_908_io_in_0 = c53_762_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_908_io_in_1 = c53_763_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_908_io_in_2 = c53_760_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_908_io_in_3 = c53_761_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_908_io_in_4 = c53_907_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_909_io_in_0 = c53_764_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_909_io_in_1 = c53_765_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_909_io_in_2 = c53_762_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_909_io_in_3 = c53_763_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_909_io_in_4 = c53_908_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_910_io_in_0 = c53_766_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_910_io_in_1 = c53_767_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_910_io_in_2 = c53_479_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_910_io_in_3 = c53_764_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_910_io_in_4 = c53_909_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_911_io_in_0 = c53_768_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_911_io_in_1 = c53_769_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_911_io_in_2 = c53_766_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_911_io_in_3 = c53_767_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_911_io_in_4 = c53_910_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_912_io_in_0 = c53_770_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_912_io_in_1 = c53_771_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_912_io_in_2 = c53_768_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_912_io_in_3 = c53_769_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_912_io_in_4 = c53_911_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_913_io_in_0 = c53_772_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_913_io_in_1 = c53_773_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_913_io_in_2 = c53_770_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_913_io_in_3 = c53_771_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_913_io_in_4 = c53_912_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_914_io_in_0 = c53_774_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_914_io_in_1 = c53_775_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_914_io_in_2 = c53_772_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_914_io_in_3 = c53_773_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_914_io_in_4 = c53_913_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_915_io_in_0 = c53_776_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_915_io_in_1 = c32_48_io_out_0; // @[Multiplier.scala 127:35]
  assign c53_915_io_in_2 = c53_775_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_915_io_in_3 = c53_774_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_915_io_in_4 = c53_914_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_916_io_in_0 = c53_777_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_916_io_in_1 = c22_64_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_916_io_in_2 = c53_776_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_916_io_in_3 = c32_48_io_out_1; // @[Multiplier.scala 128:41]
  assign c53_916_io_in_4 = c53_915_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_917_io_in_0 = c53_778_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_917_io_in_1 = c22_65_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_917_io_in_2 = c53_777_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_917_io_in_3 = c22_64_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_917_io_in_4 = c53_916_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_918_io_in_0 = c53_779_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_918_io_in_1 = c32_49_io_out_0; // @[Multiplier.scala 127:35]
  assign c53_918_io_in_2 = c53_778_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_918_io_in_3 = c22_65_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_918_io_in_4 = c53_917_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_919_io_in_0 = c53_780_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_919_io_in_1 = c22_66_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_919_io_in_2 = c53_779_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_919_io_in_3 = c32_49_io_out_1; // @[Multiplier.scala 128:41]
  assign c53_919_io_in_4 = c53_918_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_920_io_in_0 = c53_781_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_920_io_in_1 = c22_67_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_920_io_in_2 = c53_780_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_920_io_in_3 = c22_66_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_920_io_in_4 = c53_919_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_921_io_in_0 = c53_782_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_921_io_in_1 = c22_68_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_921_io_in_2 = c53_781_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_921_io_in_3 = c22_67_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_921_io_in_4 = c53_920_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_922_io_in_0 = c53_783_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_922_io_in_1 = c22_69_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_922_io_in_2 = c53_782_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_922_io_in_3 = c22_68_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_922_io_in_4 = c53_921_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_923_io_in_0 = c53_784_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_923_io_in_1 = c53_513_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_923_io_in_2 = c53_783_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_923_io_in_3 = c22_69_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_923_io_in_4 = c53_922_io_out_1; // @[Multiplier.scala 136:41]
  assign c22_113_io_in_0 = c53_785_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_113_io_in_1 = c53_784_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_114_io_in_0 = c53_786_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_114_io_in_1 = c53_785_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_62_io_in_0 = c53_787_io_out_0; // @[Multiplier.scala 135:39]
  assign c32_62_io_in_1 = c53_519_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_62_io_in_2 = c53_786_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_115_io_in_0 = c53_788_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_115_io_in_1 = c53_787_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_116_io_in_0 = c53_789_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_116_io_in_1 = c53_788_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_117_io_in_0 = c53_790_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_117_io_in_1 = c53_789_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_118_io_in_0 = c53_791_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_118_io_in_1 = c53_790_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_63_io_in_0 = c32_50_io_out_0; // @[Multiplier.scala 127:35]
  assign c32_63_io_in_1 = c53_791_io_out_1; // @[Multiplier.scala 136:41]
  assign c32_63_io_in_2 = c53_791_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_119_io_in_0 = c22_70_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_119_io_in_1 = c32_50_io_out_1; // @[Multiplier.scala 128:41]
  assign c22_120_io_in_0 = c22_71_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_120_io_in_1 = c22_70_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_121_io_in_0 = c32_51_io_out_0; // @[Multiplier.scala 127:35]
  assign c22_121_io_in_1 = c22_71_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_122_io_in_0 = c22_72_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_122_io_in_1 = c32_51_io_out_1; // @[Multiplier.scala 128:41]
  assign c22_123_io_in_0 = c22_73_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_123_io_in_1 = c22_72_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_124_io_in_0 = c22_74_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_124_io_in_1 = c22_73_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_125_io_in_0 = c22_76_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_125_io_in_1 = c22_75_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_126_io_in_0 = c22_77_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_126_io_in_1 = c22_76_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_127_io_in_0 = c22_78_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_127_io_in_1 = c22_77_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_128_io_in_0 = c22_79_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_128_io_in_1 = c22_78_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_129_io_in_0 = c22_80_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_129_io_in_1 = c22_79_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_130_io_in_0 = c22_81_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_130_io_in_1 = c22_80_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_131_io_in_0 = c22_82_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_131_io_in_1 = c22_81_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_132_io_in_0 = c22_83_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_132_io_in_1 = c22_82_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_133_io_in_0 = c22_84_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_133_io_in_1 = c22_83_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_134_io_in_0 = c22_85_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_134_io_in_1 = c22_84_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_135_io_in_0 = c22_86_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_135_io_in_1 = c22_85_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_136_io_in_0 = c32_52_io_out_0; // @[Multiplier.scala 127:35]
  assign c22_136_io_in_1 = c22_86_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_137_io_in_0 = c32_53_io_out_0; // @[Multiplier.scala 127:35]
  assign c22_137_io_in_1 = c32_52_io_out_1; // @[Multiplier.scala 128:41]
  assign c22_138_io_in_0 = c32_54_io_out_0; // @[Multiplier.scala 127:35]
  assign c22_138_io_in_1 = c32_53_io_out_1; // @[Multiplier.scala 128:41]
  assign c22_139_io_in_0 = c32_55_io_out_0; // @[Multiplier.scala 127:35]
  assign c22_139_io_in_1 = c32_54_io_out_1; // @[Multiplier.scala 128:41]
  assign c22_140_io_in_0 = c53_792_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_140_io_in_1 = c32_55_io_out_1; // @[Multiplier.scala 128:41]
  assign c22_141_io_in_0 = c53_793_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_141_io_in_1 = c53_792_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_142_io_in_0 = c53_794_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_142_io_in_1 = c53_793_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_143_io_in_0 = c53_795_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_143_io_in_1 = c53_794_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_144_io_in_0 = c53_796_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_144_io_in_1 = c53_795_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_145_io_in_0 = c53_797_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_145_io_in_1 = c53_796_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_146_io_in_0 = c53_798_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_146_io_in_1 = c53_797_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_147_io_in_0 = c53_799_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_147_io_in_1 = c53_798_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_148_io_in_0 = c53_800_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_148_io_in_1 = c53_799_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_149_io_in_0 = c53_801_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_149_io_in_1 = c53_800_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_150_io_in_0 = c53_802_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_150_io_in_1 = c53_801_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_151_io_in_0 = c53_803_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_151_io_in_1 = c53_802_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_64_io_in_0 = c53_804_io_out_0; // @[Multiplier.scala 135:39]
  assign c32_64_io_in_1 = c53_553_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_64_io_in_2 = c53_803_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_65_io_in_0 = c53_805_io_out_0; // @[Multiplier.scala 135:39]
  assign c32_65_io_in_1 = c53_555_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_65_io_in_2 = c53_804_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_66_io_in_0 = c53_806_io_out_0; // @[Multiplier.scala 135:39]
  assign c32_66_io_in_1 = c53_557_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_66_io_in_2 = c53_805_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_67_io_in_0 = c53_807_io_out_0; // @[Multiplier.scala 135:39]
  assign c32_67_io_in_1 = c53_559_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_67_io_in_2 = c53_806_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_68_io_in_0 = c53_808_io_out_0; // @[Multiplier.scala 135:39]
  assign c32_68_io_in_1 = c22_87_io_out_0; // @[Multiplier.scala 122:35]
  assign c32_68_io_in_2 = c53_807_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_924_io_in_0 = c53_809_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_924_io_in_1 = c22_88_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_924_io_in_2 = c53_808_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_924_io_in_3 = c22_87_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_924_io_in_4 = 1'h0; // @[Multiplier.scala 134:24]
  assign c53_925_io_in_0 = c53_810_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_925_io_in_1 = c22_89_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_925_io_in_2 = c53_809_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_925_io_in_3 = c22_88_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_925_io_in_4 = c53_924_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_926_io_in_0 = c53_811_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_926_io_in_1 = c22_90_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_926_io_in_2 = c53_810_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_926_io_in_3 = c22_89_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_926_io_in_4 = c53_925_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_927_io_in_0 = c53_812_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_927_io_in_1 = c22_91_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_927_io_in_2 = c53_811_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_927_io_in_3 = c22_90_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_927_io_in_4 = c53_926_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_928_io_in_0 = c53_813_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_928_io_in_1 = c22_92_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_928_io_in_2 = c53_812_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_928_io_in_3 = c22_91_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_928_io_in_4 = c53_927_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_929_io_in_0 = c53_814_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_929_io_in_1 = c22_93_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_929_io_in_2 = c53_813_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_929_io_in_3 = c22_92_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_929_io_in_4 = c53_928_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_930_io_in_0 = c53_815_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_930_io_in_1 = c22_94_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_930_io_in_2 = c53_814_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_930_io_in_3 = c22_93_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_930_io_in_4 = c53_929_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_931_io_in_0 = c53_816_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_931_io_in_1 = c22_95_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_931_io_in_2 = c53_815_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_931_io_in_3 = c22_94_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_931_io_in_4 = c53_930_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_932_io_in_0 = c53_817_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_932_io_in_1 = c22_96_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_932_io_in_2 = c53_816_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_932_io_in_3 = c22_95_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_932_io_in_4 = c53_931_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_933_io_in_0 = c53_818_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_933_io_in_1 = c22_97_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_933_io_in_2 = c53_817_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_933_io_in_3 = c22_96_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_933_io_in_4 = c53_932_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_934_io_in_0 = c53_819_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_934_io_in_1 = c22_98_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_934_io_in_2 = c53_818_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_934_io_in_3 = c22_97_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_934_io_in_4 = c53_933_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_935_io_in_0 = c53_820_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_935_io_in_1 = c32_56_io_out_0; // @[Multiplier.scala 127:35]
  assign c53_935_io_in_2 = c53_819_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_935_io_in_3 = c22_98_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_935_io_in_4 = c53_934_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_936_io_in_0 = c53_821_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_936_io_in_1 = c32_57_io_out_0; // @[Multiplier.scala 127:35]
  assign c53_936_io_in_2 = c53_820_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_936_io_in_3 = c32_56_io_out_1; // @[Multiplier.scala 128:41]
  assign c53_936_io_in_4 = c53_935_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_937_io_in_0 = c53_822_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_937_io_in_1 = c32_58_io_out_0; // @[Multiplier.scala 127:35]
  assign c53_937_io_in_2 = c53_821_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_937_io_in_3 = c32_57_io_out_1; // @[Multiplier.scala 128:41]
  assign c53_937_io_in_4 = c53_936_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_938_io_in_0 = c53_823_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_938_io_in_1 = c32_59_io_out_0; // @[Multiplier.scala 127:35]
  assign c53_938_io_in_2 = c53_822_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_938_io_in_3 = c32_58_io_out_1; // @[Multiplier.scala 128:41]
  assign c53_938_io_in_4 = c53_937_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_939_io_in_0 = c53_824_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_939_io_in_1 = c53_825_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_939_io_in_2 = c53_823_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_939_io_in_3 = c32_59_io_out_1; // @[Multiplier.scala 128:41]
  assign c53_939_io_in_4 = c53_938_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_940_io_in_0 = c53_826_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_940_io_in_1 = c53_827_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_940_io_in_2 = c53_824_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_940_io_in_3 = c53_825_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_940_io_in_4 = c53_939_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_941_io_in_0 = c53_828_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_941_io_in_1 = c53_829_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_941_io_in_2 = c53_826_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_941_io_in_3 = c53_827_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_941_io_in_4 = c53_940_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_942_io_in_0 = c53_830_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_942_io_in_1 = c53_831_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_942_io_in_2 = c53_828_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_942_io_in_3 = c53_829_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_942_io_in_4 = c53_941_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_943_io_in_0 = c53_832_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_943_io_in_1 = c53_833_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_943_io_in_2 = c53_830_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_943_io_in_3 = c53_831_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_943_io_in_4 = c53_942_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_944_io_in_0 = c53_834_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_944_io_in_1 = c53_835_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_944_io_in_2 = c53_832_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_944_io_in_3 = c53_833_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_944_io_in_4 = c53_943_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_945_io_in_0 = c53_836_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_945_io_in_1 = c53_837_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_945_io_in_2 = c53_834_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_945_io_in_3 = c53_835_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_945_io_in_4 = c53_944_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_946_io_in_0 = c53_838_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_946_io_in_1 = c53_839_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_946_io_in_2 = c53_836_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_946_io_in_3 = c53_837_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_946_io_in_4 = c53_945_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_947_io_in_0 = c53_840_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_947_io_in_1 = c53_841_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_947_io_in_2 = c53_838_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_947_io_in_3 = c53_839_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_947_io_in_4 = c53_946_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_948_io_in_0 = c53_842_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_948_io_in_1 = c53_843_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_948_io_in_2 = c53_840_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_948_io_in_3 = c53_841_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_948_io_in_4 = c53_947_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_949_io_in_0 = c53_844_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_949_io_in_1 = c53_845_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_949_io_in_2 = c53_842_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_949_io_in_3 = c53_843_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_949_io_in_4 = c53_948_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_950_io_in_0 = c53_846_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_950_io_in_1 = c53_847_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_950_io_in_2 = c53_844_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_950_io_in_3 = c53_845_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_950_io_in_4 = c53_949_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_951_io_in_0 = c53_848_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_951_io_in_1 = c53_849_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_951_io_in_2 = c53_643_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_951_io_in_3 = c53_846_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_951_io_in_4 = c53_950_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_952_io_in_0 = c53_850_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_952_io_in_1 = c53_851_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_952_io_in_2 = c53_647_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_952_io_in_3 = c53_848_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_952_io_in_4 = c53_951_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_953_io_in_0 = c53_852_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_953_io_in_1 = c53_853_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_953_io_in_2 = c53_651_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_953_io_in_3 = c53_850_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_953_io_in_4 = c53_952_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_954_io_in_0 = c53_854_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_954_io_in_1 = c53_855_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_954_io_in_2 = c53_655_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_954_io_in_3 = c53_852_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_954_io_in_4 = c53_953_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_955_io_in_0 = c53_856_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_955_io_in_1 = c53_857_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_955_io_in_2 = c53_659_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_955_io_in_3 = c53_854_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_955_io_in_4 = c53_954_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_956_io_in_0 = c53_858_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_956_io_in_1 = c53_859_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_956_io_in_2 = c53_663_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_956_io_in_3 = c53_856_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_956_io_in_4 = c53_955_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_957_io_in_0 = c53_860_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_957_io_in_1 = c53_861_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_957_io_in_2 = c53_667_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_957_io_in_3 = c53_858_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_957_io_in_4 = c53_956_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_958_io_in_0 = c53_862_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_958_io_in_1 = c53_863_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_958_io_in_2 = c53_860_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_958_io_in_3 = c53_861_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_958_io_in_4 = c53_957_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_959_io_in_0 = c53_864_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_959_io_in_1 = c53_865_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_959_io_in_2 = c53_675_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_959_io_in_3 = c53_862_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_959_io_in_4 = c53_958_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_960_io_in_0 = c53_866_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_960_io_in_1 = c53_867_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_960_io_in_2 = c53_864_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_960_io_in_3 = c53_865_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_960_io_in_4 = c53_959_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_961_io_in_0 = c53_868_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_961_io_in_1 = c53_869_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_961_io_in_2 = c53_866_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_961_io_in_3 = c53_867_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_961_io_in_4 = c53_960_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_962_io_in_0 = c53_870_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_962_io_in_1 = c53_871_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_962_io_in_2 = c53_868_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_962_io_in_3 = c53_869_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_962_io_in_4 = c53_961_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_963_io_in_0 = c53_872_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_963_io_in_1 = c53_873_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_963_io_in_2 = c53_870_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_963_io_in_3 = c53_871_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_963_io_in_4 = c53_962_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_964_io_in_0 = c53_874_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_964_io_in_1 = c53_875_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_964_io_in_2 = c53_695_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_964_io_in_3 = c53_872_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_964_io_in_4 = c53_963_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_965_io_in_0 = c53_876_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_965_io_in_1 = c53_877_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_965_io_in_2 = c53_874_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_965_io_in_3 = c53_875_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_965_io_in_4 = c53_964_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_966_io_in_0 = c53_878_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_966_io_in_1 = c53_879_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_966_io_in_2 = c53_876_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_966_io_in_3 = c53_877_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_966_io_in_4 = c53_965_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_967_io_in_0 = c53_880_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_967_io_in_1 = c53_881_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_967_io_in_2 = c53_878_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_967_io_in_3 = c53_879_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_967_io_in_4 = c53_966_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_968_io_in_0 = c53_882_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_968_io_in_1 = c53_883_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_968_io_in_2 = c53_880_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_968_io_in_3 = c53_881_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_968_io_in_4 = c53_967_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_969_io_in_0 = c53_884_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_969_io_in_1 = c53_885_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_969_io_in_2 = c53_882_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_969_io_in_3 = c53_883_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_969_io_in_4 = c53_968_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_970_io_in_0 = c53_886_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_970_io_in_1 = c53_887_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_970_io_in_2 = c53_884_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_970_io_in_3 = c53_885_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_970_io_in_4 = c53_969_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_971_io_in_0 = c53_888_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_971_io_in_1 = c53_889_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_971_io_in_2 = c53_886_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_971_io_in_3 = c53_887_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_971_io_in_4 = c53_970_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_972_io_in_0 = c53_890_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_972_io_in_1 = c53_891_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_972_io_in_2 = c53_888_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_972_io_in_3 = c53_889_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_972_io_in_4 = c53_971_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_973_io_in_0 = c53_892_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_973_io_in_1 = c22_99_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_973_io_in_2 = c53_891_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_973_io_in_3 = c53_890_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_973_io_in_4 = c53_972_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_974_io_in_0 = c53_893_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_974_io_in_1 = c22_100_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_974_io_in_2 = c53_892_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_974_io_in_3 = c22_99_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_974_io_in_4 = c53_973_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_975_io_in_0 = c53_894_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_975_io_in_1 = c32_60_io_out_0; // @[Multiplier.scala 127:35]
  assign c53_975_io_in_2 = c53_893_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_975_io_in_3 = c22_100_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_975_io_in_4 = c53_974_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_976_io_in_0 = c53_895_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_976_io_in_1 = c22_101_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_976_io_in_2 = c53_894_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_976_io_in_3 = c32_60_io_out_1; // @[Multiplier.scala 128:41]
  assign c53_976_io_in_4 = c53_975_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_977_io_in_0 = c53_896_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_977_io_in_1 = c22_102_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_977_io_in_2 = c53_895_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_977_io_in_3 = c22_101_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_977_io_in_4 = c53_976_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_978_io_in_0 = c53_897_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_978_io_in_1 = c22_103_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_978_io_in_2 = c53_896_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_978_io_in_3 = c22_102_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_978_io_in_4 = c53_977_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_979_io_in_0 = c53_898_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_979_io_in_1 = c22_104_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_979_io_in_2 = c53_897_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_979_io_in_3 = c22_103_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_979_io_in_4 = c53_978_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_980_io_in_0 = c53_899_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_980_io_in_1 = c32_61_io_out_0; // @[Multiplier.scala 127:35]
  assign c53_980_io_in_2 = c53_898_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_980_io_in_3 = c22_104_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_980_io_in_4 = c53_979_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_981_io_in_0 = c53_900_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_981_io_in_1 = c22_105_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_981_io_in_2 = c53_899_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_981_io_in_3 = c32_61_io_out_1; // @[Multiplier.scala 128:41]
  assign c53_981_io_in_4 = c53_980_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_982_io_in_0 = c53_901_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_982_io_in_1 = c22_106_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_982_io_in_2 = c53_900_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_982_io_in_3 = c22_105_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_982_io_in_4 = c53_981_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_983_io_in_0 = c53_902_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_983_io_in_1 = c22_107_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_983_io_in_2 = c53_901_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_983_io_in_3 = c22_106_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_983_io_in_4 = c53_982_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_984_io_in_0 = c53_903_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_984_io_in_1 = c22_108_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_984_io_in_2 = c53_902_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_984_io_in_3 = c22_107_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_984_io_in_4 = c53_983_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_985_io_in_0 = c53_904_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_985_io_in_1 = c22_109_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_985_io_in_2 = c53_903_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_985_io_in_3 = c22_108_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_985_io_in_4 = c53_984_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_986_io_in_0 = c53_905_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_986_io_in_1 = c22_110_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_986_io_in_2 = c53_904_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_986_io_in_3 = c22_109_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_986_io_in_4 = c53_985_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_987_io_in_0 = c53_906_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_987_io_in_1 = c22_111_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_987_io_in_2 = c53_905_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_987_io_in_3 = c22_110_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_987_io_in_4 = c53_986_io_out_1; // @[Multiplier.scala 136:41]
  assign c53_988_io_in_0 = c53_907_io_out_0; // @[Multiplier.scala 135:39]
  assign c53_988_io_in_1 = c22_112_io_out_0; // @[Multiplier.scala 122:35]
  assign c53_988_io_in_2 = c53_906_io_out_2; // @[Multiplier.scala 137:41]
  assign c53_988_io_in_3 = c22_111_io_out_1; // @[Multiplier.scala 123:41]
  assign c53_988_io_in_4 = c53_987_io_out_1; // @[Multiplier.scala 136:41]
  assign c32_69_io_in_0 = c53_908_io_out_0; // @[Multiplier.scala 135:39]
  assign c32_69_io_in_1 = c53_907_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_69_io_in_2 = c22_112_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_152_io_in_0 = c53_909_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_152_io_in_1 = c53_908_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_70_io_in_0 = c53_910_io_out_0; // @[Multiplier.scala 135:39]
  assign c32_70_io_in_1 = c53_765_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_70_io_in_2 = c53_909_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_153_io_in_0 = c53_911_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_153_io_in_1 = c53_910_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_154_io_in_0 = c53_912_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_154_io_in_1 = c53_911_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_155_io_in_0 = c53_913_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_155_io_in_1 = c53_912_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_156_io_in_0 = c53_914_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_156_io_in_1 = c53_913_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_71_io_in_0 = c53_915_io_out_0; // @[Multiplier.scala 135:39]
  assign c32_71_io_in_1 = c53_775_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_71_io_in_2 = c53_914_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_157_io_in_0 = c53_916_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_157_io_in_1 = c53_915_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_158_io_in_0 = c53_917_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_158_io_in_1 = c53_916_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_159_io_in_0 = c53_918_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_159_io_in_1 = c53_917_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_160_io_in_0 = c53_919_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_160_io_in_1 = c53_918_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_161_io_in_0 = c53_920_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_161_io_in_1 = c53_919_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_162_io_in_0 = c53_921_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_162_io_in_1 = c53_920_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_163_io_in_0 = c53_922_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_163_io_in_1 = c53_921_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_164_io_in_0 = c53_923_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_164_io_in_1 = c53_922_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_72_io_in_0 = c22_113_io_out_0; // @[Multiplier.scala 122:35]
  assign c32_72_io_in_1 = c53_923_io_out_1; // @[Multiplier.scala 136:41]
  assign c32_72_io_in_2 = c53_923_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_165_io_in_0 = c22_114_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_165_io_in_1 = c22_113_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_166_io_in_0 = c32_62_io_out_0; // @[Multiplier.scala 127:35]
  assign c22_166_io_in_1 = c22_114_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_167_io_in_0 = c22_115_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_167_io_in_1 = c32_62_io_out_1; // @[Multiplier.scala 128:41]
  assign c22_168_io_in_0 = c22_116_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_168_io_in_1 = c22_115_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_169_io_in_0 = c22_117_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_169_io_in_1 = c22_116_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_170_io_in_0 = c22_118_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_170_io_in_1 = c22_117_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_171_io_in_0 = c32_63_io_out_0; // @[Multiplier.scala 127:35]
  assign c22_171_io_in_1 = c22_118_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_172_io_in_0 = c22_119_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_172_io_in_1 = c32_63_io_out_1; // @[Multiplier.scala 128:41]
  assign c22_173_io_in_0 = c22_120_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_173_io_in_1 = c22_119_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_174_io_in_0 = c22_121_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_174_io_in_1 = c22_120_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_175_io_in_0 = c22_122_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_175_io_in_1 = c22_121_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_176_io_in_0 = c22_123_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_176_io_in_1 = c22_122_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_177_io_in_0 = c22_124_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_177_io_in_1 = c22_123_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_178_io_in_0 = c22_126_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_178_io_in_1 = c22_125_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_179_io_in_0 = c22_127_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_179_io_in_1 = c22_126_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_180_io_in_0 = c22_128_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_180_io_in_1 = c22_127_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_181_io_in_0 = c22_129_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_181_io_in_1 = c22_128_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_182_io_in_0 = c22_130_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_182_io_in_1 = c22_129_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_183_io_in_0 = c22_131_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_183_io_in_1 = c22_130_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_184_io_in_0 = c22_132_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_184_io_in_1 = c22_131_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_185_io_in_0 = c22_133_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_185_io_in_1 = c22_132_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_186_io_in_0 = c22_134_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_186_io_in_1 = c22_133_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_187_io_in_0 = c22_135_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_187_io_in_1 = c22_134_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_188_io_in_0 = c22_136_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_188_io_in_1 = c22_135_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_189_io_in_0 = c22_137_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_189_io_in_1 = c22_136_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_190_io_in_0 = c22_138_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_190_io_in_1 = c22_137_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_191_io_in_0 = c22_139_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_191_io_in_1 = c22_138_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_192_io_in_0 = c22_140_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_192_io_in_1 = c22_139_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_193_io_in_0 = c22_141_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_193_io_in_1 = c22_140_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_194_io_in_0 = c22_142_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_194_io_in_1 = c22_141_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_195_io_in_0 = c22_143_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_195_io_in_1 = c22_142_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_196_io_in_0 = c22_144_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_196_io_in_1 = c22_143_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_197_io_in_0 = c22_145_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_197_io_in_1 = c22_144_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_198_io_in_0 = c22_146_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_198_io_in_1 = c22_145_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_199_io_in_0 = c22_147_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_199_io_in_1 = c22_146_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_200_io_in_0 = c22_148_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_200_io_in_1 = c22_147_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_201_io_in_0 = c22_149_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_201_io_in_1 = c22_148_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_202_io_in_0 = c22_150_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_202_io_in_1 = c22_149_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_203_io_in_0 = c22_151_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_203_io_in_1 = c22_150_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_204_io_in_0 = c32_64_io_out_0; // @[Multiplier.scala 127:35]
  assign c22_204_io_in_1 = c22_151_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_205_io_in_0 = c32_65_io_out_0; // @[Multiplier.scala 127:35]
  assign c22_205_io_in_1 = c32_64_io_out_1; // @[Multiplier.scala 128:41]
  assign c22_206_io_in_0 = c32_66_io_out_0; // @[Multiplier.scala 127:35]
  assign c22_206_io_in_1 = c32_65_io_out_1; // @[Multiplier.scala 128:41]
  assign c22_207_io_in_0 = c32_67_io_out_0; // @[Multiplier.scala 127:35]
  assign c22_207_io_in_1 = c32_66_io_out_1; // @[Multiplier.scala 128:41]
  assign c22_208_io_in_0 = c32_68_io_out_0; // @[Multiplier.scala 127:35]
  assign c22_208_io_in_1 = c32_67_io_out_1; // @[Multiplier.scala 128:41]
  assign c22_209_io_in_0 = c53_924_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_209_io_in_1 = c32_68_io_out_1; // @[Multiplier.scala 128:41]
  assign c22_210_io_in_0 = c53_925_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_210_io_in_1 = c53_924_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_211_io_in_0 = c53_926_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_211_io_in_1 = c53_925_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_212_io_in_0 = c53_927_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_212_io_in_1 = c53_926_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_213_io_in_0 = c53_928_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_213_io_in_1 = c53_927_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_214_io_in_0 = c53_929_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_214_io_in_1 = c53_928_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_215_io_in_0 = c53_930_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_215_io_in_1 = c53_929_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_216_io_in_0 = c53_931_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_216_io_in_1 = c53_930_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_217_io_in_0 = c53_932_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_217_io_in_1 = c53_931_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_218_io_in_0 = c53_933_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_218_io_in_1 = c53_932_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_219_io_in_0 = c53_934_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_219_io_in_1 = c53_933_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_220_io_in_0 = c53_935_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_220_io_in_1 = c53_934_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_221_io_in_0 = c53_936_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_221_io_in_1 = c53_935_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_222_io_in_0 = c53_937_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_222_io_in_1 = c53_936_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_223_io_in_0 = c53_938_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_223_io_in_1 = c53_937_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_224_io_in_0 = c53_939_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_224_io_in_1 = c53_938_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_225_io_in_0 = c53_940_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_225_io_in_1 = c53_939_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_226_io_in_0 = c53_941_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_226_io_in_1 = c53_940_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_227_io_in_0 = c53_942_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_227_io_in_1 = c53_941_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_228_io_in_0 = c53_943_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_228_io_in_1 = c53_942_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_229_io_in_0 = c53_944_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_229_io_in_1 = c53_943_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_230_io_in_0 = c53_945_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_230_io_in_1 = c53_944_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_231_io_in_0 = c53_946_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_231_io_in_1 = c53_945_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_232_io_in_0 = c53_947_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_232_io_in_1 = c53_946_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_233_io_in_0 = c53_948_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_233_io_in_1 = c53_947_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_234_io_in_0 = c53_949_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_234_io_in_1 = c53_948_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_235_io_in_0 = c53_950_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_235_io_in_1 = c53_949_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_73_io_in_0 = c53_951_io_out_0; // @[Multiplier.scala 135:39]
  assign c32_73_io_in_1 = c53_847_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_73_io_in_2 = c53_950_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_74_io_in_0 = c53_952_io_out_0; // @[Multiplier.scala 135:39]
  assign c32_74_io_in_1 = c53_849_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_74_io_in_2 = c53_951_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_75_io_in_0 = c53_953_io_out_0; // @[Multiplier.scala 135:39]
  assign c32_75_io_in_1 = c53_851_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_75_io_in_2 = c53_952_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_76_io_in_0 = c53_954_io_out_0; // @[Multiplier.scala 135:39]
  assign c32_76_io_in_1 = c53_853_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_76_io_in_2 = c53_953_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_77_io_in_0 = c53_955_io_out_0; // @[Multiplier.scala 135:39]
  assign c32_77_io_in_1 = c53_855_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_77_io_in_2 = c53_954_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_78_io_in_0 = c53_956_io_out_0; // @[Multiplier.scala 135:39]
  assign c32_78_io_in_1 = c53_857_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_78_io_in_2 = c53_955_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_79_io_in_0 = c53_957_io_out_0; // @[Multiplier.scala 135:39]
  assign c32_79_io_in_1 = c53_859_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_79_io_in_2 = c53_956_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_236_io_in_0 = c53_958_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_236_io_in_1 = c53_957_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_80_io_in_0 = c53_959_io_out_0; // @[Multiplier.scala 135:39]
  assign c32_80_io_in_1 = c53_863_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_80_io_in_2 = c53_958_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_237_io_in_0 = c53_960_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_237_io_in_1 = c53_959_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_238_io_in_0 = c53_961_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_238_io_in_1 = c53_960_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_239_io_in_0 = c53_962_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_239_io_in_1 = c53_961_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_240_io_in_0 = c53_963_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_240_io_in_1 = c53_962_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_81_io_in_0 = c53_964_io_out_0; // @[Multiplier.scala 135:39]
  assign c32_81_io_in_1 = c53_873_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_81_io_in_2 = c53_963_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_241_io_in_0 = c53_965_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_241_io_in_1 = c53_964_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_242_io_in_0 = c53_966_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_242_io_in_1 = c53_965_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_243_io_in_0 = c53_967_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_243_io_in_1 = c53_966_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_244_io_in_0 = c53_968_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_244_io_in_1 = c53_967_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_245_io_in_0 = c53_969_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_245_io_in_1 = c53_968_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_246_io_in_0 = c53_970_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_246_io_in_1 = c53_969_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_247_io_in_0 = c53_971_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_247_io_in_1 = c53_970_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_248_io_in_0 = c53_972_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_248_io_in_1 = c53_971_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_82_io_in_0 = c53_973_io_out_0; // @[Multiplier.scala 135:39]
  assign c32_82_io_in_1 = c53_891_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_82_io_in_2 = c53_972_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_249_io_in_0 = c53_974_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_249_io_in_1 = c53_973_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_250_io_in_0 = c53_975_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_250_io_in_1 = c53_974_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_251_io_in_0 = c53_976_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_251_io_in_1 = c53_975_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_252_io_in_0 = c53_977_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_252_io_in_1 = c53_976_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_253_io_in_0 = c53_978_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_253_io_in_1 = c53_977_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_254_io_in_0 = c53_979_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_254_io_in_1 = c53_978_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_255_io_in_0 = c53_980_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_255_io_in_1 = c53_979_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_256_io_in_0 = c53_981_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_256_io_in_1 = c53_980_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_257_io_in_0 = c53_982_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_257_io_in_1 = c53_981_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_258_io_in_0 = c53_983_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_258_io_in_1 = c53_982_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_259_io_in_0 = c53_984_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_259_io_in_1 = c53_983_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_260_io_in_0 = c53_985_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_260_io_in_1 = c53_984_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_261_io_in_0 = c53_986_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_261_io_in_1 = c53_985_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_262_io_in_0 = c53_987_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_262_io_in_1 = c53_986_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_263_io_in_0 = c53_988_io_out_0; // @[Multiplier.scala 135:39]
  assign c22_263_io_in_1 = c53_987_io_out_2; // @[Multiplier.scala 137:41]
  assign c32_83_io_in_0 = c32_69_io_out_0; // @[Multiplier.scala 127:35]
  assign c32_83_io_in_1 = c53_988_io_out_1; // @[Multiplier.scala 136:41]
  assign c32_83_io_in_2 = c53_988_io_out_2; // @[Multiplier.scala 137:41]
  assign c22_264_io_in_0 = c22_152_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_264_io_in_1 = c32_69_io_out_1; // @[Multiplier.scala 128:41]
  assign c22_265_io_in_0 = c32_70_io_out_0; // @[Multiplier.scala 127:35]
  assign c22_265_io_in_1 = c22_152_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_266_io_in_0 = c22_153_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_266_io_in_1 = c32_70_io_out_1; // @[Multiplier.scala 128:41]
  assign c22_267_io_in_0 = c22_154_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_267_io_in_1 = c22_153_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_268_io_in_0 = c22_155_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_268_io_in_1 = c22_154_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_269_io_in_0 = c22_156_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_269_io_in_1 = c22_155_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_270_io_in_0 = c32_71_io_out_0; // @[Multiplier.scala 127:35]
  assign c22_270_io_in_1 = c22_156_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_271_io_in_0 = c22_157_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_271_io_in_1 = c32_71_io_out_1; // @[Multiplier.scala 128:41]
  assign c22_272_io_in_0 = c22_158_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_272_io_in_1 = c22_157_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_273_io_in_0 = c22_159_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_273_io_in_1 = c22_158_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_274_io_in_0 = c22_160_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_274_io_in_1 = c22_159_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_275_io_in_0 = c22_161_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_275_io_in_1 = c22_160_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_276_io_in_0 = c22_162_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_276_io_in_1 = c22_161_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_277_io_in_0 = c22_163_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_277_io_in_1 = c22_162_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_278_io_in_0 = c22_164_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_278_io_in_1 = c22_163_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_279_io_in_0 = c32_72_io_out_0; // @[Multiplier.scala 127:35]
  assign c22_279_io_in_1 = c22_164_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_280_io_in_0 = c22_165_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_280_io_in_1 = c32_72_io_out_1; // @[Multiplier.scala 128:41]
  assign c22_281_io_in_0 = c22_166_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_281_io_in_1 = c22_165_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_282_io_in_0 = c22_167_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_282_io_in_1 = c22_166_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_283_io_in_0 = c22_168_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_283_io_in_1 = c22_167_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_284_io_in_0 = c22_169_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_284_io_in_1 = c22_168_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_285_io_in_0 = c22_170_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_285_io_in_1 = c22_169_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_286_io_in_0 = c22_171_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_286_io_in_1 = c22_170_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_287_io_in_0 = c22_172_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_287_io_in_1 = c22_171_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_288_io_in_0 = c22_173_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_288_io_in_1 = c22_172_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_289_io_in_0 = c22_174_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_289_io_in_1 = c22_173_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_290_io_in_0 = c22_175_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_290_io_in_1 = c22_174_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_291_io_in_0 = c22_176_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_291_io_in_1 = c22_175_io_out_1; // @[Multiplier.scala 123:41]
  assign c22_292_io_in_0 = c22_177_io_out_0; // @[Multiplier.scala 122:35]
  assign c22_292_io_in_1 = c22_176_io_out_1; // @[Multiplier.scala 123:41]
  always @(posedge clock) begin
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r <= pp[0]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1 <= pp_1[0]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2 <= pp[1]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_3 <= pp_1[1]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_4 <= pp[2]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_5 <= pp_1[2]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_6 <= pp_2[0]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_7 <= pp[3]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_8 <= pp_1[3]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_9 <= pp_2[1]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_10 <= pp[4]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_11 <= pp_1[4]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_12 <= pp_2[2]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_13 <= pp_3[0]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_14 <= pp[5]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_15 <= pp_1[5]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_16 <= pp_2[3]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_17 <= pp_3[1]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_18 <= pp[6]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_19 <= pp_1[6]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_20 <= pp_2[4]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_21 <= pp_3[2]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_22 <= pp_4[0]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_23 <= pp[7]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_24 <= pp_1[7]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_25 <= pp_2[5]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_26 <= pp_3[3]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_27 <= pp_4[1]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_28 <= pp[8]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_29 <= pp_1[8]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_30 <= pp_2[6]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_31 <= pp_3[4]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_32 <= pp_4[2]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_33 <= pp_5[0]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_34 <= pp[9]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_35 <= pp_1[9]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_36 <= pp_2[7]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_37 <= pp_3[5]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_38 <= pp_4[3]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_39 <= pp_5[1]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_40 <= pp[10]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_41 <= pp_1[10]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_42 <= pp_2[8]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_43 <= pp_3[6]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_44 <= pp_4[4]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_45 <= pp_5[2]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_46 <= pp_6[0]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_47 <= pp[11]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_48 <= pp_1[11]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_49 <= pp_2[9]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_50 <= pp_3[7]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_51 <= pp_4[5]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_52 <= pp_5[3]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_53 <= pp_6[1]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_54 <= pp[12]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_55 <= pp_1[12]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_56 <= pp_2[10]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_57 <= pp_3[8]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_58 <= pp_4[6]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_59 <= pp_5[4]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_60 <= pp_6[2]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_61 <= pp_7[0]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_62 <= pp[13]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_63 <= pp_1[13]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_64 <= pp_2[11]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_65 <= pp_3[9]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_66 <= pp_4[7]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_67 <= pp_5[5]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_68 <= pp_6[3]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_69 <= pp_7[1]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_70 <= pp[14]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_71 <= pp_1[14]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_72 <= pp_2[12]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_73 <= pp_3[10]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_74 <= pp_4[8]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_75 <= pp_5[6]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_76 <= pp_6[4]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_77 <= pp_7[2]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_78 <= pp_8[0]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_79 <= pp[15]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_80 <= pp_1[15]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_81 <= pp_2[13]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_82 <= pp_3[11]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_83 <= pp_4[9]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_84 <= pp_5[7]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_85 <= pp_6[5]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_86 <= pp_7[3]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_87 <= pp_8[1]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_88 <= pp[16]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_89 <= pp_1[16]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_90 <= pp_2[14]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_91 <= pp_3[12]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_92 <= pp_4[10]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_93 <= pp_5[8]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_94 <= pp_6[6]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_95 <= pp_7[4]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_96 <= pp_8[2]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_97 <= pp_9[0]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_98 <= pp[17]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_99 <= pp_1[17]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_100 <= pp_2[15]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_101 <= pp_3[13]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_102 <= pp_4[11]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_103 <= pp_5[9]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_104 <= pp_6[7]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_105 <= pp_7[5]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_106 <= pp_8[3]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_107 <= pp_9[1]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_108 <= pp[18]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_109 <= pp_1[18]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_110 <= pp_2[16]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_111 <= pp_3[14]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_112 <= pp_4[12]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_113 <= pp_5[10]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_114 <= pp_6[8]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_115 <= pp_7[6]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_116 <= pp_8[4]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_117 <= pp_9[2]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_118 <= pp_10[0]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_119 <= pp[19]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_120 <= pp_1[19]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_121 <= pp_2[17]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_122 <= pp_3[15]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_123 <= pp_4[13]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_124 <= pp_5[11]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_125 <= pp_6[9]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_126 <= pp_7[7]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_127 <= pp_8[5]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_128 <= pp_9[3]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_129 <= pp_10[1]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_130 <= pp[20]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_131 <= pp_1[20]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_132 <= pp_2[18]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_133 <= pp_3[16]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_134 <= pp_4[14]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_135 <= pp_5[12]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_136 <= pp_6[10]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_137 <= pp_7[8]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_138 <= pp_8[6]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_139 <= pp_9[4]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_140 <= pp_10[2]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_141 <= pp_11[0]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_142 <= pp[21]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_143 <= pp_1[21]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_144 <= pp_2[19]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_145 <= pp_3[17]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_146 <= pp_4[15]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_147 <= pp_5[13]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_148 <= pp_6[11]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_149 <= pp_7[9]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_150 <= pp_8[7]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_151 <= pp_9[5]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_152 <= pp_10[3]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_153 <= pp_11[1]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_154 <= pp[22]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_155 <= pp_1[22]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_156 <= pp_2[20]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_157 <= pp_3[18]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_158 <= pp_4[16]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_159 <= pp_5[14]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_160 <= pp_6[12]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_161 <= pp_7[10]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_162 <= pp_8[8]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_163 <= pp_9[6]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_164 <= pp_10[4]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_165 <= pp_11[2]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_166 <= pp_12[0]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_167 <= pp[23]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_168 <= pp_1[23]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_169 <= pp_2[21]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_170 <= pp_3[19]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_171 <= pp_4[17]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_172 <= pp_5[15]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_173 <= pp_6[13]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_174 <= pp_7[11]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_175 <= pp_8[9]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_176 <= pp_9[7]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_177 <= pp_10[5]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_178 <= pp_11[3]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_179 <= pp_12[1]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_180 <= pp[24]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_181 <= pp_1[24]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_182 <= pp_2[22]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_183 <= pp_3[20]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_184 <= pp_4[18]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_185 <= pp_5[16]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_186 <= pp_6[14]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_187 <= pp_7[12]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_188 <= pp_8[10]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_189 <= pp_9[8]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_190 <= pp_10[6]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_191 <= pp_11[4]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_192 <= pp_12[2]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_193 <= pp_13[0]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_194 <= pp[25]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_195 <= pp_1[25]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_196 <= pp_2[23]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_197 <= pp_3[21]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_198 <= pp_4[19]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_199 <= pp_5[17]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_200 <= pp_6[15]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_201 <= pp_7[13]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_202 <= pp_8[11]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_203 <= pp_9[9]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_204 <= pp_10[7]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_205 <= pp_11[5]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_206 <= pp_12[3]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_207 <= pp_13[1]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_208 <= pp[26]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_209 <= pp_1[26]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_210 <= pp_2[24]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_211 <= pp_3[22]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_212 <= pp_4[20]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_213 <= pp_5[18]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_214 <= pp_6[16]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_215 <= pp_7[14]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_216 <= pp_8[12]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_217 <= pp_9[10]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_218 <= pp_10[8]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_219 <= pp_11[6]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_220 <= pp_12[4]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_221 <= pp_13[2]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_222 <= pp_14[0]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_223 <= pp[27]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_224 <= pp_1[27]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_225 <= pp_2[25]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_226 <= pp_3[23]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_227 <= pp_4[21]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_228 <= pp_5[19]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_229 <= pp_6[17]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_230 <= pp_7[15]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_231 <= pp_8[13]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_232 <= pp_9[11]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_233 <= pp_10[9]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_234 <= pp_11[7]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_235 <= pp_12[5]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_236 <= pp_13[3]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_237 <= pp_14[1]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_238 <= pp[28]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_239 <= pp_1[28]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_240 <= pp_2[26]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_241 <= pp_3[24]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_242 <= pp_4[22]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_243 <= pp_5[20]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_244 <= pp_6[18]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_245 <= pp_7[16]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_246 <= pp_8[14]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_247 <= pp_9[12]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_248 <= pp_10[10]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_249 <= pp_11[8]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_250 <= pp_12[6]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_251 <= pp_13[4]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_252 <= pp_14[2]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_253 <= pp_15[0]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_254 <= pp[29]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_255 <= pp_1[29]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_256 <= pp_2[27]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_257 <= pp_3[25]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_258 <= pp_4[23]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_259 <= pp_5[21]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_260 <= pp_6[19]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_261 <= pp_7[17]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_262 <= pp_8[15]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_263 <= pp_9[13]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_264 <= pp_10[11]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_265 <= pp_11[9]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_266 <= pp_12[7]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_267 <= pp_13[5]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_268 <= pp_14[3]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_269 <= pp_15[1]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_270 <= pp[30]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_271 <= pp_1[30]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_272 <= pp_2[28]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_273 <= pp_3[26]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_274 <= pp_4[24]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_275 <= pp_5[22]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_276 <= pp_6[20]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_277 <= pp_7[18]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_278 <= pp_8[16]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_279 <= pp_9[14]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_280 <= pp_10[12]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_281 <= pp_11[10]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_282 <= pp_12[8]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_283 <= pp_13[6]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_284 <= pp_14[4]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_285 <= pp_15[2]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_286 <= pp_16[0]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_287 <= pp[31]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_288 <= pp_1[31]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_289 <= pp_2[29]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_290 <= pp_3[27]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_291 <= pp_4[25]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_292 <= pp_5[23]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_293 <= pp_6[21]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_294 <= pp_7[19]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_295 <= pp_8[17]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_296 <= pp_9[15]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_297 <= pp_10[13]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_298 <= pp_11[11]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_299 <= pp_12[9]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_300 <= pp_13[7]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_301 <= pp_14[5]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_302 <= pp_15[3]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_303 <= pp_16[1]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_304 <= pp[32]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_305 <= pp_1[32]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_306 <= pp_2[30]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_307 <= pp_3[28]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_308 <= pp_4[26]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_309 <= pp_5[24]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_310 <= pp_6[22]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_311 <= pp_7[20]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_312 <= pp_8[18]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_313 <= pp_9[16]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_314 <= pp_10[14]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_315 <= pp_11[12]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_316 <= pp_12[10]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_317 <= pp_13[8]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_318 <= pp_14[6]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_319 <= pp_15[4]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_320 <= pp_16[2]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_321 <= pp_17[0]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_322 <= pp[33]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_323 <= pp_1[33]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_324 <= pp_2[31]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_325 <= pp_3[29]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_326 <= pp_4[27]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_327 <= pp_5[25]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_328 <= pp_6[23]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_329 <= pp_7[21]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_330 <= pp_8[19]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_331 <= pp_9[17]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_332 <= pp_10[15]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_333 <= pp_11[13]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_334 <= pp_12[11]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_335 <= pp_13[9]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_336 <= pp_14[7]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_337 <= pp_15[5]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_338 <= pp_16[3]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_339 <= pp_17[1]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_340 <= pp[34]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_341 <= pp_1[34]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_342 <= pp_2[32]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_343 <= pp_3[30]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_344 <= pp_4[28]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_345 <= pp_5[26]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_346 <= pp_6[24]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_347 <= pp_7[22]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_348 <= pp_8[20]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_349 <= pp_9[18]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_350 <= pp_10[16]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_351 <= pp_11[14]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_352 <= pp_12[12]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_353 <= pp_13[10]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_354 <= pp_14[8]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_355 <= pp_15[6]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_356 <= pp_16[4]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_357 <= pp_17[2]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_358 <= pp_18[0]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_359 <= pp[35]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_360 <= pp_1[35]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_361 <= pp_2[33]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_362 <= pp_3[31]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_363 <= pp_4[29]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_364 <= pp_5[27]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_365 <= pp_6[25]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_366 <= pp_7[23]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_367 <= pp_8[21]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_368 <= pp_9[19]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_369 <= pp_10[17]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_370 <= pp_11[15]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_371 <= pp_12[13]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_372 <= pp_13[11]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_373 <= pp_14[9]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_374 <= pp_15[7]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_375 <= pp_16[5]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_376 <= pp_17[3]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_377 <= pp_18[1]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_378 <= pp[36]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_379 <= pp_1[36]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_380 <= pp_2[34]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_381 <= pp_3[32]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_382 <= pp_4[30]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_383 <= pp_5[28]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_384 <= pp_6[26]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_385 <= pp_7[24]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_386 <= pp_8[22]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_387 <= pp_9[20]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_388 <= pp_10[18]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_389 <= pp_11[16]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_390 <= pp_12[14]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_391 <= pp_13[12]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_392 <= pp_14[10]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_393 <= pp_15[8]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_394 <= pp_16[6]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_395 <= pp_17[4]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_396 <= pp_18[2]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_397 <= pp_19[0]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_398 <= pp[37]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_399 <= pp_1[37]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_400 <= pp_2[35]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_401 <= pp_3[33]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_402 <= pp_4[31]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_403 <= pp_5[29]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_404 <= pp_6[27]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_405 <= pp_7[25]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_406 <= pp_8[23]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_407 <= pp_9[21]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_408 <= pp_10[19]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_409 <= pp_11[17]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_410 <= pp_12[15]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_411 <= pp_13[13]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_412 <= pp_14[11]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_413 <= pp_15[9]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_414 <= pp_16[7]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_415 <= pp_17[5]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_416 <= pp_18[3]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_417 <= pp_19[1]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_418 <= pp[38]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_419 <= pp_1[38]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_420 <= pp_2[36]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_421 <= pp_3[34]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_422 <= pp_4[32]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_423 <= pp_5[30]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_424 <= pp_6[28]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_425 <= pp_7[26]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_426 <= pp_8[24]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_427 <= pp_9[22]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_428 <= pp_10[20]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_429 <= pp_11[18]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_430 <= pp_12[16]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_431 <= pp_13[14]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_432 <= pp_14[12]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_433 <= pp_15[10]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_434 <= pp_16[8]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_435 <= pp_17[6]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_436 <= pp_18[4]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_437 <= pp_19[2]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_438 <= pp_20[0]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_439 <= pp[39]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_440 <= pp_1[39]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_441 <= pp_2[37]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_442 <= pp_3[35]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_443 <= pp_4[33]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_444 <= pp_5[31]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_445 <= pp_6[29]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_446 <= pp_7[27]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_447 <= pp_8[25]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_448 <= pp_9[23]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_449 <= pp_10[21]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_450 <= pp_11[19]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_451 <= pp_12[17]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_452 <= pp_13[15]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_453 <= pp_14[13]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_454 <= pp_15[11]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_455 <= pp_16[9]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_456 <= pp_17[7]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_457 <= pp_18[5]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_458 <= pp_19[3]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_459 <= pp_20[1]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_460 <= pp[40]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_461 <= pp_1[40]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_462 <= pp_2[38]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_463 <= pp_3[36]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_464 <= pp_4[34]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_465 <= pp_5[32]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_466 <= pp_6[30]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_467 <= pp_7[28]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_468 <= pp_8[26]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_469 <= pp_9[24]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_470 <= pp_10[22]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_471 <= pp_11[20]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_472 <= pp_12[18]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_473 <= pp_13[16]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_474 <= pp_14[14]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_475 <= pp_15[12]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_476 <= pp_16[10]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_477 <= pp_17[8]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_478 <= pp_18[6]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_479 <= pp_19[4]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_480 <= pp_20[2]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_481 <= pp_21[0]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_482 <= pp[41]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_483 <= pp_1[41]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_484 <= pp_2[39]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_485 <= pp_3[37]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_486 <= pp_4[35]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_487 <= pp_5[33]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_488 <= pp_6[31]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_489 <= pp_7[29]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_490 <= pp_8[27]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_491 <= pp_9[25]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_492 <= pp_10[23]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_493 <= pp_11[21]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_494 <= pp_12[19]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_495 <= pp_13[17]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_496 <= pp_14[15]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_497 <= pp_15[13]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_498 <= pp_16[11]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_499 <= pp_17[9]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_500 <= pp_18[7]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_501 <= pp_19[5]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_502 <= pp_20[3]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_503 <= pp_21[1]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_504 <= pp[42]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_505 <= pp_1[42]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_506 <= pp_2[40]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_507 <= pp_3[38]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_508 <= pp_4[36]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_509 <= pp_5[34]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_510 <= pp_6[32]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_511 <= pp_7[30]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_512 <= pp_8[28]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_513 <= pp_9[26]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_514 <= pp_10[24]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_515 <= pp_11[22]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_516 <= pp_12[20]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_517 <= pp_13[18]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_518 <= pp_14[16]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_519 <= pp_15[14]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_520 <= pp_16[12]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_521 <= pp_17[10]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_522 <= pp_18[8]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_523 <= pp_19[6]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_524 <= pp_20[4]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_525 <= pp_21[2]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_526 <= pp_22[0]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_527 <= pp[43]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_528 <= pp_1[43]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_529 <= pp_2[41]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_530 <= pp_3[39]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_531 <= pp_4[37]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_532 <= pp_5[35]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_533 <= pp_6[33]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_534 <= pp_7[31]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_535 <= pp_8[29]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_536 <= pp_9[27]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_537 <= pp_10[25]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_538 <= pp_11[23]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_539 <= pp_12[21]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_540 <= pp_13[19]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_541 <= pp_14[17]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_542 <= pp_15[15]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_543 <= pp_16[13]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_544 <= pp_17[11]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_545 <= pp_18[9]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_546 <= pp_19[7]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_547 <= pp_20[5]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_548 <= pp_21[3]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_549 <= pp_22[1]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_550 <= pp[44]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_551 <= pp_1[44]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_552 <= pp_2[42]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_553 <= pp_3[40]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_554 <= pp_4[38]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_555 <= pp_5[36]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_556 <= pp_6[34]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_557 <= pp_7[32]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_558 <= pp_8[30]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_559 <= pp_9[28]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_560 <= pp_10[26]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_561 <= pp_11[24]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_562 <= pp_12[22]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_563 <= pp_13[20]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_564 <= pp_14[18]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_565 <= pp_15[16]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_566 <= pp_16[14]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_567 <= pp_17[12]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_568 <= pp_18[10]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_569 <= pp_19[8]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_570 <= pp_20[6]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_571 <= pp_21[4]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_572 <= pp_22[2]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_573 <= pp_23[0]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_574 <= pp[45]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_575 <= pp_1[45]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_576 <= pp_2[43]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_577 <= pp_3[41]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_578 <= pp_4[39]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_579 <= pp_5[37]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_580 <= pp_6[35]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_581 <= pp_7[33]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_582 <= pp_8[31]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_583 <= pp_9[29]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_584 <= pp_10[27]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_585 <= pp_11[25]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_586 <= pp_12[23]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_587 <= pp_13[21]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_588 <= pp_14[19]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_589 <= pp_15[17]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_590 <= pp_16[15]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_591 <= pp_17[13]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_592 <= pp_18[11]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_593 <= pp_19[9]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_594 <= pp_20[7]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_595 <= pp_21[5]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_596 <= pp_22[3]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_597 <= pp_23[1]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_598 <= pp[46]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_599 <= pp_1[46]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_600 <= pp_2[44]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_601 <= pp_3[42]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_602 <= pp_4[40]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_603 <= pp_5[38]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_604 <= pp_6[36]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_605 <= pp_7[34]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_606 <= pp_8[32]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_607 <= pp_9[30]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_608 <= pp_10[28]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_609 <= pp_11[26]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_610 <= pp_12[24]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_611 <= pp_13[22]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_612 <= pp_14[20]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_613 <= pp_15[18]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_614 <= pp_16[16]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_615 <= pp_17[14]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_616 <= pp_18[12]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_617 <= pp_19[10]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_618 <= pp_20[8]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_619 <= pp_21[6]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_620 <= pp_22[4]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_621 <= pp_23[2]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_622 <= pp_24[0]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_623 <= pp[47]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_624 <= pp_1[47]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_625 <= pp_2[45]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_626 <= pp_3[43]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_627 <= pp_4[41]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_628 <= pp_5[39]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_629 <= pp_6[37]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_630 <= pp_7[35]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_631 <= pp_8[33]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_632 <= pp_9[31]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_633 <= pp_10[29]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_634 <= pp_11[27]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_635 <= pp_12[25]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_636 <= pp_13[23]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_637 <= pp_14[21]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_638 <= pp_15[19]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_639 <= pp_16[17]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_640 <= pp_17[15]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_641 <= pp_18[13]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_642 <= pp_19[11]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_643 <= pp_20[9]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_644 <= pp_21[7]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_645 <= pp_22[5]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_646 <= pp_23[3]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_647 <= pp_24[1]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_648 <= pp[48]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_649 <= pp_1[48]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_650 <= pp_2[46]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_651 <= pp_3[44]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_652 <= pp_4[42]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_653 <= pp_5[40]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_654 <= pp_6[38]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_655 <= pp_7[36]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_656 <= pp_8[34]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_657 <= pp_9[32]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_658 <= pp_10[30]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_659 <= pp_11[28]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_660 <= pp_12[26]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_661 <= pp_13[24]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_662 <= pp_14[22]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_663 <= pp_15[20]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_664 <= pp_16[18]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_665 <= pp_17[16]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_666 <= pp_18[14]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_667 <= pp_19[12]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_668 <= pp_20[10]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_669 <= pp_21[8]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_670 <= pp_22[6]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_671 <= pp_23[4]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_672 <= pp_24[2]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_673 <= pp_25[0]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_674 <= pp[49]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_675 <= pp_1[49]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_676 <= pp_2[47]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_677 <= pp_3[45]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_678 <= pp_4[43]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_679 <= pp_5[41]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_680 <= pp_6[39]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_681 <= pp_7[37]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_682 <= pp_8[35]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_683 <= pp_9[33]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_684 <= pp_10[31]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_685 <= pp_11[29]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_686 <= pp_12[27]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_687 <= pp_13[25]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_688 <= pp_14[23]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_689 <= pp_15[21]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_690 <= pp_16[19]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_691 <= pp_17[17]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_692 <= pp_18[15]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_693 <= pp_19[13]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_694 <= pp_20[11]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_695 <= pp_21[9]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_696 <= pp_22[7]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_697 <= pp_23[5]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_698 <= pp_24[3]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_699 <= pp_25[1]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_700 <= pp[50]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_701 <= pp_1[50]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_702 <= pp_2[48]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_703 <= pp_3[46]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_704 <= pp_4[44]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_705 <= pp_5[42]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_706 <= pp_6[40]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_707 <= pp_7[38]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_708 <= pp_8[36]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_709 <= pp_9[34]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_710 <= pp_10[32]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_711 <= pp_11[30]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_712 <= pp_12[28]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_713 <= pp_13[26]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_714 <= pp_14[24]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_715 <= pp_15[22]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_716 <= pp_16[20]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_717 <= pp_17[18]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_718 <= pp_18[16]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_719 <= pp_19[14]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_720 <= pp_20[12]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_721 <= pp_21[10]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_722 <= pp_22[8]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_723 <= pp_23[6]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_724 <= pp_24[4]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_725 <= pp_25[2]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_726 <= pp_26[0]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_727 <= pp[51]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_728 <= pp_1[51]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_729 <= pp_2[49]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_730 <= pp_3[47]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_731 <= pp_4[45]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_732 <= pp_5[43]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_733 <= pp_6[41]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_734 <= pp_7[39]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_735 <= pp_8[37]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_736 <= pp_9[35]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_737 <= pp_10[33]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_738 <= pp_11[31]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_739 <= pp_12[29]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_740 <= pp_13[27]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_741 <= pp_14[25]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_742 <= pp_15[23]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_743 <= pp_16[21]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_744 <= pp_17[19]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_745 <= pp_18[17]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_746 <= pp_19[15]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_747 <= pp_20[13]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_748 <= pp_21[11]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_749 <= pp_22[9]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_750 <= pp_23[7]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_751 <= pp_24[5]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_752 <= pp_25[3]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_753 <= pp_26[1]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_754 <= pp[52]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_755 <= pp_1[52]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_756 <= pp_2[50]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_757 <= pp_3[48]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_758 <= pp_4[46]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_759 <= pp_5[44]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_760 <= pp_6[42]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_761 <= pp_7[40]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_762 <= pp_8[38]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_763 <= pp_9[36]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_764 <= pp_10[34]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_765 <= pp_11[32]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_766 <= pp_12[30]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_767 <= pp_13[28]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_768 <= pp_14[26]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_769 <= pp_15[24]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_770 <= pp_16[22]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_771 <= pp_17[20]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_772 <= pp_18[18]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_773 <= pp_19[16]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_774 <= pp_20[14]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_775 <= pp_21[12]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_776 <= pp_22[10]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_777 <= pp_23[8]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_778 <= pp_24[6]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_779 <= pp_25[4]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_780 <= pp_26[2]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_781 <= pp_27[0]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_782 <= pp[53]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_783 <= pp_1[53]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_784 <= pp_2[51]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_785 <= pp_3[49]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_786 <= pp_4[47]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_787 <= pp_5[45]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_788 <= pp_6[43]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_789 <= pp_7[41]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_790 <= pp_8[39]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_791 <= pp_9[37]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_792 <= pp_10[35]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_793 <= pp_11[33]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_794 <= pp_12[31]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_795 <= pp_13[29]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_796 <= pp_14[27]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_797 <= pp_15[25]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_798 <= pp_16[23]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_799 <= pp_17[21]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_800 <= pp_18[19]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_801 <= pp_19[17]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_802 <= pp_20[15]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_803 <= pp_21[13]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_804 <= pp_22[11]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_805 <= pp_23[9]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_806 <= pp_24[7]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_807 <= pp_25[5]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_808 <= pp_26[3]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_809 <= pp_27[1]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_810 <= pp[54]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_811 <= pp_1[54]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_812 <= pp_2[52]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_813 <= pp_3[50]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_814 <= pp_4[48]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_815 <= pp_5[46]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_816 <= pp_6[44]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_817 <= pp_7[42]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_818 <= pp_8[40]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_819 <= pp_9[38]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_820 <= pp_10[36]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_821 <= pp_11[34]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_822 <= pp_12[32]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_823 <= pp_13[30]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_824 <= pp_14[28]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_825 <= pp_15[26]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_826 <= pp_16[24]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_827 <= pp_17[22]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_828 <= pp_18[20]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_829 <= pp_19[18]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_830 <= pp_20[16]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_831 <= pp_21[14]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_832 <= pp_22[12]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_833 <= pp_23[10]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_834 <= pp_24[8]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_835 <= pp_25[6]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_836 <= pp_26[4]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_837 <= pp_27[2]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_838 <= pp_28[0]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_839 <= pp[55]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_840 <= pp_1[55]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_841 <= pp_2[53]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_842 <= pp_3[51]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_843 <= pp_4[49]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_844 <= pp_5[47]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_845 <= pp_6[45]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_846 <= pp_7[43]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_847 <= pp_8[41]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_848 <= pp_9[39]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_849 <= pp_10[37]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_850 <= pp_11[35]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_851 <= pp_12[33]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_852 <= pp_13[31]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_853 <= pp_14[29]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_854 <= pp_15[27]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_855 <= pp_16[25]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_856 <= pp_17[23]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_857 <= pp_18[21]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_858 <= pp_19[19]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_859 <= pp_20[17]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_860 <= pp_21[15]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_861 <= pp_22[13]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_862 <= pp_23[11]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_863 <= pp_24[9]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_864 <= pp_25[7]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_865 <= pp_26[5]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_866 <= pp_27[3]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_867 <= pp_28[1]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_868 <= pp[56]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_869 <= pp_1[56]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_870 <= pp_2[54]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_871 <= pp_3[52]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_872 <= pp_4[50]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_873 <= pp_5[48]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_874 <= pp_6[46]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_875 <= pp_7[44]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_876 <= pp_8[42]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_877 <= pp_9[40]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_878 <= pp_10[38]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_879 <= pp_11[36]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_880 <= pp_12[34]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_881 <= pp_13[32]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_882 <= pp_14[30]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_883 <= pp_15[28]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_884 <= pp_16[26]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_885 <= pp_17[24]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_886 <= pp_18[22]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_887 <= pp_19[20]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_888 <= pp_20[18]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_889 <= pp_21[16]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_890 <= pp_22[14]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_891 <= pp_23[12]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_892 <= pp_24[10]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_893 <= pp_25[8]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_894 <= pp_26[6]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_895 <= pp_27[4]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_896 <= pp_28[2]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_897 <= pp_29[0]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_898 <= pp[57]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_899 <= pp_1[57]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_900 <= pp_2[55]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_901 <= pp_3[53]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_902 <= pp_4[51]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_903 <= pp_5[49]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_904 <= pp_6[47]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_905 <= pp_7[45]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_906 <= pp_8[43]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_907 <= pp_9[41]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_908 <= pp_10[39]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_909 <= pp_11[37]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_910 <= pp_12[35]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_911 <= pp_13[33]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_912 <= pp_14[31]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_913 <= pp_15[29]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_914 <= pp_16[27]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_915 <= pp_17[25]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_916 <= pp_18[23]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_917 <= pp_19[21]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_918 <= pp_20[19]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_919 <= pp_21[17]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_920 <= pp_22[15]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_921 <= pp_23[13]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_922 <= pp_24[11]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_923 <= pp_25[9]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_924 <= pp_26[7]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_925 <= pp_27[5]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_926 <= pp_28[3]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_927 <= pp_29[1]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_928 <= pp[58]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_929 <= pp_1[58]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_930 <= pp_2[56]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_931 <= pp_3[54]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_932 <= pp_4[52]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_933 <= pp_5[50]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_934 <= pp_6[48]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_935 <= pp_7[46]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_936 <= pp_8[44]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_937 <= pp_9[42]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_938 <= pp_10[40]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_939 <= pp_11[38]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_940 <= pp_12[36]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_941 <= pp_13[34]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_942 <= pp_14[32]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_943 <= pp_15[30]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_944 <= pp_16[28]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_945 <= pp_17[26]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_946 <= pp_18[24]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_947 <= pp_19[22]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_948 <= pp_20[20]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_949 <= pp_21[18]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_950 <= pp_22[16]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_951 <= pp_23[14]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_952 <= pp_24[12]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_953 <= pp_25[10]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_954 <= pp_26[8]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_955 <= pp_27[6]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_956 <= pp_28[4]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_957 <= pp_29[2]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_958 <= pp_30[0]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_959 <= pp[59]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_960 <= pp_1[59]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_961 <= pp_2[57]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_962 <= pp_3[55]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_963 <= pp_4[53]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_964 <= pp_5[51]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_965 <= pp_6[49]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_966 <= pp_7[47]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_967 <= pp_8[45]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_968 <= pp_9[43]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_969 <= pp_10[41]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_970 <= pp_11[39]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_971 <= pp_12[37]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_972 <= pp_13[35]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_973 <= pp_14[33]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_974 <= pp_15[31]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_975 <= pp_16[29]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_976 <= pp_17[27]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_977 <= pp_18[25]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_978 <= pp_19[23]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_979 <= pp_20[21]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_980 <= pp_21[19]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_981 <= pp_22[17]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_982 <= pp_23[15]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_983 <= pp_24[13]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_984 <= pp_25[11]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_985 <= pp_26[9]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_986 <= pp_27[7]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_987 <= pp_28[5]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_988 <= pp_29[3]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_989 <= pp_30[1]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_990 <= pp[60]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_991 <= pp_1[60]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_992 <= pp_2[58]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_993 <= pp_3[56]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_994 <= pp_4[54]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_995 <= pp_5[52]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_996 <= pp_6[50]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_997 <= pp_7[48]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_998 <= pp_8[46]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_999 <= pp_9[44]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1000 <= pp_10[42]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1001 <= pp_11[40]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1002 <= pp_12[38]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1003 <= pp_13[36]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1004 <= pp_14[34]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1005 <= pp_15[32]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1006 <= pp_16[30]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1007 <= pp_17[28]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1008 <= pp_18[26]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1009 <= pp_19[24]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1010 <= pp_20[22]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1011 <= pp_21[20]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1012 <= pp_22[18]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1013 <= pp_23[16]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1014 <= pp_24[14]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1015 <= pp_25[12]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1016 <= pp_26[10]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1017 <= pp_27[8]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1018 <= pp_28[6]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1019 <= pp_29[4]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1020 <= pp_30[2]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1021 <= pp_31[0]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1022 <= pp[61]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1023 <= pp_1[61]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1024 <= pp_2[59]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1025 <= pp_3[57]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1026 <= pp_4[55]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1027 <= pp_5[53]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1028 <= pp_6[51]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1029 <= pp_7[49]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1030 <= pp_8[47]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1031 <= pp_9[45]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1032 <= pp_10[43]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1033 <= pp_11[41]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1034 <= pp_12[39]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1035 <= pp_13[37]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1036 <= pp_14[35]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1037 <= pp_15[33]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1038 <= pp_16[31]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1039 <= pp_17[29]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1040 <= pp_18[27]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1041 <= pp_19[25]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1042 <= pp_20[23]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1043 <= pp_21[21]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1044 <= pp_22[19]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1045 <= pp_23[17]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1046 <= pp_24[15]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1047 <= pp_25[13]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1048 <= pp_26[11]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1049 <= pp_27[9]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1050 <= pp_28[7]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1051 <= pp_29[5]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1052 <= pp_30[3]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1053 <= pp_31[1]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1054 <= pp[62]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1055 <= pp_1[62]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1056 <= pp_2[60]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1057 <= pp_3[58]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1058 <= pp_4[56]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1059 <= pp_5[54]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1060 <= pp_6[52]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1061 <= pp_7[50]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1062 <= pp_8[48]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1063 <= pp_9[46]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1064 <= pp_10[44]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1065 <= pp_11[42]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1066 <= pp_12[40]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1067 <= pp_13[38]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1068 <= pp_14[36]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1069 <= pp_15[34]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1070 <= pp_16[32]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1071 <= pp_17[30]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1072 <= pp_18[28]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1073 <= pp_19[26]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1074 <= pp_20[24]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1075 <= pp_21[22]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1076 <= pp_22[20]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1077 <= pp_23[18]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1078 <= pp_24[16]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1079 <= pp_25[14]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1080 <= pp_26[12]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1081 <= pp_27[10]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1082 <= pp_28[8]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1083 <= pp_29[6]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1084 <= pp_30[4]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1085 <= pp_31[2]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1086 <= pp_32[0]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1087 <= pp[63]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1088 <= pp_1[63]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1089 <= pp_2[61]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1090 <= pp_3[59]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1091 <= pp_4[57]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1092 <= pp_5[55]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1093 <= pp_6[53]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1094 <= pp_7[51]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1095 <= pp_8[49]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1096 <= pp_9[47]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1097 <= pp_10[45]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1098 <= pp_11[43]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1099 <= pp_12[41]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1100 <= pp_13[39]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1101 <= pp_14[37]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1102 <= pp_15[35]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1103 <= pp_16[33]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1104 <= pp_17[31]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1105 <= pp_18[29]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1106 <= pp_19[27]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1107 <= pp_20[25]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1108 <= pp_21[23]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1109 <= pp_22[21]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1110 <= pp_23[19]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1111 <= pp_24[17]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1112 <= pp_25[15]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1113 <= pp_26[13]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1114 <= pp_27[11]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1115 <= pp_28[9]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1116 <= pp_29[7]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1117 <= pp_30[5]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1118 <= pp_31[3]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1119 <= pp_32[1]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1120 <= pp[64]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1121 <= pp_1[64]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1122 <= pp_2[62]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1123 <= pp_3[60]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1124 <= pp_4[58]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1125 <= pp_5[56]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1126 <= pp_6[54]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1127 <= pp_7[52]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1128 <= pp_8[50]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1129 <= pp_9[48]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1130 <= pp_10[46]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1131 <= pp_11[44]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1132 <= pp_12[42]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1133 <= pp_13[40]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1134 <= pp_14[38]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1135 <= pp_15[36]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1136 <= pp_16[34]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1137 <= pp_17[32]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1138 <= pp_18[30]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1139 <= pp_19[28]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1140 <= pp_20[26]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1141 <= pp_21[24]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1142 <= pp_22[22]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1143 <= pp_23[20]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1144 <= pp_24[18]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1145 <= pp_25[16]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1146 <= pp_26[14]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1147 <= pp_27[12]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1148 <= pp_28[10]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1149 <= pp_29[8]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1150 <= pp_30[6]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1151 <= pp_31[4]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1152 <= pp_32[2]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1153 <= pp[65]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1154 <= pp_1[65]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1155 <= pp_2[63]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1156 <= pp_3[61]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1157 <= pp_4[59]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1158 <= pp_5[57]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1159 <= pp_6[55]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1160 <= pp_7[53]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1161 <= pp_8[51]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1162 <= pp_9[49]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1163 <= pp_10[47]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1164 <= pp_11[45]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1165 <= pp_12[43]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1166 <= pp_13[41]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1167 <= pp_14[39]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1168 <= pp_15[37]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1169 <= pp_16[35]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1170 <= pp_17[33]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1171 <= pp_18[31]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1172 <= pp_19[29]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1173 <= pp_20[27]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1174 <= pp_21[25]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1175 <= pp_22[23]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1176 <= pp_23[21]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1177 <= pp_24[19]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1178 <= pp_25[17]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1179 <= pp_26[15]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1180 <= pp_27[13]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1181 <= pp_28[11]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1182 <= pp_29[9]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1183 <= pp_30[7]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1184 <= pp_31[5]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1185 <= pp_32[3]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1186 <= pp[66]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1187 <= pp_1[66]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1188 <= pp_2[64]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1189 <= pp_3[62]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1190 <= pp_4[60]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1191 <= pp_5[58]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1192 <= pp_6[56]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1193 <= pp_7[54]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1194 <= pp_8[52]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1195 <= pp_9[50]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1196 <= pp_10[48]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1197 <= pp_11[46]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1198 <= pp_12[44]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1199 <= pp_13[42]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1200 <= pp_14[40]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1201 <= pp_15[38]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1202 <= pp_16[36]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1203 <= pp_17[34]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1204 <= pp_18[32]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1205 <= pp_19[30]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1206 <= pp_20[28]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1207 <= pp_21[26]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1208 <= pp_22[24]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1209 <= pp_23[22]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1210 <= pp_24[20]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1211 <= pp_25[18]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1212 <= pp_26[16]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1213 <= pp_27[14]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1214 <= pp_28[12]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1215 <= pp_29[10]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1216 <= pp_30[8]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1217 <= pp_31[6]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1218 <= pp_32[4]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1219 <= pp[67]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1220 <= pp_1[67]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1221 <= pp_2[65]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1222 <= pp_3[63]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1223 <= pp_4[61]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1224 <= pp_5[59]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1225 <= pp_6[57]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1226 <= pp_7[55]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1227 <= pp_8[53]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1228 <= pp_9[51]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1229 <= pp_10[49]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1230 <= pp_11[47]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1231 <= pp_12[45]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1232 <= pp_13[43]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1233 <= pp_14[41]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1234 <= pp_15[39]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1235 <= pp_16[37]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1236 <= pp_17[35]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1237 <= pp_18[33]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1238 <= pp_19[31]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1239 <= pp_20[29]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1240 <= pp_21[27]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1241 <= pp_22[25]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1242 <= pp_23[23]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1243 <= pp_24[21]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1244 <= pp_25[19]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1245 <= pp_26[17]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1246 <= pp_27[15]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1247 <= pp_28[13]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1248 <= pp_29[11]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1249 <= pp_30[9]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1250 <= pp_31[7]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1251 <= pp_32[5]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1252 <= pp[68]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1253 <= pp_1[68]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1254 <= pp_2[66]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1255 <= pp_3[64]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1256 <= pp_4[62]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1257 <= pp_5[60]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1258 <= pp_6[58]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1259 <= pp_7[56]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1260 <= pp_8[54]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1261 <= pp_9[52]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1262 <= pp_10[50]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1263 <= pp_11[48]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1264 <= pp_12[46]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1265 <= pp_13[44]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1266 <= pp_14[42]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1267 <= pp_15[40]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1268 <= pp_16[38]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1269 <= pp_17[36]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1270 <= pp_18[34]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1271 <= pp_19[32]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1272 <= pp_20[30]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1273 <= pp_21[28]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1274 <= pp_22[26]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1275 <= pp_23[24]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1276 <= pp_24[22]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1277 <= pp_25[20]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1278 <= pp_26[18]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1279 <= pp_27[16]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1280 <= pp_28[14]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1281 <= pp_29[12]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1282 <= pp_30[10]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1283 <= pp_31[8]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1284 <= pp_32[6]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1285 <= pp_1[69]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1286 <= pp_2[67]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1287 <= pp_3[65]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1288 <= pp_4[63]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1289 <= pp_5[61]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1290 <= pp_6[59]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1291 <= pp_7[57]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1292 <= pp_8[55]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1293 <= pp_9[53]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1294 <= pp_10[51]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1295 <= pp_11[49]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1296 <= pp_12[47]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1297 <= pp_13[45]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1298 <= pp_14[43]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1299 <= pp_15[41]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1300 <= pp_16[39]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1301 <= pp_17[37]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1302 <= pp_18[35]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1303 <= pp_19[33]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1304 <= pp_20[31]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1305 <= pp_21[29]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1306 <= pp_22[27]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1307 <= pp_23[25]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1308 <= pp_24[23]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1309 <= pp_25[21]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1310 <= pp_26[19]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1311 <= pp_27[17]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1312 <= pp_28[15]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1313 <= pp_29[13]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1314 <= pp_30[11]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1315 <= pp_31[9]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1316 <= pp_32[7]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1317 <= pp_2[68]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1318 <= pp_3[66]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1319 <= pp_4[64]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1320 <= pp_5[62]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1321 <= pp_6[60]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1322 <= pp_7[58]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1323 <= pp_8[56]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1324 <= pp_9[54]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1325 <= pp_10[52]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1326 <= pp_11[50]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1327 <= pp_12[48]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1328 <= pp_13[46]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1329 <= pp_14[44]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1330 <= pp_15[42]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1331 <= pp_16[40]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1332 <= pp_17[38]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1333 <= pp_18[36]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1334 <= pp_19[34]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1335 <= pp_20[32]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1336 <= pp_21[30]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1337 <= pp_22[28]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1338 <= pp_23[26]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1339 <= pp_24[24]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1340 <= pp_25[22]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1341 <= pp_26[20]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1342 <= pp_27[18]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1343 <= pp_28[16]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1344 <= pp_29[14]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1345 <= pp_30[12]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1346 <= pp_31[10]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1347 <= pp_32[8]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1348 <= pp_2[69]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1349 <= pp_3[67]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1350 <= pp_4[65]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1351 <= pp_5[63]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1352 <= pp_6[61]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1353 <= pp_7[59]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1354 <= pp_8[57]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1355 <= pp_9[55]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1356 <= pp_10[53]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1357 <= pp_11[51]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1358 <= pp_12[49]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1359 <= pp_13[47]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1360 <= pp_14[45]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1361 <= pp_15[43]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1362 <= pp_16[41]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1363 <= pp_17[39]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1364 <= pp_18[37]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1365 <= pp_19[35]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1366 <= pp_20[33]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1367 <= pp_21[31]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1368 <= pp_22[29]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1369 <= pp_23[27]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1370 <= pp_24[25]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1371 <= pp_25[23]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1372 <= pp_26[21]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1373 <= pp_27[19]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1374 <= pp_28[17]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1375 <= pp_29[15]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1376 <= pp_30[13]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1377 <= pp_31[11]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1378 <= pp_32[9]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1379 <= pp_3[68]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1380 <= pp_4[66]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1381 <= pp_5[64]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1382 <= pp_6[62]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1383 <= pp_7[60]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1384 <= pp_8[58]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1385 <= pp_9[56]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1386 <= pp_10[54]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1387 <= pp_11[52]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1388 <= pp_12[50]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1389 <= pp_13[48]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1390 <= pp_14[46]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1391 <= pp_15[44]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1392 <= pp_16[42]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1393 <= pp_17[40]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1394 <= pp_18[38]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1395 <= pp_19[36]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1396 <= pp_20[34]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1397 <= pp_21[32]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1398 <= pp_22[30]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1399 <= pp_23[28]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1400 <= pp_24[26]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1401 <= pp_25[24]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1402 <= pp_26[22]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1403 <= pp_27[20]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1404 <= pp_28[18]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1405 <= pp_29[16]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1406 <= pp_30[14]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1407 <= pp_31[12]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1408 <= pp_32[10]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1409 <= pp_3[69]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1410 <= pp_4[67]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1411 <= pp_5[65]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1412 <= pp_6[63]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1413 <= pp_7[61]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1414 <= pp_8[59]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1415 <= pp_9[57]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1416 <= pp_10[55]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1417 <= pp_11[53]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1418 <= pp_12[51]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1419 <= pp_13[49]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1420 <= pp_14[47]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1421 <= pp_15[45]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1422 <= pp_16[43]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1423 <= pp_17[41]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1424 <= pp_18[39]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1425 <= pp_19[37]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1426 <= pp_20[35]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1427 <= pp_21[33]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1428 <= pp_22[31]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1429 <= pp_23[29]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1430 <= pp_24[27]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1431 <= pp_25[25]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1432 <= pp_26[23]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1433 <= pp_27[21]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1434 <= pp_28[19]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1435 <= pp_29[17]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1436 <= pp_30[15]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1437 <= pp_31[13]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1438 <= pp_32[11]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1439 <= pp_4[68]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1440 <= pp_5[66]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1441 <= pp_6[64]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1442 <= pp_7[62]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1443 <= pp_8[60]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1444 <= pp_9[58]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1445 <= pp_10[56]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1446 <= pp_11[54]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1447 <= pp_12[52]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1448 <= pp_13[50]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1449 <= pp_14[48]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1450 <= pp_15[46]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1451 <= pp_16[44]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1452 <= pp_17[42]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1453 <= pp_18[40]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1454 <= pp_19[38]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1455 <= pp_20[36]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1456 <= pp_21[34]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1457 <= pp_22[32]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1458 <= pp_23[30]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1459 <= pp_24[28]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1460 <= pp_25[26]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1461 <= pp_26[24]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1462 <= pp_27[22]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1463 <= pp_28[20]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1464 <= pp_29[18]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1465 <= pp_30[16]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1466 <= pp_31[14]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1467 <= pp_32[12]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1468 <= pp_4[69]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1469 <= pp_5[67]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1470 <= pp_6[65]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1471 <= pp_7[63]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1472 <= pp_8[61]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1473 <= pp_9[59]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1474 <= pp_10[57]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1475 <= pp_11[55]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1476 <= pp_12[53]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1477 <= pp_13[51]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1478 <= pp_14[49]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1479 <= pp_15[47]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1480 <= pp_16[45]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1481 <= pp_17[43]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1482 <= pp_18[41]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1483 <= pp_19[39]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1484 <= pp_20[37]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1485 <= pp_21[35]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1486 <= pp_22[33]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1487 <= pp_23[31]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1488 <= pp_24[29]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1489 <= pp_25[27]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1490 <= pp_26[25]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1491 <= pp_27[23]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1492 <= pp_28[21]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1493 <= pp_29[19]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1494 <= pp_30[17]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1495 <= pp_31[15]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1496 <= pp_32[13]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1497 <= pp_5[68]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1498 <= pp_6[66]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1499 <= pp_7[64]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1500 <= pp_8[62]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1501 <= pp_9[60]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1502 <= pp_10[58]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1503 <= pp_11[56]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1504 <= pp_12[54]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1505 <= pp_13[52]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1506 <= pp_14[50]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1507 <= pp_15[48]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1508 <= pp_16[46]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1509 <= pp_17[44]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1510 <= pp_18[42]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1511 <= pp_19[40]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1512 <= pp_20[38]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1513 <= pp_21[36]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1514 <= pp_22[34]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1515 <= pp_23[32]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1516 <= pp_24[30]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1517 <= pp_25[28]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1518 <= pp_26[26]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1519 <= pp_27[24]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1520 <= pp_28[22]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1521 <= pp_29[20]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1522 <= pp_30[18]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1523 <= pp_31[16]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1524 <= pp_32[14]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1525 <= pp_5[69]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1526 <= pp_6[67]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1527 <= pp_7[65]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1528 <= pp_8[63]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1529 <= pp_9[61]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1530 <= pp_10[59]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1531 <= pp_11[57]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1532 <= pp_12[55]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1533 <= pp_13[53]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1534 <= pp_14[51]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1535 <= pp_15[49]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1536 <= pp_16[47]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1537 <= pp_17[45]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1538 <= pp_18[43]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1539 <= pp_19[41]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1540 <= pp_20[39]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1541 <= pp_21[37]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1542 <= pp_22[35]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1543 <= pp_23[33]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1544 <= pp_24[31]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1545 <= pp_25[29]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1546 <= pp_26[27]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1547 <= pp_27[25]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1548 <= pp_28[23]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1549 <= pp_29[21]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1550 <= pp_30[19]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1551 <= pp_31[17]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1552 <= pp_32[15]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1553 <= pp_6[68]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1554 <= pp_7[66]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1555 <= pp_8[64]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1556 <= pp_9[62]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1557 <= pp_10[60]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1558 <= pp_11[58]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1559 <= pp_12[56]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1560 <= pp_13[54]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1561 <= pp_14[52]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1562 <= pp_15[50]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1563 <= pp_16[48]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1564 <= pp_17[46]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1565 <= pp_18[44]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1566 <= pp_19[42]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1567 <= pp_20[40]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1568 <= pp_21[38]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1569 <= pp_22[36]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1570 <= pp_23[34]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1571 <= pp_24[32]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1572 <= pp_25[30]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1573 <= pp_26[28]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1574 <= pp_27[26]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1575 <= pp_28[24]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1576 <= pp_29[22]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1577 <= pp_30[20]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1578 <= pp_31[18]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1579 <= pp_32[16]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1580 <= pp_6[69]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1581 <= pp_7[67]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1582 <= pp_8[65]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1583 <= pp_9[63]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1584 <= pp_10[61]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1585 <= pp_11[59]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1586 <= pp_12[57]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1587 <= pp_13[55]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1588 <= pp_14[53]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1589 <= pp_15[51]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1590 <= pp_16[49]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1591 <= pp_17[47]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1592 <= pp_18[45]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1593 <= pp_19[43]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1594 <= pp_20[41]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1595 <= pp_21[39]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1596 <= pp_22[37]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1597 <= pp_23[35]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1598 <= pp_24[33]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1599 <= pp_25[31]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1600 <= pp_26[29]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1601 <= pp_27[27]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1602 <= pp_28[25]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1603 <= pp_29[23]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1604 <= pp_30[21]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1605 <= pp_31[19]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1606 <= pp_32[17]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1607 <= pp_7[68]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1608 <= pp_8[66]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1609 <= pp_9[64]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1610 <= pp_10[62]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1611 <= pp_11[60]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1612 <= pp_12[58]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1613 <= pp_13[56]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1614 <= pp_14[54]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1615 <= pp_15[52]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1616 <= pp_16[50]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1617 <= pp_17[48]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1618 <= pp_18[46]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1619 <= pp_19[44]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1620 <= pp_20[42]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1621 <= pp_21[40]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1622 <= pp_22[38]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1623 <= pp_23[36]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1624 <= pp_24[34]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1625 <= pp_25[32]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1626 <= pp_26[30]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1627 <= pp_27[28]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1628 <= pp_28[26]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1629 <= pp_29[24]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1630 <= pp_30[22]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1631 <= pp_31[20]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1632 <= pp_32[18]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1633 <= pp_7[69]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1634 <= pp_8[67]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1635 <= pp_9[65]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1636 <= pp_10[63]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1637 <= pp_11[61]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1638 <= pp_12[59]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1639 <= pp_13[57]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1640 <= pp_14[55]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1641 <= pp_15[53]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1642 <= pp_16[51]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1643 <= pp_17[49]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1644 <= pp_18[47]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1645 <= pp_19[45]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1646 <= pp_20[43]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1647 <= pp_21[41]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1648 <= pp_22[39]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1649 <= pp_23[37]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1650 <= pp_24[35]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1651 <= pp_25[33]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1652 <= pp_26[31]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1653 <= pp_27[29]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1654 <= pp_28[27]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1655 <= pp_29[25]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1656 <= pp_30[23]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1657 <= pp_31[21]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1658 <= pp_32[19]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1659 <= pp_8[68]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1660 <= pp_9[66]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1661 <= pp_10[64]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1662 <= pp_11[62]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1663 <= pp_12[60]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1664 <= pp_13[58]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1665 <= pp_14[56]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1666 <= pp_15[54]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1667 <= pp_16[52]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1668 <= pp_17[50]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1669 <= pp_18[48]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1670 <= pp_19[46]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1671 <= pp_20[44]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1672 <= pp_21[42]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1673 <= pp_22[40]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1674 <= pp_23[38]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1675 <= pp_24[36]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1676 <= pp_25[34]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1677 <= pp_26[32]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1678 <= pp_27[30]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1679 <= pp_28[28]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1680 <= pp_29[26]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1681 <= pp_30[24]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1682 <= pp_31[22]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1683 <= pp_32[20]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1684 <= pp_8[69]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1685 <= pp_9[67]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1686 <= pp_10[65]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1687 <= pp_11[63]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1688 <= pp_12[61]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1689 <= pp_13[59]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1690 <= pp_14[57]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1691 <= pp_15[55]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1692 <= pp_16[53]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1693 <= pp_17[51]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1694 <= pp_18[49]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1695 <= pp_19[47]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1696 <= pp_20[45]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1697 <= pp_21[43]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1698 <= pp_22[41]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1699 <= pp_23[39]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1700 <= pp_24[37]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1701 <= pp_25[35]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1702 <= pp_26[33]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1703 <= pp_27[31]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1704 <= pp_28[29]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1705 <= pp_29[27]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1706 <= pp_30[25]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1707 <= pp_31[23]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1708 <= pp_32[21]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1709 <= pp_9[68]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1710 <= pp_10[66]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1711 <= pp_11[64]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1712 <= pp_12[62]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1713 <= pp_13[60]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1714 <= pp_14[58]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1715 <= pp_15[56]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1716 <= pp_16[54]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1717 <= pp_17[52]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1718 <= pp_18[50]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1719 <= pp_19[48]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1720 <= pp_20[46]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1721 <= pp_21[44]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1722 <= pp_22[42]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1723 <= pp_23[40]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1724 <= pp_24[38]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1725 <= pp_25[36]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1726 <= pp_26[34]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1727 <= pp_27[32]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1728 <= pp_28[30]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1729 <= pp_29[28]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1730 <= pp_30[26]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1731 <= pp_31[24]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1732 <= pp_32[22]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1733 <= pp_9[69]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1734 <= pp_10[67]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1735 <= pp_11[65]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1736 <= pp_12[63]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1737 <= pp_13[61]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1738 <= pp_14[59]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1739 <= pp_15[57]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1740 <= pp_16[55]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1741 <= pp_17[53]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1742 <= pp_18[51]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1743 <= pp_19[49]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1744 <= pp_20[47]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1745 <= pp_21[45]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1746 <= pp_22[43]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1747 <= pp_23[41]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1748 <= pp_24[39]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1749 <= pp_25[37]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1750 <= pp_26[35]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1751 <= pp_27[33]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1752 <= pp_28[31]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1753 <= pp_29[29]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1754 <= pp_30[27]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1755 <= pp_31[25]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1756 <= pp_32[23]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1757 <= pp_10[68]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1758 <= pp_11[66]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1759 <= pp_12[64]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1760 <= pp_13[62]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1761 <= pp_14[60]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1762 <= pp_15[58]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1763 <= pp_16[56]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1764 <= pp_17[54]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1765 <= pp_18[52]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1766 <= pp_19[50]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1767 <= pp_20[48]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1768 <= pp_21[46]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1769 <= pp_22[44]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1770 <= pp_23[42]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1771 <= pp_24[40]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1772 <= pp_25[38]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1773 <= pp_26[36]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1774 <= pp_27[34]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1775 <= pp_28[32]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1776 <= pp_29[30]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1777 <= pp_30[28]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1778 <= pp_31[26]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1779 <= pp_32[24]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1780 <= pp_10[69]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1781 <= pp_11[67]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1782 <= pp_12[65]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1783 <= pp_13[63]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1784 <= pp_14[61]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1785 <= pp_15[59]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1786 <= pp_16[57]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1787 <= pp_17[55]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1788 <= pp_18[53]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1789 <= pp_19[51]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1790 <= pp_20[49]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1791 <= pp_21[47]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1792 <= pp_22[45]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1793 <= pp_23[43]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1794 <= pp_24[41]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1795 <= pp_25[39]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1796 <= pp_26[37]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1797 <= pp_27[35]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1798 <= pp_28[33]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1799 <= pp_29[31]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1800 <= pp_30[29]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1801 <= pp_31[27]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1802 <= pp_32[25]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1803 <= pp_11[68]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1804 <= pp_12[66]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1805 <= pp_13[64]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1806 <= pp_14[62]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1807 <= pp_15[60]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1808 <= pp_16[58]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1809 <= pp_17[56]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1810 <= pp_18[54]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1811 <= pp_19[52]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1812 <= pp_20[50]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1813 <= pp_21[48]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1814 <= pp_22[46]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1815 <= pp_23[44]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1816 <= pp_24[42]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1817 <= pp_25[40]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1818 <= pp_26[38]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1819 <= pp_27[36]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1820 <= pp_28[34]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1821 <= pp_29[32]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1822 <= pp_30[30]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1823 <= pp_31[28]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1824 <= pp_32[26]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1825 <= pp_11[69]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1826 <= pp_12[67]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1827 <= pp_13[65]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1828 <= pp_14[63]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1829 <= pp_15[61]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1830 <= pp_16[59]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1831 <= pp_17[57]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1832 <= pp_18[55]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1833 <= pp_19[53]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1834 <= pp_20[51]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1835 <= pp_21[49]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1836 <= pp_22[47]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1837 <= pp_23[45]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1838 <= pp_24[43]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1839 <= pp_25[41]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1840 <= pp_26[39]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1841 <= pp_27[37]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1842 <= pp_28[35]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1843 <= pp_29[33]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1844 <= pp_30[31]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1845 <= pp_31[29]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1846 <= pp_32[27]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1847 <= pp_12[68]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1848 <= pp_13[66]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1849 <= pp_14[64]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1850 <= pp_15[62]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1851 <= pp_16[60]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1852 <= pp_17[58]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1853 <= pp_18[56]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1854 <= pp_19[54]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1855 <= pp_20[52]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1856 <= pp_21[50]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1857 <= pp_22[48]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1858 <= pp_23[46]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1859 <= pp_24[44]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1860 <= pp_25[42]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1861 <= pp_26[40]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1862 <= pp_27[38]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1863 <= pp_28[36]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1864 <= pp_29[34]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1865 <= pp_30[32]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1866 <= pp_31[30]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1867 <= pp_32[28]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1868 <= pp_12[69]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1869 <= pp_13[67]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1870 <= pp_14[65]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1871 <= pp_15[63]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1872 <= pp_16[61]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1873 <= pp_17[59]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1874 <= pp_18[57]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1875 <= pp_19[55]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1876 <= pp_20[53]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1877 <= pp_21[51]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1878 <= pp_22[49]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1879 <= pp_23[47]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1880 <= pp_24[45]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1881 <= pp_25[43]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1882 <= pp_26[41]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1883 <= pp_27[39]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1884 <= pp_28[37]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1885 <= pp_29[35]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1886 <= pp_30[33]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1887 <= pp_31[31]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1888 <= pp_32[29]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1889 <= pp_13[68]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1890 <= pp_14[66]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1891 <= pp_15[64]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1892 <= pp_16[62]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1893 <= pp_17[60]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1894 <= pp_18[58]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1895 <= pp_19[56]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1896 <= pp_20[54]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1897 <= pp_21[52]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1898 <= pp_22[50]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1899 <= pp_23[48]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1900 <= pp_24[46]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1901 <= pp_25[44]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1902 <= pp_26[42]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1903 <= pp_27[40]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1904 <= pp_28[38]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1905 <= pp_29[36]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1906 <= pp_30[34]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1907 <= pp_31[32]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1908 <= pp_32[30]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1909 <= pp_13[69]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1910 <= pp_14[67]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1911 <= pp_15[65]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1912 <= pp_16[63]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1913 <= pp_17[61]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1914 <= pp_18[59]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1915 <= pp_19[57]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1916 <= pp_20[55]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1917 <= pp_21[53]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1918 <= pp_22[51]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1919 <= pp_23[49]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1920 <= pp_24[47]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1921 <= pp_25[45]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1922 <= pp_26[43]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1923 <= pp_27[41]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1924 <= pp_28[39]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1925 <= pp_29[37]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1926 <= pp_30[35]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1927 <= pp_31[33]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1928 <= pp_32[31]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1929 <= pp_14[68]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1930 <= pp_15[66]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1931 <= pp_16[64]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1932 <= pp_17[62]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1933 <= pp_18[60]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1934 <= pp_19[58]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1935 <= pp_20[56]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1936 <= pp_21[54]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1937 <= pp_22[52]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1938 <= pp_23[50]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1939 <= pp_24[48]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1940 <= pp_25[46]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1941 <= pp_26[44]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1942 <= pp_27[42]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1943 <= pp_28[40]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1944 <= pp_29[38]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1945 <= pp_30[36]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1946 <= pp_31[34]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1947 <= pp_32[32]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1948 <= pp_14[69]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1949 <= pp_15[67]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1950 <= pp_16[65]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1951 <= pp_17[63]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1952 <= pp_18[61]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1953 <= pp_19[59]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1954 <= pp_20[57]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1955 <= pp_21[55]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1956 <= pp_22[53]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1957 <= pp_23[51]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1958 <= pp_24[49]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1959 <= pp_25[47]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1960 <= pp_26[45]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1961 <= pp_27[43]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1962 <= pp_28[41]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1963 <= pp_29[39]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1964 <= pp_30[37]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1965 <= pp_31[35]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1966 <= pp_32[33]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1967 <= pp_15[68]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1968 <= pp_16[66]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1969 <= pp_17[64]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1970 <= pp_18[62]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1971 <= pp_19[60]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1972 <= pp_20[58]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1973 <= pp_21[56]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1974 <= pp_22[54]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1975 <= pp_23[52]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1976 <= pp_24[50]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1977 <= pp_25[48]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1978 <= pp_26[46]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1979 <= pp_27[44]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1980 <= pp_28[42]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1981 <= pp_29[40]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1982 <= pp_30[38]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1983 <= pp_31[36]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1984 <= pp_32[34]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1985 <= pp_15[69]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1986 <= pp_16[67]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1987 <= pp_17[65]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1988 <= pp_18[63]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1989 <= pp_19[61]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1990 <= pp_20[59]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1991 <= pp_21[57]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1992 <= pp_22[55]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1993 <= pp_23[53]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1994 <= pp_24[51]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1995 <= pp_25[49]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1996 <= pp_26[47]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1997 <= pp_27[45]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1998 <= pp_28[43]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1999 <= pp_29[41]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2000 <= pp_30[39]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2001 <= pp_31[37]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2002 <= pp_32[35]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2003 <= pp_16[68]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2004 <= pp_17[66]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2005 <= pp_18[64]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2006 <= pp_19[62]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2007 <= pp_20[60]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2008 <= pp_21[58]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2009 <= pp_22[56]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2010 <= pp_23[54]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2011 <= pp_24[52]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2012 <= pp_25[50]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2013 <= pp_26[48]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2014 <= pp_27[46]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2015 <= pp_28[44]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2016 <= pp_29[42]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2017 <= pp_30[40]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2018 <= pp_31[38]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2019 <= pp_32[36]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2020 <= pp_16[69]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2021 <= pp_17[67]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2022 <= pp_18[65]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2023 <= pp_19[63]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2024 <= pp_20[61]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2025 <= pp_21[59]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2026 <= pp_22[57]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2027 <= pp_23[55]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2028 <= pp_24[53]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2029 <= pp_25[51]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2030 <= pp_26[49]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2031 <= pp_27[47]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2032 <= pp_28[45]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2033 <= pp_29[43]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2034 <= pp_30[41]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2035 <= pp_31[39]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2036 <= pp_32[37]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2037 <= pp_17[68]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2038 <= pp_18[66]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2039 <= pp_19[64]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2040 <= pp_20[62]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2041 <= pp_21[60]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2042 <= pp_22[58]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2043 <= pp_23[56]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2044 <= pp_24[54]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2045 <= pp_25[52]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2046 <= pp_26[50]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2047 <= pp_27[48]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2048 <= pp_28[46]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2049 <= pp_29[44]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2050 <= pp_30[42]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2051 <= pp_31[40]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2052 <= pp_32[38]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2053 <= pp_17[69]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2054 <= pp_18[67]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2055 <= pp_19[65]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2056 <= pp_20[63]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2057 <= pp_21[61]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2058 <= pp_22[59]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2059 <= pp_23[57]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2060 <= pp_24[55]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2061 <= pp_25[53]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2062 <= pp_26[51]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2063 <= pp_27[49]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2064 <= pp_28[47]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2065 <= pp_29[45]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2066 <= pp_30[43]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2067 <= pp_31[41]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2068 <= pp_32[39]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2069 <= pp_18[68]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2070 <= pp_19[66]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2071 <= pp_20[64]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2072 <= pp_21[62]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2073 <= pp_22[60]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2074 <= pp_23[58]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2075 <= pp_24[56]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2076 <= pp_25[54]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2077 <= pp_26[52]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2078 <= pp_27[50]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2079 <= pp_28[48]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2080 <= pp_29[46]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2081 <= pp_30[44]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2082 <= pp_31[42]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2083 <= pp_32[40]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2084 <= pp_18[69]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2085 <= pp_19[67]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2086 <= pp_20[65]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2087 <= pp_21[63]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2088 <= pp_22[61]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2089 <= pp_23[59]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2090 <= pp_24[57]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2091 <= pp_25[55]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2092 <= pp_26[53]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2093 <= pp_27[51]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2094 <= pp_28[49]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2095 <= pp_29[47]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2096 <= pp_30[45]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2097 <= pp_31[43]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2098 <= pp_32[41]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2099 <= pp_19[68]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2100 <= pp_20[66]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2101 <= pp_21[64]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2102 <= pp_22[62]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2103 <= pp_23[60]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2104 <= pp_24[58]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2105 <= pp_25[56]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2106 <= pp_26[54]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2107 <= pp_27[52]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2108 <= pp_28[50]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2109 <= pp_29[48]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2110 <= pp_30[46]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2111 <= pp_31[44]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2112 <= pp_32[42]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2113 <= pp_19[69]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2114 <= pp_20[67]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2115 <= pp_21[65]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2116 <= pp_22[63]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2117 <= pp_23[61]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2118 <= pp_24[59]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2119 <= pp_25[57]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2120 <= pp_26[55]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2121 <= pp_27[53]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2122 <= pp_28[51]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2123 <= pp_29[49]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2124 <= pp_30[47]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2125 <= pp_31[45]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2126 <= pp_32[43]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2127 <= pp_20[68]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2128 <= pp_21[66]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2129 <= pp_22[64]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2130 <= pp_23[62]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2131 <= pp_24[60]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2132 <= pp_25[58]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2133 <= pp_26[56]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2134 <= pp_27[54]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2135 <= pp_28[52]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2136 <= pp_29[50]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2137 <= pp_30[48]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2138 <= pp_31[46]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2139 <= pp_32[44]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2140 <= pp_20[69]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2141 <= pp_21[67]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2142 <= pp_22[65]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2143 <= pp_23[63]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2144 <= pp_24[61]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2145 <= pp_25[59]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2146 <= pp_26[57]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2147 <= pp_27[55]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2148 <= pp_28[53]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2149 <= pp_29[51]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2150 <= pp_30[49]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2151 <= pp_31[47]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2152 <= pp_32[45]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2153 <= pp_21[68]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2154 <= pp_22[66]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2155 <= pp_23[64]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2156 <= pp_24[62]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2157 <= pp_25[60]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2158 <= pp_26[58]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2159 <= pp_27[56]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2160 <= pp_28[54]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2161 <= pp_29[52]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2162 <= pp_30[50]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2163 <= pp_31[48]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2164 <= pp_32[46]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2165 <= pp_21[69]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2166 <= pp_22[67]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2167 <= pp_23[65]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2168 <= pp_24[63]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2169 <= pp_25[61]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2170 <= pp_26[59]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2171 <= pp_27[57]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2172 <= pp_28[55]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2173 <= pp_29[53]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2174 <= pp_30[51]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2175 <= pp_31[49]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2176 <= pp_32[47]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2177 <= pp_22[68]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2178 <= pp_23[66]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2179 <= pp_24[64]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2180 <= pp_25[62]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2181 <= pp_26[60]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2182 <= pp_27[58]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2183 <= pp_28[56]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2184 <= pp_29[54]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2185 <= pp_30[52]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2186 <= pp_31[50]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2187 <= pp_32[48]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2188 <= pp_22[69]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2189 <= pp_23[67]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2190 <= pp_24[65]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2191 <= pp_25[63]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2192 <= pp_26[61]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2193 <= pp_27[59]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2194 <= pp_28[57]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2195 <= pp_29[55]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2196 <= pp_30[53]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2197 <= pp_31[51]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2198 <= pp_32[49]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2199 <= pp_23[68]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2200 <= pp_24[66]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2201 <= pp_25[64]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2202 <= pp_26[62]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2203 <= pp_27[60]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2204 <= pp_28[58]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2205 <= pp_29[56]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2206 <= pp_30[54]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2207 <= pp_31[52]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2208 <= pp_32[50]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2209 <= pp_23[69]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2210 <= pp_24[67]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2211 <= pp_25[65]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2212 <= pp_26[63]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2213 <= pp_27[61]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2214 <= pp_28[59]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2215 <= pp_29[57]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2216 <= pp_30[55]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2217 <= pp_31[53]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2218 <= pp_32[51]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2219 <= pp_24[68]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2220 <= pp_25[66]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2221 <= pp_26[64]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2222 <= pp_27[62]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2223 <= pp_28[60]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2224 <= pp_29[58]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2225 <= pp_30[56]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2226 <= pp_31[54]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2227 <= pp_32[52]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2228 <= pp_24[69]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2229 <= pp_25[67]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2230 <= pp_26[65]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2231 <= pp_27[63]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2232 <= pp_28[61]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2233 <= pp_29[59]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2234 <= pp_30[57]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2235 <= pp_31[55]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2236 <= pp_32[53]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2237 <= pp_25[68]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2238 <= pp_26[66]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2239 <= pp_27[64]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2240 <= pp_28[62]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2241 <= pp_29[60]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2242 <= pp_30[58]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2243 <= pp_31[56]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2244 <= pp_32[54]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2245 <= pp_25[69]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2246 <= pp_26[67]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2247 <= pp_27[65]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2248 <= pp_28[63]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2249 <= pp_29[61]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2250 <= pp_30[59]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2251 <= pp_31[57]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2252 <= pp_32[55]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2253 <= pp_26[68]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2254 <= pp_27[66]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2255 <= pp_28[64]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2256 <= pp_29[62]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2257 <= pp_30[60]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2258 <= pp_31[58]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2259 <= pp_32[56]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2260 <= pp_26[69]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2261 <= pp_27[67]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2262 <= pp_28[65]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2263 <= pp_29[63]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2264 <= pp_30[61]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2265 <= pp_31[59]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2266 <= pp_32[57]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2267 <= pp_27[68]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2268 <= pp_28[66]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2269 <= pp_29[64]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2270 <= pp_30[62]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2271 <= pp_31[60]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2272 <= pp_32[58]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2273 <= pp_27[69]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2274 <= pp_28[67]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2275 <= pp_29[65]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2276 <= pp_30[63]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2277 <= pp_31[61]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2278 <= pp_32[59]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2279 <= pp_28[68]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2280 <= pp_29[66]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2281 <= pp_30[64]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2282 <= pp_31[62]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2283 <= pp_32[60]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2284 <= pp_28[69]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2285 <= pp_29[67]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2286 <= pp_30[65]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2287 <= pp_31[63]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2288 <= pp_32[61]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2289 <= pp_29[68]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2290 <= pp_30[66]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2291 <= pp_31[64]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2292 <= pp_32[62]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2293 <= pp_29[69]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2294 <= pp_30[67]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2295 <= pp_31[65]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2296 <= pp_32[63]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2297 <= pp_30[68]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2298 <= pp_31[66]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2299 <= pp_32[64]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2300 <= pp_30[69]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2301 <= pp_31[67]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2302 <= pp_32[65]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2303 <= pp_31[68]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2304 <= pp_32[66]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2305 <= pp_31[69]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2306 <= pp_32[67]; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2307 <= s_0; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2308 <= s_0_130; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2309 <= s_0_259; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2310 <= s_0_387; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2311 <= s_0_514; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2312 <= s_0_515; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2313 <= c2_0_514; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2314 <= s_0_516; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2315 <= c2_0_515; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2316 <= s_0_517; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2317 <= c2_0_516; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2318 <= s_0_518; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2319 <= c2_0_517; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2320 <= s_0_519; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2321 <= c2_0_518; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2322 <= s_0_520; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2323 <= c2_0_519; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2324 <= s_0_521; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2325 <= c2_0_520; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2326 <= s_0_522; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2327 <= c2_0_521; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2328 <= s_0_523; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2329 <= c2_0_522; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2330 <= s_0_524; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2331 <= c2_0_523; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2332 <= s_0_525; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2333 <= c2_0_524; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2334 <= s_0_526; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2335 <= c2_0_525; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2336 <= s_0_527; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2337 <= c2_0_526; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2338 <= s_0_528; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2339 <= c2_0_527; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2340 <= s_0_529; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2341 <= c2_0_528; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2342 <= s_0_530; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2343 <= c2_0_529; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2344 <= s_0_531; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2345 <= c2_0_530; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2346 <= s_0_532; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2347 <= c2_0_531; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2348 <= s_0_533; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2349 <= c2_0_532; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2350 <= s_0_534; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2351 <= c2_0_533; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2352 <= s_0_535; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2353 <= c2_0_534; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2354 <= s_0_536; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2355 <= c2_0_535; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2356 <= s_0_537; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2357 <= c2_0_536; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2358 <= s_0_538; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2359 <= c2_0_537; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2360 <= s_0_539; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2361 <= c2_0_538; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2362 <= s_0_540; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2363 <= c2_0_539; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2364 <= s_0_541; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2365 <= c2_0_540; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2366 <= s_0_542; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2367 <= c2_0_541; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2368 <= s_0_543; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2369 <= c2_0_542; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2370 <= s_0_544; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2371 <= c2_0_543; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2372 <= s_0_545; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2373 <= c2_0_544; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2374 <= s_0_546; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2375 <= c2_0_545; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2376 <= s_0_547; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2377 <= c2_0_546; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2378 <= s_0_548; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2379 <= c2_0_547; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2380 <= s_0_549; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2381 <= c2_0_548; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2382 <= s_0_550; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2383 <= c2_0_549; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2384 <= s_0_551; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2385 <= c2_0_550; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2386 <= s_0_552; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2387 <= c2_0_551; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2388 <= s_0_553; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2389 <= c2_0_552; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2390 <= s_0_554; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2391 <= c2_0_553; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2392 <= s_0_555; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2393 <= c2_0_554; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2394 <= s_0_556; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2395 <= c2_0_555; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2396 <= s_0_557; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2397 <= c2_0_556; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2398 <= s_0_558; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2399 <= c2_0_557; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2400 <= s_0_559; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2401 <= c2_0_558; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2402 <= s_0_560; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2403 <= c2_0_559; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2404 <= s_0_561; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2405 <= c2_0_560; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2406 <= s_0_562; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2407 <= c2_0_561; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2408 <= s_0_563; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2409 <= c2_0_562; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2410 <= s_0_564; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2411 <= c2_0_563; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2412 <= s_0_565; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2413 <= c2_0_564; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2414 <= s_0_566; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2415 <= c2_0_565; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2416 <= s_0_567; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2417 <= c2_0_566; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2418 <= s_0_568; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2419 <= c2_0_567; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2420 <= s_0_569; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2421 <= c2_0_568; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2422 <= s_0_570; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2423 <= c2_0_569; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2424 <= s_0_571; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2425 <= c2_0_570; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2426 <= s_0_572; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2427 <= c2_0_571; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2428 <= s_0_573; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2429 <= c2_0_572; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2430 <= s_0_574; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2431 <= c2_0_573; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2432 <= s_0_575; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2433 <= c2_0_574; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2434 <= s_0_576; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2435 <= c2_0_575; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2436 <= s_0_577; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2437 <= c2_0_576; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2438 <= s_0_578; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2439 <= c2_0_577; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2440 <= s_0_579; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2441 <= c2_0_578; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2442 <= s_0_580; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2443 <= c2_0_579; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2444 <= s_0_581; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2445 <= c2_0_580; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2446 <= s_0_582; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2447 <= c2_0_581; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2448 <= s_0_583; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2449 <= c2_0_582; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2450 <= s_0_584; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2451 <= c2_0_583; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2452 <= s_0_585; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2453 <= c2_0_584; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2454 <= s_0_586; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2455 <= c2_0_585; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2456 <= s_0_587; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2457 <= c2_0_586; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2458 <= s_0_588; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2459 <= c2_0_587; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2460 <= s_0_589; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2461 <= c2_0_588; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2462 <= s_0_590; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2463 <= c2_0_589; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2464 <= s_0_591; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2465 <= c2_0_590; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2466 <= s_0_592; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2467 <= c2_0_591; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2468 <= s_0_593; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2469 <= c2_0_592; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2470 <= s_0_594; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2471 <= c2_0_593; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2472 <= s_0_595; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2473 <= c2_0_594; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2474 <= s_0_596; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2475 <= c2_0_595; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2476 <= s_0_597; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2477 <= c2_0_596; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2478 <= s_0_598; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2479 <= c2_0_597; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2480 <= s_0_599; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2481 <= c2_0_598; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2482 <= s_0_600; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2483 <= c2_0_599; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2484 <= s_0_601; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2485 <= c2_0_600; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2486 <= s_0_602; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2487 <= c2_0_601; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2488 <= s_0_603; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2489 <= c2_0_602; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2490 <= s_0_604; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2491 <= c2_0_603; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2492 <= s_0_605; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2493 <= c2_0_604; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2494 <= s_0_606; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2495 <= c2_0_605; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2496 <= s_0_607; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2497 <= c2_0_606; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2498 <= s_0_608; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2499 <= c2_0_607; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2500 <= s_0_609; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2501 <= c2_0_608; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2502 <= s_0_610; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2503 <= c2_0_609; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2504 <= s_0_611; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2505 <= c2_0_610; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2506 <= s_0_612; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2507 <= c2_0_611; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2508 <= s_0_613; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2509 <= c2_0_612; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2510 <= s_0_614; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2511 <= c2_0_613; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2512 <= s_0_615; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2513 <= c2_0_614; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2514 <= s_0_616; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2515 <= c2_0_615; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2516 <= s_0_617; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2517 <= c2_0_616; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2518 <= s_0_618; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2519 <= c2_0_617; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2520 <= s_0_619; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2521 <= c2_0_618; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2522 <= s_0_620; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2523 <= c2_0_619; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2524 <= s_0_621; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2525 <= c2_0_620; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2526 <= s_0_622; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2527 <= c2_0_621; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2528 <= s_0_623; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2529 <= c2_0_622; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2530 <= s_0_624; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2531 <= c2_0_623; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2532 <= s_0_625; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2533 <= c2_0_624; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2534 <= s_0_626; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2535 <= c2_0_625; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2536 <= s_0_627; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2537 <= c2_0_626; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2538 <= s_0_628; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2539 <= c2_0_627; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2540 <= s_0_629; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2541 <= c2_0_628; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2542 <= s_0_630; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2543 <= c2_0_629; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2544 <= s_0_631; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2545 <= c2_0_630; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2546 <= s_0_632; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2547 <= c2_0_631; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2548 <= s_0_633; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2549 <= c2_0_632; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2550 <= s_0_634; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2551 <= c2_0_633; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2552 <= s_0_635; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2553 <= c2_0_634; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2554 <= s_0_636; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2555 <= c2_0_635; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2556 <= s_0_637; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2557 <= c2_0_636; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2558 <= s_0_638; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2559 <= c2_0_637; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2560 <= s_0_639; // @[Reg.scala 17:22]
    end
    if (io_regEnables_1) begin // @[Reg.scala 17:18]
      r_2561 <= c2_0_638; // @[Reg.scala 17:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  r_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  r_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  r_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  r_4 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  r_5 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  r_6 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  r_7 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  r_8 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  r_9 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  r_10 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  r_11 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  r_12 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  r_13 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  r_14 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  r_15 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  r_16 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  r_17 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  r_18 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  r_19 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  r_20 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  r_21 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  r_22 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  r_23 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  r_24 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  r_25 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  r_26 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  r_27 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  r_28 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  r_29 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  r_30 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  r_31 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  r_32 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  r_33 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  r_34 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  r_35 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  r_36 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  r_37 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  r_38 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  r_39 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  r_40 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  r_41 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  r_42 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  r_43 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  r_44 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  r_45 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  r_46 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  r_47 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  r_48 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  r_49 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  r_50 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  r_51 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  r_52 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  r_53 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  r_54 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  r_55 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  r_56 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  r_57 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  r_58 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  r_59 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  r_60 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  r_61 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  r_62 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  r_63 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  r_64 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  r_65 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  r_66 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  r_67 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  r_68 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  r_69 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  r_70 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  r_71 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  r_72 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  r_73 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  r_74 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  r_75 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  r_76 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  r_77 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  r_78 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  r_79 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  r_80 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  r_81 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  r_82 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  r_83 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  r_84 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  r_85 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  r_86 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  r_87 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  r_88 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  r_89 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  r_90 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  r_91 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  r_92 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  r_93 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  r_94 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  r_95 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  r_96 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  r_97 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  r_98 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  r_99 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  r_100 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  r_101 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  r_102 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  r_103 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  r_104 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  r_105 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  r_106 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  r_107 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  r_108 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  r_109 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  r_110 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  r_111 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  r_112 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  r_113 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  r_114 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  r_115 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  r_116 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  r_117 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  r_118 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  r_119 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  r_120 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  r_121 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  r_122 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  r_123 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  r_124 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  r_125 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  r_126 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  r_127 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  r_128 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  r_129 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  r_130 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  r_131 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  r_132 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  r_133 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  r_134 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  r_135 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  r_136 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  r_137 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  r_138 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  r_139 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  r_140 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  r_141 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  r_142 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  r_143 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  r_144 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  r_145 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  r_146 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  r_147 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  r_148 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  r_149 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  r_150 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  r_151 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  r_152 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  r_153 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  r_154 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  r_155 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  r_156 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  r_157 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  r_158 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  r_159 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  r_160 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  r_161 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  r_162 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  r_163 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  r_164 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  r_165 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  r_166 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  r_167 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  r_168 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  r_169 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  r_170 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  r_171 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  r_172 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  r_173 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  r_174 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  r_175 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  r_176 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  r_177 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  r_178 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  r_179 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  r_180 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  r_181 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  r_182 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  r_183 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  r_184 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  r_185 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  r_186 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  r_187 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  r_188 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  r_189 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  r_190 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  r_191 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  r_192 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  r_193 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  r_194 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  r_195 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  r_196 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  r_197 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  r_198 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  r_199 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  r_200 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  r_201 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  r_202 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  r_203 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  r_204 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  r_205 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  r_206 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  r_207 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  r_208 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  r_209 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  r_210 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  r_211 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  r_212 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  r_213 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  r_214 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  r_215 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  r_216 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  r_217 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  r_218 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  r_219 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  r_220 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  r_221 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  r_222 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  r_223 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  r_224 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  r_225 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  r_226 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  r_227 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  r_228 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  r_229 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  r_230 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  r_231 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  r_232 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  r_233 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  r_234 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  r_235 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  r_236 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  r_237 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  r_238 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  r_239 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  r_240 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  r_241 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  r_242 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  r_243 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  r_244 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  r_245 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  r_246 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  r_247 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  r_248 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  r_249 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  r_250 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  r_251 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  r_252 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  r_253 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  r_254 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  r_255 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  r_256 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  r_257 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  r_258 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  r_259 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  r_260 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  r_261 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  r_262 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  r_263 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  r_264 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  r_265 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  r_266 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  r_267 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  r_268 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  r_269 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  r_270 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  r_271 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  r_272 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  r_273 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  r_274 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  r_275 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  r_276 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  r_277 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  r_278 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  r_279 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  r_280 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  r_281 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  r_282 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  r_283 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  r_284 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  r_285 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  r_286 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  r_287 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  r_288 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  r_289 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  r_290 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  r_291 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  r_292 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  r_293 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  r_294 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  r_295 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  r_296 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  r_297 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  r_298 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  r_299 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  r_300 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  r_301 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  r_302 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  r_303 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  r_304 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  r_305 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  r_306 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  r_307 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  r_308 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  r_309 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  r_310 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  r_311 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  r_312 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  r_313 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  r_314 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  r_315 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  r_316 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  r_317 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  r_318 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  r_319 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  r_320 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  r_321 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  r_322 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  r_323 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  r_324 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  r_325 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  r_326 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  r_327 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  r_328 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  r_329 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  r_330 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  r_331 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  r_332 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  r_333 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  r_334 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  r_335 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  r_336 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  r_337 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  r_338 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  r_339 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  r_340 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  r_341 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  r_342 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  r_343 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  r_344 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  r_345 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  r_346 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  r_347 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  r_348 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  r_349 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  r_350 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  r_351 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  r_352 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  r_353 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  r_354 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  r_355 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  r_356 = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  r_357 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  r_358 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  r_359 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  r_360 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  r_361 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  r_362 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  r_363 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  r_364 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  r_365 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  r_366 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  r_367 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  r_368 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  r_369 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  r_370 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  r_371 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  r_372 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  r_373 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  r_374 = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  r_375 = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  r_376 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  r_377 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  r_378 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  r_379 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  r_380 = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  r_381 = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  r_382 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  r_383 = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  r_384 = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  r_385 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  r_386 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  r_387 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  r_388 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  r_389 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  r_390 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  r_391 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  r_392 = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  r_393 = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  r_394 = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  r_395 = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  r_396 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  r_397 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  r_398 = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  r_399 = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  r_400 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  r_401 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  r_402 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  r_403 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  r_404 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  r_405 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  r_406 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  r_407 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  r_408 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  r_409 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  r_410 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  r_411 = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  r_412 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  r_413 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  r_414 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  r_415 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  r_416 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  r_417 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  r_418 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  r_419 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  r_420 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  r_421 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  r_422 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  r_423 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  r_424 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  r_425 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  r_426 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  r_427 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  r_428 = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  r_429 = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  r_430 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  r_431 = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  r_432 = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  r_433 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  r_434 = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  r_435 = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  r_436 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  r_437 = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  r_438 = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  r_439 = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  r_440 = _RAND_440[0:0];
  _RAND_441 = {1{`RANDOM}};
  r_441 = _RAND_441[0:0];
  _RAND_442 = {1{`RANDOM}};
  r_442 = _RAND_442[0:0];
  _RAND_443 = {1{`RANDOM}};
  r_443 = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  r_444 = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  r_445 = _RAND_445[0:0];
  _RAND_446 = {1{`RANDOM}};
  r_446 = _RAND_446[0:0];
  _RAND_447 = {1{`RANDOM}};
  r_447 = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  r_448 = _RAND_448[0:0];
  _RAND_449 = {1{`RANDOM}};
  r_449 = _RAND_449[0:0];
  _RAND_450 = {1{`RANDOM}};
  r_450 = _RAND_450[0:0];
  _RAND_451 = {1{`RANDOM}};
  r_451 = _RAND_451[0:0];
  _RAND_452 = {1{`RANDOM}};
  r_452 = _RAND_452[0:0];
  _RAND_453 = {1{`RANDOM}};
  r_453 = _RAND_453[0:0];
  _RAND_454 = {1{`RANDOM}};
  r_454 = _RAND_454[0:0];
  _RAND_455 = {1{`RANDOM}};
  r_455 = _RAND_455[0:0];
  _RAND_456 = {1{`RANDOM}};
  r_456 = _RAND_456[0:0];
  _RAND_457 = {1{`RANDOM}};
  r_457 = _RAND_457[0:0];
  _RAND_458 = {1{`RANDOM}};
  r_458 = _RAND_458[0:0];
  _RAND_459 = {1{`RANDOM}};
  r_459 = _RAND_459[0:0];
  _RAND_460 = {1{`RANDOM}};
  r_460 = _RAND_460[0:0];
  _RAND_461 = {1{`RANDOM}};
  r_461 = _RAND_461[0:0];
  _RAND_462 = {1{`RANDOM}};
  r_462 = _RAND_462[0:0];
  _RAND_463 = {1{`RANDOM}};
  r_463 = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  r_464 = _RAND_464[0:0];
  _RAND_465 = {1{`RANDOM}};
  r_465 = _RAND_465[0:0];
  _RAND_466 = {1{`RANDOM}};
  r_466 = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  r_467 = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  r_468 = _RAND_468[0:0];
  _RAND_469 = {1{`RANDOM}};
  r_469 = _RAND_469[0:0];
  _RAND_470 = {1{`RANDOM}};
  r_470 = _RAND_470[0:0];
  _RAND_471 = {1{`RANDOM}};
  r_471 = _RAND_471[0:0];
  _RAND_472 = {1{`RANDOM}};
  r_472 = _RAND_472[0:0];
  _RAND_473 = {1{`RANDOM}};
  r_473 = _RAND_473[0:0];
  _RAND_474 = {1{`RANDOM}};
  r_474 = _RAND_474[0:0];
  _RAND_475 = {1{`RANDOM}};
  r_475 = _RAND_475[0:0];
  _RAND_476 = {1{`RANDOM}};
  r_476 = _RAND_476[0:0];
  _RAND_477 = {1{`RANDOM}};
  r_477 = _RAND_477[0:0];
  _RAND_478 = {1{`RANDOM}};
  r_478 = _RAND_478[0:0];
  _RAND_479 = {1{`RANDOM}};
  r_479 = _RAND_479[0:0];
  _RAND_480 = {1{`RANDOM}};
  r_480 = _RAND_480[0:0];
  _RAND_481 = {1{`RANDOM}};
  r_481 = _RAND_481[0:0];
  _RAND_482 = {1{`RANDOM}};
  r_482 = _RAND_482[0:0];
  _RAND_483 = {1{`RANDOM}};
  r_483 = _RAND_483[0:0];
  _RAND_484 = {1{`RANDOM}};
  r_484 = _RAND_484[0:0];
  _RAND_485 = {1{`RANDOM}};
  r_485 = _RAND_485[0:0];
  _RAND_486 = {1{`RANDOM}};
  r_486 = _RAND_486[0:0];
  _RAND_487 = {1{`RANDOM}};
  r_487 = _RAND_487[0:0];
  _RAND_488 = {1{`RANDOM}};
  r_488 = _RAND_488[0:0];
  _RAND_489 = {1{`RANDOM}};
  r_489 = _RAND_489[0:0];
  _RAND_490 = {1{`RANDOM}};
  r_490 = _RAND_490[0:0];
  _RAND_491 = {1{`RANDOM}};
  r_491 = _RAND_491[0:0];
  _RAND_492 = {1{`RANDOM}};
  r_492 = _RAND_492[0:0];
  _RAND_493 = {1{`RANDOM}};
  r_493 = _RAND_493[0:0];
  _RAND_494 = {1{`RANDOM}};
  r_494 = _RAND_494[0:0];
  _RAND_495 = {1{`RANDOM}};
  r_495 = _RAND_495[0:0];
  _RAND_496 = {1{`RANDOM}};
  r_496 = _RAND_496[0:0];
  _RAND_497 = {1{`RANDOM}};
  r_497 = _RAND_497[0:0];
  _RAND_498 = {1{`RANDOM}};
  r_498 = _RAND_498[0:0];
  _RAND_499 = {1{`RANDOM}};
  r_499 = _RAND_499[0:0];
  _RAND_500 = {1{`RANDOM}};
  r_500 = _RAND_500[0:0];
  _RAND_501 = {1{`RANDOM}};
  r_501 = _RAND_501[0:0];
  _RAND_502 = {1{`RANDOM}};
  r_502 = _RAND_502[0:0];
  _RAND_503 = {1{`RANDOM}};
  r_503 = _RAND_503[0:0];
  _RAND_504 = {1{`RANDOM}};
  r_504 = _RAND_504[0:0];
  _RAND_505 = {1{`RANDOM}};
  r_505 = _RAND_505[0:0];
  _RAND_506 = {1{`RANDOM}};
  r_506 = _RAND_506[0:0];
  _RAND_507 = {1{`RANDOM}};
  r_507 = _RAND_507[0:0];
  _RAND_508 = {1{`RANDOM}};
  r_508 = _RAND_508[0:0];
  _RAND_509 = {1{`RANDOM}};
  r_509 = _RAND_509[0:0];
  _RAND_510 = {1{`RANDOM}};
  r_510 = _RAND_510[0:0];
  _RAND_511 = {1{`RANDOM}};
  r_511 = _RAND_511[0:0];
  _RAND_512 = {1{`RANDOM}};
  r_512 = _RAND_512[0:0];
  _RAND_513 = {1{`RANDOM}};
  r_513 = _RAND_513[0:0];
  _RAND_514 = {1{`RANDOM}};
  r_514 = _RAND_514[0:0];
  _RAND_515 = {1{`RANDOM}};
  r_515 = _RAND_515[0:0];
  _RAND_516 = {1{`RANDOM}};
  r_516 = _RAND_516[0:0];
  _RAND_517 = {1{`RANDOM}};
  r_517 = _RAND_517[0:0];
  _RAND_518 = {1{`RANDOM}};
  r_518 = _RAND_518[0:0];
  _RAND_519 = {1{`RANDOM}};
  r_519 = _RAND_519[0:0];
  _RAND_520 = {1{`RANDOM}};
  r_520 = _RAND_520[0:0];
  _RAND_521 = {1{`RANDOM}};
  r_521 = _RAND_521[0:0];
  _RAND_522 = {1{`RANDOM}};
  r_522 = _RAND_522[0:0];
  _RAND_523 = {1{`RANDOM}};
  r_523 = _RAND_523[0:0];
  _RAND_524 = {1{`RANDOM}};
  r_524 = _RAND_524[0:0];
  _RAND_525 = {1{`RANDOM}};
  r_525 = _RAND_525[0:0];
  _RAND_526 = {1{`RANDOM}};
  r_526 = _RAND_526[0:0];
  _RAND_527 = {1{`RANDOM}};
  r_527 = _RAND_527[0:0];
  _RAND_528 = {1{`RANDOM}};
  r_528 = _RAND_528[0:0];
  _RAND_529 = {1{`RANDOM}};
  r_529 = _RAND_529[0:0];
  _RAND_530 = {1{`RANDOM}};
  r_530 = _RAND_530[0:0];
  _RAND_531 = {1{`RANDOM}};
  r_531 = _RAND_531[0:0];
  _RAND_532 = {1{`RANDOM}};
  r_532 = _RAND_532[0:0];
  _RAND_533 = {1{`RANDOM}};
  r_533 = _RAND_533[0:0];
  _RAND_534 = {1{`RANDOM}};
  r_534 = _RAND_534[0:0];
  _RAND_535 = {1{`RANDOM}};
  r_535 = _RAND_535[0:0];
  _RAND_536 = {1{`RANDOM}};
  r_536 = _RAND_536[0:0];
  _RAND_537 = {1{`RANDOM}};
  r_537 = _RAND_537[0:0];
  _RAND_538 = {1{`RANDOM}};
  r_538 = _RAND_538[0:0];
  _RAND_539 = {1{`RANDOM}};
  r_539 = _RAND_539[0:0];
  _RAND_540 = {1{`RANDOM}};
  r_540 = _RAND_540[0:0];
  _RAND_541 = {1{`RANDOM}};
  r_541 = _RAND_541[0:0];
  _RAND_542 = {1{`RANDOM}};
  r_542 = _RAND_542[0:0];
  _RAND_543 = {1{`RANDOM}};
  r_543 = _RAND_543[0:0];
  _RAND_544 = {1{`RANDOM}};
  r_544 = _RAND_544[0:0];
  _RAND_545 = {1{`RANDOM}};
  r_545 = _RAND_545[0:0];
  _RAND_546 = {1{`RANDOM}};
  r_546 = _RAND_546[0:0];
  _RAND_547 = {1{`RANDOM}};
  r_547 = _RAND_547[0:0];
  _RAND_548 = {1{`RANDOM}};
  r_548 = _RAND_548[0:0];
  _RAND_549 = {1{`RANDOM}};
  r_549 = _RAND_549[0:0];
  _RAND_550 = {1{`RANDOM}};
  r_550 = _RAND_550[0:0];
  _RAND_551 = {1{`RANDOM}};
  r_551 = _RAND_551[0:0];
  _RAND_552 = {1{`RANDOM}};
  r_552 = _RAND_552[0:0];
  _RAND_553 = {1{`RANDOM}};
  r_553 = _RAND_553[0:0];
  _RAND_554 = {1{`RANDOM}};
  r_554 = _RAND_554[0:0];
  _RAND_555 = {1{`RANDOM}};
  r_555 = _RAND_555[0:0];
  _RAND_556 = {1{`RANDOM}};
  r_556 = _RAND_556[0:0];
  _RAND_557 = {1{`RANDOM}};
  r_557 = _RAND_557[0:0];
  _RAND_558 = {1{`RANDOM}};
  r_558 = _RAND_558[0:0];
  _RAND_559 = {1{`RANDOM}};
  r_559 = _RAND_559[0:0];
  _RAND_560 = {1{`RANDOM}};
  r_560 = _RAND_560[0:0];
  _RAND_561 = {1{`RANDOM}};
  r_561 = _RAND_561[0:0];
  _RAND_562 = {1{`RANDOM}};
  r_562 = _RAND_562[0:0];
  _RAND_563 = {1{`RANDOM}};
  r_563 = _RAND_563[0:0];
  _RAND_564 = {1{`RANDOM}};
  r_564 = _RAND_564[0:0];
  _RAND_565 = {1{`RANDOM}};
  r_565 = _RAND_565[0:0];
  _RAND_566 = {1{`RANDOM}};
  r_566 = _RAND_566[0:0];
  _RAND_567 = {1{`RANDOM}};
  r_567 = _RAND_567[0:0];
  _RAND_568 = {1{`RANDOM}};
  r_568 = _RAND_568[0:0];
  _RAND_569 = {1{`RANDOM}};
  r_569 = _RAND_569[0:0];
  _RAND_570 = {1{`RANDOM}};
  r_570 = _RAND_570[0:0];
  _RAND_571 = {1{`RANDOM}};
  r_571 = _RAND_571[0:0];
  _RAND_572 = {1{`RANDOM}};
  r_572 = _RAND_572[0:0];
  _RAND_573 = {1{`RANDOM}};
  r_573 = _RAND_573[0:0];
  _RAND_574 = {1{`RANDOM}};
  r_574 = _RAND_574[0:0];
  _RAND_575 = {1{`RANDOM}};
  r_575 = _RAND_575[0:0];
  _RAND_576 = {1{`RANDOM}};
  r_576 = _RAND_576[0:0];
  _RAND_577 = {1{`RANDOM}};
  r_577 = _RAND_577[0:0];
  _RAND_578 = {1{`RANDOM}};
  r_578 = _RAND_578[0:0];
  _RAND_579 = {1{`RANDOM}};
  r_579 = _RAND_579[0:0];
  _RAND_580 = {1{`RANDOM}};
  r_580 = _RAND_580[0:0];
  _RAND_581 = {1{`RANDOM}};
  r_581 = _RAND_581[0:0];
  _RAND_582 = {1{`RANDOM}};
  r_582 = _RAND_582[0:0];
  _RAND_583 = {1{`RANDOM}};
  r_583 = _RAND_583[0:0];
  _RAND_584 = {1{`RANDOM}};
  r_584 = _RAND_584[0:0];
  _RAND_585 = {1{`RANDOM}};
  r_585 = _RAND_585[0:0];
  _RAND_586 = {1{`RANDOM}};
  r_586 = _RAND_586[0:0];
  _RAND_587 = {1{`RANDOM}};
  r_587 = _RAND_587[0:0];
  _RAND_588 = {1{`RANDOM}};
  r_588 = _RAND_588[0:0];
  _RAND_589 = {1{`RANDOM}};
  r_589 = _RAND_589[0:0];
  _RAND_590 = {1{`RANDOM}};
  r_590 = _RAND_590[0:0];
  _RAND_591 = {1{`RANDOM}};
  r_591 = _RAND_591[0:0];
  _RAND_592 = {1{`RANDOM}};
  r_592 = _RAND_592[0:0];
  _RAND_593 = {1{`RANDOM}};
  r_593 = _RAND_593[0:0];
  _RAND_594 = {1{`RANDOM}};
  r_594 = _RAND_594[0:0];
  _RAND_595 = {1{`RANDOM}};
  r_595 = _RAND_595[0:0];
  _RAND_596 = {1{`RANDOM}};
  r_596 = _RAND_596[0:0];
  _RAND_597 = {1{`RANDOM}};
  r_597 = _RAND_597[0:0];
  _RAND_598 = {1{`RANDOM}};
  r_598 = _RAND_598[0:0];
  _RAND_599 = {1{`RANDOM}};
  r_599 = _RAND_599[0:0];
  _RAND_600 = {1{`RANDOM}};
  r_600 = _RAND_600[0:0];
  _RAND_601 = {1{`RANDOM}};
  r_601 = _RAND_601[0:0];
  _RAND_602 = {1{`RANDOM}};
  r_602 = _RAND_602[0:0];
  _RAND_603 = {1{`RANDOM}};
  r_603 = _RAND_603[0:0];
  _RAND_604 = {1{`RANDOM}};
  r_604 = _RAND_604[0:0];
  _RAND_605 = {1{`RANDOM}};
  r_605 = _RAND_605[0:0];
  _RAND_606 = {1{`RANDOM}};
  r_606 = _RAND_606[0:0];
  _RAND_607 = {1{`RANDOM}};
  r_607 = _RAND_607[0:0];
  _RAND_608 = {1{`RANDOM}};
  r_608 = _RAND_608[0:0];
  _RAND_609 = {1{`RANDOM}};
  r_609 = _RAND_609[0:0];
  _RAND_610 = {1{`RANDOM}};
  r_610 = _RAND_610[0:0];
  _RAND_611 = {1{`RANDOM}};
  r_611 = _RAND_611[0:0];
  _RAND_612 = {1{`RANDOM}};
  r_612 = _RAND_612[0:0];
  _RAND_613 = {1{`RANDOM}};
  r_613 = _RAND_613[0:0];
  _RAND_614 = {1{`RANDOM}};
  r_614 = _RAND_614[0:0];
  _RAND_615 = {1{`RANDOM}};
  r_615 = _RAND_615[0:0];
  _RAND_616 = {1{`RANDOM}};
  r_616 = _RAND_616[0:0];
  _RAND_617 = {1{`RANDOM}};
  r_617 = _RAND_617[0:0];
  _RAND_618 = {1{`RANDOM}};
  r_618 = _RAND_618[0:0];
  _RAND_619 = {1{`RANDOM}};
  r_619 = _RAND_619[0:0];
  _RAND_620 = {1{`RANDOM}};
  r_620 = _RAND_620[0:0];
  _RAND_621 = {1{`RANDOM}};
  r_621 = _RAND_621[0:0];
  _RAND_622 = {1{`RANDOM}};
  r_622 = _RAND_622[0:0];
  _RAND_623 = {1{`RANDOM}};
  r_623 = _RAND_623[0:0];
  _RAND_624 = {1{`RANDOM}};
  r_624 = _RAND_624[0:0];
  _RAND_625 = {1{`RANDOM}};
  r_625 = _RAND_625[0:0];
  _RAND_626 = {1{`RANDOM}};
  r_626 = _RAND_626[0:0];
  _RAND_627 = {1{`RANDOM}};
  r_627 = _RAND_627[0:0];
  _RAND_628 = {1{`RANDOM}};
  r_628 = _RAND_628[0:0];
  _RAND_629 = {1{`RANDOM}};
  r_629 = _RAND_629[0:0];
  _RAND_630 = {1{`RANDOM}};
  r_630 = _RAND_630[0:0];
  _RAND_631 = {1{`RANDOM}};
  r_631 = _RAND_631[0:0];
  _RAND_632 = {1{`RANDOM}};
  r_632 = _RAND_632[0:0];
  _RAND_633 = {1{`RANDOM}};
  r_633 = _RAND_633[0:0];
  _RAND_634 = {1{`RANDOM}};
  r_634 = _RAND_634[0:0];
  _RAND_635 = {1{`RANDOM}};
  r_635 = _RAND_635[0:0];
  _RAND_636 = {1{`RANDOM}};
  r_636 = _RAND_636[0:0];
  _RAND_637 = {1{`RANDOM}};
  r_637 = _RAND_637[0:0];
  _RAND_638 = {1{`RANDOM}};
  r_638 = _RAND_638[0:0];
  _RAND_639 = {1{`RANDOM}};
  r_639 = _RAND_639[0:0];
  _RAND_640 = {1{`RANDOM}};
  r_640 = _RAND_640[0:0];
  _RAND_641 = {1{`RANDOM}};
  r_641 = _RAND_641[0:0];
  _RAND_642 = {1{`RANDOM}};
  r_642 = _RAND_642[0:0];
  _RAND_643 = {1{`RANDOM}};
  r_643 = _RAND_643[0:0];
  _RAND_644 = {1{`RANDOM}};
  r_644 = _RAND_644[0:0];
  _RAND_645 = {1{`RANDOM}};
  r_645 = _RAND_645[0:0];
  _RAND_646 = {1{`RANDOM}};
  r_646 = _RAND_646[0:0];
  _RAND_647 = {1{`RANDOM}};
  r_647 = _RAND_647[0:0];
  _RAND_648 = {1{`RANDOM}};
  r_648 = _RAND_648[0:0];
  _RAND_649 = {1{`RANDOM}};
  r_649 = _RAND_649[0:0];
  _RAND_650 = {1{`RANDOM}};
  r_650 = _RAND_650[0:0];
  _RAND_651 = {1{`RANDOM}};
  r_651 = _RAND_651[0:0];
  _RAND_652 = {1{`RANDOM}};
  r_652 = _RAND_652[0:0];
  _RAND_653 = {1{`RANDOM}};
  r_653 = _RAND_653[0:0];
  _RAND_654 = {1{`RANDOM}};
  r_654 = _RAND_654[0:0];
  _RAND_655 = {1{`RANDOM}};
  r_655 = _RAND_655[0:0];
  _RAND_656 = {1{`RANDOM}};
  r_656 = _RAND_656[0:0];
  _RAND_657 = {1{`RANDOM}};
  r_657 = _RAND_657[0:0];
  _RAND_658 = {1{`RANDOM}};
  r_658 = _RAND_658[0:0];
  _RAND_659 = {1{`RANDOM}};
  r_659 = _RAND_659[0:0];
  _RAND_660 = {1{`RANDOM}};
  r_660 = _RAND_660[0:0];
  _RAND_661 = {1{`RANDOM}};
  r_661 = _RAND_661[0:0];
  _RAND_662 = {1{`RANDOM}};
  r_662 = _RAND_662[0:0];
  _RAND_663 = {1{`RANDOM}};
  r_663 = _RAND_663[0:0];
  _RAND_664 = {1{`RANDOM}};
  r_664 = _RAND_664[0:0];
  _RAND_665 = {1{`RANDOM}};
  r_665 = _RAND_665[0:0];
  _RAND_666 = {1{`RANDOM}};
  r_666 = _RAND_666[0:0];
  _RAND_667 = {1{`RANDOM}};
  r_667 = _RAND_667[0:0];
  _RAND_668 = {1{`RANDOM}};
  r_668 = _RAND_668[0:0];
  _RAND_669 = {1{`RANDOM}};
  r_669 = _RAND_669[0:0];
  _RAND_670 = {1{`RANDOM}};
  r_670 = _RAND_670[0:0];
  _RAND_671 = {1{`RANDOM}};
  r_671 = _RAND_671[0:0];
  _RAND_672 = {1{`RANDOM}};
  r_672 = _RAND_672[0:0];
  _RAND_673 = {1{`RANDOM}};
  r_673 = _RAND_673[0:0];
  _RAND_674 = {1{`RANDOM}};
  r_674 = _RAND_674[0:0];
  _RAND_675 = {1{`RANDOM}};
  r_675 = _RAND_675[0:0];
  _RAND_676 = {1{`RANDOM}};
  r_676 = _RAND_676[0:0];
  _RAND_677 = {1{`RANDOM}};
  r_677 = _RAND_677[0:0];
  _RAND_678 = {1{`RANDOM}};
  r_678 = _RAND_678[0:0];
  _RAND_679 = {1{`RANDOM}};
  r_679 = _RAND_679[0:0];
  _RAND_680 = {1{`RANDOM}};
  r_680 = _RAND_680[0:0];
  _RAND_681 = {1{`RANDOM}};
  r_681 = _RAND_681[0:0];
  _RAND_682 = {1{`RANDOM}};
  r_682 = _RAND_682[0:0];
  _RAND_683 = {1{`RANDOM}};
  r_683 = _RAND_683[0:0];
  _RAND_684 = {1{`RANDOM}};
  r_684 = _RAND_684[0:0];
  _RAND_685 = {1{`RANDOM}};
  r_685 = _RAND_685[0:0];
  _RAND_686 = {1{`RANDOM}};
  r_686 = _RAND_686[0:0];
  _RAND_687 = {1{`RANDOM}};
  r_687 = _RAND_687[0:0];
  _RAND_688 = {1{`RANDOM}};
  r_688 = _RAND_688[0:0];
  _RAND_689 = {1{`RANDOM}};
  r_689 = _RAND_689[0:0];
  _RAND_690 = {1{`RANDOM}};
  r_690 = _RAND_690[0:0];
  _RAND_691 = {1{`RANDOM}};
  r_691 = _RAND_691[0:0];
  _RAND_692 = {1{`RANDOM}};
  r_692 = _RAND_692[0:0];
  _RAND_693 = {1{`RANDOM}};
  r_693 = _RAND_693[0:0];
  _RAND_694 = {1{`RANDOM}};
  r_694 = _RAND_694[0:0];
  _RAND_695 = {1{`RANDOM}};
  r_695 = _RAND_695[0:0];
  _RAND_696 = {1{`RANDOM}};
  r_696 = _RAND_696[0:0];
  _RAND_697 = {1{`RANDOM}};
  r_697 = _RAND_697[0:0];
  _RAND_698 = {1{`RANDOM}};
  r_698 = _RAND_698[0:0];
  _RAND_699 = {1{`RANDOM}};
  r_699 = _RAND_699[0:0];
  _RAND_700 = {1{`RANDOM}};
  r_700 = _RAND_700[0:0];
  _RAND_701 = {1{`RANDOM}};
  r_701 = _RAND_701[0:0];
  _RAND_702 = {1{`RANDOM}};
  r_702 = _RAND_702[0:0];
  _RAND_703 = {1{`RANDOM}};
  r_703 = _RAND_703[0:0];
  _RAND_704 = {1{`RANDOM}};
  r_704 = _RAND_704[0:0];
  _RAND_705 = {1{`RANDOM}};
  r_705 = _RAND_705[0:0];
  _RAND_706 = {1{`RANDOM}};
  r_706 = _RAND_706[0:0];
  _RAND_707 = {1{`RANDOM}};
  r_707 = _RAND_707[0:0];
  _RAND_708 = {1{`RANDOM}};
  r_708 = _RAND_708[0:0];
  _RAND_709 = {1{`RANDOM}};
  r_709 = _RAND_709[0:0];
  _RAND_710 = {1{`RANDOM}};
  r_710 = _RAND_710[0:0];
  _RAND_711 = {1{`RANDOM}};
  r_711 = _RAND_711[0:0];
  _RAND_712 = {1{`RANDOM}};
  r_712 = _RAND_712[0:0];
  _RAND_713 = {1{`RANDOM}};
  r_713 = _RAND_713[0:0];
  _RAND_714 = {1{`RANDOM}};
  r_714 = _RAND_714[0:0];
  _RAND_715 = {1{`RANDOM}};
  r_715 = _RAND_715[0:0];
  _RAND_716 = {1{`RANDOM}};
  r_716 = _RAND_716[0:0];
  _RAND_717 = {1{`RANDOM}};
  r_717 = _RAND_717[0:0];
  _RAND_718 = {1{`RANDOM}};
  r_718 = _RAND_718[0:0];
  _RAND_719 = {1{`RANDOM}};
  r_719 = _RAND_719[0:0];
  _RAND_720 = {1{`RANDOM}};
  r_720 = _RAND_720[0:0];
  _RAND_721 = {1{`RANDOM}};
  r_721 = _RAND_721[0:0];
  _RAND_722 = {1{`RANDOM}};
  r_722 = _RAND_722[0:0];
  _RAND_723 = {1{`RANDOM}};
  r_723 = _RAND_723[0:0];
  _RAND_724 = {1{`RANDOM}};
  r_724 = _RAND_724[0:0];
  _RAND_725 = {1{`RANDOM}};
  r_725 = _RAND_725[0:0];
  _RAND_726 = {1{`RANDOM}};
  r_726 = _RAND_726[0:0];
  _RAND_727 = {1{`RANDOM}};
  r_727 = _RAND_727[0:0];
  _RAND_728 = {1{`RANDOM}};
  r_728 = _RAND_728[0:0];
  _RAND_729 = {1{`RANDOM}};
  r_729 = _RAND_729[0:0];
  _RAND_730 = {1{`RANDOM}};
  r_730 = _RAND_730[0:0];
  _RAND_731 = {1{`RANDOM}};
  r_731 = _RAND_731[0:0];
  _RAND_732 = {1{`RANDOM}};
  r_732 = _RAND_732[0:0];
  _RAND_733 = {1{`RANDOM}};
  r_733 = _RAND_733[0:0];
  _RAND_734 = {1{`RANDOM}};
  r_734 = _RAND_734[0:0];
  _RAND_735 = {1{`RANDOM}};
  r_735 = _RAND_735[0:0];
  _RAND_736 = {1{`RANDOM}};
  r_736 = _RAND_736[0:0];
  _RAND_737 = {1{`RANDOM}};
  r_737 = _RAND_737[0:0];
  _RAND_738 = {1{`RANDOM}};
  r_738 = _RAND_738[0:0];
  _RAND_739 = {1{`RANDOM}};
  r_739 = _RAND_739[0:0];
  _RAND_740 = {1{`RANDOM}};
  r_740 = _RAND_740[0:0];
  _RAND_741 = {1{`RANDOM}};
  r_741 = _RAND_741[0:0];
  _RAND_742 = {1{`RANDOM}};
  r_742 = _RAND_742[0:0];
  _RAND_743 = {1{`RANDOM}};
  r_743 = _RAND_743[0:0];
  _RAND_744 = {1{`RANDOM}};
  r_744 = _RAND_744[0:0];
  _RAND_745 = {1{`RANDOM}};
  r_745 = _RAND_745[0:0];
  _RAND_746 = {1{`RANDOM}};
  r_746 = _RAND_746[0:0];
  _RAND_747 = {1{`RANDOM}};
  r_747 = _RAND_747[0:0];
  _RAND_748 = {1{`RANDOM}};
  r_748 = _RAND_748[0:0];
  _RAND_749 = {1{`RANDOM}};
  r_749 = _RAND_749[0:0];
  _RAND_750 = {1{`RANDOM}};
  r_750 = _RAND_750[0:0];
  _RAND_751 = {1{`RANDOM}};
  r_751 = _RAND_751[0:0];
  _RAND_752 = {1{`RANDOM}};
  r_752 = _RAND_752[0:0];
  _RAND_753 = {1{`RANDOM}};
  r_753 = _RAND_753[0:0];
  _RAND_754 = {1{`RANDOM}};
  r_754 = _RAND_754[0:0];
  _RAND_755 = {1{`RANDOM}};
  r_755 = _RAND_755[0:0];
  _RAND_756 = {1{`RANDOM}};
  r_756 = _RAND_756[0:0];
  _RAND_757 = {1{`RANDOM}};
  r_757 = _RAND_757[0:0];
  _RAND_758 = {1{`RANDOM}};
  r_758 = _RAND_758[0:0];
  _RAND_759 = {1{`RANDOM}};
  r_759 = _RAND_759[0:0];
  _RAND_760 = {1{`RANDOM}};
  r_760 = _RAND_760[0:0];
  _RAND_761 = {1{`RANDOM}};
  r_761 = _RAND_761[0:0];
  _RAND_762 = {1{`RANDOM}};
  r_762 = _RAND_762[0:0];
  _RAND_763 = {1{`RANDOM}};
  r_763 = _RAND_763[0:0];
  _RAND_764 = {1{`RANDOM}};
  r_764 = _RAND_764[0:0];
  _RAND_765 = {1{`RANDOM}};
  r_765 = _RAND_765[0:0];
  _RAND_766 = {1{`RANDOM}};
  r_766 = _RAND_766[0:0];
  _RAND_767 = {1{`RANDOM}};
  r_767 = _RAND_767[0:0];
  _RAND_768 = {1{`RANDOM}};
  r_768 = _RAND_768[0:0];
  _RAND_769 = {1{`RANDOM}};
  r_769 = _RAND_769[0:0];
  _RAND_770 = {1{`RANDOM}};
  r_770 = _RAND_770[0:0];
  _RAND_771 = {1{`RANDOM}};
  r_771 = _RAND_771[0:0];
  _RAND_772 = {1{`RANDOM}};
  r_772 = _RAND_772[0:0];
  _RAND_773 = {1{`RANDOM}};
  r_773 = _RAND_773[0:0];
  _RAND_774 = {1{`RANDOM}};
  r_774 = _RAND_774[0:0];
  _RAND_775 = {1{`RANDOM}};
  r_775 = _RAND_775[0:0];
  _RAND_776 = {1{`RANDOM}};
  r_776 = _RAND_776[0:0];
  _RAND_777 = {1{`RANDOM}};
  r_777 = _RAND_777[0:0];
  _RAND_778 = {1{`RANDOM}};
  r_778 = _RAND_778[0:0];
  _RAND_779 = {1{`RANDOM}};
  r_779 = _RAND_779[0:0];
  _RAND_780 = {1{`RANDOM}};
  r_780 = _RAND_780[0:0];
  _RAND_781 = {1{`RANDOM}};
  r_781 = _RAND_781[0:0];
  _RAND_782 = {1{`RANDOM}};
  r_782 = _RAND_782[0:0];
  _RAND_783 = {1{`RANDOM}};
  r_783 = _RAND_783[0:0];
  _RAND_784 = {1{`RANDOM}};
  r_784 = _RAND_784[0:0];
  _RAND_785 = {1{`RANDOM}};
  r_785 = _RAND_785[0:0];
  _RAND_786 = {1{`RANDOM}};
  r_786 = _RAND_786[0:0];
  _RAND_787 = {1{`RANDOM}};
  r_787 = _RAND_787[0:0];
  _RAND_788 = {1{`RANDOM}};
  r_788 = _RAND_788[0:0];
  _RAND_789 = {1{`RANDOM}};
  r_789 = _RAND_789[0:0];
  _RAND_790 = {1{`RANDOM}};
  r_790 = _RAND_790[0:0];
  _RAND_791 = {1{`RANDOM}};
  r_791 = _RAND_791[0:0];
  _RAND_792 = {1{`RANDOM}};
  r_792 = _RAND_792[0:0];
  _RAND_793 = {1{`RANDOM}};
  r_793 = _RAND_793[0:0];
  _RAND_794 = {1{`RANDOM}};
  r_794 = _RAND_794[0:0];
  _RAND_795 = {1{`RANDOM}};
  r_795 = _RAND_795[0:0];
  _RAND_796 = {1{`RANDOM}};
  r_796 = _RAND_796[0:0];
  _RAND_797 = {1{`RANDOM}};
  r_797 = _RAND_797[0:0];
  _RAND_798 = {1{`RANDOM}};
  r_798 = _RAND_798[0:0];
  _RAND_799 = {1{`RANDOM}};
  r_799 = _RAND_799[0:0];
  _RAND_800 = {1{`RANDOM}};
  r_800 = _RAND_800[0:0];
  _RAND_801 = {1{`RANDOM}};
  r_801 = _RAND_801[0:0];
  _RAND_802 = {1{`RANDOM}};
  r_802 = _RAND_802[0:0];
  _RAND_803 = {1{`RANDOM}};
  r_803 = _RAND_803[0:0];
  _RAND_804 = {1{`RANDOM}};
  r_804 = _RAND_804[0:0];
  _RAND_805 = {1{`RANDOM}};
  r_805 = _RAND_805[0:0];
  _RAND_806 = {1{`RANDOM}};
  r_806 = _RAND_806[0:0];
  _RAND_807 = {1{`RANDOM}};
  r_807 = _RAND_807[0:0];
  _RAND_808 = {1{`RANDOM}};
  r_808 = _RAND_808[0:0];
  _RAND_809 = {1{`RANDOM}};
  r_809 = _RAND_809[0:0];
  _RAND_810 = {1{`RANDOM}};
  r_810 = _RAND_810[0:0];
  _RAND_811 = {1{`RANDOM}};
  r_811 = _RAND_811[0:0];
  _RAND_812 = {1{`RANDOM}};
  r_812 = _RAND_812[0:0];
  _RAND_813 = {1{`RANDOM}};
  r_813 = _RAND_813[0:0];
  _RAND_814 = {1{`RANDOM}};
  r_814 = _RAND_814[0:0];
  _RAND_815 = {1{`RANDOM}};
  r_815 = _RAND_815[0:0];
  _RAND_816 = {1{`RANDOM}};
  r_816 = _RAND_816[0:0];
  _RAND_817 = {1{`RANDOM}};
  r_817 = _RAND_817[0:0];
  _RAND_818 = {1{`RANDOM}};
  r_818 = _RAND_818[0:0];
  _RAND_819 = {1{`RANDOM}};
  r_819 = _RAND_819[0:0];
  _RAND_820 = {1{`RANDOM}};
  r_820 = _RAND_820[0:0];
  _RAND_821 = {1{`RANDOM}};
  r_821 = _RAND_821[0:0];
  _RAND_822 = {1{`RANDOM}};
  r_822 = _RAND_822[0:0];
  _RAND_823 = {1{`RANDOM}};
  r_823 = _RAND_823[0:0];
  _RAND_824 = {1{`RANDOM}};
  r_824 = _RAND_824[0:0];
  _RAND_825 = {1{`RANDOM}};
  r_825 = _RAND_825[0:0];
  _RAND_826 = {1{`RANDOM}};
  r_826 = _RAND_826[0:0];
  _RAND_827 = {1{`RANDOM}};
  r_827 = _RAND_827[0:0];
  _RAND_828 = {1{`RANDOM}};
  r_828 = _RAND_828[0:0];
  _RAND_829 = {1{`RANDOM}};
  r_829 = _RAND_829[0:0];
  _RAND_830 = {1{`RANDOM}};
  r_830 = _RAND_830[0:0];
  _RAND_831 = {1{`RANDOM}};
  r_831 = _RAND_831[0:0];
  _RAND_832 = {1{`RANDOM}};
  r_832 = _RAND_832[0:0];
  _RAND_833 = {1{`RANDOM}};
  r_833 = _RAND_833[0:0];
  _RAND_834 = {1{`RANDOM}};
  r_834 = _RAND_834[0:0];
  _RAND_835 = {1{`RANDOM}};
  r_835 = _RAND_835[0:0];
  _RAND_836 = {1{`RANDOM}};
  r_836 = _RAND_836[0:0];
  _RAND_837 = {1{`RANDOM}};
  r_837 = _RAND_837[0:0];
  _RAND_838 = {1{`RANDOM}};
  r_838 = _RAND_838[0:0];
  _RAND_839 = {1{`RANDOM}};
  r_839 = _RAND_839[0:0];
  _RAND_840 = {1{`RANDOM}};
  r_840 = _RAND_840[0:0];
  _RAND_841 = {1{`RANDOM}};
  r_841 = _RAND_841[0:0];
  _RAND_842 = {1{`RANDOM}};
  r_842 = _RAND_842[0:0];
  _RAND_843 = {1{`RANDOM}};
  r_843 = _RAND_843[0:0];
  _RAND_844 = {1{`RANDOM}};
  r_844 = _RAND_844[0:0];
  _RAND_845 = {1{`RANDOM}};
  r_845 = _RAND_845[0:0];
  _RAND_846 = {1{`RANDOM}};
  r_846 = _RAND_846[0:0];
  _RAND_847 = {1{`RANDOM}};
  r_847 = _RAND_847[0:0];
  _RAND_848 = {1{`RANDOM}};
  r_848 = _RAND_848[0:0];
  _RAND_849 = {1{`RANDOM}};
  r_849 = _RAND_849[0:0];
  _RAND_850 = {1{`RANDOM}};
  r_850 = _RAND_850[0:0];
  _RAND_851 = {1{`RANDOM}};
  r_851 = _RAND_851[0:0];
  _RAND_852 = {1{`RANDOM}};
  r_852 = _RAND_852[0:0];
  _RAND_853 = {1{`RANDOM}};
  r_853 = _RAND_853[0:0];
  _RAND_854 = {1{`RANDOM}};
  r_854 = _RAND_854[0:0];
  _RAND_855 = {1{`RANDOM}};
  r_855 = _RAND_855[0:0];
  _RAND_856 = {1{`RANDOM}};
  r_856 = _RAND_856[0:0];
  _RAND_857 = {1{`RANDOM}};
  r_857 = _RAND_857[0:0];
  _RAND_858 = {1{`RANDOM}};
  r_858 = _RAND_858[0:0];
  _RAND_859 = {1{`RANDOM}};
  r_859 = _RAND_859[0:0];
  _RAND_860 = {1{`RANDOM}};
  r_860 = _RAND_860[0:0];
  _RAND_861 = {1{`RANDOM}};
  r_861 = _RAND_861[0:0];
  _RAND_862 = {1{`RANDOM}};
  r_862 = _RAND_862[0:0];
  _RAND_863 = {1{`RANDOM}};
  r_863 = _RAND_863[0:0];
  _RAND_864 = {1{`RANDOM}};
  r_864 = _RAND_864[0:0];
  _RAND_865 = {1{`RANDOM}};
  r_865 = _RAND_865[0:0];
  _RAND_866 = {1{`RANDOM}};
  r_866 = _RAND_866[0:0];
  _RAND_867 = {1{`RANDOM}};
  r_867 = _RAND_867[0:0];
  _RAND_868 = {1{`RANDOM}};
  r_868 = _RAND_868[0:0];
  _RAND_869 = {1{`RANDOM}};
  r_869 = _RAND_869[0:0];
  _RAND_870 = {1{`RANDOM}};
  r_870 = _RAND_870[0:0];
  _RAND_871 = {1{`RANDOM}};
  r_871 = _RAND_871[0:0];
  _RAND_872 = {1{`RANDOM}};
  r_872 = _RAND_872[0:0];
  _RAND_873 = {1{`RANDOM}};
  r_873 = _RAND_873[0:0];
  _RAND_874 = {1{`RANDOM}};
  r_874 = _RAND_874[0:0];
  _RAND_875 = {1{`RANDOM}};
  r_875 = _RAND_875[0:0];
  _RAND_876 = {1{`RANDOM}};
  r_876 = _RAND_876[0:0];
  _RAND_877 = {1{`RANDOM}};
  r_877 = _RAND_877[0:0];
  _RAND_878 = {1{`RANDOM}};
  r_878 = _RAND_878[0:0];
  _RAND_879 = {1{`RANDOM}};
  r_879 = _RAND_879[0:0];
  _RAND_880 = {1{`RANDOM}};
  r_880 = _RAND_880[0:0];
  _RAND_881 = {1{`RANDOM}};
  r_881 = _RAND_881[0:0];
  _RAND_882 = {1{`RANDOM}};
  r_882 = _RAND_882[0:0];
  _RAND_883 = {1{`RANDOM}};
  r_883 = _RAND_883[0:0];
  _RAND_884 = {1{`RANDOM}};
  r_884 = _RAND_884[0:0];
  _RAND_885 = {1{`RANDOM}};
  r_885 = _RAND_885[0:0];
  _RAND_886 = {1{`RANDOM}};
  r_886 = _RAND_886[0:0];
  _RAND_887 = {1{`RANDOM}};
  r_887 = _RAND_887[0:0];
  _RAND_888 = {1{`RANDOM}};
  r_888 = _RAND_888[0:0];
  _RAND_889 = {1{`RANDOM}};
  r_889 = _RAND_889[0:0];
  _RAND_890 = {1{`RANDOM}};
  r_890 = _RAND_890[0:0];
  _RAND_891 = {1{`RANDOM}};
  r_891 = _RAND_891[0:0];
  _RAND_892 = {1{`RANDOM}};
  r_892 = _RAND_892[0:0];
  _RAND_893 = {1{`RANDOM}};
  r_893 = _RAND_893[0:0];
  _RAND_894 = {1{`RANDOM}};
  r_894 = _RAND_894[0:0];
  _RAND_895 = {1{`RANDOM}};
  r_895 = _RAND_895[0:0];
  _RAND_896 = {1{`RANDOM}};
  r_896 = _RAND_896[0:0];
  _RAND_897 = {1{`RANDOM}};
  r_897 = _RAND_897[0:0];
  _RAND_898 = {1{`RANDOM}};
  r_898 = _RAND_898[0:0];
  _RAND_899 = {1{`RANDOM}};
  r_899 = _RAND_899[0:0];
  _RAND_900 = {1{`RANDOM}};
  r_900 = _RAND_900[0:0];
  _RAND_901 = {1{`RANDOM}};
  r_901 = _RAND_901[0:0];
  _RAND_902 = {1{`RANDOM}};
  r_902 = _RAND_902[0:0];
  _RAND_903 = {1{`RANDOM}};
  r_903 = _RAND_903[0:0];
  _RAND_904 = {1{`RANDOM}};
  r_904 = _RAND_904[0:0];
  _RAND_905 = {1{`RANDOM}};
  r_905 = _RAND_905[0:0];
  _RAND_906 = {1{`RANDOM}};
  r_906 = _RAND_906[0:0];
  _RAND_907 = {1{`RANDOM}};
  r_907 = _RAND_907[0:0];
  _RAND_908 = {1{`RANDOM}};
  r_908 = _RAND_908[0:0];
  _RAND_909 = {1{`RANDOM}};
  r_909 = _RAND_909[0:0];
  _RAND_910 = {1{`RANDOM}};
  r_910 = _RAND_910[0:0];
  _RAND_911 = {1{`RANDOM}};
  r_911 = _RAND_911[0:0];
  _RAND_912 = {1{`RANDOM}};
  r_912 = _RAND_912[0:0];
  _RAND_913 = {1{`RANDOM}};
  r_913 = _RAND_913[0:0];
  _RAND_914 = {1{`RANDOM}};
  r_914 = _RAND_914[0:0];
  _RAND_915 = {1{`RANDOM}};
  r_915 = _RAND_915[0:0];
  _RAND_916 = {1{`RANDOM}};
  r_916 = _RAND_916[0:0];
  _RAND_917 = {1{`RANDOM}};
  r_917 = _RAND_917[0:0];
  _RAND_918 = {1{`RANDOM}};
  r_918 = _RAND_918[0:0];
  _RAND_919 = {1{`RANDOM}};
  r_919 = _RAND_919[0:0];
  _RAND_920 = {1{`RANDOM}};
  r_920 = _RAND_920[0:0];
  _RAND_921 = {1{`RANDOM}};
  r_921 = _RAND_921[0:0];
  _RAND_922 = {1{`RANDOM}};
  r_922 = _RAND_922[0:0];
  _RAND_923 = {1{`RANDOM}};
  r_923 = _RAND_923[0:0];
  _RAND_924 = {1{`RANDOM}};
  r_924 = _RAND_924[0:0];
  _RAND_925 = {1{`RANDOM}};
  r_925 = _RAND_925[0:0];
  _RAND_926 = {1{`RANDOM}};
  r_926 = _RAND_926[0:0];
  _RAND_927 = {1{`RANDOM}};
  r_927 = _RAND_927[0:0];
  _RAND_928 = {1{`RANDOM}};
  r_928 = _RAND_928[0:0];
  _RAND_929 = {1{`RANDOM}};
  r_929 = _RAND_929[0:0];
  _RAND_930 = {1{`RANDOM}};
  r_930 = _RAND_930[0:0];
  _RAND_931 = {1{`RANDOM}};
  r_931 = _RAND_931[0:0];
  _RAND_932 = {1{`RANDOM}};
  r_932 = _RAND_932[0:0];
  _RAND_933 = {1{`RANDOM}};
  r_933 = _RAND_933[0:0];
  _RAND_934 = {1{`RANDOM}};
  r_934 = _RAND_934[0:0];
  _RAND_935 = {1{`RANDOM}};
  r_935 = _RAND_935[0:0];
  _RAND_936 = {1{`RANDOM}};
  r_936 = _RAND_936[0:0];
  _RAND_937 = {1{`RANDOM}};
  r_937 = _RAND_937[0:0];
  _RAND_938 = {1{`RANDOM}};
  r_938 = _RAND_938[0:0];
  _RAND_939 = {1{`RANDOM}};
  r_939 = _RAND_939[0:0];
  _RAND_940 = {1{`RANDOM}};
  r_940 = _RAND_940[0:0];
  _RAND_941 = {1{`RANDOM}};
  r_941 = _RAND_941[0:0];
  _RAND_942 = {1{`RANDOM}};
  r_942 = _RAND_942[0:0];
  _RAND_943 = {1{`RANDOM}};
  r_943 = _RAND_943[0:0];
  _RAND_944 = {1{`RANDOM}};
  r_944 = _RAND_944[0:0];
  _RAND_945 = {1{`RANDOM}};
  r_945 = _RAND_945[0:0];
  _RAND_946 = {1{`RANDOM}};
  r_946 = _RAND_946[0:0];
  _RAND_947 = {1{`RANDOM}};
  r_947 = _RAND_947[0:0];
  _RAND_948 = {1{`RANDOM}};
  r_948 = _RAND_948[0:0];
  _RAND_949 = {1{`RANDOM}};
  r_949 = _RAND_949[0:0];
  _RAND_950 = {1{`RANDOM}};
  r_950 = _RAND_950[0:0];
  _RAND_951 = {1{`RANDOM}};
  r_951 = _RAND_951[0:0];
  _RAND_952 = {1{`RANDOM}};
  r_952 = _RAND_952[0:0];
  _RAND_953 = {1{`RANDOM}};
  r_953 = _RAND_953[0:0];
  _RAND_954 = {1{`RANDOM}};
  r_954 = _RAND_954[0:0];
  _RAND_955 = {1{`RANDOM}};
  r_955 = _RAND_955[0:0];
  _RAND_956 = {1{`RANDOM}};
  r_956 = _RAND_956[0:0];
  _RAND_957 = {1{`RANDOM}};
  r_957 = _RAND_957[0:0];
  _RAND_958 = {1{`RANDOM}};
  r_958 = _RAND_958[0:0];
  _RAND_959 = {1{`RANDOM}};
  r_959 = _RAND_959[0:0];
  _RAND_960 = {1{`RANDOM}};
  r_960 = _RAND_960[0:0];
  _RAND_961 = {1{`RANDOM}};
  r_961 = _RAND_961[0:0];
  _RAND_962 = {1{`RANDOM}};
  r_962 = _RAND_962[0:0];
  _RAND_963 = {1{`RANDOM}};
  r_963 = _RAND_963[0:0];
  _RAND_964 = {1{`RANDOM}};
  r_964 = _RAND_964[0:0];
  _RAND_965 = {1{`RANDOM}};
  r_965 = _RAND_965[0:0];
  _RAND_966 = {1{`RANDOM}};
  r_966 = _RAND_966[0:0];
  _RAND_967 = {1{`RANDOM}};
  r_967 = _RAND_967[0:0];
  _RAND_968 = {1{`RANDOM}};
  r_968 = _RAND_968[0:0];
  _RAND_969 = {1{`RANDOM}};
  r_969 = _RAND_969[0:0];
  _RAND_970 = {1{`RANDOM}};
  r_970 = _RAND_970[0:0];
  _RAND_971 = {1{`RANDOM}};
  r_971 = _RAND_971[0:0];
  _RAND_972 = {1{`RANDOM}};
  r_972 = _RAND_972[0:0];
  _RAND_973 = {1{`RANDOM}};
  r_973 = _RAND_973[0:0];
  _RAND_974 = {1{`RANDOM}};
  r_974 = _RAND_974[0:0];
  _RAND_975 = {1{`RANDOM}};
  r_975 = _RAND_975[0:0];
  _RAND_976 = {1{`RANDOM}};
  r_976 = _RAND_976[0:0];
  _RAND_977 = {1{`RANDOM}};
  r_977 = _RAND_977[0:0];
  _RAND_978 = {1{`RANDOM}};
  r_978 = _RAND_978[0:0];
  _RAND_979 = {1{`RANDOM}};
  r_979 = _RAND_979[0:0];
  _RAND_980 = {1{`RANDOM}};
  r_980 = _RAND_980[0:0];
  _RAND_981 = {1{`RANDOM}};
  r_981 = _RAND_981[0:0];
  _RAND_982 = {1{`RANDOM}};
  r_982 = _RAND_982[0:0];
  _RAND_983 = {1{`RANDOM}};
  r_983 = _RAND_983[0:0];
  _RAND_984 = {1{`RANDOM}};
  r_984 = _RAND_984[0:0];
  _RAND_985 = {1{`RANDOM}};
  r_985 = _RAND_985[0:0];
  _RAND_986 = {1{`RANDOM}};
  r_986 = _RAND_986[0:0];
  _RAND_987 = {1{`RANDOM}};
  r_987 = _RAND_987[0:0];
  _RAND_988 = {1{`RANDOM}};
  r_988 = _RAND_988[0:0];
  _RAND_989 = {1{`RANDOM}};
  r_989 = _RAND_989[0:0];
  _RAND_990 = {1{`RANDOM}};
  r_990 = _RAND_990[0:0];
  _RAND_991 = {1{`RANDOM}};
  r_991 = _RAND_991[0:0];
  _RAND_992 = {1{`RANDOM}};
  r_992 = _RAND_992[0:0];
  _RAND_993 = {1{`RANDOM}};
  r_993 = _RAND_993[0:0];
  _RAND_994 = {1{`RANDOM}};
  r_994 = _RAND_994[0:0];
  _RAND_995 = {1{`RANDOM}};
  r_995 = _RAND_995[0:0];
  _RAND_996 = {1{`RANDOM}};
  r_996 = _RAND_996[0:0];
  _RAND_997 = {1{`RANDOM}};
  r_997 = _RAND_997[0:0];
  _RAND_998 = {1{`RANDOM}};
  r_998 = _RAND_998[0:0];
  _RAND_999 = {1{`RANDOM}};
  r_999 = _RAND_999[0:0];
  _RAND_1000 = {1{`RANDOM}};
  r_1000 = _RAND_1000[0:0];
  _RAND_1001 = {1{`RANDOM}};
  r_1001 = _RAND_1001[0:0];
  _RAND_1002 = {1{`RANDOM}};
  r_1002 = _RAND_1002[0:0];
  _RAND_1003 = {1{`RANDOM}};
  r_1003 = _RAND_1003[0:0];
  _RAND_1004 = {1{`RANDOM}};
  r_1004 = _RAND_1004[0:0];
  _RAND_1005 = {1{`RANDOM}};
  r_1005 = _RAND_1005[0:0];
  _RAND_1006 = {1{`RANDOM}};
  r_1006 = _RAND_1006[0:0];
  _RAND_1007 = {1{`RANDOM}};
  r_1007 = _RAND_1007[0:0];
  _RAND_1008 = {1{`RANDOM}};
  r_1008 = _RAND_1008[0:0];
  _RAND_1009 = {1{`RANDOM}};
  r_1009 = _RAND_1009[0:0];
  _RAND_1010 = {1{`RANDOM}};
  r_1010 = _RAND_1010[0:0];
  _RAND_1011 = {1{`RANDOM}};
  r_1011 = _RAND_1011[0:0];
  _RAND_1012 = {1{`RANDOM}};
  r_1012 = _RAND_1012[0:0];
  _RAND_1013 = {1{`RANDOM}};
  r_1013 = _RAND_1013[0:0];
  _RAND_1014 = {1{`RANDOM}};
  r_1014 = _RAND_1014[0:0];
  _RAND_1015 = {1{`RANDOM}};
  r_1015 = _RAND_1015[0:0];
  _RAND_1016 = {1{`RANDOM}};
  r_1016 = _RAND_1016[0:0];
  _RAND_1017 = {1{`RANDOM}};
  r_1017 = _RAND_1017[0:0];
  _RAND_1018 = {1{`RANDOM}};
  r_1018 = _RAND_1018[0:0];
  _RAND_1019 = {1{`RANDOM}};
  r_1019 = _RAND_1019[0:0];
  _RAND_1020 = {1{`RANDOM}};
  r_1020 = _RAND_1020[0:0];
  _RAND_1021 = {1{`RANDOM}};
  r_1021 = _RAND_1021[0:0];
  _RAND_1022 = {1{`RANDOM}};
  r_1022 = _RAND_1022[0:0];
  _RAND_1023 = {1{`RANDOM}};
  r_1023 = _RAND_1023[0:0];
  _RAND_1024 = {1{`RANDOM}};
  r_1024 = _RAND_1024[0:0];
  _RAND_1025 = {1{`RANDOM}};
  r_1025 = _RAND_1025[0:0];
  _RAND_1026 = {1{`RANDOM}};
  r_1026 = _RAND_1026[0:0];
  _RAND_1027 = {1{`RANDOM}};
  r_1027 = _RAND_1027[0:0];
  _RAND_1028 = {1{`RANDOM}};
  r_1028 = _RAND_1028[0:0];
  _RAND_1029 = {1{`RANDOM}};
  r_1029 = _RAND_1029[0:0];
  _RAND_1030 = {1{`RANDOM}};
  r_1030 = _RAND_1030[0:0];
  _RAND_1031 = {1{`RANDOM}};
  r_1031 = _RAND_1031[0:0];
  _RAND_1032 = {1{`RANDOM}};
  r_1032 = _RAND_1032[0:0];
  _RAND_1033 = {1{`RANDOM}};
  r_1033 = _RAND_1033[0:0];
  _RAND_1034 = {1{`RANDOM}};
  r_1034 = _RAND_1034[0:0];
  _RAND_1035 = {1{`RANDOM}};
  r_1035 = _RAND_1035[0:0];
  _RAND_1036 = {1{`RANDOM}};
  r_1036 = _RAND_1036[0:0];
  _RAND_1037 = {1{`RANDOM}};
  r_1037 = _RAND_1037[0:0];
  _RAND_1038 = {1{`RANDOM}};
  r_1038 = _RAND_1038[0:0];
  _RAND_1039 = {1{`RANDOM}};
  r_1039 = _RAND_1039[0:0];
  _RAND_1040 = {1{`RANDOM}};
  r_1040 = _RAND_1040[0:0];
  _RAND_1041 = {1{`RANDOM}};
  r_1041 = _RAND_1041[0:0];
  _RAND_1042 = {1{`RANDOM}};
  r_1042 = _RAND_1042[0:0];
  _RAND_1043 = {1{`RANDOM}};
  r_1043 = _RAND_1043[0:0];
  _RAND_1044 = {1{`RANDOM}};
  r_1044 = _RAND_1044[0:0];
  _RAND_1045 = {1{`RANDOM}};
  r_1045 = _RAND_1045[0:0];
  _RAND_1046 = {1{`RANDOM}};
  r_1046 = _RAND_1046[0:0];
  _RAND_1047 = {1{`RANDOM}};
  r_1047 = _RAND_1047[0:0];
  _RAND_1048 = {1{`RANDOM}};
  r_1048 = _RAND_1048[0:0];
  _RAND_1049 = {1{`RANDOM}};
  r_1049 = _RAND_1049[0:0];
  _RAND_1050 = {1{`RANDOM}};
  r_1050 = _RAND_1050[0:0];
  _RAND_1051 = {1{`RANDOM}};
  r_1051 = _RAND_1051[0:0];
  _RAND_1052 = {1{`RANDOM}};
  r_1052 = _RAND_1052[0:0];
  _RAND_1053 = {1{`RANDOM}};
  r_1053 = _RAND_1053[0:0];
  _RAND_1054 = {1{`RANDOM}};
  r_1054 = _RAND_1054[0:0];
  _RAND_1055 = {1{`RANDOM}};
  r_1055 = _RAND_1055[0:0];
  _RAND_1056 = {1{`RANDOM}};
  r_1056 = _RAND_1056[0:0];
  _RAND_1057 = {1{`RANDOM}};
  r_1057 = _RAND_1057[0:0];
  _RAND_1058 = {1{`RANDOM}};
  r_1058 = _RAND_1058[0:0];
  _RAND_1059 = {1{`RANDOM}};
  r_1059 = _RAND_1059[0:0];
  _RAND_1060 = {1{`RANDOM}};
  r_1060 = _RAND_1060[0:0];
  _RAND_1061 = {1{`RANDOM}};
  r_1061 = _RAND_1061[0:0];
  _RAND_1062 = {1{`RANDOM}};
  r_1062 = _RAND_1062[0:0];
  _RAND_1063 = {1{`RANDOM}};
  r_1063 = _RAND_1063[0:0];
  _RAND_1064 = {1{`RANDOM}};
  r_1064 = _RAND_1064[0:0];
  _RAND_1065 = {1{`RANDOM}};
  r_1065 = _RAND_1065[0:0];
  _RAND_1066 = {1{`RANDOM}};
  r_1066 = _RAND_1066[0:0];
  _RAND_1067 = {1{`RANDOM}};
  r_1067 = _RAND_1067[0:0];
  _RAND_1068 = {1{`RANDOM}};
  r_1068 = _RAND_1068[0:0];
  _RAND_1069 = {1{`RANDOM}};
  r_1069 = _RAND_1069[0:0];
  _RAND_1070 = {1{`RANDOM}};
  r_1070 = _RAND_1070[0:0];
  _RAND_1071 = {1{`RANDOM}};
  r_1071 = _RAND_1071[0:0];
  _RAND_1072 = {1{`RANDOM}};
  r_1072 = _RAND_1072[0:0];
  _RAND_1073 = {1{`RANDOM}};
  r_1073 = _RAND_1073[0:0];
  _RAND_1074 = {1{`RANDOM}};
  r_1074 = _RAND_1074[0:0];
  _RAND_1075 = {1{`RANDOM}};
  r_1075 = _RAND_1075[0:0];
  _RAND_1076 = {1{`RANDOM}};
  r_1076 = _RAND_1076[0:0];
  _RAND_1077 = {1{`RANDOM}};
  r_1077 = _RAND_1077[0:0];
  _RAND_1078 = {1{`RANDOM}};
  r_1078 = _RAND_1078[0:0];
  _RAND_1079 = {1{`RANDOM}};
  r_1079 = _RAND_1079[0:0];
  _RAND_1080 = {1{`RANDOM}};
  r_1080 = _RAND_1080[0:0];
  _RAND_1081 = {1{`RANDOM}};
  r_1081 = _RAND_1081[0:0];
  _RAND_1082 = {1{`RANDOM}};
  r_1082 = _RAND_1082[0:0];
  _RAND_1083 = {1{`RANDOM}};
  r_1083 = _RAND_1083[0:0];
  _RAND_1084 = {1{`RANDOM}};
  r_1084 = _RAND_1084[0:0];
  _RAND_1085 = {1{`RANDOM}};
  r_1085 = _RAND_1085[0:0];
  _RAND_1086 = {1{`RANDOM}};
  r_1086 = _RAND_1086[0:0];
  _RAND_1087 = {1{`RANDOM}};
  r_1087 = _RAND_1087[0:0];
  _RAND_1088 = {1{`RANDOM}};
  r_1088 = _RAND_1088[0:0];
  _RAND_1089 = {1{`RANDOM}};
  r_1089 = _RAND_1089[0:0];
  _RAND_1090 = {1{`RANDOM}};
  r_1090 = _RAND_1090[0:0];
  _RAND_1091 = {1{`RANDOM}};
  r_1091 = _RAND_1091[0:0];
  _RAND_1092 = {1{`RANDOM}};
  r_1092 = _RAND_1092[0:0];
  _RAND_1093 = {1{`RANDOM}};
  r_1093 = _RAND_1093[0:0];
  _RAND_1094 = {1{`RANDOM}};
  r_1094 = _RAND_1094[0:0];
  _RAND_1095 = {1{`RANDOM}};
  r_1095 = _RAND_1095[0:0];
  _RAND_1096 = {1{`RANDOM}};
  r_1096 = _RAND_1096[0:0];
  _RAND_1097 = {1{`RANDOM}};
  r_1097 = _RAND_1097[0:0];
  _RAND_1098 = {1{`RANDOM}};
  r_1098 = _RAND_1098[0:0];
  _RAND_1099 = {1{`RANDOM}};
  r_1099 = _RAND_1099[0:0];
  _RAND_1100 = {1{`RANDOM}};
  r_1100 = _RAND_1100[0:0];
  _RAND_1101 = {1{`RANDOM}};
  r_1101 = _RAND_1101[0:0];
  _RAND_1102 = {1{`RANDOM}};
  r_1102 = _RAND_1102[0:0];
  _RAND_1103 = {1{`RANDOM}};
  r_1103 = _RAND_1103[0:0];
  _RAND_1104 = {1{`RANDOM}};
  r_1104 = _RAND_1104[0:0];
  _RAND_1105 = {1{`RANDOM}};
  r_1105 = _RAND_1105[0:0];
  _RAND_1106 = {1{`RANDOM}};
  r_1106 = _RAND_1106[0:0];
  _RAND_1107 = {1{`RANDOM}};
  r_1107 = _RAND_1107[0:0];
  _RAND_1108 = {1{`RANDOM}};
  r_1108 = _RAND_1108[0:0];
  _RAND_1109 = {1{`RANDOM}};
  r_1109 = _RAND_1109[0:0];
  _RAND_1110 = {1{`RANDOM}};
  r_1110 = _RAND_1110[0:0];
  _RAND_1111 = {1{`RANDOM}};
  r_1111 = _RAND_1111[0:0];
  _RAND_1112 = {1{`RANDOM}};
  r_1112 = _RAND_1112[0:0];
  _RAND_1113 = {1{`RANDOM}};
  r_1113 = _RAND_1113[0:0];
  _RAND_1114 = {1{`RANDOM}};
  r_1114 = _RAND_1114[0:0];
  _RAND_1115 = {1{`RANDOM}};
  r_1115 = _RAND_1115[0:0];
  _RAND_1116 = {1{`RANDOM}};
  r_1116 = _RAND_1116[0:0];
  _RAND_1117 = {1{`RANDOM}};
  r_1117 = _RAND_1117[0:0];
  _RAND_1118 = {1{`RANDOM}};
  r_1118 = _RAND_1118[0:0];
  _RAND_1119 = {1{`RANDOM}};
  r_1119 = _RAND_1119[0:0];
  _RAND_1120 = {1{`RANDOM}};
  r_1120 = _RAND_1120[0:0];
  _RAND_1121 = {1{`RANDOM}};
  r_1121 = _RAND_1121[0:0];
  _RAND_1122 = {1{`RANDOM}};
  r_1122 = _RAND_1122[0:0];
  _RAND_1123 = {1{`RANDOM}};
  r_1123 = _RAND_1123[0:0];
  _RAND_1124 = {1{`RANDOM}};
  r_1124 = _RAND_1124[0:0];
  _RAND_1125 = {1{`RANDOM}};
  r_1125 = _RAND_1125[0:0];
  _RAND_1126 = {1{`RANDOM}};
  r_1126 = _RAND_1126[0:0];
  _RAND_1127 = {1{`RANDOM}};
  r_1127 = _RAND_1127[0:0];
  _RAND_1128 = {1{`RANDOM}};
  r_1128 = _RAND_1128[0:0];
  _RAND_1129 = {1{`RANDOM}};
  r_1129 = _RAND_1129[0:0];
  _RAND_1130 = {1{`RANDOM}};
  r_1130 = _RAND_1130[0:0];
  _RAND_1131 = {1{`RANDOM}};
  r_1131 = _RAND_1131[0:0];
  _RAND_1132 = {1{`RANDOM}};
  r_1132 = _RAND_1132[0:0];
  _RAND_1133 = {1{`RANDOM}};
  r_1133 = _RAND_1133[0:0];
  _RAND_1134 = {1{`RANDOM}};
  r_1134 = _RAND_1134[0:0];
  _RAND_1135 = {1{`RANDOM}};
  r_1135 = _RAND_1135[0:0];
  _RAND_1136 = {1{`RANDOM}};
  r_1136 = _RAND_1136[0:0];
  _RAND_1137 = {1{`RANDOM}};
  r_1137 = _RAND_1137[0:0];
  _RAND_1138 = {1{`RANDOM}};
  r_1138 = _RAND_1138[0:0];
  _RAND_1139 = {1{`RANDOM}};
  r_1139 = _RAND_1139[0:0];
  _RAND_1140 = {1{`RANDOM}};
  r_1140 = _RAND_1140[0:0];
  _RAND_1141 = {1{`RANDOM}};
  r_1141 = _RAND_1141[0:0];
  _RAND_1142 = {1{`RANDOM}};
  r_1142 = _RAND_1142[0:0];
  _RAND_1143 = {1{`RANDOM}};
  r_1143 = _RAND_1143[0:0];
  _RAND_1144 = {1{`RANDOM}};
  r_1144 = _RAND_1144[0:0];
  _RAND_1145 = {1{`RANDOM}};
  r_1145 = _RAND_1145[0:0];
  _RAND_1146 = {1{`RANDOM}};
  r_1146 = _RAND_1146[0:0];
  _RAND_1147 = {1{`RANDOM}};
  r_1147 = _RAND_1147[0:0];
  _RAND_1148 = {1{`RANDOM}};
  r_1148 = _RAND_1148[0:0];
  _RAND_1149 = {1{`RANDOM}};
  r_1149 = _RAND_1149[0:0];
  _RAND_1150 = {1{`RANDOM}};
  r_1150 = _RAND_1150[0:0];
  _RAND_1151 = {1{`RANDOM}};
  r_1151 = _RAND_1151[0:0];
  _RAND_1152 = {1{`RANDOM}};
  r_1152 = _RAND_1152[0:0];
  _RAND_1153 = {1{`RANDOM}};
  r_1153 = _RAND_1153[0:0];
  _RAND_1154 = {1{`RANDOM}};
  r_1154 = _RAND_1154[0:0];
  _RAND_1155 = {1{`RANDOM}};
  r_1155 = _RAND_1155[0:0];
  _RAND_1156 = {1{`RANDOM}};
  r_1156 = _RAND_1156[0:0];
  _RAND_1157 = {1{`RANDOM}};
  r_1157 = _RAND_1157[0:0];
  _RAND_1158 = {1{`RANDOM}};
  r_1158 = _RAND_1158[0:0];
  _RAND_1159 = {1{`RANDOM}};
  r_1159 = _RAND_1159[0:0];
  _RAND_1160 = {1{`RANDOM}};
  r_1160 = _RAND_1160[0:0];
  _RAND_1161 = {1{`RANDOM}};
  r_1161 = _RAND_1161[0:0];
  _RAND_1162 = {1{`RANDOM}};
  r_1162 = _RAND_1162[0:0];
  _RAND_1163 = {1{`RANDOM}};
  r_1163 = _RAND_1163[0:0];
  _RAND_1164 = {1{`RANDOM}};
  r_1164 = _RAND_1164[0:0];
  _RAND_1165 = {1{`RANDOM}};
  r_1165 = _RAND_1165[0:0];
  _RAND_1166 = {1{`RANDOM}};
  r_1166 = _RAND_1166[0:0];
  _RAND_1167 = {1{`RANDOM}};
  r_1167 = _RAND_1167[0:0];
  _RAND_1168 = {1{`RANDOM}};
  r_1168 = _RAND_1168[0:0];
  _RAND_1169 = {1{`RANDOM}};
  r_1169 = _RAND_1169[0:0];
  _RAND_1170 = {1{`RANDOM}};
  r_1170 = _RAND_1170[0:0];
  _RAND_1171 = {1{`RANDOM}};
  r_1171 = _RAND_1171[0:0];
  _RAND_1172 = {1{`RANDOM}};
  r_1172 = _RAND_1172[0:0];
  _RAND_1173 = {1{`RANDOM}};
  r_1173 = _RAND_1173[0:0];
  _RAND_1174 = {1{`RANDOM}};
  r_1174 = _RAND_1174[0:0];
  _RAND_1175 = {1{`RANDOM}};
  r_1175 = _RAND_1175[0:0];
  _RAND_1176 = {1{`RANDOM}};
  r_1176 = _RAND_1176[0:0];
  _RAND_1177 = {1{`RANDOM}};
  r_1177 = _RAND_1177[0:0];
  _RAND_1178 = {1{`RANDOM}};
  r_1178 = _RAND_1178[0:0];
  _RAND_1179 = {1{`RANDOM}};
  r_1179 = _RAND_1179[0:0];
  _RAND_1180 = {1{`RANDOM}};
  r_1180 = _RAND_1180[0:0];
  _RAND_1181 = {1{`RANDOM}};
  r_1181 = _RAND_1181[0:0];
  _RAND_1182 = {1{`RANDOM}};
  r_1182 = _RAND_1182[0:0];
  _RAND_1183 = {1{`RANDOM}};
  r_1183 = _RAND_1183[0:0];
  _RAND_1184 = {1{`RANDOM}};
  r_1184 = _RAND_1184[0:0];
  _RAND_1185 = {1{`RANDOM}};
  r_1185 = _RAND_1185[0:0];
  _RAND_1186 = {1{`RANDOM}};
  r_1186 = _RAND_1186[0:0];
  _RAND_1187 = {1{`RANDOM}};
  r_1187 = _RAND_1187[0:0];
  _RAND_1188 = {1{`RANDOM}};
  r_1188 = _RAND_1188[0:0];
  _RAND_1189 = {1{`RANDOM}};
  r_1189 = _RAND_1189[0:0];
  _RAND_1190 = {1{`RANDOM}};
  r_1190 = _RAND_1190[0:0];
  _RAND_1191 = {1{`RANDOM}};
  r_1191 = _RAND_1191[0:0];
  _RAND_1192 = {1{`RANDOM}};
  r_1192 = _RAND_1192[0:0];
  _RAND_1193 = {1{`RANDOM}};
  r_1193 = _RAND_1193[0:0];
  _RAND_1194 = {1{`RANDOM}};
  r_1194 = _RAND_1194[0:0];
  _RAND_1195 = {1{`RANDOM}};
  r_1195 = _RAND_1195[0:0];
  _RAND_1196 = {1{`RANDOM}};
  r_1196 = _RAND_1196[0:0];
  _RAND_1197 = {1{`RANDOM}};
  r_1197 = _RAND_1197[0:0];
  _RAND_1198 = {1{`RANDOM}};
  r_1198 = _RAND_1198[0:0];
  _RAND_1199 = {1{`RANDOM}};
  r_1199 = _RAND_1199[0:0];
  _RAND_1200 = {1{`RANDOM}};
  r_1200 = _RAND_1200[0:0];
  _RAND_1201 = {1{`RANDOM}};
  r_1201 = _RAND_1201[0:0];
  _RAND_1202 = {1{`RANDOM}};
  r_1202 = _RAND_1202[0:0];
  _RAND_1203 = {1{`RANDOM}};
  r_1203 = _RAND_1203[0:0];
  _RAND_1204 = {1{`RANDOM}};
  r_1204 = _RAND_1204[0:0];
  _RAND_1205 = {1{`RANDOM}};
  r_1205 = _RAND_1205[0:0];
  _RAND_1206 = {1{`RANDOM}};
  r_1206 = _RAND_1206[0:0];
  _RAND_1207 = {1{`RANDOM}};
  r_1207 = _RAND_1207[0:0];
  _RAND_1208 = {1{`RANDOM}};
  r_1208 = _RAND_1208[0:0];
  _RAND_1209 = {1{`RANDOM}};
  r_1209 = _RAND_1209[0:0];
  _RAND_1210 = {1{`RANDOM}};
  r_1210 = _RAND_1210[0:0];
  _RAND_1211 = {1{`RANDOM}};
  r_1211 = _RAND_1211[0:0];
  _RAND_1212 = {1{`RANDOM}};
  r_1212 = _RAND_1212[0:0];
  _RAND_1213 = {1{`RANDOM}};
  r_1213 = _RAND_1213[0:0];
  _RAND_1214 = {1{`RANDOM}};
  r_1214 = _RAND_1214[0:0];
  _RAND_1215 = {1{`RANDOM}};
  r_1215 = _RAND_1215[0:0];
  _RAND_1216 = {1{`RANDOM}};
  r_1216 = _RAND_1216[0:0];
  _RAND_1217 = {1{`RANDOM}};
  r_1217 = _RAND_1217[0:0];
  _RAND_1218 = {1{`RANDOM}};
  r_1218 = _RAND_1218[0:0];
  _RAND_1219 = {1{`RANDOM}};
  r_1219 = _RAND_1219[0:0];
  _RAND_1220 = {1{`RANDOM}};
  r_1220 = _RAND_1220[0:0];
  _RAND_1221 = {1{`RANDOM}};
  r_1221 = _RAND_1221[0:0];
  _RAND_1222 = {1{`RANDOM}};
  r_1222 = _RAND_1222[0:0];
  _RAND_1223 = {1{`RANDOM}};
  r_1223 = _RAND_1223[0:0];
  _RAND_1224 = {1{`RANDOM}};
  r_1224 = _RAND_1224[0:0];
  _RAND_1225 = {1{`RANDOM}};
  r_1225 = _RAND_1225[0:0];
  _RAND_1226 = {1{`RANDOM}};
  r_1226 = _RAND_1226[0:0];
  _RAND_1227 = {1{`RANDOM}};
  r_1227 = _RAND_1227[0:0];
  _RAND_1228 = {1{`RANDOM}};
  r_1228 = _RAND_1228[0:0];
  _RAND_1229 = {1{`RANDOM}};
  r_1229 = _RAND_1229[0:0];
  _RAND_1230 = {1{`RANDOM}};
  r_1230 = _RAND_1230[0:0];
  _RAND_1231 = {1{`RANDOM}};
  r_1231 = _RAND_1231[0:0];
  _RAND_1232 = {1{`RANDOM}};
  r_1232 = _RAND_1232[0:0];
  _RAND_1233 = {1{`RANDOM}};
  r_1233 = _RAND_1233[0:0];
  _RAND_1234 = {1{`RANDOM}};
  r_1234 = _RAND_1234[0:0];
  _RAND_1235 = {1{`RANDOM}};
  r_1235 = _RAND_1235[0:0];
  _RAND_1236 = {1{`RANDOM}};
  r_1236 = _RAND_1236[0:0];
  _RAND_1237 = {1{`RANDOM}};
  r_1237 = _RAND_1237[0:0];
  _RAND_1238 = {1{`RANDOM}};
  r_1238 = _RAND_1238[0:0];
  _RAND_1239 = {1{`RANDOM}};
  r_1239 = _RAND_1239[0:0];
  _RAND_1240 = {1{`RANDOM}};
  r_1240 = _RAND_1240[0:0];
  _RAND_1241 = {1{`RANDOM}};
  r_1241 = _RAND_1241[0:0];
  _RAND_1242 = {1{`RANDOM}};
  r_1242 = _RAND_1242[0:0];
  _RAND_1243 = {1{`RANDOM}};
  r_1243 = _RAND_1243[0:0];
  _RAND_1244 = {1{`RANDOM}};
  r_1244 = _RAND_1244[0:0];
  _RAND_1245 = {1{`RANDOM}};
  r_1245 = _RAND_1245[0:0];
  _RAND_1246 = {1{`RANDOM}};
  r_1246 = _RAND_1246[0:0];
  _RAND_1247 = {1{`RANDOM}};
  r_1247 = _RAND_1247[0:0];
  _RAND_1248 = {1{`RANDOM}};
  r_1248 = _RAND_1248[0:0];
  _RAND_1249 = {1{`RANDOM}};
  r_1249 = _RAND_1249[0:0];
  _RAND_1250 = {1{`RANDOM}};
  r_1250 = _RAND_1250[0:0];
  _RAND_1251 = {1{`RANDOM}};
  r_1251 = _RAND_1251[0:0];
  _RAND_1252 = {1{`RANDOM}};
  r_1252 = _RAND_1252[0:0];
  _RAND_1253 = {1{`RANDOM}};
  r_1253 = _RAND_1253[0:0];
  _RAND_1254 = {1{`RANDOM}};
  r_1254 = _RAND_1254[0:0];
  _RAND_1255 = {1{`RANDOM}};
  r_1255 = _RAND_1255[0:0];
  _RAND_1256 = {1{`RANDOM}};
  r_1256 = _RAND_1256[0:0];
  _RAND_1257 = {1{`RANDOM}};
  r_1257 = _RAND_1257[0:0];
  _RAND_1258 = {1{`RANDOM}};
  r_1258 = _RAND_1258[0:0];
  _RAND_1259 = {1{`RANDOM}};
  r_1259 = _RAND_1259[0:0];
  _RAND_1260 = {1{`RANDOM}};
  r_1260 = _RAND_1260[0:0];
  _RAND_1261 = {1{`RANDOM}};
  r_1261 = _RAND_1261[0:0];
  _RAND_1262 = {1{`RANDOM}};
  r_1262 = _RAND_1262[0:0];
  _RAND_1263 = {1{`RANDOM}};
  r_1263 = _RAND_1263[0:0];
  _RAND_1264 = {1{`RANDOM}};
  r_1264 = _RAND_1264[0:0];
  _RAND_1265 = {1{`RANDOM}};
  r_1265 = _RAND_1265[0:0];
  _RAND_1266 = {1{`RANDOM}};
  r_1266 = _RAND_1266[0:0];
  _RAND_1267 = {1{`RANDOM}};
  r_1267 = _RAND_1267[0:0];
  _RAND_1268 = {1{`RANDOM}};
  r_1268 = _RAND_1268[0:0];
  _RAND_1269 = {1{`RANDOM}};
  r_1269 = _RAND_1269[0:0];
  _RAND_1270 = {1{`RANDOM}};
  r_1270 = _RAND_1270[0:0];
  _RAND_1271 = {1{`RANDOM}};
  r_1271 = _RAND_1271[0:0];
  _RAND_1272 = {1{`RANDOM}};
  r_1272 = _RAND_1272[0:0];
  _RAND_1273 = {1{`RANDOM}};
  r_1273 = _RAND_1273[0:0];
  _RAND_1274 = {1{`RANDOM}};
  r_1274 = _RAND_1274[0:0];
  _RAND_1275 = {1{`RANDOM}};
  r_1275 = _RAND_1275[0:0];
  _RAND_1276 = {1{`RANDOM}};
  r_1276 = _RAND_1276[0:0];
  _RAND_1277 = {1{`RANDOM}};
  r_1277 = _RAND_1277[0:0];
  _RAND_1278 = {1{`RANDOM}};
  r_1278 = _RAND_1278[0:0];
  _RAND_1279 = {1{`RANDOM}};
  r_1279 = _RAND_1279[0:0];
  _RAND_1280 = {1{`RANDOM}};
  r_1280 = _RAND_1280[0:0];
  _RAND_1281 = {1{`RANDOM}};
  r_1281 = _RAND_1281[0:0];
  _RAND_1282 = {1{`RANDOM}};
  r_1282 = _RAND_1282[0:0];
  _RAND_1283 = {1{`RANDOM}};
  r_1283 = _RAND_1283[0:0];
  _RAND_1284 = {1{`RANDOM}};
  r_1284 = _RAND_1284[0:0];
  _RAND_1285 = {1{`RANDOM}};
  r_1285 = _RAND_1285[0:0];
  _RAND_1286 = {1{`RANDOM}};
  r_1286 = _RAND_1286[0:0];
  _RAND_1287 = {1{`RANDOM}};
  r_1287 = _RAND_1287[0:0];
  _RAND_1288 = {1{`RANDOM}};
  r_1288 = _RAND_1288[0:0];
  _RAND_1289 = {1{`RANDOM}};
  r_1289 = _RAND_1289[0:0];
  _RAND_1290 = {1{`RANDOM}};
  r_1290 = _RAND_1290[0:0];
  _RAND_1291 = {1{`RANDOM}};
  r_1291 = _RAND_1291[0:0];
  _RAND_1292 = {1{`RANDOM}};
  r_1292 = _RAND_1292[0:0];
  _RAND_1293 = {1{`RANDOM}};
  r_1293 = _RAND_1293[0:0];
  _RAND_1294 = {1{`RANDOM}};
  r_1294 = _RAND_1294[0:0];
  _RAND_1295 = {1{`RANDOM}};
  r_1295 = _RAND_1295[0:0];
  _RAND_1296 = {1{`RANDOM}};
  r_1296 = _RAND_1296[0:0];
  _RAND_1297 = {1{`RANDOM}};
  r_1297 = _RAND_1297[0:0];
  _RAND_1298 = {1{`RANDOM}};
  r_1298 = _RAND_1298[0:0];
  _RAND_1299 = {1{`RANDOM}};
  r_1299 = _RAND_1299[0:0];
  _RAND_1300 = {1{`RANDOM}};
  r_1300 = _RAND_1300[0:0];
  _RAND_1301 = {1{`RANDOM}};
  r_1301 = _RAND_1301[0:0];
  _RAND_1302 = {1{`RANDOM}};
  r_1302 = _RAND_1302[0:0];
  _RAND_1303 = {1{`RANDOM}};
  r_1303 = _RAND_1303[0:0];
  _RAND_1304 = {1{`RANDOM}};
  r_1304 = _RAND_1304[0:0];
  _RAND_1305 = {1{`RANDOM}};
  r_1305 = _RAND_1305[0:0];
  _RAND_1306 = {1{`RANDOM}};
  r_1306 = _RAND_1306[0:0];
  _RAND_1307 = {1{`RANDOM}};
  r_1307 = _RAND_1307[0:0];
  _RAND_1308 = {1{`RANDOM}};
  r_1308 = _RAND_1308[0:0];
  _RAND_1309 = {1{`RANDOM}};
  r_1309 = _RAND_1309[0:0];
  _RAND_1310 = {1{`RANDOM}};
  r_1310 = _RAND_1310[0:0];
  _RAND_1311 = {1{`RANDOM}};
  r_1311 = _RAND_1311[0:0];
  _RAND_1312 = {1{`RANDOM}};
  r_1312 = _RAND_1312[0:0];
  _RAND_1313 = {1{`RANDOM}};
  r_1313 = _RAND_1313[0:0];
  _RAND_1314 = {1{`RANDOM}};
  r_1314 = _RAND_1314[0:0];
  _RAND_1315 = {1{`RANDOM}};
  r_1315 = _RAND_1315[0:0];
  _RAND_1316 = {1{`RANDOM}};
  r_1316 = _RAND_1316[0:0];
  _RAND_1317 = {1{`RANDOM}};
  r_1317 = _RAND_1317[0:0];
  _RAND_1318 = {1{`RANDOM}};
  r_1318 = _RAND_1318[0:0];
  _RAND_1319 = {1{`RANDOM}};
  r_1319 = _RAND_1319[0:0];
  _RAND_1320 = {1{`RANDOM}};
  r_1320 = _RAND_1320[0:0];
  _RAND_1321 = {1{`RANDOM}};
  r_1321 = _RAND_1321[0:0];
  _RAND_1322 = {1{`RANDOM}};
  r_1322 = _RAND_1322[0:0];
  _RAND_1323 = {1{`RANDOM}};
  r_1323 = _RAND_1323[0:0];
  _RAND_1324 = {1{`RANDOM}};
  r_1324 = _RAND_1324[0:0];
  _RAND_1325 = {1{`RANDOM}};
  r_1325 = _RAND_1325[0:0];
  _RAND_1326 = {1{`RANDOM}};
  r_1326 = _RAND_1326[0:0];
  _RAND_1327 = {1{`RANDOM}};
  r_1327 = _RAND_1327[0:0];
  _RAND_1328 = {1{`RANDOM}};
  r_1328 = _RAND_1328[0:0];
  _RAND_1329 = {1{`RANDOM}};
  r_1329 = _RAND_1329[0:0];
  _RAND_1330 = {1{`RANDOM}};
  r_1330 = _RAND_1330[0:0];
  _RAND_1331 = {1{`RANDOM}};
  r_1331 = _RAND_1331[0:0];
  _RAND_1332 = {1{`RANDOM}};
  r_1332 = _RAND_1332[0:0];
  _RAND_1333 = {1{`RANDOM}};
  r_1333 = _RAND_1333[0:0];
  _RAND_1334 = {1{`RANDOM}};
  r_1334 = _RAND_1334[0:0];
  _RAND_1335 = {1{`RANDOM}};
  r_1335 = _RAND_1335[0:0];
  _RAND_1336 = {1{`RANDOM}};
  r_1336 = _RAND_1336[0:0];
  _RAND_1337 = {1{`RANDOM}};
  r_1337 = _RAND_1337[0:0];
  _RAND_1338 = {1{`RANDOM}};
  r_1338 = _RAND_1338[0:0];
  _RAND_1339 = {1{`RANDOM}};
  r_1339 = _RAND_1339[0:0];
  _RAND_1340 = {1{`RANDOM}};
  r_1340 = _RAND_1340[0:0];
  _RAND_1341 = {1{`RANDOM}};
  r_1341 = _RAND_1341[0:0];
  _RAND_1342 = {1{`RANDOM}};
  r_1342 = _RAND_1342[0:0];
  _RAND_1343 = {1{`RANDOM}};
  r_1343 = _RAND_1343[0:0];
  _RAND_1344 = {1{`RANDOM}};
  r_1344 = _RAND_1344[0:0];
  _RAND_1345 = {1{`RANDOM}};
  r_1345 = _RAND_1345[0:0];
  _RAND_1346 = {1{`RANDOM}};
  r_1346 = _RAND_1346[0:0];
  _RAND_1347 = {1{`RANDOM}};
  r_1347 = _RAND_1347[0:0];
  _RAND_1348 = {1{`RANDOM}};
  r_1348 = _RAND_1348[0:0];
  _RAND_1349 = {1{`RANDOM}};
  r_1349 = _RAND_1349[0:0];
  _RAND_1350 = {1{`RANDOM}};
  r_1350 = _RAND_1350[0:0];
  _RAND_1351 = {1{`RANDOM}};
  r_1351 = _RAND_1351[0:0];
  _RAND_1352 = {1{`RANDOM}};
  r_1352 = _RAND_1352[0:0];
  _RAND_1353 = {1{`RANDOM}};
  r_1353 = _RAND_1353[0:0];
  _RAND_1354 = {1{`RANDOM}};
  r_1354 = _RAND_1354[0:0];
  _RAND_1355 = {1{`RANDOM}};
  r_1355 = _RAND_1355[0:0];
  _RAND_1356 = {1{`RANDOM}};
  r_1356 = _RAND_1356[0:0];
  _RAND_1357 = {1{`RANDOM}};
  r_1357 = _RAND_1357[0:0];
  _RAND_1358 = {1{`RANDOM}};
  r_1358 = _RAND_1358[0:0];
  _RAND_1359 = {1{`RANDOM}};
  r_1359 = _RAND_1359[0:0];
  _RAND_1360 = {1{`RANDOM}};
  r_1360 = _RAND_1360[0:0];
  _RAND_1361 = {1{`RANDOM}};
  r_1361 = _RAND_1361[0:0];
  _RAND_1362 = {1{`RANDOM}};
  r_1362 = _RAND_1362[0:0];
  _RAND_1363 = {1{`RANDOM}};
  r_1363 = _RAND_1363[0:0];
  _RAND_1364 = {1{`RANDOM}};
  r_1364 = _RAND_1364[0:0];
  _RAND_1365 = {1{`RANDOM}};
  r_1365 = _RAND_1365[0:0];
  _RAND_1366 = {1{`RANDOM}};
  r_1366 = _RAND_1366[0:0];
  _RAND_1367 = {1{`RANDOM}};
  r_1367 = _RAND_1367[0:0];
  _RAND_1368 = {1{`RANDOM}};
  r_1368 = _RAND_1368[0:0];
  _RAND_1369 = {1{`RANDOM}};
  r_1369 = _RAND_1369[0:0];
  _RAND_1370 = {1{`RANDOM}};
  r_1370 = _RAND_1370[0:0];
  _RAND_1371 = {1{`RANDOM}};
  r_1371 = _RAND_1371[0:0];
  _RAND_1372 = {1{`RANDOM}};
  r_1372 = _RAND_1372[0:0];
  _RAND_1373 = {1{`RANDOM}};
  r_1373 = _RAND_1373[0:0];
  _RAND_1374 = {1{`RANDOM}};
  r_1374 = _RAND_1374[0:0];
  _RAND_1375 = {1{`RANDOM}};
  r_1375 = _RAND_1375[0:0];
  _RAND_1376 = {1{`RANDOM}};
  r_1376 = _RAND_1376[0:0];
  _RAND_1377 = {1{`RANDOM}};
  r_1377 = _RAND_1377[0:0];
  _RAND_1378 = {1{`RANDOM}};
  r_1378 = _RAND_1378[0:0];
  _RAND_1379 = {1{`RANDOM}};
  r_1379 = _RAND_1379[0:0];
  _RAND_1380 = {1{`RANDOM}};
  r_1380 = _RAND_1380[0:0];
  _RAND_1381 = {1{`RANDOM}};
  r_1381 = _RAND_1381[0:0];
  _RAND_1382 = {1{`RANDOM}};
  r_1382 = _RAND_1382[0:0];
  _RAND_1383 = {1{`RANDOM}};
  r_1383 = _RAND_1383[0:0];
  _RAND_1384 = {1{`RANDOM}};
  r_1384 = _RAND_1384[0:0];
  _RAND_1385 = {1{`RANDOM}};
  r_1385 = _RAND_1385[0:0];
  _RAND_1386 = {1{`RANDOM}};
  r_1386 = _RAND_1386[0:0];
  _RAND_1387 = {1{`RANDOM}};
  r_1387 = _RAND_1387[0:0];
  _RAND_1388 = {1{`RANDOM}};
  r_1388 = _RAND_1388[0:0];
  _RAND_1389 = {1{`RANDOM}};
  r_1389 = _RAND_1389[0:0];
  _RAND_1390 = {1{`RANDOM}};
  r_1390 = _RAND_1390[0:0];
  _RAND_1391 = {1{`RANDOM}};
  r_1391 = _RAND_1391[0:0];
  _RAND_1392 = {1{`RANDOM}};
  r_1392 = _RAND_1392[0:0];
  _RAND_1393 = {1{`RANDOM}};
  r_1393 = _RAND_1393[0:0];
  _RAND_1394 = {1{`RANDOM}};
  r_1394 = _RAND_1394[0:0];
  _RAND_1395 = {1{`RANDOM}};
  r_1395 = _RAND_1395[0:0];
  _RAND_1396 = {1{`RANDOM}};
  r_1396 = _RAND_1396[0:0];
  _RAND_1397 = {1{`RANDOM}};
  r_1397 = _RAND_1397[0:0];
  _RAND_1398 = {1{`RANDOM}};
  r_1398 = _RAND_1398[0:0];
  _RAND_1399 = {1{`RANDOM}};
  r_1399 = _RAND_1399[0:0];
  _RAND_1400 = {1{`RANDOM}};
  r_1400 = _RAND_1400[0:0];
  _RAND_1401 = {1{`RANDOM}};
  r_1401 = _RAND_1401[0:0];
  _RAND_1402 = {1{`RANDOM}};
  r_1402 = _RAND_1402[0:0];
  _RAND_1403 = {1{`RANDOM}};
  r_1403 = _RAND_1403[0:0];
  _RAND_1404 = {1{`RANDOM}};
  r_1404 = _RAND_1404[0:0];
  _RAND_1405 = {1{`RANDOM}};
  r_1405 = _RAND_1405[0:0];
  _RAND_1406 = {1{`RANDOM}};
  r_1406 = _RAND_1406[0:0];
  _RAND_1407 = {1{`RANDOM}};
  r_1407 = _RAND_1407[0:0];
  _RAND_1408 = {1{`RANDOM}};
  r_1408 = _RAND_1408[0:0];
  _RAND_1409 = {1{`RANDOM}};
  r_1409 = _RAND_1409[0:0];
  _RAND_1410 = {1{`RANDOM}};
  r_1410 = _RAND_1410[0:0];
  _RAND_1411 = {1{`RANDOM}};
  r_1411 = _RAND_1411[0:0];
  _RAND_1412 = {1{`RANDOM}};
  r_1412 = _RAND_1412[0:0];
  _RAND_1413 = {1{`RANDOM}};
  r_1413 = _RAND_1413[0:0];
  _RAND_1414 = {1{`RANDOM}};
  r_1414 = _RAND_1414[0:0];
  _RAND_1415 = {1{`RANDOM}};
  r_1415 = _RAND_1415[0:0];
  _RAND_1416 = {1{`RANDOM}};
  r_1416 = _RAND_1416[0:0];
  _RAND_1417 = {1{`RANDOM}};
  r_1417 = _RAND_1417[0:0];
  _RAND_1418 = {1{`RANDOM}};
  r_1418 = _RAND_1418[0:0];
  _RAND_1419 = {1{`RANDOM}};
  r_1419 = _RAND_1419[0:0];
  _RAND_1420 = {1{`RANDOM}};
  r_1420 = _RAND_1420[0:0];
  _RAND_1421 = {1{`RANDOM}};
  r_1421 = _RAND_1421[0:0];
  _RAND_1422 = {1{`RANDOM}};
  r_1422 = _RAND_1422[0:0];
  _RAND_1423 = {1{`RANDOM}};
  r_1423 = _RAND_1423[0:0];
  _RAND_1424 = {1{`RANDOM}};
  r_1424 = _RAND_1424[0:0];
  _RAND_1425 = {1{`RANDOM}};
  r_1425 = _RAND_1425[0:0];
  _RAND_1426 = {1{`RANDOM}};
  r_1426 = _RAND_1426[0:0];
  _RAND_1427 = {1{`RANDOM}};
  r_1427 = _RAND_1427[0:0];
  _RAND_1428 = {1{`RANDOM}};
  r_1428 = _RAND_1428[0:0];
  _RAND_1429 = {1{`RANDOM}};
  r_1429 = _RAND_1429[0:0];
  _RAND_1430 = {1{`RANDOM}};
  r_1430 = _RAND_1430[0:0];
  _RAND_1431 = {1{`RANDOM}};
  r_1431 = _RAND_1431[0:0];
  _RAND_1432 = {1{`RANDOM}};
  r_1432 = _RAND_1432[0:0];
  _RAND_1433 = {1{`RANDOM}};
  r_1433 = _RAND_1433[0:0];
  _RAND_1434 = {1{`RANDOM}};
  r_1434 = _RAND_1434[0:0];
  _RAND_1435 = {1{`RANDOM}};
  r_1435 = _RAND_1435[0:0];
  _RAND_1436 = {1{`RANDOM}};
  r_1436 = _RAND_1436[0:0];
  _RAND_1437 = {1{`RANDOM}};
  r_1437 = _RAND_1437[0:0];
  _RAND_1438 = {1{`RANDOM}};
  r_1438 = _RAND_1438[0:0];
  _RAND_1439 = {1{`RANDOM}};
  r_1439 = _RAND_1439[0:0];
  _RAND_1440 = {1{`RANDOM}};
  r_1440 = _RAND_1440[0:0];
  _RAND_1441 = {1{`RANDOM}};
  r_1441 = _RAND_1441[0:0];
  _RAND_1442 = {1{`RANDOM}};
  r_1442 = _RAND_1442[0:0];
  _RAND_1443 = {1{`RANDOM}};
  r_1443 = _RAND_1443[0:0];
  _RAND_1444 = {1{`RANDOM}};
  r_1444 = _RAND_1444[0:0];
  _RAND_1445 = {1{`RANDOM}};
  r_1445 = _RAND_1445[0:0];
  _RAND_1446 = {1{`RANDOM}};
  r_1446 = _RAND_1446[0:0];
  _RAND_1447 = {1{`RANDOM}};
  r_1447 = _RAND_1447[0:0];
  _RAND_1448 = {1{`RANDOM}};
  r_1448 = _RAND_1448[0:0];
  _RAND_1449 = {1{`RANDOM}};
  r_1449 = _RAND_1449[0:0];
  _RAND_1450 = {1{`RANDOM}};
  r_1450 = _RAND_1450[0:0];
  _RAND_1451 = {1{`RANDOM}};
  r_1451 = _RAND_1451[0:0];
  _RAND_1452 = {1{`RANDOM}};
  r_1452 = _RAND_1452[0:0];
  _RAND_1453 = {1{`RANDOM}};
  r_1453 = _RAND_1453[0:0];
  _RAND_1454 = {1{`RANDOM}};
  r_1454 = _RAND_1454[0:0];
  _RAND_1455 = {1{`RANDOM}};
  r_1455 = _RAND_1455[0:0];
  _RAND_1456 = {1{`RANDOM}};
  r_1456 = _RAND_1456[0:0];
  _RAND_1457 = {1{`RANDOM}};
  r_1457 = _RAND_1457[0:0];
  _RAND_1458 = {1{`RANDOM}};
  r_1458 = _RAND_1458[0:0];
  _RAND_1459 = {1{`RANDOM}};
  r_1459 = _RAND_1459[0:0];
  _RAND_1460 = {1{`RANDOM}};
  r_1460 = _RAND_1460[0:0];
  _RAND_1461 = {1{`RANDOM}};
  r_1461 = _RAND_1461[0:0];
  _RAND_1462 = {1{`RANDOM}};
  r_1462 = _RAND_1462[0:0];
  _RAND_1463 = {1{`RANDOM}};
  r_1463 = _RAND_1463[0:0];
  _RAND_1464 = {1{`RANDOM}};
  r_1464 = _RAND_1464[0:0];
  _RAND_1465 = {1{`RANDOM}};
  r_1465 = _RAND_1465[0:0];
  _RAND_1466 = {1{`RANDOM}};
  r_1466 = _RAND_1466[0:0];
  _RAND_1467 = {1{`RANDOM}};
  r_1467 = _RAND_1467[0:0];
  _RAND_1468 = {1{`RANDOM}};
  r_1468 = _RAND_1468[0:0];
  _RAND_1469 = {1{`RANDOM}};
  r_1469 = _RAND_1469[0:0];
  _RAND_1470 = {1{`RANDOM}};
  r_1470 = _RAND_1470[0:0];
  _RAND_1471 = {1{`RANDOM}};
  r_1471 = _RAND_1471[0:0];
  _RAND_1472 = {1{`RANDOM}};
  r_1472 = _RAND_1472[0:0];
  _RAND_1473 = {1{`RANDOM}};
  r_1473 = _RAND_1473[0:0];
  _RAND_1474 = {1{`RANDOM}};
  r_1474 = _RAND_1474[0:0];
  _RAND_1475 = {1{`RANDOM}};
  r_1475 = _RAND_1475[0:0];
  _RAND_1476 = {1{`RANDOM}};
  r_1476 = _RAND_1476[0:0];
  _RAND_1477 = {1{`RANDOM}};
  r_1477 = _RAND_1477[0:0];
  _RAND_1478 = {1{`RANDOM}};
  r_1478 = _RAND_1478[0:0];
  _RAND_1479 = {1{`RANDOM}};
  r_1479 = _RAND_1479[0:0];
  _RAND_1480 = {1{`RANDOM}};
  r_1480 = _RAND_1480[0:0];
  _RAND_1481 = {1{`RANDOM}};
  r_1481 = _RAND_1481[0:0];
  _RAND_1482 = {1{`RANDOM}};
  r_1482 = _RAND_1482[0:0];
  _RAND_1483 = {1{`RANDOM}};
  r_1483 = _RAND_1483[0:0];
  _RAND_1484 = {1{`RANDOM}};
  r_1484 = _RAND_1484[0:0];
  _RAND_1485 = {1{`RANDOM}};
  r_1485 = _RAND_1485[0:0];
  _RAND_1486 = {1{`RANDOM}};
  r_1486 = _RAND_1486[0:0];
  _RAND_1487 = {1{`RANDOM}};
  r_1487 = _RAND_1487[0:0];
  _RAND_1488 = {1{`RANDOM}};
  r_1488 = _RAND_1488[0:0];
  _RAND_1489 = {1{`RANDOM}};
  r_1489 = _RAND_1489[0:0];
  _RAND_1490 = {1{`RANDOM}};
  r_1490 = _RAND_1490[0:0];
  _RAND_1491 = {1{`RANDOM}};
  r_1491 = _RAND_1491[0:0];
  _RAND_1492 = {1{`RANDOM}};
  r_1492 = _RAND_1492[0:0];
  _RAND_1493 = {1{`RANDOM}};
  r_1493 = _RAND_1493[0:0];
  _RAND_1494 = {1{`RANDOM}};
  r_1494 = _RAND_1494[0:0];
  _RAND_1495 = {1{`RANDOM}};
  r_1495 = _RAND_1495[0:0];
  _RAND_1496 = {1{`RANDOM}};
  r_1496 = _RAND_1496[0:0];
  _RAND_1497 = {1{`RANDOM}};
  r_1497 = _RAND_1497[0:0];
  _RAND_1498 = {1{`RANDOM}};
  r_1498 = _RAND_1498[0:0];
  _RAND_1499 = {1{`RANDOM}};
  r_1499 = _RAND_1499[0:0];
  _RAND_1500 = {1{`RANDOM}};
  r_1500 = _RAND_1500[0:0];
  _RAND_1501 = {1{`RANDOM}};
  r_1501 = _RAND_1501[0:0];
  _RAND_1502 = {1{`RANDOM}};
  r_1502 = _RAND_1502[0:0];
  _RAND_1503 = {1{`RANDOM}};
  r_1503 = _RAND_1503[0:0];
  _RAND_1504 = {1{`RANDOM}};
  r_1504 = _RAND_1504[0:0];
  _RAND_1505 = {1{`RANDOM}};
  r_1505 = _RAND_1505[0:0];
  _RAND_1506 = {1{`RANDOM}};
  r_1506 = _RAND_1506[0:0];
  _RAND_1507 = {1{`RANDOM}};
  r_1507 = _RAND_1507[0:0];
  _RAND_1508 = {1{`RANDOM}};
  r_1508 = _RAND_1508[0:0];
  _RAND_1509 = {1{`RANDOM}};
  r_1509 = _RAND_1509[0:0];
  _RAND_1510 = {1{`RANDOM}};
  r_1510 = _RAND_1510[0:0];
  _RAND_1511 = {1{`RANDOM}};
  r_1511 = _RAND_1511[0:0];
  _RAND_1512 = {1{`RANDOM}};
  r_1512 = _RAND_1512[0:0];
  _RAND_1513 = {1{`RANDOM}};
  r_1513 = _RAND_1513[0:0];
  _RAND_1514 = {1{`RANDOM}};
  r_1514 = _RAND_1514[0:0];
  _RAND_1515 = {1{`RANDOM}};
  r_1515 = _RAND_1515[0:0];
  _RAND_1516 = {1{`RANDOM}};
  r_1516 = _RAND_1516[0:0];
  _RAND_1517 = {1{`RANDOM}};
  r_1517 = _RAND_1517[0:0];
  _RAND_1518 = {1{`RANDOM}};
  r_1518 = _RAND_1518[0:0];
  _RAND_1519 = {1{`RANDOM}};
  r_1519 = _RAND_1519[0:0];
  _RAND_1520 = {1{`RANDOM}};
  r_1520 = _RAND_1520[0:0];
  _RAND_1521 = {1{`RANDOM}};
  r_1521 = _RAND_1521[0:0];
  _RAND_1522 = {1{`RANDOM}};
  r_1522 = _RAND_1522[0:0];
  _RAND_1523 = {1{`RANDOM}};
  r_1523 = _RAND_1523[0:0];
  _RAND_1524 = {1{`RANDOM}};
  r_1524 = _RAND_1524[0:0];
  _RAND_1525 = {1{`RANDOM}};
  r_1525 = _RAND_1525[0:0];
  _RAND_1526 = {1{`RANDOM}};
  r_1526 = _RAND_1526[0:0];
  _RAND_1527 = {1{`RANDOM}};
  r_1527 = _RAND_1527[0:0];
  _RAND_1528 = {1{`RANDOM}};
  r_1528 = _RAND_1528[0:0];
  _RAND_1529 = {1{`RANDOM}};
  r_1529 = _RAND_1529[0:0];
  _RAND_1530 = {1{`RANDOM}};
  r_1530 = _RAND_1530[0:0];
  _RAND_1531 = {1{`RANDOM}};
  r_1531 = _RAND_1531[0:0];
  _RAND_1532 = {1{`RANDOM}};
  r_1532 = _RAND_1532[0:0];
  _RAND_1533 = {1{`RANDOM}};
  r_1533 = _RAND_1533[0:0];
  _RAND_1534 = {1{`RANDOM}};
  r_1534 = _RAND_1534[0:0];
  _RAND_1535 = {1{`RANDOM}};
  r_1535 = _RAND_1535[0:0];
  _RAND_1536 = {1{`RANDOM}};
  r_1536 = _RAND_1536[0:0];
  _RAND_1537 = {1{`RANDOM}};
  r_1537 = _RAND_1537[0:0];
  _RAND_1538 = {1{`RANDOM}};
  r_1538 = _RAND_1538[0:0];
  _RAND_1539 = {1{`RANDOM}};
  r_1539 = _RAND_1539[0:0];
  _RAND_1540 = {1{`RANDOM}};
  r_1540 = _RAND_1540[0:0];
  _RAND_1541 = {1{`RANDOM}};
  r_1541 = _RAND_1541[0:0];
  _RAND_1542 = {1{`RANDOM}};
  r_1542 = _RAND_1542[0:0];
  _RAND_1543 = {1{`RANDOM}};
  r_1543 = _RAND_1543[0:0];
  _RAND_1544 = {1{`RANDOM}};
  r_1544 = _RAND_1544[0:0];
  _RAND_1545 = {1{`RANDOM}};
  r_1545 = _RAND_1545[0:0];
  _RAND_1546 = {1{`RANDOM}};
  r_1546 = _RAND_1546[0:0];
  _RAND_1547 = {1{`RANDOM}};
  r_1547 = _RAND_1547[0:0];
  _RAND_1548 = {1{`RANDOM}};
  r_1548 = _RAND_1548[0:0];
  _RAND_1549 = {1{`RANDOM}};
  r_1549 = _RAND_1549[0:0];
  _RAND_1550 = {1{`RANDOM}};
  r_1550 = _RAND_1550[0:0];
  _RAND_1551 = {1{`RANDOM}};
  r_1551 = _RAND_1551[0:0];
  _RAND_1552 = {1{`RANDOM}};
  r_1552 = _RAND_1552[0:0];
  _RAND_1553 = {1{`RANDOM}};
  r_1553 = _RAND_1553[0:0];
  _RAND_1554 = {1{`RANDOM}};
  r_1554 = _RAND_1554[0:0];
  _RAND_1555 = {1{`RANDOM}};
  r_1555 = _RAND_1555[0:0];
  _RAND_1556 = {1{`RANDOM}};
  r_1556 = _RAND_1556[0:0];
  _RAND_1557 = {1{`RANDOM}};
  r_1557 = _RAND_1557[0:0];
  _RAND_1558 = {1{`RANDOM}};
  r_1558 = _RAND_1558[0:0];
  _RAND_1559 = {1{`RANDOM}};
  r_1559 = _RAND_1559[0:0];
  _RAND_1560 = {1{`RANDOM}};
  r_1560 = _RAND_1560[0:0];
  _RAND_1561 = {1{`RANDOM}};
  r_1561 = _RAND_1561[0:0];
  _RAND_1562 = {1{`RANDOM}};
  r_1562 = _RAND_1562[0:0];
  _RAND_1563 = {1{`RANDOM}};
  r_1563 = _RAND_1563[0:0];
  _RAND_1564 = {1{`RANDOM}};
  r_1564 = _RAND_1564[0:0];
  _RAND_1565 = {1{`RANDOM}};
  r_1565 = _RAND_1565[0:0];
  _RAND_1566 = {1{`RANDOM}};
  r_1566 = _RAND_1566[0:0];
  _RAND_1567 = {1{`RANDOM}};
  r_1567 = _RAND_1567[0:0];
  _RAND_1568 = {1{`RANDOM}};
  r_1568 = _RAND_1568[0:0];
  _RAND_1569 = {1{`RANDOM}};
  r_1569 = _RAND_1569[0:0];
  _RAND_1570 = {1{`RANDOM}};
  r_1570 = _RAND_1570[0:0];
  _RAND_1571 = {1{`RANDOM}};
  r_1571 = _RAND_1571[0:0];
  _RAND_1572 = {1{`RANDOM}};
  r_1572 = _RAND_1572[0:0];
  _RAND_1573 = {1{`RANDOM}};
  r_1573 = _RAND_1573[0:0];
  _RAND_1574 = {1{`RANDOM}};
  r_1574 = _RAND_1574[0:0];
  _RAND_1575 = {1{`RANDOM}};
  r_1575 = _RAND_1575[0:0];
  _RAND_1576 = {1{`RANDOM}};
  r_1576 = _RAND_1576[0:0];
  _RAND_1577 = {1{`RANDOM}};
  r_1577 = _RAND_1577[0:0];
  _RAND_1578 = {1{`RANDOM}};
  r_1578 = _RAND_1578[0:0];
  _RAND_1579 = {1{`RANDOM}};
  r_1579 = _RAND_1579[0:0];
  _RAND_1580 = {1{`RANDOM}};
  r_1580 = _RAND_1580[0:0];
  _RAND_1581 = {1{`RANDOM}};
  r_1581 = _RAND_1581[0:0];
  _RAND_1582 = {1{`RANDOM}};
  r_1582 = _RAND_1582[0:0];
  _RAND_1583 = {1{`RANDOM}};
  r_1583 = _RAND_1583[0:0];
  _RAND_1584 = {1{`RANDOM}};
  r_1584 = _RAND_1584[0:0];
  _RAND_1585 = {1{`RANDOM}};
  r_1585 = _RAND_1585[0:0];
  _RAND_1586 = {1{`RANDOM}};
  r_1586 = _RAND_1586[0:0];
  _RAND_1587 = {1{`RANDOM}};
  r_1587 = _RAND_1587[0:0];
  _RAND_1588 = {1{`RANDOM}};
  r_1588 = _RAND_1588[0:0];
  _RAND_1589 = {1{`RANDOM}};
  r_1589 = _RAND_1589[0:0];
  _RAND_1590 = {1{`RANDOM}};
  r_1590 = _RAND_1590[0:0];
  _RAND_1591 = {1{`RANDOM}};
  r_1591 = _RAND_1591[0:0];
  _RAND_1592 = {1{`RANDOM}};
  r_1592 = _RAND_1592[0:0];
  _RAND_1593 = {1{`RANDOM}};
  r_1593 = _RAND_1593[0:0];
  _RAND_1594 = {1{`RANDOM}};
  r_1594 = _RAND_1594[0:0];
  _RAND_1595 = {1{`RANDOM}};
  r_1595 = _RAND_1595[0:0];
  _RAND_1596 = {1{`RANDOM}};
  r_1596 = _RAND_1596[0:0];
  _RAND_1597 = {1{`RANDOM}};
  r_1597 = _RAND_1597[0:0];
  _RAND_1598 = {1{`RANDOM}};
  r_1598 = _RAND_1598[0:0];
  _RAND_1599 = {1{`RANDOM}};
  r_1599 = _RAND_1599[0:0];
  _RAND_1600 = {1{`RANDOM}};
  r_1600 = _RAND_1600[0:0];
  _RAND_1601 = {1{`RANDOM}};
  r_1601 = _RAND_1601[0:0];
  _RAND_1602 = {1{`RANDOM}};
  r_1602 = _RAND_1602[0:0];
  _RAND_1603 = {1{`RANDOM}};
  r_1603 = _RAND_1603[0:0];
  _RAND_1604 = {1{`RANDOM}};
  r_1604 = _RAND_1604[0:0];
  _RAND_1605 = {1{`RANDOM}};
  r_1605 = _RAND_1605[0:0];
  _RAND_1606 = {1{`RANDOM}};
  r_1606 = _RAND_1606[0:0];
  _RAND_1607 = {1{`RANDOM}};
  r_1607 = _RAND_1607[0:0];
  _RAND_1608 = {1{`RANDOM}};
  r_1608 = _RAND_1608[0:0];
  _RAND_1609 = {1{`RANDOM}};
  r_1609 = _RAND_1609[0:0];
  _RAND_1610 = {1{`RANDOM}};
  r_1610 = _RAND_1610[0:0];
  _RAND_1611 = {1{`RANDOM}};
  r_1611 = _RAND_1611[0:0];
  _RAND_1612 = {1{`RANDOM}};
  r_1612 = _RAND_1612[0:0];
  _RAND_1613 = {1{`RANDOM}};
  r_1613 = _RAND_1613[0:0];
  _RAND_1614 = {1{`RANDOM}};
  r_1614 = _RAND_1614[0:0];
  _RAND_1615 = {1{`RANDOM}};
  r_1615 = _RAND_1615[0:0];
  _RAND_1616 = {1{`RANDOM}};
  r_1616 = _RAND_1616[0:0];
  _RAND_1617 = {1{`RANDOM}};
  r_1617 = _RAND_1617[0:0];
  _RAND_1618 = {1{`RANDOM}};
  r_1618 = _RAND_1618[0:0];
  _RAND_1619 = {1{`RANDOM}};
  r_1619 = _RAND_1619[0:0];
  _RAND_1620 = {1{`RANDOM}};
  r_1620 = _RAND_1620[0:0];
  _RAND_1621 = {1{`RANDOM}};
  r_1621 = _RAND_1621[0:0];
  _RAND_1622 = {1{`RANDOM}};
  r_1622 = _RAND_1622[0:0];
  _RAND_1623 = {1{`RANDOM}};
  r_1623 = _RAND_1623[0:0];
  _RAND_1624 = {1{`RANDOM}};
  r_1624 = _RAND_1624[0:0];
  _RAND_1625 = {1{`RANDOM}};
  r_1625 = _RAND_1625[0:0];
  _RAND_1626 = {1{`RANDOM}};
  r_1626 = _RAND_1626[0:0];
  _RAND_1627 = {1{`RANDOM}};
  r_1627 = _RAND_1627[0:0];
  _RAND_1628 = {1{`RANDOM}};
  r_1628 = _RAND_1628[0:0];
  _RAND_1629 = {1{`RANDOM}};
  r_1629 = _RAND_1629[0:0];
  _RAND_1630 = {1{`RANDOM}};
  r_1630 = _RAND_1630[0:0];
  _RAND_1631 = {1{`RANDOM}};
  r_1631 = _RAND_1631[0:0];
  _RAND_1632 = {1{`RANDOM}};
  r_1632 = _RAND_1632[0:0];
  _RAND_1633 = {1{`RANDOM}};
  r_1633 = _RAND_1633[0:0];
  _RAND_1634 = {1{`RANDOM}};
  r_1634 = _RAND_1634[0:0];
  _RAND_1635 = {1{`RANDOM}};
  r_1635 = _RAND_1635[0:0];
  _RAND_1636 = {1{`RANDOM}};
  r_1636 = _RAND_1636[0:0];
  _RAND_1637 = {1{`RANDOM}};
  r_1637 = _RAND_1637[0:0];
  _RAND_1638 = {1{`RANDOM}};
  r_1638 = _RAND_1638[0:0];
  _RAND_1639 = {1{`RANDOM}};
  r_1639 = _RAND_1639[0:0];
  _RAND_1640 = {1{`RANDOM}};
  r_1640 = _RAND_1640[0:0];
  _RAND_1641 = {1{`RANDOM}};
  r_1641 = _RAND_1641[0:0];
  _RAND_1642 = {1{`RANDOM}};
  r_1642 = _RAND_1642[0:0];
  _RAND_1643 = {1{`RANDOM}};
  r_1643 = _RAND_1643[0:0];
  _RAND_1644 = {1{`RANDOM}};
  r_1644 = _RAND_1644[0:0];
  _RAND_1645 = {1{`RANDOM}};
  r_1645 = _RAND_1645[0:0];
  _RAND_1646 = {1{`RANDOM}};
  r_1646 = _RAND_1646[0:0];
  _RAND_1647 = {1{`RANDOM}};
  r_1647 = _RAND_1647[0:0];
  _RAND_1648 = {1{`RANDOM}};
  r_1648 = _RAND_1648[0:0];
  _RAND_1649 = {1{`RANDOM}};
  r_1649 = _RAND_1649[0:0];
  _RAND_1650 = {1{`RANDOM}};
  r_1650 = _RAND_1650[0:0];
  _RAND_1651 = {1{`RANDOM}};
  r_1651 = _RAND_1651[0:0];
  _RAND_1652 = {1{`RANDOM}};
  r_1652 = _RAND_1652[0:0];
  _RAND_1653 = {1{`RANDOM}};
  r_1653 = _RAND_1653[0:0];
  _RAND_1654 = {1{`RANDOM}};
  r_1654 = _RAND_1654[0:0];
  _RAND_1655 = {1{`RANDOM}};
  r_1655 = _RAND_1655[0:0];
  _RAND_1656 = {1{`RANDOM}};
  r_1656 = _RAND_1656[0:0];
  _RAND_1657 = {1{`RANDOM}};
  r_1657 = _RAND_1657[0:0];
  _RAND_1658 = {1{`RANDOM}};
  r_1658 = _RAND_1658[0:0];
  _RAND_1659 = {1{`RANDOM}};
  r_1659 = _RAND_1659[0:0];
  _RAND_1660 = {1{`RANDOM}};
  r_1660 = _RAND_1660[0:0];
  _RAND_1661 = {1{`RANDOM}};
  r_1661 = _RAND_1661[0:0];
  _RAND_1662 = {1{`RANDOM}};
  r_1662 = _RAND_1662[0:0];
  _RAND_1663 = {1{`RANDOM}};
  r_1663 = _RAND_1663[0:0];
  _RAND_1664 = {1{`RANDOM}};
  r_1664 = _RAND_1664[0:0];
  _RAND_1665 = {1{`RANDOM}};
  r_1665 = _RAND_1665[0:0];
  _RAND_1666 = {1{`RANDOM}};
  r_1666 = _RAND_1666[0:0];
  _RAND_1667 = {1{`RANDOM}};
  r_1667 = _RAND_1667[0:0];
  _RAND_1668 = {1{`RANDOM}};
  r_1668 = _RAND_1668[0:0];
  _RAND_1669 = {1{`RANDOM}};
  r_1669 = _RAND_1669[0:0];
  _RAND_1670 = {1{`RANDOM}};
  r_1670 = _RAND_1670[0:0];
  _RAND_1671 = {1{`RANDOM}};
  r_1671 = _RAND_1671[0:0];
  _RAND_1672 = {1{`RANDOM}};
  r_1672 = _RAND_1672[0:0];
  _RAND_1673 = {1{`RANDOM}};
  r_1673 = _RAND_1673[0:0];
  _RAND_1674 = {1{`RANDOM}};
  r_1674 = _RAND_1674[0:0];
  _RAND_1675 = {1{`RANDOM}};
  r_1675 = _RAND_1675[0:0];
  _RAND_1676 = {1{`RANDOM}};
  r_1676 = _RAND_1676[0:0];
  _RAND_1677 = {1{`RANDOM}};
  r_1677 = _RAND_1677[0:0];
  _RAND_1678 = {1{`RANDOM}};
  r_1678 = _RAND_1678[0:0];
  _RAND_1679 = {1{`RANDOM}};
  r_1679 = _RAND_1679[0:0];
  _RAND_1680 = {1{`RANDOM}};
  r_1680 = _RAND_1680[0:0];
  _RAND_1681 = {1{`RANDOM}};
  r_1681 = _RAND_1681[0:0];
  _RAND_1682 = {1{`RANDOM}};
  r_1682 = _RAND_1682[0:0];
  _RAND_1683 = {1{`RANDOM}};
  r_1683 = _RAND_1683[0:0];
  _RAND_1684 = {1{`RANDOM}};
  r_1684 = _RAND_1684[0:0];
  _RAND_1685 = {1{`RANDOM}};
  r_1685 = _RAND_1685[0:0];
  _RAND_1686 = {1{`RANDOM}};
  r_1686 = _RAND_1686[0:0];
  _RAND_1687 = {1{`RANDOM}};
  r_1687 = _RAND_1687[0:0];
  _RAND_1688 = {1{`RANDOM}};
  r_1688 = _RAND_1688[0:0];
  _RAND_1689 = {1{`RANDOM}};
  r_1689 = _RAND_1689[0:0];
  _RAND_1690 = {1{`RANDOM}};
  r_1690 = _RAND_1690[0:0];
  _RAND_1691 = {1{`RANDOM}};
  r_1691 = _RAND_1691[0:0];
  _RAND_1692 = {1{`RANDOM}};
  r_1692 = _RAND_1692[0:0];
  _RAND_1693 = {1{`RANDOM}};
  r_1693 = _RAND_1693[0:0];
  _RAND_1694 = {1{`RANDOM}};
  r_1694 = _RAND_1694[0:0];
  _RAND_1695 = {1{`RANDOM}};
  r_1695 = _RAND_1695[0:0];
  _RAND_1696 = {1{`RANDOM}};
  r_1696 = _RAND_1696[0:0];
  _RAND_1697 = {1{`RANDOM}};
  r_1697 = _RAND_1697[0:0];
  _RAND_1698 = {1{`RANDOM}};
  r_1698 = _RAND_1698[0:0];
  _RAND_1699 = {1{`RANDOM}};
  r_1699 = _RAND_1699[0:0];
  _RAND_1700 = {1{`RANDOM}};
  r_1700 = _RAND_1700[0:0];
  _RAND_1701 = {1{`RANDOM}};
  r_1701 = _RAND_1701[0:0];
  _RAND_1702 = {1{`RANDOM}};
  r_1702 = _RAND_1702[0:0];
  _RAND_1703 = {1{`RANDOM}};
  r_1703 = _RAND_1703[0:0];
  _RAND_1704 = {1{`RANDOM}};
  r_1704 = _RAND_1704[0:0];
  _RAND_1705 = {1{`RANDOM}};
  r_1705 = _RAND_1705[0:0];
  _RAND_1706 = {1{`RANDOM}};
  r_1706 = _RAND_1706[0:0];
  _RAND_1707 = {1{`RANDOM}};
  r_1707 = _RAND_1707[0:0];
  _RAND_1708 = {1{`RANDOM}};
  r_1708 = _RAND_1708[0:0];
  _RAND_1709 = {1{`RANDOM}};
  r_1709 = _RAND_1709[0:0];
  _RAND_1710 = {1{`RANDOM}};
  r_1710 = _RAND_1710[0:0];
  _RAND_1711 = {1{`RANDOM}};
  r_1711 = _RAND_1711[0:0];
  _RAND_1712 = {1{`RANDOM}};
  r_1712 = _RAND_1712[0:0];
  _RAND_1713 = {1{`RANDOM}};
  r_1713 = _RAND_1713[0:0];
  _RAND_1714 = {1{`RANDOM}};
  r_1714 = _RAND_1714[0:0];
  _RAND_1715 = {1{`RANDOM}};
  r_1715 = _RAND_1715[0:0];
  _RAND_1716 = {1{`RANDOM}};
  r_1716 = _RAND_1716[0:0];
  _RAND_1717 = {1{`RANDOM}};
  r_1717 = _RAND_1717[0:0];
  _RAND_1718 = {1{`RANDOM}};
  r_1718 = _RAND_1718[0:0];
  _RAND_1719 = {1{`RANDOM}};
  r_1719 = _RAND_1719[0:0];
  _RAND_1720 = {1{`RANDOM}};
  r_1720 = _RAND_1720[0:0];
  _RAND_1721 = {1{`RANDOM}};
  r_1721 = _RAND_1721[0:0];
  _RAND_1722 = {1{`RANDOM}};
  r_1722 = _RAND_1722[0:0];
  _RAND_1723 = {1{`RANDOM}};
  r_1723 = _RAND_1723[0:0];
  _RAND_1724 = {1{`RANDOM}};
  r_1724 = _RAND_1724[0:0];
  _RAND_1725 = {1{`RANDOM}};
  r_1725 = _RAND_1725[0:0];
  _RAND_1726 = {1{`RANDOM}};
  r_1726 = _RAND_1726[0:0];
  _RAND_1727 = {1{`RANDOM}};
  r_1727 = _RAND_1727[0:0];
  _RAND_1728 = {1{`RANDOM}};
  r_1728 = _RAND_1728[0:0];
  _RAND_1729 = {1{`RANDOM}};
  r_1729 = _RAND_1729[0:0];
  _RAND_1730 = {1{`RANDOM}};
  r_1730 = _RAND_1730[0:0];
  _RAND_1731 = {1{`RANDOM}};
  r_1731 = _RAND_1731[0:0];
  _RAND_1732 = {1{`RANDOM}};
  r_1732 = _RAND_1732[0:0];
  _RAND_1733 = {1{`RANDOM}};
  r_1733 = _RAND_1733[0:0];
  _RAND_1734 = {1{`RANDOM}};
  r_1734 = _RAND_1734[0:0];
  _RAND_1735 = {1{`RANDOM}};
  r_1735 = _RAND_1735[0:0];
  _RAND_1736 = {1{`RANDOM}};
  r_1736 = _RAND_1736[0:0];
  _RAND_1737 = {1{`RANDOM}};
  r_1737 = _RAND_1737[0:0];
  _RAND_1738 = {1{`RANDOM}};
  r_1738 = _RAND_1738[0:0];
  _RAND_1739 = {1{`RANDOM}};
  r_1739 = _RAND_1739[0:0];
  _RAND_1740 = {1{`RANDOM}};
  r_1740 = _RAND_1740[0:0];
  _RAND_1741 = {1{`RANDOM}};
  r_1741 = _RAND_1741[0:0];
  _RAND_1742 = {1{`RANDOM}};
  r_1742 = _RAND_1742[0:0];
  _RAND_1743 = {1{`RANDOM}};
  r_1743 = _RAND_1743[0:0];
  _RAND_1744 = {1{`RANDOM}};
  r_1744 = _RAND_1744[0:0];
  _RAND_1745 = {1{`RANDOM}};
  r_1745 = _RAND_1745[0:0];
  _RAND_1746 = {1{`RANDOM}};
  r_1746 = _RAND_1746[0:0];
  _RAND_1747 = {1{`RANDOM}};
  r_1747 = _RAND_1747[0:0];
  _RAND_1748 = {1{`RANDOM}};
  r_1748 = _RAND_1748[0:0];
  _RAND_1749 = {1{`RANDOM}};
  r_1749 = _RAND_1749[0:0];
  _RAND_1750 = {1{`RANDOM}};
  r_1750 = _RAND_1750[0:0];
  _RAND_1751 = {1{`RANDOM}};
  r_1751 = _RAND_1751[0:0];
  _RAND_1752 = {1{`RANDOM}};
  r_1752 = _RAND_1752[0:0];
  _RAND_1753 = {1{`RANDOM}};
  r_1753 = _RAND_1753[0:0];
  _RAND_1754 = {1{`RANDOM}};
  r_1754 = _RAND_1754[0:0];
  _RAND_1755 = {1{`RANDOM}};
  r_1755 = _RAND_1755[0:0];
  _RAND_1756 = {1{`RANDOM}};
  r_1756 = _RAND_1756[0:0];
  _RAND_1757 = {1{`RANDOM}};
  r_1757 = _RAND_1757[0:0];
  _RAND_1758 = {1{`RANDOM}};
  r_1758 = _RAND_1758[0:0];
  _RAND_1759 = {1{`RANDOM}};
  r_1759 = _RAND_1759[0:0];
  _RAND_1760 = {1{`RANDOM}};
  r_1760 = _RAND_1760[0:0];
  _RAND_1761 = {1{`RANDOM}};
  r_1761 = _RAND_1761[0:0];
  _RAND_1762 = {1{`RANDOM}};
  r_1762 = _RAND_1762[0:0];
  _RAND_1763 = {1{`RANDOM}};
  r_1763 = _RAND_1763[0:0];
  _RAND_1764 = {1{`RANDOM}};
  r_1764 = _RAND_1764[0:0];
  _RAND_1765 = {1{`RANDOM}};
  r_1765 = _RAND_1765[0:0];
  _RAND_1766 = {1{`RANDOM}};
  r_1766 = _RAND_1766[0:0];
  _RAND_1767 = {1{`RANDOM}};
  r_1767 = _RAND_1767[0:0];
  _RAND_1768 = {1{`RANDOM}};
  r_1768 = _RAND_1768[0:0];
  _RAND_1769 = {1{`RANDOM}};
  r_1769 = _RAND_1769[0:0];
  _RAND_1770 = {1{`RANDOM}};
  r_1770 = _RAND_1770[0:0];
  _RAND_1771 = {1{`RANDOM}};
  r_1771 = _RAND_1771[0:0];
  _RAND_1772 = {1{`RANDOM}};
  r_1772 = _RAND_1772[0:0];
  _RAND_1773 = {1{`RANDOM}};
  r_1773 = _RAND_1773[0:0];
  _RAND_1774 = {1{`RANDOM}};
  r_1774 = _RAND_1774[0:0];
  _RAND_1775 = {1{`RANDOM}};
  r_1775 = _RAND_1775[0:0];
  _RAND_1776 = {1{`RANDOM}};
  r_1776 = _RAND_1776[0:0];
  _RAND_1777 = {1{`RANDOM}};
  r_1777 = _RAND_1777[0:0];
  _RAND_1778 = {1{`RANDOM}};
  r_1778 = _RAND_1778[0:0];
  _RAND_1779 = {1{`RANDOM}};
  r_1779 = _RAND_1779[0:0];
  _RAND_1780 = {1{`RANDOM}};
  r_1780 = _RAND_1780[0:0];
  _RAND_1781 = {1{`RANDOM}};
  r_1781 = _RAND_1781[0:0];
  _RAND_1782 = {1{`RANDOM}};
  r_1782 = _RAND_1782[0:0];
  _RAND_1783 = {1{`RANDOM}};
  r_1783 = _RAND_1783[0:0];
  _RAND_1784 = {1{`RANDOM}};
  r_1784 = _RAND_1784[0:0];
  _RAND_1785 = {1{`RANDOM}};
  r_1785 = _RAND_1785[0:0];
  _RAND_1786 = {1{`RANDOM}};
  r_1786 = _RAND_1786[0:0];
  _RAND_1787 = {1{`RANDOM}};
  r_1787 = _RAND_1787[0:0];
  _RAND_1788 = {1{`RANDOM}};
  r_1788 = _RAND_1788[0:0];
  _RAND_1789 = {1{`RANDOM}};
  r_1789 = _RAND_1789[0:0];
  _RAND_1790 = {1{`RANDOM}};
  r_1790 = _RAND_1790[0:0];
  _RAND_1791 = {1{`RANDOM}};
  r_1791 = _RAND_1791[0:0];
  _RAND_1792 = {1{`RANDOM}};
  r_1792 = _RAND_1792[0:0];
  _RAND_1793 = {1{`RANDOM}};
  r_1793 = _RAND_1793[0:0];
  _RAND_1794 = {1{`RANDOM}};
  r_1794 = _RAND_1794[0:0];
  _RAND_1795 = {1{`RANDOM}};
  r_1795 = _RAND_1795[0:0];
  _RAND_1796 = {1{`RANDOM}};
  r_1796 = _RAND_1796[0:0];
  _RAND_1797 = {1{`RANDOM}};
  r_1797 = _RAND_1797[0:0];
  _RAND_1798 = {1{`RANDOM}};
  r_1798 = _RAND_1798[0:0];
  _RAND_1799 = {1{`RANDOM}};
  r_1799 = _RAND_1799[0:0];
  _RAND_1800 = {1{`RANDOM}};
  r_1800 = _RAND_1800[0:0];
  _RAND_1801 = {1{`RANDOM}};
  r_1801 = _RAND_1801[0:0];
  _RAND_1802 = {1{`RANDOM}};
  r_1802 = _RAND_1802[0:0];
  _RAND_1803 = {1{`RANDOM}};
  r_1803 = _RAND_1803[0:0];
  _RAND_1804 = {1{`RANDOM}};
  r_1804 = _RAND_1804[0:0];
  _RAND_1805 = {1{`RANDOM}};
  r_1805 = _RAND_1805[0:0];
  _RAND_1806 = {1{`RANDOM}};
  r_1806 = _RAND_1806[0:0];
  _RAND_1807 = {1{`RANDOM}};
  r_1807 = _RAND_1807[0:0];
  _RAND_1808 = {1{`RANDOM}};
  r_1808 = _RAND_1808[0:0];
  _RAND_1809 = {1{`RANDOM}};
  r_1809 = _RAND_1809[0:0];
  _RAND_1810 = {1{`RANDOM}};
  r_1810 = _RAND_1810[0:0];
  _RAND_1811 = {1{`RANDOM}};
  r_1811 = _RAND_1811[0:0];
  _RAND_1812 = {1{`RANDOM}};
  r_1812 = _RAND_1812[0:0];
  _RAND_1813 = {1{`RANDOM}};
  r_1813 = _RAND_1813[0:0];
  _RAND_1814 = {1{`RANDOM}};
  r_1814 = _RAND_1814[0:0];
  _RAND_1815 = {1{`RANDOM}};
  r_1815 = _RAND_1815[0:0];
  _RAND_1816 = {1{`RANDOM}};
  r_1816 = _RAND_1816[0:0];
  _RAND_1817 = {1{`RANDOM}};
  r_1817 = _RAND_1817[0:0];
  _RAND_1818 = {1{`RANDOM}};
  r_1818 = _RAND_1818[0:0];
  _RAND_1819 = {1{`RANDOM}};
  r_1819 = _RAND_1819[0:0];
  _RAND_1820 = {1{`RANDOM}};
  r_1820 = _RAND_1820[0:0];
  _RAND_1821 = {1{`RANDOM}};
  r_1821 = _RAND_1821[0:0];
  _RAND_1822 = {1{`RANDOM}};
  r_1822 = _RAND_1822[0:0];
  _RAND_1823 = {1{`RANDOM}};
  r_1823 = _RAND_1823[0:0];
  _RAND_1824 = {1{`RANDOM}};
  r_1824 = _RAND_1824[0:0];
  _RAND_1825 = {1{`RANDOM}};
  r_1825 = _RAND_1825[0:0];
  _RAND_1826 = {1{`RANDOM}};
  r_1826 = _RAND_1826[0:0];
  _RAND_1827 = {1{`RANDOM}};
  r_1827 = _RAND_1827[0:0];
  _RAND_1828 = {1{`RANDOM}};
  r_1828 = _RAND_1828[0:0];
  _RAND_1829 = {1{`RANDOM}};
  r_1829 = _RAND_1829[0:0];
  _RAND_1830 = {1{`RANDOM}};
  r_1830 = _RAND_1830[0:0];
  _RAND_1831 = {1{`RANDOM}};
  r_1831 = _RAND_1831[0:0];
  _RAND_1832 = {1{`RANDOM}};
  r_1832 = _RAND_1832[0:0];
  _RAND_1833 = {1{`RANDOM}};
  r_1833 = _RAND_1833[0:0];
  _RAND_1834 = {1{`RANDOM}};
  r_1834 = _RAND_1834[0:0];
  _RAND_1835 = {1{`RANDOM}};
  r_1835 = _RAND_1835[0:0];
  _RAND_1836 = {1{`RANDOM}};
  r_1836 = _RAND_1836[0:0];
  _RAND_1837 = {1{`RANDOM}};
  r_1837 = _RAND_1837[0:0];
  _RAND_1838 = {1{`RANDOM}};
  r_1838 = _RAND_1838[0:0];
  _RAND_1839 = {1{`RANDOM}};
  r_1839 = _RAND_1839[0:0];
  _RAND_1840 = {1{`RANDOM}};
  r_1840 = _RAND_1840[0:0];
  _RAND_1841 = {1{`RANDOM}};
  r_1841 = _RAND_1841[0:0];
  _RAND_1842 = {1{`RANDOM}};
  r_1842 = _RAND_1842[0:0];
  _RAND_1843 = {1{`RANDOM}};
  r_1843 = _RAND_1843[0:0];
  _RAND_1844 = {1{`RANDOM}};
  r_1844 = _RAND_1844[0:0];
  _RAND_1845 = {1{`RANDOM}};
  r_1845 = _RAND_1845[0:0];
  _RAND_1846 = {1{`RANDOM}};
  r_1846 = _RAND_1846[0:0];
  _RAND_1847 = {1{`RANDOM}};
  r_1847 = _RAND_1847[0:0];
  _RAND_1848 = {1{`RANDOM}};
  r_1848 = _RAND_1848[0:0];
  _RAND_1849 = {1{`RANDOM}};
  r_1849 = _RAND_1849[0:0];
  _RAND_1850 = {1{`RANDOM}};
  r_1850 = _RAND_1850[0:0];
  _RAND_1851 = {1{`RANDOM}};
  r_1851 = _RAND_1851[0:0];
  _RAND_1852 = {1{`RANDOM}};
  r_1852 = _RAND_1852[0:0];
  _RAND_1853 = {1{`RANDOM}};
  r_1853 = _RAND_1853[0:0];
  _RAND_1854 = {1{`RANDOM}};
  r_1854 = _RAND_1854[0:0];
  _RAND_1855 = {1{`RANDOM}};
  r_1855 = _RAND_1855[0:0];
  _RAND_1856 = {1{`RANDOM}};
  r_1856 = _RAND_1856[0:0];
  _RAND_1857 = {1{`RANDOM}};
  r_1857 = _RAND_1857[0:0];
  _RAND_1858 = {1{`RANDOM}};
  r_1858 = _RAND_1858[0:0];
  _RAND_1859 = {1{`RANDOM}};
  r_1859 = _RAND_1859[0:0];
  _RAND_1860 = {1{`RANDOM}};
  r_1860 = _RAND_1860[0:0];
  _RAND_1861 = {1{`RANDOM}};
  r_1861 = _RAND_1861[0:0];
  _RAND_1862 = {1{`RANDOM}};
  r_1862 = _RAND_1862[0:0];
  _RAND_1863 = {1{`RANDOM}};
  r_1863 = _RAND_1863[0:0];
  _RAND_1864 = {1{`RANDOM}};
  r_1864 = _RAND_1864[0:0];
  _RAND_1865 = {1{`RANDOM}};
  r_1865 = _RAND_1865[0:0];
  _RAND_1866 = {1{`RANDOM}};
  r_1866 = _RAND_1866[0:0];
  _RAND_1867 = {1{`RANDOM}};
  r_1867 = _RAND_1867[0:0];
  _RAND_1868 = {1{`RANDOM}};
  r_1868 = _RAND_1868[0:0];
  _RAND_1869 = {1{`RANDOM}};
  r_1869 = _RAND_1869[0:0];
  _RAND_1870 = {1{`RANDOM}};
  r_1870 = _RAND_1870[0:0];
  _RAND_1871 = {1{`RANDOM}};
  r_1871 = _RAND_1871[0:0];
  _RAND_1872 = {1{`RANDOM}};
  r_1872 = _RAND_1872[0:0];
  _RAND_1873 = {1{`RANDOM}};
  r_1873 = _RAND_1873[0:0];
  _RAND_1874 = {1{`RANDOM}};
  r_1874 = _RAND_1874[0:0];
  _RAND_1875 = {1{`RANDOM}};
  r_1875 = _RAND_1875[0:0];
  _RAND_1876 = {1{`RANDOM}};
  r_1876 = _RAND_1876[0:0];
  _RAND_1877 = {1{`RANDOM}};
  r_1877 = _RAND_1877[0:0];
  _RAND_1878 = {1{`RANDOM}};
  r_1878 = _RAND_1878[0:0];
  _RAND_1879 = {1{`RANDOM}};
  r_1879 = _RAND_1879[0:0];
  _RAND_1880 = {1{`RANDOM}};
  r_1880 = _RAND_1880[0:0];
  _RAND_1881 = {1{`RANDOM}};
  r_1881 = _RAND_1881[0:0];
  _RAND_1882 = {1{`RANDOM}};
  r_1882 = _RAND_1882[0:0];
  _RAND_1883 = {1{`RANDOM}};
  r_1883 = _RAND_1883[0:0];
  _RAND_1884 = {1{`RANDOM}};
  r_1884 = _RAND_1884[0:0];
  _RAND_1885 = {1{`RANDOM}};
  r_1885 = _RAND_1885[0:0];
  _RAND_1886 = {1{`RANDOM}};
  r_1886 = _RAND_1886[0:0];
  _RAND_1887 = {1{`RANDOM}};
  r_1887 = _RAND_1887[0:0];
  _RAND_1888 = {1{`RANDOM}};
  r_1888 = _RAND_1888[0:0];
  _RAND_1889 = {1{`RANDOM}};
  r_1889 = _RAND_1889[0:0];
  _RAND_1890 = {1{`RANDOM}};
  r_1890 = _RAND_1890[0:0];
  _RAND_1891 = {1{`RANDOM}};
  r_1891 = _RAND_1891[0:0];
  _RAND_1892 = {1{`RANDOM}};
  r_1892 = _RAND_1892[0:0];
  _RAND_1893 = {1{`RANDOM}};
  r_1893 = _RAND_1893[0:0];
  _RAND_1894 = {1{`RANDOM}};
  r_1894 = _RAND_1894[0:0];
  _RAND_1895 = {1{`RANDOM}};
  r_1895 = _RAND_1895[0:0];
  _RAND_1896 = {1{`RANDOM}};
  r_1896 = _RAND_1896[0:0];
  _RAND_1897 = {1{`RANDOM}};
  r_1897 = _RAND_1897[0:0];
  _RAND_1898 = {1{`RANDOM}};
  r_1898 = _RAND_1898[0:0];
  _RAND_1899 = {1{`RANDOM}};
  r_1899 = _RAND_1899[0:0];
  _RAND_1900 = {1{`RANDOM}};
  r_1900 = _RAND_1900[0:0];
  _RAND_1901 = {1{`RANDOM}};
  r_1901 = _RAND_1901[0:0];
  _RAND_1902 = {1{`RANDOM}};
  r_1902 = _RAND_1902[0:0];
  _RAND_1903 = {1{`RANDOM}};
  r_1903 = _RAND_1903[0:0];
  _RAND_1904 = {1{`RANDOM}};
  r_1904 = _RAND_1904[0:0];
  _RAND_1905 = {1{`RANDOM}};
  r_1905 = _RAND_1905[0:0];
  _RAND_1906 = {1{`RANDOM}};
  r_1906 = _RAND_1906[0:0];
  _RAND_1907 = {1{`RANDOM}};
  r_1907 = _RAND_1907[0:0];
  _RAND_1908 = {1{`RANDOM}};
  r_1908 = _RAND_1908[0:0];
  _RAND_1909 = {1{`RANDOM}};
  r_1909 = _RAND_1909[0:0];
  _RAND_1910 = {1{`RANDOM}};
  r_1910 = _RAND_1910[0:0];
  _RAND_1911 = {1{`RANDOM}};
  r_1911 = _RAND_1911[0:0];
  _RAND_1912 = {1{`RANDOM}};
  r_1912 = _RAND_1912[0:0];
  _RAND_1913 = {1{`RANDOM}};
  r_1913 = _RAND_1913[0:0];
  _RAND_1914 = {1{`RANDOM}};
  r_1914 = _RAND_1914[0:0];
  _RAND_1915 = {1{`RANDOM}};
  r_1915 = _RAND_1915[0:0];
  _RAND_1916 = {1{`RANDOM}};
  r_1916 = _RAND_1916[0:0];
  _RAND_1917 = {1{`RANDOM}};
  r_1917 = _RAND_1917[0:0];
  _RAND_1918 = {1{`RANDOM}};
  r_1918 = _RAND_1918[0:0];
  _RAND_1919 = {1{`RANDOM}};
  r_1919 = _RAND_1919[0:0];
  _RAND_1920 = {1{`RANDOM}};
  r_1920 = _RAND_1920[0:0];
  _RAND_1921 = {1{`RANDOM}};
  r_1921 = _RAND_1921[0:0];
  _RAND_1922 = {1{`RANDOM}};
  r_1922 = _RAND_1922[0:0];
  _RAND_1923 = {1{`RANDOM}};
  r_1923 = _RAND_1923[0:0];
  _RAND_1924 = {1{`RANDOM}};
  r_1924 = _RAND_1924[0:0];
  _RAND_1925 = {1{`RANDOM}};
  r_1925 = _RAND_1925[0:0];
  _RAND_1926 = {1{`RANDOM}};
  r_1926 = _RAND_1926[0:0];
  _RAND_1927 = {1{`RANDOM}};
  r_1927 = _RAND_1927[0:0];
  _RAND_1928 = {1{`RANDOM}};
  r_1928 = _RAND_1928[0:0];
  _RAND_1929 = {1{`RANDOM}};
  r_1929 = _RAND_1929[0:0];
  _RAND_1930 = {1{`RANDOM}};
  r_1930 = _RAND_1930[0:0];
  _RAND_1931 = {1{`RANDOM}};
  r_1931 = _RAND_1931[0:0];
  _RAND_1932 = {1{`RANDOM}};
  r_1932 = _RAND_1932[0:0];
  _RAND_1933 = {1{`RANDOM}};
  r_1933 = _RAND_1933[0:0];
  _RAND_1934 = {1{`RANDOM}};
  r_1934 = _RAND_1934[0:0];
  _RAND_1935 = {1{`RANDOM}};
  r_1935 = _RAND_1935[0:0];
  _RAND_1936 = {1{`RANDOM}};
  r_1936 = _RAND_1936[0:0];
  _RAND_1937 = {1{`RANDOM}};
  r_1937 = _RAND_1937[0:0];
  _RAND_1938 = {1{`RANDOM}};
  r_1938 = _RAND_1938[0:0];
  _RAND_1939 = {1{`RANDOM}};
  r_1939 = _RAND_1939[0:0];
  _RAND_1940 = {1{`RANDOM}};
  r_1940 = _RAND_1940[0:0];
  _RAND_1941 = {1{`RANDOM}};
  r_1941 = _RAND_1941[0:0];
  _RAND_1942 = {1{`RANDOM}};
  r_1942 = _RAND_1942[0:0];
  _RAND_1943 = {1{`RANDOM}};
  r_1943 = _RAND_1943[0:0];
  _RAND_1944 = {1{`RANDOM}};
  r_1944 = _RAND_1944[0:0];
  _RAND_1945 = {1{`RANDOM}};
  r_1945 = _RAND_1945[0:0];
  _RAND_1946 = {1{`RANDOM}};
  r_1946 = _RAND_1946[0:0];
  _RAND_1947 = {1{`RANDOM}};
  r_1947 = _RAND_1947[0:0];
  _RAND_1948 = {1{`RANDOM}};
  r_1948 = _RAND_1948[0:0];
  _RAND_1949 = {1{`RANDOM}};
  r_1949 = _RAND_1949[0:0];
  _RAND_1950 = {1{`RANDOM}};
  r_1950 = _RAND_1950[0:0];
  _RAND_1951 = {1{`RANDOM}};
  r_1951 = _RAND_1951[0:0];
  _RAND_1952 = {1{`RANDOM}};
  r_1952 = _RAND_1952[0:0];
  _RAND_1953 = {1{`RANDOM}};
  r_1953 = _RAND_1953[0:0];
  _RAND_1954 = {1{`RANDOM}};
  r_1954 = _RAND_1954[0:0];
  _RAND_1955 = {1{`RANDOM}};
  r_1955 = _RAND_1955[0:0];
  _RAND_1956 = {1{`RANDOM}};
  r_1956 = _RAND_1956[0:0];
  _RAND_1957 = {1{`RANDOM}};
  r_1957 = _RAND_1957[0:0];
  _RAND_1958 = {1{`RANDOM}};
  r_1958 = _RAND_1958[0:0];
  _RAND_1959 = {1{`RANDOM}};
  r_1959 = _RAND_1959[0:0];
  _RAND_1960 = {1{`RANDOM}};
  r_1960 = _RAND_1960[0:0];
  _RAND_1961 = {1{`RANDOM}};
  r_1961 = _RAND_1961[0:0];
  _RAND_1962 = {1{`RANDOM}};
  r_1962 = _RAND_1962[0:0];
  _RAND_1963 = {1{`RANDOM}};
  r_1963 = _RAND_1963[0:0];
  _RAND_1964 = {1{`RANDOM}};
  r_1964 = _RAND_1964[0:0];
  _RAND_1965 = {1{`RANDOM}};
  r_1965 = _RAND_1965[0:0];
  _RAND_1966 = {1{`RANDOM}};
  r_1966 = _RAND_1966[0:0];
  _RAND_1967 = {1{`RANDOM}};
  r_1967 = _RAND_1967[0:0];
  _RAND_1968 = {1{`RANDOM}};
  r_1968 = _RAND_1968[0:0];
  _RAND_1969 = {1{`RANDOM}};
  r_1969 = _RAND_1969[0:0];
  _RAND_1970 = {1{`RANDOM}};
  r_1970 = _RAND_1970[0:0];
  _RAND_1971 = {1{`RANDOM}};
  r_1971 = _RAND_1971[0:0];
  _RAND_1972 = {1{`RANDOM}};
  r_1972 = _RAND_1972[0:0];
  _RAND_1973 = {1{`RANDOM}};
  r_1973 = _RAND_1973[0:0];
  _RAND_1974 = {1{`RANDOM}};
  r_1974 = _RAND_1974[0:0];
  _RAND_1975 = {1{`RANDOM}};
  r_1975 = _RAND_1975[0:0];
  _RAND_1976 = {1{`RANDOM}};
  r_1976 = _RAND_1976[0:0];
  _RAND_1977 = {1{`RANDOM}};
  r_1977 = _RAND_1977[0:0];
  _RAND_1978 = {1{`RANDOM}};
  r_1978 = _RAND_1978[0:0];
  _RAND_1979 = {1{`RANDOM}};
  r_1979 = _RAND_1979[0:0];
  _RAND_1980 = {1{`RANDOM}};
  r_1980 = _RAND_1980[0:0];
  _RAND_1981 = {1{`RANDOM}};
  r_1981 = _RAND_1981[0:0];
  _RAND_1982 = {1{`RANDOM}};
  r_1982 = _RAND_1982[0:0];
  _RAND_1983 = {1{`RANDOM}};
  r_1983 = _RAND_1983[0:0];
  _RAND_1984 = {1{`RANDOM}};
  r_1984 = _RAND_1984[0:0];
  _RAND_1985 = {1{`RANDOM}};
  r_1985 = _RAND_1985[0:0];
  _RAND_1986 = {1{`RANDOM}};
  r_1986 = _RAND_1986[0:0];
  _RAND_1987 = {1{`RANDOM}};
  r_1987 = _RAND_1987[0:0];
  _RAND_1988 = {1{`RANDOM}};
  r_1988 = _RAND_1988[0:0];
  _RAND_1989 = {1{`RANDOM}};
  r_1989 = _RAND_1989[0:0];
  _RAND_1990 = {1{`RANDOM}};
  r_1990 = _RAND_1990[0:0];
  _RAND_1991 = {1{`RANDOM}};
  r_1991 = _RAND_1991[0:0];
  _RAND_1992 = {1{`RANDOM}};
  r_1992 = _RAND_1992[0:0];
  _RAND_1993 = {1{`RANDOM}};
  r_1993 = _RAND_1993[0:0];
  _RAND_1994 = {1{`RANDOM}};
  r_1994 = _RAND_1994[0:0];
  _RAND_1995 = {1{`RANDOM}};
  r_1995 = _RAND_1995[0:0];
  _RAND_1996 = {1{`RANDOM}};
  r_1996 = _RAND_1996[0:0];
  _RAND_1997 = {1{`RANDOM}};
  r_1997 = _RAND_1997[0:0];
  _RAND_1998 = {1{`RANDOM}};
  r_1998 = _RAND_1998[0:0];
  _RAND_1999 = {1{`RANDOM}};
  r_1999 = _RAND_1999[0:0];
  _RAND_2000 = {1{`RANDOM}};
  r_2000 = _RAND_2000[0:0];
  _RAND_2001 = {1{`RANDOM}};
  r_2001 = _RAND_2001[0:0];
  _RAND_2002 = {1{`RANDOM}};
  r_2002 = _RAND_2002[0:0];
  _RAND_2003 = {1{`RANDOM}};
  r_2003 = _RAND_2003[0:0];
  _RAND_2004 = {1{`RANDOM}};
  r_2004 = _RAND_2004[0:0];
  _RAND_2005 = {1{`RANDOM}};
  r_2005 = _RAND_2005[0:0];
  _RAND_2006 = {1{`RANDOM}};
  r_2006 = _RAND_2006[0:0];
  _RAND_2007 = {1{`RANDOM}};
  r_2007 = _RAND_2007[0:0];
  _RAND_2008 = {1{`RANDOM}};
  r_2008 = _RAND_2008[0:0];
  _RAND_2009 = {1{`RANDOM}};
  r_2009 = _RAND_2009[0:0];
  _RAND_2010 = {1{`RANDOM}};
  r_2010 = _RAND_2010[0:0];
  _RAND_2011 = {1{`RANDOM}};
  r_2011 = _RAND_2011[0:0];
  _RAND_2012 = {1{`RANDOM}};
  r_2012 = _RAND_2012[0:0];
  _RAND_2013 = {1{`RANDOM}};
  r_2013 = _RAND_2013[0:0];
  _RAND_2014 = {1{`RANDOM}};
  r_2014 = _RAND_2014[0:0];
  _RAND_2015 = {1{`RANDOM}};
  r_2015 = _RAND_2015[0:0];
  _RAND_2016 = {1{`RANDOM}};
  r_2016 = _RAND_2016[0:0];
  _RAND_2017 = {1{`RANDOM}};
  r_2017 = _RAND_2017[0:0];
  _RAND_2018 = {1{`RANDOM}};
  r_2018 = _RAND_2018[0:0];
  _RAND_2019 = {1{`RANDOM}};
  r_2019 = _RAND_2019[0:0];
  _RAND_2020 = {1{`RANDOM}};
  r_2020 = _RAND_2020[0:0];
  _RAND_2021 = {1{`RANDOM}};
  r_2021 = _RAND_2021[0:0];
  _RAND_2022 = {1{`RANDOM}};
  r_2022 = _RAND_2022[0:0];
  _RAND_2023 = {1{`RANDOM}};
  r_2023 = _RAND_2023[0:0];
  _RAND_2024 = {1{`RANDOM}};
  r_2024 = _RAND_2024[0:0];
  _RAND_2025 = {1{`RANDOM}};
  r_2025 = _RAND_2025[0:0];
  _RAND_2026 = {1{`RANDOM}};
  r_2026 = _RAND_2026[0:0];
  _RAND_2027 = {1{`RANDOM}};
  r_2027 = _RAND_2027[0:0];
  _RAND_2028 = {1{`RANDOM}};
  r_2028 = _RAND_2028[0:0];
  _RAND_2029 = {1{`RANDOM}};
  r_2029 = _RAND_2029[0:0];
  _RAND_2030 = {1{`RANDOM}};
  r_2030 = _RAND_2030[0:0];
  _RAND_2031 = {1{`RANDOM}};
  r_2031 = _RAND_2031[0:0];
  _RAND_2032 = {1{`RANDOM}};
  r_2032 = _RAND_2032[0:0];
  _RAND_2033 = {1{`RANDOM}};
  r_2033 = _RAND_2033[0:0];
  _RAND_2034 = {1{`RANDOM}};
  r_2034 = _RAND_2034[0:0];
  _RAND_2035 = {1{`RANDOM}};
  r_2035 = _RAND_2035[0:0];
  _RAND_2036 = {1{`RANDOM}};
  r_2036 = _RAND_2036[0:0];
  _RAND_2037 = {1{`RANDOM}};
  r_2037 = _RAND_2037[0:0];
  _RAND_2038 = {1{`RANDOM}};
  r_2038 = _RAND_2038[0:0];
  _RAND_2039 = {1{`RANDOM}};
  r_2039 = _RAND_2039[0:0];
  _RAND_2040 = {1{`RANDOM}};
  r_2040 = _RAND_2040[0:0];
  _RAND_2041 = {1{`RANDOM}};
  r_2041 = _RAND_2041[0:0];
  _RAND_2042 = {1{`RANDOM}};
  r_2042 = _RAND_2042[0:0];
  _RAND_2043 = {1{`RANDOM}};
  r_2043 = _RAND_2043[0:0];
  _RAND_2044 = {1{`RANDOM}};
  r_2044 = _RAND_2044[0:0];
  _RAND_2045 = {1{`RANDOM}};
  r_2045 = _RAND_2045[0:0];
  _RAND_2046 = {1{`RANDOM}};
  r_2046 = _RAND_2046[0:0];
  _RAND_2047 = {1{`RANDOM}};
  r_2047 = _RAND_2047[0:0];
  _RAND_2048 = {1{`RANDOM}};
  r_2048 = _RAND_2048[0:0];
  _RAND_2049 = {1{`RANDOM}};
  r_2049 = _RAND_2049[0:0];
  _RAND_2050 = {1{`RANDOM}};
  r_2050 = _RAND_2050[0:0];
  _RAND_2051 = {1{`RANDOM}};
  r_2051 = _RAND_2051[0:0];
  _RAND_2052 = {1{`RANDOM}};
  r_2052 = _RAND_2052[0:0];
  _RAND_2053 = {1{`RANDOM}};
  r_2053 = _RAND_2053[0:0];
  _RAND_2054 = {1{`RANDOM}};
  r_2054 = _RAND_2054[0:0];
  _RAND_2055 = {1{`RANDOM}};
  r_2055 = _RAND_2055[0:0];
  _RAND_2056 = {1{`RANDOM}};
  r_2056 = _RAND_2056[0:0];
  _RAND_2057 = {1{`RANDOM}};
  r_2057 = _RAND_2057[0:0];
  _RAND_2058 = {1{`RANDOM}};
  r_2058 = _RAND_2058[0:0];
  _RAND_2059 = {1{`RANDOM}};
  r_2059 = _RAND_2059[0:0];
  _RAND_2060 = {1{`RANDOM}};
  r_2060 = _RAND_2060[0:0];
  _RAND_2061 = {1{`RANDOM}};
  r_2061 = _RAND_2061[0:0];
  _RAND_2062 = {1{`RANDOM}};
  r_2062 = _RAND_2062[0:0];
  _RAND_2063 = {1{`RANDOM}};
  r_2063 = _RAND_2063[0:0];
  _RAND_2064 = {1{`RANDOM}};
  r_2064 = _RAND_2064[0:0];
  _RAND_2065 = {1{`RANDOM}};
  r_2065 = _RAND_2065[0:0];
  _RAND_2066 = {1{`RANDOM}};
  r_2066 = _RAND_2066[0:0];
  _RAND_2067 = {1{`RANDOM}};
  r_2067 = _RAND_2067[0:0];
  _RAND_2068 = {1{`RANDOM}};
  r_2068 = _RAND_2068[0:0];
  _RAND_2069 = {1{`RANDOM}};
  r_2069 = _RAND_2069[0:0];
  _RAND_2070 = {1{`RANDOM}};
  r_2070 = _RAND_2070[0:0];
  _RAND_2071 = {1{`RANDOM}};
  r_2071 = _RAND_2071[0:0];
  _RAND_2072 = {1{`RANDOM}};
  r_2072 = _RAND_2072[0:0];
  _RAND_2073 = {1{`RANDOM}};
  r_2073 = _RAND_2073[0:0];
  _RAND_2074 = {1{`RANDOM}};
  r_2074 = _RAND_2074[0:0];
  _RAND_2075 = {1{`RANDOM}};
  r_2075 = _RAND_2075[0:0];
  _RAND_2076 = {1{`RANDOM}};
  r_2076 = _RAND_2076[0:0];
  _RAND_2077 = {1{`RANDOM}};
  r_2077 = _RAND_2077[0:0];
  _RAND_2078 = {1{`RANDOM}};
  r_2078 = _RAND_2078[0:0];
  _RAND_2079 = {1{`RANDOM}};
  r_2079 = _RAND_2079[0:0];
  _RAND_2080 = {1{`RANDOM}};
  r_2080 = _RAND_2080[0:0];
  _RAND_2081 = {1{`RANDOM}};
  r_2081 = _RAND_2081[0:0];
  _RAND_2082 = {1{`RANDOM}};
  r_2082 = _RAND_2082[0:0];
  _RAND_2083 = {1{`RANDOM}};
  r_2083 = _RAND_2083[0:0];
  _RAND_2084 = {1{`RANDOM}};
  r_2084 = _RAND_2084[0:0];
  _RAND_2085 = {1{`RANDOM}};
  r_2085 = _RAND_2085[0:0];
  _RAND_2086 = {1{`RANDOM}};
  r_2086 = _RAND_2086[0:0];
  _RAND_2087 = {1{`RANDOM}};
  r_2087 = _RAND_2087[0:0];
  _RAND_2088 = {1{`RANDOM}};
  r_2088 = _RAND_2088[0:0];
  _RAND_2089 = {1{`RANDOM}};
  r_2089 = _RAND_2089[0:0];
  _RAND_2090 = {1{`RANDOM}};
  r_2090 = _RAND_2090[0:0];
  _RAND_2091 = {1{`RANDOM}};
  r_2091 = _RAND_2091[0:0];
  _RAND_2092 = {1{`RANDOM}};
  r_2092 = _RAND_2092[0:0];
  _RAND_2093 = {1{`RANDOM}};
  r_2093 = _RAND_2093[0:0];
  _RAND_2094 = {1{`RANDOM}};
  r_2094 = _RAND_2094[0:0];
  _RAND_2095 = {1{`RANDOM}};
  r_2095 = _RAND_2095[0:0];
  _RAND_2096 = {1{`RANDOM}};
  r_2096 = _RAND_2096[0:0];
  _RAND_2097 = {1{`RANDOM}};
  r_2097 = _RAND_2097[0:0];
  _RAND_2098 = {1{`RANDOM}};
  r_2098 = _RAND_2098[0:0];
  _RAND_2099 = {1{`RANDOM}};
  r_2099 = _RAND_2099[0:0];
  _RAND_2100 = {1{`RANDOM}};
  r_2100 = _RAND_2100[0:0];
  _RAND_2101 = {1{`RANDOM}};
  r_2101 = _RAND_2101[0:0];
  _RAND_2102 = {1{`RANDOM}};
  r_2102 = _RAND_2102[0:0];
  _RAND_2103 = {1{`RANDOM}};
  r_2103 = _RAND_2103[0:0];
  _RAND_2104 = {1{`RANDOM}};
  r_2104 = _RAND_2104[0:0];
  _RAND_2105 = {1{`RANDOM}};
  r_2105 = _RAND_2105[0:0];
  _RAND_2106 = {1{`RANDOM}};
  r_2106 = _RAND_2106[0:0];
  _RAND_2107 = {1{`RANDOM}};
  r_2107 = _RAND_2107[0:0];
  _RAND_2108 = {1{`RANDOM}};
  r_2108 = _RAND_2108[0:0];
  _RAND_2109 = {1{`RANDOM}};
  r_2109 = _RAND_2109[0:0];
  _RAND_2110 = {1{`RANDOM}};
  r_2110 = _RAND_2110[0:0];
  _RAND_2111 = {1{`RANDOM}};
  r_2111 = _RAND_2111[0:0];
  _RAND_2112 = {1{`RANDOM}};
  r_2112 = _RAND_2112[0:0];
  _RAND_2113 = {1{`RANDOM}};
  r_2113 = _RAND_2113[0:0];
  _RAND_2114 = {1{`RANDOM}};
  r_2114 = _RAND_2114[0:0];
  _RAND_2115 = {1{`RANDOM}};
  r_2115 = _RAND_2115[0:0];
  _RAND_2116 = {1{`RANDOM}};
  r_2116 = _RAND_2116[0:0];
  _RAND_2117 = {1{`RANDOM}};
  r_2117 = _RAND_2117[0:0];
  _RAND_2118 = {1{`RANDOM}};
  r_2118 = _RAND_2118[0:0];
  _RAND_2119 = {1{`RANDOM}};
  r_2119 = _RAND_2119[0:0];
  _RAND_2120 = {1{`RANDOM}};
  r_2120 = _RAND_2120[0:0];
  _RAND_2121 = {1{`RANDOM}};
  r_2121 = _RAND_2121[0:0];
  _RAND_2122 = {1{`RANDOM}};
  r_2122 = _RAND_2122[0:0];
  _RAND_2123 = {1{`RANDOM}};
  r_2123 = _RAND_2123[0:0];
  _RAND_2124 = {1{`RANDOM}};
  r_2124 = _RAND_2124[0:0];
  _RAND_2125 = {1{`RANDOM}};
  r_2125 = _RAND_2125[0:0];
  _RAND_2126 = {1{`RANDOM}};
  r_2126 = _RAND_2126[0:0];
  _RAND_2127 = {1{`RANDOM}};
  r_2127 = _RAND_2127[0:0];
  _RAND_2128 = {1{`RANDOM}};
  r_2128 = _RAND_2128[0:0];
  _RAND_2129 = {1{`RANDOM}};
  r_2129 = _RAND_2129[0:0];
  _RAND_2130 = {1{`RANDOM}};
  r_2130 = _RAND_2130[0:0];
  _RAND_2131 = {1{`RANDOM}};
  r_2131 = _RAND_2131[0:0];
  _RAND_2132 = {1{`RANDOM}};
  r_2132 = _RAND_2132[0:0];
  _RAND_2133 = {1{`RANDOM}};
  r_2133 = _RAND_2133[0:0];
  _RAND_2134 = {1{`RANDOM}};
  r_2134 = _RAND_2134[0:0];
  _RAND_2135 = {1{`RANDOM}};
  r_2135 = _RAND_2135[0:0];
  _RAND_2136 = {1{`RANDOM}};
  r_2136 = _RAND_2136[0:0];
  _RAND_2137 = {1{`RANDOM}};
  r_2137 = _RAND_2137[0:0];
  _RAND_2138 = {1{`RANDOM}};
  r_2138 = _RAND_2138[0:0];
  _RAND_2139 = {1{`RANDOM}};
  r_2139 = _RAND_2139[0:0];
  _RAND_2140 = {1{`RANDOM}};
  r_2140 = _RAND_2140[0:0];
  _RAND_2141 = {1{`RANDOM}};
  r_2141 = _RAND_2141[0:0];
  _RAND_2142 = {1{`RANDOM}};
  r_2142 = _RAND_2142[0:0];
  _RAND_2143 = {1{`RANDOM}};
  r_2143 = _RAND_2143[0:0];
  _RAND_2144 = {1{`RANDOM}};
  r_2144 = _RAND_2144[0:0];
  _RAND_2145 = {1{`RANDOM}};
  r_2145 = _RAND_2145[0:0];
  _RAND_2146 = {1{`RANDOM}};
  r_2146 = _RAND_2146[0:0];
  _RAND_2147 = {1{`RANDOM}};
  r_2147 = _RAND_2147[0:0];
  _RAND_2148 = {1{`RANDOM}};
  r_2148 = _RAND_2148[0:0];
  _RAND_2149 = {1{`RANDOM}};
  r_2149 = _RAND_2149[0:0];
  _RAND_2150 = {1{`RANDOM}};
  r_2150 = _RAND_2150[0:0];
  _RAND_2151 = {1{`RANDOM}};
  r_2151 = _RAND_2151[0:0];
  _RAND_2152 = {1{`RANDOM}};
  r_2152 = _RAND_2152[0:0];
  _RAND_2153 = {1{`RANDOM}};
  r_2153 = _RAND_2153[0:0];
  _RAND_2154 = {1{`RANDOM}};
  r_2154 = _RAND_2154[0:0];
  _RAND_2155 = {1{`RANDOM}};
  r_2155 = _RAND_2155[0:0];
  _RAND_2156 = {1{`RANDOM}};
  r_2156 = _RAND_2156[0:0];
  _RAND_2157 = {1{`RANDOM}};
  r_2157 = _RAND_2157[0:0];
  _RAND_2158 = {1{`RANDOM}};
  r_2158 = _RAND_2158[0:0];
  _RAND_2159 = {1{`RANDOM}};
  r_2159 = _RAND_2159[0:0];
  _RAND_2160 = {1{`RANDOM}};
  r_2160 = _RAND_2160[0:0];
  _RAND_2161 = {1{`RANDOM}};
  r_2161 = _RAND_2161[0:0];
  _RAND_2162 = {1{`RANDOM}};
  r_2162 = _RAND_2162[0:0];
  _RAND_2163 = {1{`RANDOM}};
  r_2163 = _RAND_2163[0:0];
  _RAND_2164 = {1{`RANDOM}};
  r_2164 = _RAND_2164[0:0];
  _RAND_2165 = {1{`RANDOM}};
  r_2165 = _RAND_2165[0:0];
  _RAND_2166 = {1{`RANDOM}};
  r_2166 = _RAND_2166[0:0];
  _RAND_2167 = {1{`RANDOM}};
  r_2167 = _RAND_2167[0:0];
  _RAND_2168 = {1{`RANDOM}};
  r_2168 = _RAND_2168[0:0];
  _RAND_2169 = {1{`RANDOM}};
  r_2169 = _RAND_2169[0:0];
  _RAND_2170 = {1{`RANDOM}};
  r_2170 = _RAND_2170[0:0];
  _RAND_2171 = {1{`RANDOM}};
  r_2171 = _RAND_2171[0:0];
  _RAND_2172 = {1{`RANDOM}};
  r_2172 = _RAND_2172[0:0];
  _RAND_2173 = {1{`RANDOM}};
  r_2173 = _RAND_2173[0:0];
  _RAND_2174 = {1{`RANDOM}};
  r_2174 = _RAND_2174[0:0];
  _RAND_2175 = {1{`RANDOM}};
  r_2175 = _RAND_2175[0:0];
  _RAND_2176 = {1{`RANDOM}};
  r_2176 = _RAND_2176[0:0];
  _RAND_2177 = {1{`RANDOM}};
  r_2177 = _RAND_2177[0:0];
  _RAND_2178 = {1{`RANDOM}};
  r_2178 = _RAND_2178[0:0];
  _RAND_2179 = {1{`RANDOM}};
  r_2179 = _RAND_2179[0:0];
  _RAND_2180 = {1{`RANDOM}};
  r_2180 = _RAND_2180[0:0];
  _RAND_2181 = {1{`RANDOM}};
  r_2181 = _RAND_2181[0:0];
  _RAND_2182 = {1{`RANDOM}};
  r_2182 = _RAND_2182[0:0];
  _RAND_2183 = {1{`RANDOM}};
  r_2183 = _RAND_2183[0:0];
  _RAND_2184 = {1{`RANDOM}};
  r_2184 = _RAND_2184[0:0];
  _RAND_2185 = {1{`RANDOM}};
  r_2185 = _RAND_2185[0:0];
  _RAND_2186 = {1{`RANDOM}};
  r_2186 = _RAND_2186[0:0];
  _RAND_2187 = {1{`RANDOM}};
  r_2187 = _RAND_2187[0:0];
  _RAND_2188 = {1{`RANDOM}};
  r_2188 = _RAND_2188[0:0];
  _RAND_2189 = {1{`RANDOM}};
  r_2189 = _RAND_2189[0:0];
  _RAND_2190 = {1{`RANDOM}};
  r_2190 = _RAND_2190[0:0];
  _RAND_2191 = {1{`RANDOM}};
  r_2191 = _RAND_2191[0:0];
  _RAND_2192 = {1{`RANDOM}};
  r_2192 = _RAND_2192[0:0];
  _RAND_2193 = {1{`RANDOM}};
  r_2193 = _RAND_2193[0:0];
  _RAND_2194 = {1{`RANDOM}};
  r_2194 = _RAND_2194[0:0];
  _RAND_2195 = {1{`RANDOM}};
  r_2195 = _RAND_2195[0:0];
  _RAND_2196 = {1{`RANDOM}};
  r_2196 = _RAND_2196[0:0];
  _RAND_2197 = {1{`RANDOM}};
  r_2197 = _RAND_2197[0:0];
  _RAND_2198 = {1{`RANDOM}};
  r_2198 = _RAND_2198[0:0];
  _RAND_2199 = {1{`RANDOM}};
  r_2199 = _RAND_2199[0:0];
  _RAND_2200 = {1{`RANDOM}};
  r_2200 = _RAND_2200[0:0];
  _RAND_2201 = {1{`RANDOM}};
  r_2201 = _RAND_2201[0:0];
  _RAND_2202 = {1{`RANDOM}};
  r_2202 = _RAND_2202[0:0];
  _RAND_2203 = {1{`RANDOM}};
  r_2203 = _RAND_2203[0:0];
  _RAND_2204 = {1{`RANDOM}};
  r_2204 = _RAND_2204[0:0];
  _RAND_2205 = {1{`RANDOM}};
  r_2205 = _RAND_2205[0:0];
  _RAND_2206 = {1{`RANDOM}};
  r_2206 = _RAND_2206[0:0];
  _RAND_2207 = {1{`RANDOM}};
  r_2207 = _RAND_2207[0:0];
  _RAND_2208 = {1{`RANDOM}};
  r_2208 = _RAND_2208[0:0];
  _RAND_2209 = {1{`RANDOM}};
  r_2209 = _RAND_2209[0:0];
  _RAND_2210 = {1{`RANDOM}};
  r_2210 = _RAND_2210[0:0];
  _RAND_2211 = {1{`RANDOM}};
  r_2211 = _RAND_2211[0:0];
  _RAND_2212 = {1{`RANDOM}};
  r_2212 = _RAND_2212[0:0];
  _RAND_2213 = {1{`RANDOM}};
  r_2213 = _RAND_2213[0:0];
  _RAND_2214 = {1{`RANDOM}};
  r_2214 = _RAND_2214[0:0];
  _RAND_2215 = {1{`RANDOM}};
  r_2215 = _RAND_2215[0:0];
  _RAND_2216 = {1{`RANDOM}};
  r_2216 = _RAND_2216[0:0];
  _RAND_2217 = {1{`RANDOM}};
  r_2217 = _RAND_2217[0:0];
  _RAND_2218 = {1{`RANDOM}};
  r_2218 = _RAND_2218[0:0];
  _RAND_2219 = {1{`RANDOM}};
  r_2219 = _RAND_2219[0:0];
  _RAND_2220 = {1{`RANDOM}};
  r_2220 = _RAND_2220[0:0];
  _RAND_2221 = {1{`RANDOM}};
  r_2221 = _RAND_2221[0:0];
  _RAND_2222 = {1{`RANDOM}};
  r_2222 = _RAND_2222[0:0];
  _RAND_2223 = {1{`RANDOM}};
  r_2223 = _RAND_2223[0:0];
  _RAND_2224 = {1{`RANDOM}};
  r_2224 = _RAND_2224[0:0];
  _RAND_2225 = {1{`RANDOM}};
  r_2225 = _RAND_2225[0:0];
  _RAND_2226 = {1{`RANDOM}};
  r_2226 = _RAND_2226[0:0];
  _RAND_2227 = {1{`RANDOM}};
  r_2227 = _RAND_2227[0:0];
  _RAND_2228 = {1{`RANDOM}};
  r_2228 = _RAND_2228[0:0];
  _RAND_2229 = {1{`RANDOM}};
  r_2229 = _RAND_2229[0:0];
  _RAND_2230 = {1{`RANDOM}};
  r_2230 = _RAND_2230[0:0];
  _RAND_2231 = {1{`RANDOM}};
  r_2231 = _RAND_2231[0:0];
  _RAND_2232 = {1{`RANDOM}};
  r_2232 = _RAND_2232[0:0];
  _RAND_2233 = {1{`RANDOM}};
  r_2233 = _RAND_2233[0:0];
  _RAND_2234 = {1{`RANDOM}};
  r_2234 = _RAND_2234[0:0];
  _RAND_2235 = {1{`RANDOM}};
  r_2235 = _RAND_2235[0:0];
  _RAND_2236 = {1{`RANDOM}};
  r_2236 = _RAND_2236[0:0];
  _RAND_2237 = {1{`RANDOM}};
  r_2237 = _RAND_2237[0:0];
  _RAND_2238 = {1{`RANDOM}};
  r_2238 = _RAND_2238[0:0];
  _RAND_2239 = {1{`RANDOM}};
  r_2239 = _RAND_2239[0:0];
  _RAND_2240 = {1{`RANDOM}};
  r_2240 = _RAND_2240[0:0];
  _RAND_2241 = {1{`RANDOM}};
  r_2241 = _RAND_2241[0:0];
  _RAND_2242 = {1{`RANDOM}};
  r_2242 = _RAND_2242[0:0];
  _RAND_2243 = {1{`RANDOM}};
  r_2243 = _RAND_2243[0:0];
  _RAND_2244 = {1{`RANDOM}};
  r_2244 = _RAND_2244[0:0];
  _RAND_2245 = {1{`RANDOM}};
  r_2245 = _RAND_2245[0:0];
  _RAND_2246 = {1{`RANDOM}};
  r_2246 = _RAND_2246[0:0];
  _RAND_2247 = {1{`RANDOM}};
  r_2247 = _RAND_2247[0:0];
  _RAND_2248 = {1{`RANDOM}};
  r_2248 = _RAND_2248[0:0];
  _RAND_2249 = {1{`RANDOM}};
  r_2249 = _RAND_2249[0:0];
  _RAND_2250 = {1{`RANDOM}};
  r_2250 = _RAND_2250[0:0];
  _RAND_2251 = {1{`RANDOM}};
  r_2251 = _RAND_2251[0:0];
  _RAND_2252 = {1{`RANDOM}};
  r_2252 = _RAND_2252[0:0];
  _RAND_2253 = {1{`RANDOM}};
  r_2253 = _RAND_2253[0:0];
  _RAND_2254 = {1{`RANDOM}};
  r_2254 = _RAND_2254[0:0];
  _RAND_2255 = {1{`RANDOM}};
  r_2255 = _RAND_2255[0:0];
  _RAND_2256 = {1{`RANDOM}};
  r_2256 = _RAND_2256[0:0];
  _RAND_2257 = {1{`RANDOM}};
  r_2257 = _RAND_2257[0:0];
  _RAND_2258 = {1{`RANDOM}};
  r_2258 = _RAND_2258[0:0];
  _RAND_2259 = {1{`RANDOM}};
  r_2259 = _RAND_2259[0:0];
  _RAND_2260 = {1{`RANDOM}};
  r_2260 = _RAND_2260[0:0];
  _RAND_2261 = {1{`RANDOM}};
  r_2261 = _RAND_2261[0:0];
  _RAND_2262 = {1{`RANDOM}};
  r_2262 = _RAND_2262[0:0];
  _RAND_2263 = {1{`RANDOM}};
  r_2263 = _RAND_2263[0:0];
  _RAND_2264 = {1{`RANDOM}};
  r_2264 = _RAND_2264[0:0];
  _RAND_2265 = {1{`RANDOM}};
  r_2265 = _RAND_2265[0:0];
  _RAND_2266 = {1{`RANDOM}};
  r_2266 = _RAND_2266[0:0];
  _RAND_2267 = {1{`RANDOM}};
  r_2267 = _RAND_2267[0:0];
  _RAND_2268 = {1{`RANDOM}};
  r_2268 = _RAND_2268[0:0];
  _RAND_2269 = {1{`RANDOM}};
  r_2269 = _RAND_2269[0:0];
  _RAND_2270 = {1{`RANDOM}};
  r_2270 = _RAND_2270[0:0];
  _RAND_2271 = {1{`RANDOM}};
  r_2271 = _RAND_2271[0:0];
  _RAND_2272 = {1{`RANDOM}};
  r_2272 = _RAND_2272[0:0];
  _RAND_2273 = {1{`RANDOM}};
  r_2273 = _RAND_2273[0:0];
  _RAND_2274 = {1{`RANDOM}};
  r_2274 = _RAND_2274[0:0];
  _RAND_2275 = {1{`RANDOM}};
  r_2275 = _RAND_2275[0:0];
  _RAND_2276 = {1{`RANDOM}};
  r_2276 = _RAND_2276[0:0];
  _RAND_2277 = {1{`RANDOM}};
  r_2277 = _RAND_2277[0:0];
  _RAND_2278 = {1{`RANDOM}};
  r_2278 = _RAND_2278[0:0];
  _RAND_2279 = {1{`RANDOM}};
  r_2279 = _RAND_2279[0:0];
  _RAND_2280 = {1{`RANDOM}};
  r_2280 = _RAND_2280[0:0];
  _RAND_2281 = {1{`RANDOM}};
  r_2281 = _RAND_2281[0:0];
  _RAND_2282 = {1{`RANDOM}};
  r_2282 = _RAND_2282[0:0];
  _RAND_2283 = {1{`RANDOM}};
  r_2283 = _RAND_2283[0:0];
  _RAND_2284 = {1{`RANDOM}};
  r_2284 = _RAND_2284[0:0];
  _RAND_2285 = {1{`RANDOM}};
  r_2285 = _RAND_2285[0:0];
  _RAND_2286 = {1{`RANDOM}};
  r_2286 = _RAND_2286[0:0];
  _RAND_2287 = {1{`RANDOM}};
  r_2287 = _RAND_2287[0:0];
  _RAND_2288 = {1{`RANDOM}};
  r_2288 = _RAND_2288[0:0];
  _RAND_2289 = {1{`RANDOM}};
  r_2289 = _RAND_2289[0:0];
  _RAND_2290 = {1{`RANDOM}};
  r_2290 = _RAND_2290[0:0];
  _RAND_2291 = {1{`RANDOM}};
  r_2291 = _RAND_2291[0:0];
  _RAND_2292 = {1{`RANDOM}};
  r_2292 = _RAND_2292[0:0];
  _RAND_2293 = {1{`RANDOM}};
  r_2293 = _RAND_2293[0:0];
  _RAND_2294 = {1{`RANDOM}};
  r_2294 = _RAND_2294[0:0];
  _RAND_2295 = {1{`RANDOM}};
  r_2295 = _RAND_2295[0:0];
  _RAND_2296 = {1{`RANDOM}};
  r_2296 = _RAND_2296[0:0];
  _RAND_2297 = {1{`RANDOM}};
  r_2297 = _RAND_2297[0:0];
  _RAND_2298 = {1{`RANDOM}};
  r_2298 = _RAND_2298[0:0];
  _RAND_2299 = {1{`RANDOM}};
  r_2299 = _RAND_2299[0:0];
  _RAND_2300 = {1{`RANDOM}};
  r_2300 = _RAND_2300[0:0];
  _RAND_2301 = {1{`RANDOM}};
  r_2301 = _RAND_2301[0:0];
  _RAND_2302 = {1{`RANDOM}};
  r_2302 = _RAND_2302[0:0];
  _RAND_2303 = {1{`RANDOM}};
  r_2303 = _RAND_2303[0:0];
  _RAND_2304 = {1{`RANDOM}};
  r_2304 = _RAND_2304[0:0];
  _RAND_2305 = {1{`RANDOM}};
  r_2305 = _RAND_2305[0:0];
  _RAND_2306 = {1{`RANDOM}};
  r_2306 = _RAND_2306[0:0];
  _RAND_2307 = {1{`RANDOM}};
  r_2307 = _RAND_2307[0:0];
  _RAND_2308 = {1{`RANDOM}};
  r_2308 = _RAND_2308[0:0];
  _RAND_2309 = {1{`RANDOM}};
  r_2309 = _RAND_2309[0:0];
  _RAND_2310 = {1{`RANDOM}};
  r_2310 = _RAND_2310[0:0];
  _RAND_2311 = {1{`RANDOM}};
  r_2311 = _RAND_2311[0:0];
  _RAND_2312 = {1{`RANDOM}};
  r_2312 = _RAND_2312[0:0];
  _RAND_2313 = {1{`RANDOM}};
  r_2313 = _RAND_2313[0:0];
  _RAND_2314 = {1{`RANDOM}};
  r_2314 = _RAND_2314[0:0];
  _RAND_2315 = {1{`RANDOM}};
  r_2315 = _RAND_2315[0:0];
  _RAND_2316 = {1{`RANDOM}};
  r_2316 = _RAND_2316[0:0];
  _RAND_2317 = {1{`RANDOM}};
  r_2317 = _RAND_2317[0:0];
  _RAND_2318 = {1{`RANDOM}};
  r_2318 = _RAND_2318[0:0];
  _RAND_2319 = {1{`RANDOM}};
  r_2319 = _RAND_2319[0:0];
  _RAND_2320 = {1{`RANDOM}};
  r_2320 = _RAND_2320[0:0];
  _RAND_2321 = {1{`RANDOM}};
  r_2321 = _RAND_2321[0:0];
  _RAND_2322 = {1{`RANDOM}};
  r_2322 = _RAND_2322[0:0];
  _RAND_2323 = {1{`RANDOM}};
  r_2323 = _RAND_2323[0:0];
  _RAND_2324 = {1{`RANDOM}};
  r_2324 = _RAND_2324[0:0];
  _RAND_2325 = {1{`RANDOM}};
  r_2325 = _RAND_2325[0:0];
  _RAND_2326 = {1{`RANDOM}};
  r_2326 = _RAND_2326[0:0];
  _RAND_2327 = {1{`RANDOM}};
  r_2327 = _RAND_2327[0:0];
  _RAND_2328 = {1{`RANDOM}};
  r_2328 = _RAND_2328[0:0];
  _RAND_2329 = {1{`RANDOM}};
  r_2329 = _RAND_2329[0:0];
  _RAND_2330 = {1{`RANDOM}};
  r_2330 = _RAND_2330[0:0];
  _RAND_2331 = {1{`RANDOM}};
  r_2331 = _RAND_2331[0:0];
  _RAND_2332 = {1{`RANDOM}};
  r_2332 = _RAND_2332[0:0];
  _RAND_2333 = {1{`RANDOM}};
  r_2333 = _RAND_2333[0:0];
  _RAND_2334 = {1{`RANDOM}};
  r_2334 = _RAND_2334[0:0];
  _RAND_2335 = {1{`RANDOM}};
  r_2335 = _RAND_2335[0:0];
  _RAND_2336 = {1{`RANDOM}};
  r_2336 = _RAND_2336[0:0];
  _RAND_2337 = {1{`RANDOM}};
  r_2337 = _RAND_2337[0:0];
  _RAND_2338 = {1{`RANDOM}};
  r_2338 = _RAND_2338[0:0];
  _RAND_2339 = {1{`RANDOM}};
  r_2339 = _RAND_2339[0:0];
  _RAND_2340 = {1{`RANDOM}};
  r_2340 = _RAND_2340[0:0];
  _RAND_2341 = {1{`RANDOM}};
  r_2341 = _RAND_2341[0:0];
  _RAND_2342 = {1{`RANDOM}};
  r_2342 = _RAND_2342[0:0];
  _RAND_2343 = {1{`RANDOM}};
  r_2343 = _RAND_2343[0:0];
  _RAND_2344 = {1{`RANDOM}};
  r_2344 = _RAND_2344[0:0];
  _RAND_2345 = {1{`RANDOM}};
  r_2345 = _RAND_2345[0:0];
  _RAND_2346 = {1{`RANDOM}};
  r_2346 = _RAND_2346[0:0];
  _RAND_2347 = {1{`RANDOM}};
  r_2347 = _RAND_2347[0:0];
  _RAND_2348 = {1{`RANDOM}};
  r_2348 = _RAND_2348[0:0];
  _RAND_2349 = {1{`RANDOM}};
  r_2349 = _RAND_2349[0:0];
  _RAND_2350 = {1{`RANDOM}};
  r_2350 = _RAND_2350[0:0];
  _RAND_2351 = {1{`RANDOM}};
  r_2351 = _RAND_2351[0:0];
  _RAND_2352 = {1{`RANDOM}};
  r_2352 = _RAND_2352[0:0];
  _RAND_2353 = {1{`RANDOM}};
  r_2353 = _RAND_2353[0:0];
  _RAND_2354 = {1{`RANDOM}};
  r_2354 = _RAND_2354[0:0];
  _RAND_2355 = {1{`RANDOM}};
  r_2355 = _RAND_2355[0:0];
  _RAND_2356 = {1{`RANDOM}};
  r_2356 = _RAND_2356[0:0];
  _RAND_2357 = {1{`RANDOM}};
  r_2357 = _RAND_2357[0:0];
  _RAND_2358 = {1{`RANDOM}};
  r_2358 = _RAND_2358[0:0];
  _RAND_2359 = {1{`RANDOM}};
  r_2359 = _RAND_2359[0:0];
  _RAND_2360 = {1{`RANDOM}};
  r_2360 = _RAND_2360[0:0];
  _RAND_2361 = {1{`RANDOM}};
  r_2361 = _RAND_2361[0:0];
  _RAND_2362 = {1{`RANDOM}};
  r_2362 = _RAND_2362[0:0];
  _RAND_2363 = {1{`RANDOM}};
  r_2363 = _RAND_2363[0:0];
  _RAND_2364 = {1{`RANDOM}};
  r_2364 = _RAND_2364[0:0];
  _RAND_2365 = {1{`RANDOM}};
  r_2365 = _RAND_2365[0:0];
  _RAND_2366 = {1{`RANDOM}};
  r_2366 = _RAND_2366[0:0];
  _RAND_2367 = {1{`RANDOM}};
  r_2367 = _RAND_2367[0:0];
  _RAND_2368 = {1{`RANDOM}};
  r_2368 = _RAND_2368[0:0];
  _RAND_2369 = {1{`RANDOM}};
  r_2369 = _RAND_2369[0:0];
  _RAND_2370 = {1{`RANDOM}};
  r_2370 = _RAND_2370[0:0];
  _RAND_2371 = {1{`RANDOM}};
  r_2371 = _RAND_2371[0:0];
  _RAND_2372 = {1{`RANDOM}};
  r_2372 = _RAND_2372[0:0];
  _RAND_2373 = {1{`RANDOM}};
  r_2373 = _RAND_2373[0:0];
  _RAND_2374 = {1{`RANDOM}};
  r_2374 = _RAND_2374[0:0];
  _RAND_2375 = {1{`RANDOM}};
  r_2375 = _RAND_2375[0:0];
  _RAND_2376 = {1{`RANDOM}};
  r_2376 = _RAND_2376[0:0];
  _RAND_2377 = {1{`RANDOM}};
  r_2377 = _RAND_2377[0:0];
  _RAND_2378 = {1{`RANDOM}};
  r_2378 = _RAND_2378[0:0];
  _RAND_2379 = {1{`RANDOM}};
  r_2379 = _RAND_2379[0:0];
  _RAND_2380 = {1{`RANDOM}};
  r_2380 = _RAND_2380[0:0];
  _RAND_2381 = {1{`RANDOM}};
  r_2381 = _RAND_2381[0:0];
  _RAND_2382 = {1{`RANDOM}};
  r_2382 = _RAND_2382[0:0];
  _RAND_2383 = {1{`RANDOM}};
  r_2383 = _RAND_2383[0:0];
  _RAND_2384 = {1{`RANDOM}};
  r_2384 = _RAND_2384[0:0];
  _RAND_2385 = {1{`RANDOM}};
  r_2385 = _RAND_2385[0:0];
  _RAND_2386 = {1{`RANDOM}};
  r_2386 = _RAND_2386[0:0];
  _RAND_2387 = {1{`RANDOM}};
  r_2387 = _RAND_2387[0:0];
  _RAND_2388 = {1{`RANDOM}};
  r_2388 = _RAND_2388[0:0];
  _RAND_2389 = {1{`RANDOM}};
  r_2389 = _RAND_2389[0:0];
  _RAND_2390 = {1{`RANDOM}};
  r_2390 = _RAND_2390[0:0];
  _RAND_2391 = {1{`RANDOM}};
  r_2391 = _RAND_2391[0:0];
  _RAND_2392 = {1{`RANDOM}};
  r_2392 = _RAND_2392[0:0];
  _RAND_2393 = {1{`RANDOM}};
  r_2393 = _RAND_2393[0:0];
  _RAND_2394 = {1{`RANDOM}};
  r_2394 = _RAND_2394[0:0];
  _RAND_2395 = {1{`RANDOM}};
  r_2395 = _RAND_2395[0:0];
  _RAND_2396 = {1{`RANDOM}};
  r_2396 = _RAND_2396[0:0];
  _RAND_2397 = {1{`RANDOM}};
  r_2397 = _RAND_2397[0:0];
  _RAND_2398 = {1{`RANDOM}};
  r_2398 = _RAND_2398[0:0];
  _RAND_2399 = {1{`RANDOM}};
  r_2399 = _RAND_2399[0:0];
  _RAND_2400 = {1{`RANDOM}};
  r_2400 = _RAND_2400[0:0];
  _RAND_2401 = {1{`RANDOM}};
  r_2401 = _RAND_2401[0:0];
  _RAND_2402 = {1{`RANDOM}};
  r_2402 = _RAND_2402[0:0];
  _RAND_2403 = {1{`RANDOM}};
  r_2403 = _RAND_2403[0:0];
  _RAND_2404 = {1{`RANDOM}};
  r_2404 = _RAND_2404[0:0];
  _RAND_2405 = {1{`RANDOM}};
  r_2405 = _RAND_2405[0:0];
  _RAND_2406 = {1{`RANDOM}};
  r_2406 = _RAND_2406[0:0];
  _RAND_2407 = {1{`RANDOM}};
  r_2407 = _RAND_2407[0:0];
  _RAND_2408 = {1{`RANDOM}};
  r_2408 = _RAND_2408[0:0];
  _RAND_2409 = {1{`RANDOM}};
  r_2409 = _RAND_2409[0:0];
  _RAND_2410 = {1{`RANDOM}};
  r_2410 = _RAND_2410[0:0];
  _RAND_2411 = {1{`RANDOM}};
  r_2411 = _RAND_2411[0:0];
  _RAND_2412 = {1{`RANDOM}};
  r_2412 = _RAND_2412[0:0];
  _RAND_2413 = {1{`RANDOM}};
  r_2413 = _RAND_2413[0:0];
  _RAND_2414 = {1{`RANDOM}};
  r_2414 = _RAND_2414[0:0];
  _RAND_2415 = {1{`RANDOM}};
  r_2415 = _RAND_2415[0:0];
  _RAND_2416 = {1{`RANDOM}};
  r_2416 = _RAND_2416[0:0];
  _RAND_2417 = {1{`RANDOM}};
  r_2417 = _RAND_2417[0:0];
  _RAND_2418 = {1{`RANDOM}};
  r_2418 = _RAND_2418[0:0];
  _RAND_2419 = {1{`RANDOM}};
  r_2419 = _RAND_2419[0:0];
  _RAND_2420 = {1{`RANDOM}};
  r_2420 = _RAND_2420[0:0];
  _RAND_2421 = {1{`RANDOM}};
  r_2421 = _RAND_2421[0:0];
  _RAND_2422 = {1{`RANDOM}};
  r_2422 = _RAND_2422[0:0];
  _RAND_2423 = {1{`RANDOM}};
  r_2423 = _RAND_2423[0:0];
  _RAND_2424 = {1{`RANDOM}};
  r_2424 = _RAND_2424[0:0];
  _RAND_2425 = {1{`RANDOM}};
  r_2425 = _RAND_2425[0:0];
  _RAND_2426 = {1{`RANDOM}};
  r_2426 = _RAND_2426[0:0];
  _RAND_2427 = {1{`RANDOM}};
  r_2427 = _RAND_2427[0:0];
  _RAND_2428 = {1{`RANDOM}};
  r_2428 = _RAND_2428[0:0];
  _RAND_2429 = {1{`RANDOM}};
  r_2429 = _RAND_2429[0:0];
  _RAND_2430 = {1{`RANDOM}};
  r_2430 = _RAND_2430[0:0];
  _RAND_2431 = {1{`RANDOM}};
  r_2431 = _RAND_2431[0:0];
  _RAND_2432 = {1{`RANDOM}};
  r_2432 = _RAND_2432[0:0];
  _RAND_2433 = {1{`RANDOM}};
  r_2433 = _RAND_2433[0:0];
  _RAND_2434 = {1{`RANDOM}};
  r_2434 = _RAND_2434[0:0];
  _RAND_2435 = {1{`RANDOM}};
  r_2435 = _RAND_2435[0:0];
  _RAND_2436 = {1{`RANDOM}};
  r_2436 = _RAND_2436[0:0];
  _RAND_2437 = {1{`RANDOM}};
  r_2437 = _RAND_2437[0:0];
  _RAND_2438 = {1{`RANDOM}};
  r_2438 = _RAND_2438[0:0];
  _RAND_2439 = {1{`RANDOM}};
  r_2439 = _RAND_2439[0:0];
  _RAND_2440 = {1{`RANDOM}};
  r_2440 = _RAND_2440[0:0];
  _RAND_2441 = {1{`RANDOM}};
  r_2441 = _RAND_2441[0:0];
  _RAND_2442 = {1{`RANDOM}};
  r_2442 = _RAND_2442[0:0];
  _RAND_2443 = {1{`RANDOM}};
  r_2443 = _RAND_2443[0:0];
  _RAND_2444 = {1{`RANDOM}};
  r_2444 = _RAND_2444[0:0];
  _RAND_2445 = {1{`RANDOM}};
  r_2445 = _RAND_2445[0:0];
  _RAND_2446 = {1{`RANDOM}};
  r_2446 = _RAND_2446[0:0];
  _RAND_2447 = {1{`RANDOM}};
  r_2447 = _RAND_2447[0:0];
  _RAND_2448 = {1{`RANDOM}};
  r_2448 = _RAND_2448[0:0];
  _RAND_2449 = {1{`RANDOM}};
  r_2449 = _RAND_2449[0:0];
  _RAND_2450 = {1{`RANDOM}};
  r_2450 = _RAND_2450[0:0];
  _RAND_2451 = {1{`RANDOM}};
  r_2451 = _RAND_2451[0:0];
  _RAND_2452 = {1{`RANDOM}};
  r_2452 = _RAND_2452[0:0];
  _RAND_2453 = {1{`RANDOM}};
  r_2453 = _RAND_2453[0:0];
  _RAND_2454 = {1{`RANDOM}};
  r_2454 = _RAND_2454[0:0];
  _RAND_2455 = {1{`RANDOM}};
  r_2455 = _RAND_2455[0:0];
  _RAND_2456 = {1{`RANDOM}};
  r_2456 = _RAND_2456[0:0];
  _RAND_2457 = {1{`RANDOM}};
  r_2457 = _RAND_2457[0:0];
  _RAND_2458 = {1{`RANDOM}};
  r_2458 = _RAND_2458[0:0];
  _RAND_2459 = {1{`RANDOM}};
  r_2459 = _RAND_2459[0:0];
  _RAND_2460 = {1{`RANDOM}};
  r_2460 = _RAND_2460[0:0];
  _RAND_2461 = {1{`RANDOM}};
  r_2461 = _RAND_2461[0:0];
  _RAND_2462 = {1{`RANDOM}};
  r_2462 = _RAND_2462[0:0];
  _RAND_2463 = {1{`RANDOM}};
  r_2463 = _RAND_2463[0:0];
  _RAND_2464 = {1{`RANDOM}};
  r_2464 = _RAND_2464[0:0];
  _RAND_2465 = {1{`RANDOM}};
  r_2465 = _RAND_2465[0:0];
  _RAND_2466 = {1{`RANDOM}};
  r_2466 = _RAND_2466[0:0];
  _RAND_2467 = {1{`RANDOM}};
  r_2467 = _RAND_2467[0:0];
  _RAND_2468 = {1{`RANDOM}};
  r_2468 = _RAND_2468[0:0];
  _RAND_2469 = {1{`RANDOM}};
  r_2469 = _RAND_2469[0:0];
  _RAND_2470 = {1{`RANDOM}};
  r_2470 = _RAND_2470[0:0];
  _RAND_2471 = {1{`RANDOM}};
  r_2471 = _RAND_2471[0:0];
  _RAND_2472 = {1{`RANDOM}};
  r_2472 = _RAND_2472[0:0];
  _RAND_2473 = {1{`RANDOM}};
  r_2473 = _RAND_2473[0:0];
  _RAND_2474 = {1{`RANDOM}};
  r_2474 = _RAND_2474[0:0];
  _RAND_2475 = {1{`RANDOM}};
  r_2475 = _RAND_2475[0:0];
  _RAND_2476 = {1{`RANDOM}};
  r_2476 = _RAND_2476[0:0];
  _RAND_2477 = {1{`RANDOM}};
  r_2477 = _RAND_2477[0:0];
  _RAND_2478 = {1{`RANDOM}};
  r_2478 = _RAND_2478[0:0];
  _RAND_2479 = {1{`RANDOM}};
  r_2479 = _RAND_2479[0:0];
  _RAND_2480 = {1{`RANDOM}};
  r_2480 = _RAND_2480[0:0];
  _RAND_2481 = {1{`RANDOM}};
  r_2481 = _RAND_2481[0:0];
  _RAND_2482 = {1{`RANDOM}};
  r_2482 = _RAND_2482[0:0];
  _RAND_2483 = {1{`RANDOM}};
  r_2483 = _RAND_2483[0:0];
  _RAND_2484 = {1{`RANDOM}};
  r_2484 = _RAND_2484[0:0];
  _RAND_2485 = {1{`RANDOM}};
  r_2485 = _RAND_2485[0:0];
  _RAND_2486 = {1{`RANDOM}};
  r_2486 = _RAND_2486[0:0];
  _RAND_2487 = {1{`RANDOM}};
  r_2487 = _RAND_2487[0:0];
  _RAND_2488 = {1{`RANDOM}};
  r_2488 = _RAND_2488[0:0];
  _RAND_2489 = {1{`RANDOM}};
  r_2489 = _RAND_2489[0:0];
  _RAND_2490 = {1{`RANDOM}};
  r_2490 = _RAND_2490[0:0];
  _RAND_2491 = {1{`RANDOM}};
  r_2491 = _RAND_2491[0:0];
  _RAND_2492 = {1{`RANDOM}};
  r_2492 = _RAND_2492[0:0];
  _RAND_2493 = {1{`RANDOM}};
  r_2493 = _RAND_2493[0:0];
  _RAND_2494 = {1{`RANDOM}};
  r_2494 = _RAND_2494[0:0];
  _RAND_2495 = {1{`RANDOM}};
  r_2495 = _RAND_2495[0:0];
  _RAND_2496 = {1{`RANDOM}};
  r_2496 = _RAND_2496[0:0];
  _RAND_2497 = {1{`RANDOM}};
  r_2497 = _RAND_2497[0:0];
  _RAND_2498 = {1{`RANDOM}};
  r_2498 = _RAND_2498[0:0];
  _RAND_2499 = {1{`RANDOM}};
  r_2499 = _RAND_2499[0:0];
  _RAND_2500 = {1{`RANDOM}};
  r_2500 = _RAND_2500[0:0];
  _RAND_2501 = {1{`RANDOM}};
  r_2501 = _RAND_2501[0:0];
  _RAND_2502 = {1{`RANDOM}};
  r_2502 = _RAND_2502[0:0];
  _RAND_2503 = {1{`RANDOM}};
  r_2503 = _RAND_2503[0:0];
  _RAND_2504 = {1{`RANDOM}};
  r_2504 = _RAND_2504[0:0];
  _RAND_2505 = {1{`RANDOM}};
  r_2505 = _RAND_2505[0:0];
  _RAND_2506 = {1{`RANDOM}};
  r_2506 = _RAND_2506[0:0];
  _RAND_2507 = {1{`RANDOM}};
  r_2507 = _RAND_2507[0:0];
  _RAND_2508 = {1{`RANDOM}};
  r_2508 = _RAND_2508[0:0];
  _RAND_2509 = {1{`RANDOM}};
  r_2509 = _RAND_2509[0:0];
  _RAND_2510 = {1{`RANDOM}};
  r_2510 = _RAND_2510[0:0];
  _RAND_2511 = {1{`RANDOM}};
  r_2511 = _RAND_2511[0:0];
  _RAND_2512 = {1{`RANDOM}};
  r_2512 = _RAND_2512[0:0];
  _RAND_2513 = {1{`RANDOM}};
  r_2513 = _RAND_2513[0:0];
  _RAND_2514 = {1{`RANDOM}};
  r_2514 = _RAND_2514[0:0];
  _RAND_2515 = {1{`RANDOM}};
  r_2515 = _RAND_2515[0:0];
  _RAND_2516 = {1{`RANDOM}};
  r_2516 = _RAND_2516[0:0];
  _RAND_2517 = {1{`RANDOM}};
  r_2517 = _RAND_2517[0:0];
  _RAND_2518 = {1{`RANDOM}};
  r_2518 = _RAND_2518[0:0];
  _RAND_2519 = {1{`RANDOM}};
  r_2519 = _RAND_2519[0:0];
  _RAND_2520 = {1{`RANDOM}};
  r_2520 = _RAND_2520[0:0];
  _RAND_2521 = {1{`RANDOM}};
  r_2521 = _RAND_2521[0:0];
  _RAND_2522 = {1{`RANDOM}};
  r_2522 = _RAND_2522[0:0];
  _RAND_2523 = {1{`RANDOM}};
  r_2523 = _RAND_2523[0:0];
  _RAND_2524 = {1{`RANDOM}};
  r_2524 = _RAND_2524[0:0];
  _RAND_2525 = {1{`RANDOM}};
  r_2525 = _RAND_2525[0:0];
  _RAND_2526 = {1{`RANDOM}};
  r_2526 = _RAND_2526[0:0];
  _RAND_2527 = {1{`RANDOM}};
  r_2527 = _RAND_2527[0:0];
  _RAND_2528 = {1{`RANDOM}};
  r_2528 = _RAND_2528[0:0];
  _RAND_2529 = {1{`RANDOM}};
  r_2529 = _RAND_2529[0:0];
  _RAND_2530 = {1{`RANDOM}};
  r_2530 = _RAND_2530[0:0];
  _RAND_2531 = {1{`RANDOM}};
  r_2531 = _RAND_2531[0:0];
  _RAND_2532 = {1{`RANDOM}};
  r_2532 = _RAND_2532[0:0];
  _RAND_2533 = {1{`RANDOM}};
  r_2533 = _RAND_2533[0:0];
  _RAND_2534 = {1{`RANDOM}};
  r_2534 = _RAND_2534[0:0];
  _RAND_2535 = {1{`RANDOM}};
  r_2535 = _RAND_2535[0:0];
  _RAND_2536 = {1{`RANDOM}};
  r_2536 = _RAND_2536[0:0];
  _RAND_2537 = {1{`RANDOM}};
  r_2537 = _RAND_2537[0:0];
  _RAND_2538 = {1{`RANDOM}};
  r_2538 = _RAND_2538[0:0];
  _RAND_2539 = {1{`RANDOM}};
  r_2539 = _RAND_2539[0:0];
  _RAND_2540 = {1{`RANDOM}};
  r_2540 = _RAND_2540[0:0];
  _RAND_2541 = {1{`RANDOM}};
  r_2541 = _RAND_2541[0:0];
  _RAND_2542 = {1{`RANDOM}};
  r_2542 = _RAND_2542[0:0];
  _RAND_2543 = {1{`RANDOM}};
  r_2543 = _RAND_2543[0:0];
  _RAND_2544 = {1{`RANDOM}};
  r_2544 = _RAND_2544[0:0];
  _RAND_2545 = {1{`RANDOM}};
  r_2545 = _RAND_2545[0:0];
  _RAND_2546 = {1{`RANDOM}};
  r_2546 = _RAND_2546[0:0];
  _RAND_2547 = {1{`RANDOM}};
  r_2547 = _RAND_2547[0:0];
  _RAND_2548 = {1{`RANDOM}};
  r_2548 = _RAND_2548[0:0];
  _RAND_2549 = {1{`RANDOM}};
  r_2549 = _RAND_2549[0:0];
  _RAND_2550 = {1{`RANDOM}};
  r_2550 = _RAND_2550[0:0];
  _RAND_2551 = {1{`RANDOM}};
  r_2551 = _RAND_2551[0:0];
  _RAND_2552 = {1{`RANDOM}};
  r_2552 = _RAND_2552[0:0];
  _RAND_2553 = {1{`RANDOM}};
  r_2553 = _RAND_2553[0:0];
  _RAND_2554 = {1{`RANDOM}};
  r_2554 = _RAND_2554[0:0];
  _RAND_2555 = {1{`RANDOM}};
  r_2555 = _RAND_2555[0:0];
  _RAND_2556 = {1{`RANDOM}};
  r_2556 = _RAND_2556[0:0];
  _RAND_2557 = {1{`RANDOM}};
  r_2557 = _RAND_2557[0:0];
  _RAND_2558 = {1{`RANDOM}};
  r_2558 = _RAND_2558[0:0];
  _RAND_2559 = {1{`RANDOM}};
  r_2559 = _RAND_2559[0:0];
  _RAND_2560 = {1{`RANDOM}};
  r_2560 = _RAND_2560[0:0];
  _RAND_2561 = {1{`RANDOM}};
  r_2561 = _RAND_2561[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule

