module OldestSelection_1(
  input   io_oldest_valid,
  output  io_isOverrided_0
);
  assign io_isOverrided_0 = io_oldest_valid; // @[SelectPolicy.scala 99:29]
endmodule

