module NewIFU(
  input          clock,
  input          reset,
  output         io_ftqInter_fromFtq_req_ready,
  input          io_ftqInter_fromFtq_req_valid,
  input  [38:0]  io_ftqInter_fromFtq_req_bits_startAddr,
  input  [38:0]  io_ftqInter_fromFtq_req_bits_nextlineStart,
  input  [38:0]  io_ftqInter_fromFtq_req_bits_nextStartAddr,
  input          io_ftqInter_fromFtq_req_bits_ftqIdx_flag,
  input  [2:0]   io_ftqInter_fromFtq_req_bits_ftqIdx_value,
  input          io_ftqInter_fromFtq_req_bits_ftqOffset_valid,
  input  [2:0]   io_ftqInter_fromFtq_req_bits_ftqOffset_bits,
  input          io_ftqInter_fromFtq_redirect_valid,
  input          io_ftqInter_fromFtq_redirect_bits_ftqIdx_flag,
  input  [2:0]   io_ftqInter_fromFtq_redirect_bits_ftqIdx_value,
  input  [2:0]   io_ftqInter_fromFtq_redirect_bits_ftqOffset,
  input          io_ftqInter_fromFtq_redirect_bits_level,
  input          io_ftqInter_fromFtq_flushFromBpu_s2_valid,
  input          io_ftqInter_fromFtq_flushFromBpu_s2_bits_flag,
  input  [2:0]   io_ftqInter_fromFtq_flushFromBpu_s2_bits_value,
  input          io_ftqInter_fromFtq_flushFromBpu_s3_valid,
  input          io_ftqInter_fromFtq_flushFromBpu_s3_bits_flag,
  input  [2:0]   io_ftqInter_fromFtq_flushFromBpu_s3_bits_value,
  output         io_ftqInter_toFtq_pdWb_valid,
  output [38:0]  io_ftqInter_toFtq_pdWb_bits_pc_0,
  output [38:0]  io_ftqInter_toFtq_pdWb_bits_pc_1,
  output [38:0]  io_ftqInter_toFtq_pdWb_bits_pc_2,
  output [38:0]  io_ftqInter_toFtq_pdWb_bits_pc_3,
  output [38:0]  io_ftqInter_toFtq_pdWb_bits_pc_4,
  output [38:0]  io_ftqInter_toFtq_pdWb_bits_pc_5,
  output [38:0]  io_ftqInter_toFtq_pdWb_bits_pc_6,
  output [38:0]  io_ftqInter_toFtq_pdWb_bits_pc_7,
  output         io_ftqInter_toFtq_pdWb_bits_pd_0_valid,
  output         io_ftqInter_toFtq_pdWb_bits_pd_0_isRVC,
  output [1:0]   io_ftqInter_toFtq_pdWb_bits_pd_0_brType,
  output         io_ftqInter_toFtq_pdWb_bits_pd_0_isCall,
  output         io_ftqInter_toFtq_pdWb_bits_pd_0_isRet,
  output         io_ftqInter_toFtq_pdWb_bits_pd_1_valid,
  output         io_ftqInter_toFtq_pdWb_bits_pd_1_isRVC,
  output [1:0]   io_ftqInter_toFtq_pdWb_bits_pd_1_brType,
  output         io_ftqInter_toFtq_pdWb_bits_pd_1_isCall,
  output         io_ftqInter_toFtq_pdWb_bits_pd_1_isRet,
  output         io_ftqInter_toFtq_pdWb_bits_pd_2_valid,
  output         io_ftqInter_toFtq_pdWb_bits_pd_2_isRVC,
  output [1:0]   io_ftqInter_toFtq_pdWb_bits_pd_2_brType,
  output         io_ftqInter_toFtq_pdWb_bits_pd_2_isCall,
  output         io_ftqInter_toFtq_pdWb_bits_pd_2_isRet,
  output         io_ftqInter_toFtq_pdWb_bits_pd_3_valid,
  output         io_ftqInter_toFtq_pdWb_bits_pd_3_isRVC,
  output [1:0]   io_ftqInter_toFtq_pdWb_bits_pd_3_brType,
  output         io_ftqInter_toFtq_pdWb_bits_pd_3_isCall,
  output         io_ftqInter_toFtq_pdWb_bits_pd_3_isRet,
  output         io_ftqInter_toFtq_pdWb_bits_pd_4_valid,
  output         io_ftqInter_toFtq_pdWb_bits_pd_4_isRVC,
  output [1:0]   io_ftqInter_toFtq_pdWb_bits_pd_4_brType,
  output         io_ftqInter_toFtq_pdWb_bits_pd_4_isCall,
  output         io_ftqInter_toFtq_pdWb_bits_pd_4_isRet,
  output         io_ftqInter_toFtq_pdWb_bits_pd_5_valid,
  output         io_ftqInter_toFtq_pdWb_bits_pd_5_isRVC,
  output [1:0]   io_ftqInter_toFtq_pdWb_bits_pd_5_brType,
  output         io_ftqInter_toFtq_pdWb_bits_pd_5_isCall,
  output         io_ftqInter_toFtq_pdWb_bits_pd_5_isRet,
  output         io_ftqInter_toFtq_pdWb_bits_pd_6_valid,
  output         io_ftqInter_toFtq_pdWb_bits_pd_6_isRVC,
  output [1:0]   io_ftqInter_toFtq_pdWb_bits_pd_6_brType,
  output         io_ftqInter_toFtq_pdWb_bits_pd_6_isCall,
  output         io_ftqInter_toFtq_pdWb_bits_pd_6_isRet,
  output         io_ftqInter_toFtq_pdWb_bits_pd_7_valid,
  output         io_ftqInter_toFtq_pdWb_bits_pd_7_isRVC,
  output [1:0]   io_ftqInter_toFtq_pdWb_bits_pd_7_brType,
  output         io_ftqInter_toFtq_pdWb_bits_pd_7_isCall,
  output         io_ftqInter_toFtq_pdWb_bits_pd_7_isRet,
  output         io_ftqInter_toFtq_pdWb_bits_ftqIdx_flag,
  output [2:0]   io_ftqInter_toFtq_pdWb_bits_ftqIdx_value,
  output         io_ftqInter_toFtq_pdWb_bits_misOffset_valid,
  output [2:0]   io_ftqInter_toFtq_pdWb_bits_misOffset_bits,
  output         io_ftqInter_toFtq_pdWb_bits_cfiOffset_valid,
  output [38:0]  io_ftqInter_toFtq_pdWb_bits_target,
  output [38:0]  io_ftqInter_toFtq_pdWb_bits_jalTarget,
  output         io_ftqInter_toFtq_pdWb_bits_instrRange_0,
  output         io_ftqInter_toFtq_pdWb_bits_instrRange_1,
  output         io_ftqInter_toFtq_pdWb_bits_instrRange_2,
  output         io_ftqInter_toFtq_pdWb_bits_instrRange_3,
  output         io_ftqInter_toFtq_pdWb_bits_instrRange_4,
  output         io_ftqInter_toFtq_pdWb_bits_instrRange_5,
  output         io_ftqInter_toFtq_pdWb_bits_instrRange_6,
  output         io_ftqInter_toFtq_pdWb_bits_instrRange_7,
  input          io_icacheInter_icacheReady,
  input          io_icacheInter_resp_0_valid,
  input  [38:0]  io_icacheInter_resp_0_bits_vaddr,
  input  [511:0] io_icacheInter_resp_0_bits_registerData,
  input  [511:0] io_icacheInter_resp_0_bits_sramData,
  input          io_icacheInter_resp_0_bits_select,
  input  [35:0]  io_icacheInter_resp_0_bits_paddr,
  input          io_icacheInter_resp_0_bits_tlbExcp_pageFault,
  input          io_icacheInter_resp_0_bits_tlbExcp_accessFault,
  input          io_icacheInter_resp_0_bits_tlbExcp_mmio,
  input          io_icacheInter_resp_1_valid,
  input  [38:0]  io_icacheInter_resp_1_bits_vaddr,
  input  [511:0] io_icacheInter_resp_1_bits_registerData,
  input  [511:0] io_icacheInter_resp_1_bits_sramData,
  input          io_icacheInter_resp_1_bits_select,
  input          io_icacheInter_resp_1_bits_tlbExcp_pageFault,
  input          io_icacheInter_resp_1_bits_tlbExcp_accessFault,
  output         io_icacheStop,
  input          io_icachePerfInfo_only_0_hit,
  input          io_icachePerfInfo_only_0_miss,
  input          io_icachePerfInfo_hit_0_hit_1,
  input          io_icachePerfInfo_hit_0_miss_1,
  input          io_icachePerfInfo_miss_0_hit_1,
  input          io_icachePerfInfo_miss_0_miss_1,
  input          io_icachePerfInfo_hit_0_except_1,
  input          io_icachePerfInfo_miss_0_except_1,
  input          io_icachePerfInfo_except_0,
  input          io_icachePerfInfo_bank_hit_1,
  input          io_icachePerfInfo_hit,
  input          io_toIbuffer_ready,
  output         io_toIbuffer_valid,
  output [31:0]  io_toIbuffer_bits_instrs_0,
  output [31:0]  io_toIbuffer_bits_instrs_1,
  output [31:0]  io_toIbuffer_bits_instrs_2,
  output [31:0]  io_toIbuffer_bits_instrs_3,
  output [31:0]  io_toIbuffer_bits_instrs_4,
  output [31:0]  io_toIbuffer_bits_instrs_5,
  output [31:0]  io_toIbuffer_bits_instrs_6,
  output [31:0]  io_toIbuffer_bits_instrs_7,
  output [7:0]   io_toIbuffer_bits_valid,
  output [7:0]   io_toIbuffer_bits_enqEnable,
  output         io_toIbuffer_bits_pd_0_isRVC,
  output [1:0]   io_toIbuffer_bits_pd_0_brType,
  output         io_toIbuffer_bits_pd_0_isCall,
  output         io_toIbuffer_bits_pd_0_isRet,
  output         io_toIbuffer_bits_pd_1_isRVC,
  output [1:0]   io_toIbuffer_bits_pd_1_brType,
  output         io_toIbuffer_bits_pd_1_isCall,
  output         io_toIbuffer_bits_pd_1_isRet,
  output         io_toIbuffer_bits_pd_2_isRVC,
  output [1:0]   io_toIbuffer_bits_pd_2_brType,
  output         io_toIbuffer_bits_pd_2_isCall,
  output         io_toIbuffer_bits_pd_2_isRet,
  output         io_toIbuffer_bits_pd_3_isRVC,
  output [1:0]   io_toIbuffer_bits_pd_3_brType,
  output         io_toIbuffer_bits_pd_3_isCall,
  output         io_toIbuffer_bits_pd_3_isRet,
  output         io_toIbuffer_bits_pd_4_isRVC,
  output [1:0]   io_toIbuffer_bits_pd_4_brType,
  output         io_toIbuffer_bits_pd_4_isCall,
  output         io_toIbuffer_bits_pd_4_isRet,
  output         io_toIbuffer_bits_pd_5_isRVC,
  output [1:0]   io_toIbuffer_bits_pd_5_brType,
  output         io_toIbuffer_bits_pd_5_isCall,
  output         io_toIbuffer_bits_pd_5_isRet,
  output         io_toIbuffer_bits_pd_6_isRVC,
  output [1:0]   io_toIbuffer_bits_pd_6_brType,
  output         io_toIbuffer_bits_pd_6_isCall,
  output         io_toIbuffer_bits_pd_6_isRet,
  output         io_toIbuffer_bits_pd_7_isRVC,
  output [1:0]   io_toIbuffer_bits_pd_7_brType,
  output         io_toIbuffer_bits_pd_7_isCall,
  output         io_toIbuffer_bits_pd_7_isRet,
  output [9:0]   io_toIbuffer_bits_foldpc_0,
  output [9:0]   io_toIbuffer_bits_foldpc_1,
  output [9:0]   io_toIbuffer_bits_foldpc_2,
  output [9:0]   io_toIbuffer_bits_foldpc_3,
  output [9:0]   io_toIbuffer_bits_foldpc_4,
  output [9:0]   io_toIbuffer_bits_foldpc_5,
  output [9:0]   io_toIbuffer_bits_foldpc_6,
  output [9:0]   io_toIbuffer_bits_foldpc_7,
  output         io_toIbuffer_bits_ftqPtr_flag,
  output [2:0]   io_toIbuffer_bits_ftqPtr_value,
  output         io_toIbuffer_bits_ftqOffset_0_valid,
  output         io_toIbuffer_bits_ftqOffset_1_valid,
  output         io_toIbuffer_bits_ftqOffset_2_valid,
  output         io_toIbuffer_bits_ftqOffset_3_valid,
  output         io_toIbuffer_bits_ftqOffset_4_valid,
  output         io_toIbuffer_bits_ftqOffset_5_valid,
  output         io_toIbuffer_bits_ftqOffset_6_valid,
  output         io_toIbuffer_bits_ftqOffset_7_valid,
  output         io_toIbuffer_bits_ipf_0,
  output         io_toIbuffer_bits_ipf_1,
  output         io_toIbuffer_bits_ipf_2,
  output         io_toIbuffer_bits_ipf_3,
  output         io_toIbuffer_bits_ipf_4,
  output         io_toIbuffer_bits_ipf_5,
  output         io_toIbuffer_bits_ipf_6,
  output         io_toIbuffer_bits_ipf_7,
  output         io_toIbuffer_bits_acf_0,
  output         io_toIbuffer_bits_acf_1,
  output         io_toIbuffer_bits_acf_2,
  output         io_toIbuffer_bits_acf_3,
  output         io_toIbuffer_bits_acf_4,
  output         io_toIbuffer_bits_acf_5,
  output         io_toIbuffer_bits_acf_6,
  output         io_toIbuffer_bits_acf_7,
  output         io_toIbuffer_bits_crossPageIPFFix_0,
  output         io_toIbuffer_bits_crossPageIPFFix_1,
  output         io_toIbuffer_bits_crossPageIPFFix_2,
  output         io_toIbuffer_bits_crossPageIPFFix_3,
  output         io_toIbuffer_bits_crossPageIPFFix_4,
  output         io_toIbuffer_bits_crossPageIPFFix_5,
  output         io_toIbuffer_bits_crossPageIPFFix_6,
  output         io_toIbuffer_bits_crossPageIPFFix_7,
  output         io_toIbuffer_bits_triggered_0_frontendHit_0,
  output         io_toIbuffer_bits_triggered_0_frontendHit_1,
  output         io_toIbuffer_bits_triggered_0_frontendHit_2,
  output         io_toIbuffer_bits_triggered_0_frontendHit_3,
  output         io_toIbuffer_bits_triggered_0_backendEn_0,
  output         io_toIbuffer_bits_triggered_0_backendEn_1,
  output         io_toIbuffer_bits_triggered_1_frontendHit_0,
  output         io_toIbuffer_bits_triggered_1_frontendHit_1,
  output         io_toIbuffer_bits_triggered_1_frontendHit_2,
  output         io_toIbuffer_bits_triggered_1_frontendHit_3,
  output         io_toIbuffer_bits_triggered_1_backendEn_0,
  output         io_toIbuffer_bits_triggered_1_backendEn_1,
  output         io_toIbuffer_bits_triggered_2_frontendHit_0,
  output         io_toIbuffer_bits_triggered_2_frontendHit_1,
  output         io_toIbuffer_bits_triggered_2_frontendHit_2,
  output         io_toIbuffer_bits_triggered_2_frontendHit_3,
  output         io_toIbuffer_bits_triggered_2_backendEn_0,
  output         io_toIbuffer_bits_triggered_2_backendEn_1,
  output         io_toIbuffer_bits_triggered_3_frontendHit_0,
  output         io_toIbuffer_bits_triggered_3_frontendHit_1,
  output         io_toIbuffer_bits_triggered_3_frontendHit_2,
  output         io_toIbuffer_bits_triggered_3_frontendHit_3,
  output         io_toIbuffer_bits_triggered_3_backendEn_0,
  output         io_toIbuffer_bits_triggered_3_backendEn_1,
  output         io_toIbuffer_bits_triggered_4_frontendHit_0,
  output         io_toIbuffer_bits_triggered_4_frontendHit_1,
  output         io_toIbuffer_bits_triggered_4_frontendHit_2,
  output         io_toIbuffer_bits_triggered_4_frontendHit_3,
  output         io_toIbuffer_bits_triggered_4_backendEn_0,
  output         io_toIbuffer_bits_triggered_4_backendEn_1,
  output         io_toIbuffer_bits_triggered_5_frontendHit_0,
  output         io_toIbuffer_bits_triggered_5_frontendHit_1,
  output         io_toIbuffer_bits_triggered_5_frontendHit_2,
  output         io_toIbuffer_bits_triggered_5_frontendHit_3,
  output         io_toIbuffer_bits_triggered_5_backendEn_0,
  output         io_toIbuffer_bits_triggered_5_backendEn_1,
  output         io_toIbuffer_bits_triggered_6_frontendHit_0,
  output         io_toIbuffer_bits_triggered_6_frontendHit_1,
  output         io_toIbuffer_bits_triggered_6_frontendHit_2,
  output         io_toIbuffer_bits_triggered_6_frontendHit_3,
  output         io_toIbuffer_bits_triggered_6_backendEn_0,
  output         io_toIbuffer_bits_triggered_6_backendEn_1,
  output         io_toIbuffer_bits_triggered_7_frontendHit_0,
  output         io_toIbuffer_bits_triggered_7_frontendHit_1,
  output         io_toIbuffer_bits_triggered_7_frontendHit_2,
  output         io_toIbuffer_bits_triggered_7_frontendHit_3,
  output         io_toIbuffer_bits_triggered_7_backendEn_0,
  output         io_toIbuffer_bits_triggered_7_backendEn_1,
  output         io_uncacheInter_fromUncache_ready,
  input          io_uncacheInter_fromUncache_valid,
  input  [31:0]  io_uncacheInter_fromUncache_bits_data,
  input          io_uncacheInter_toUncache_ready,
  output         io_uncacheInter_toUncache_valid,
  output [35:0]  io_uncacheInter_toUncache_bits_addr,
  input          io_frontendTrigger_t_valid,
  input  [1:0]   io_frontendTrigger_t_bits_addr,
  input  [1:0]   io_frontendTrigger_t_bits_tdata_matchType,
  input          io_frontendTrigger_t_bits_tdata_select,
  input          io_frontendTrigger_t_bits_tdata_timing,
  input          io_frontendTrigger_t_bits_tdata_chain,
  input  [63:0]  io_frontendTrigger_t_bits_tdata_tdata2,
  input          io_csrTriggerEnable_0,
  input          io_csrTriggerEnable_1,
  input          io_csrTriggerEnable_2,
  input          io_csrTriggerEnable_3,
  input          io_rob_commits_0_valid,
  input          io_rob_commits_0_bits_ftqIdx_flag,
  input  [2:0]   io_rob_commits_0_bits_ftqIdx_value,
  input  [2:0]   io_rob_commits_0_bits_ftqOffset,
  input          io_rob_commits_1_valid,
  input          io_rob_commits_1_bits_ftqIdx_flag,
  input  [2:0]   io_rob_commits_1_bits_ftqIdx_value,
  input  [2:0]   io_rob_commits_1_bits_ftqOffset,
  output         io_iTLBInter_req_valid,
  output [38:0]  io_iTLBInter_req_bits_vaddr,
  input  [35:0]  io_iTLBInter_resp_bits_paddr_0,
  input          io_iTLBInter_resp_bits_miss,
  input          io_iTLBInter_resp_bits_excp_0_pf_instr,
  input          io_iTLBInter_resp_bits_excp_0_af_instr,
  output [35:0]  io_pmp_req_bits_addr,
  input          io_pmp_resp_instr,
  input          io_pmp_resp_mmio,
  output         io_mmioCommitRead_mmioFtqPtr_flag,
  output [2:0]   io_mmioCommitRead_mmioFtqPtr_value,
  input          io_mmioCommitRead_mmioLastCommit,
  output [5:0]   io_perf_0_value,
  output [5:0]   io_perf_1_value,
  output [5:0]   io_perf_2_value,
  output [5:0]   io_perf_3_value,
  output [5:0]   io_perf_4_value,
  output [5:0]   io_perf_5_value,
  output [5:0]   io_perf_6_value,
  output [5:0]   io_perf_7_value,
  output [5:0]   io_perf_8_value,
  output [5:0]   io_perf_9_value,
  output [5:0]   io_perf_10_value,
  output [5:0]   io_perf_11_value,
  output [5:0]   io_perf_12_value
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [63:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [63:0] _RAND_39;
  reg [63:0] _RAND_40;
  reg [63:0] _RAND_41;
  reg [63:0] _RAND_42;
  reg [63:0] _RAND_43;
  reg [63:0] _RAND_44;
  reg [63:0] _RAND_45;
  reg [63:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [63:0] _RAND_56;
  reg [63:0] _RAND_57;
  reg [63:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [63:0] _RAND_119;
  reg [63:0] _RAND_120;
  reg [63:0] _RAND_121;
  reg [63:0] _RAND_122;
  reg [63:0] _RAND_123;
  reg [63:0] _RAND_124;
  reg [63:0] _RAND_125;
  reg [63:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [63:0] _RAND_143;
  reg [63:0] _RAND_144;
  reg [63:0] _RAND_145;
  reg [63:0] _RAND_146;
  reg [63:0] _RAND_147;
  reg [63:0] _RAND_148;
  reg [63:0] _RAND_149;
  reg [63:0] _RAND_150;
  reg [63:0] _RAND_151;
  reg [63:0] _RAND_152;
  reg [63:0] _RAND_153;
  reg [63:0] _RAND_154;
  reg [63:0] _RAND_155;
  reg [63:0] _RAND_156;
  reg [63:0] _RAND_157;
  reg [63:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [63:0] _RAND_183;
  reg [63:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [63:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [63:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [63:0] _RAND_216;
  reg [63:0] _RAND_217;
  reg [63:0] _RAND_218;
  reg [63:0] _RAND_219;
  reg [63:0] _RAND_220;
  reg [63:0] _RAND_221;
  reg [63:0] _RAND_222;
  reg [63:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [63:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [63:0] _RAND_305;
  reg [63:0] _RAND_306;
`endif // RANDOMIZE_REG_INIT
  wire [15:0] preDecoders_0_io_in_data_0; // @[IFU.scala 142:46]
  wire [15:0] preDecoders_0_io_in_data_1; // @[IFU.scala 142:46]
  wire [15:0] preDecoders_0_io_in_data_2; // @[IFU.scala 142:46]
  wire [15:0] preDecoders_0_io_in_data_3; // @[IFU.scala 142:46]
  wire [15:0] preDecoders_0_io_in_data_4; // @[IFU.scala 142:46]
  wire [15:0] preDecoders_0_io_in_data_5; // @[IFU.scala 142:46]
  wire [15:0] preDecoders_0_io_in_data_6; // @[IFU.scala 142:46]
  wire [15:0] preDecoders_0_io_in_data_7; // @[IFU.scala 142:46]
  wire [15:0] preDecoders_0_io_in_data_8; // @[IFU.scala 142:46]
  wire  preDecoders_0_io_out_pd_0_isRVC; // @[IFU.scala 142:46]
  wire [1:0] preDecoders_0_io_out_pd_0_brType; // @[IFU.scala 142:46]
  wire  preDecoders_0_io_out_pd_0_isCall; // @[IFU.scala 142:46]
  wire  preDecoders_0_io_out_pd_0_isRet; // @[IFU.scala 142:46]
  wire  preDecoders_0_io_out_pd_1_valid; // @[IFU.scala 142:46]
  wire  preDecoders_0_io_out_pd_1_isRVC; // @[IFU.scala 142:46]
  wire [1:0] preDecoders_0_io_out_pd_1_brType; // @[IFU.scala 142:46]
  wire  preDecoders_0_io_out_pd_1_isCall; // @[IFU.scala 142:46]
  wire  preDecoders_0_io_out_pd_1_isRet; // @[IFU.scala 142:46]
  wire  preDecoders_0_io_out_pd_2_valid; // @[IFU.scala 142:46]
  wire  preDecoders_0_io_out_pd_2_isRVC; // @[IFU.scala 142:46]
  wire [1:0] preDecoders_0_io_out_pd_2_brType; // @[IFU.scala 142:46]
  wire  preDecoders_0_io_out_pd_2_isCall; // @[IFU.scala 142:46]
  wire  preDecoders_0_io_out_pd_2_isRet; // @[IFU.scala 142:46]
  wire  preDecoders_0_io_out_pd_3_valid; // @[IFU.scala 142:46]
  wire  preDecoders_0_io_out_pd_3_isRVC; // @[IFU.scala 142:46]
  wire [1:0] preDecoders_0_io_out_pd_3_brType; // @[IFU.scala 142:46]
  wire  preDecoders_0_io_out_pd_3_isCall; // @[IFU.scala 142:46]
  wire  preDecoders_0_io_out_pd_3_isRet; // @[IFU.scala 142:46]
  wire  preDecoders_0_io_out_pd_4_valid; // @[IFU.scala 142:46]
  wire  preDecoders_0_io_out_pd_4_isRVC; // @[IFU.scala 142:46]
  wire [1:0] preDecoders_0_io_out_pd_4_brType; // @[IFU.scala 142:46]
  wire  preDecoders_0_io_out_pd_4_isCall; // @[IFU.scala 142:46]
  wire  preDecoders_0_io_out_pd_4_isRet; // @[IFU.scala 142:46]
  wire  preDecoders_0_io_out_pd_5_valid; // @[IFU.scala 142:46]
  wire  preDecoders_0_io_out_pd_5_isRVC; // @[IFU.scala 142:46]
  wire [1:0] preDecoders_0_io_out_pd_5_brType; // @[IFU.scala 142:46]
  wire  preDecoders_0_io_out_pd_5_isCall; // @[IFU.scala 142:46]
  wire  preDecoders_0_io_out_pd_5_isRet; // @[IFU.scala 142:46]
  wire  preDecoders_0_io_out_pd_6_valid; // @[IFU.scala 142:46]
  wire  preDecoders_0_io_out_pd_6_isRVC; // @[IFU.scala 142:46]
  wire [1:0] preDecoders_0_io_out_pd_6_brType; // @[IFU.scala 142:46]
  wire  preDecoders_0_io_out_pd_6_isCall; // @[IFU.scala 142:46]
  wire  preDecoders_0_io_out_pd_6_isRet; // @[IFU.scala 142:46]
  wire  preDecoders_0_io_out_pd_7_valid; // @[IFU.scala 142:46]
  wire  preDecoders_0_io_out_pd_7_isRVC; // @[IFU.scala 142:46]
  wire [1:0] preDecoders_0_io_out_pd_7_brType; // @[IFU.scala 142:46]
  wire  preDecoders_0_io_out_pd_7_isCall; // @[IFU.scala 142:46]
  wire  preDecoders_0_io_out_pd_7_isRet; // @[IFU.scala 142:46]
  wire  preDecoders_0_io_out_hasHalfValid_2; // @[IFU.scala 142:46]
  wire  preDecoders_0_io_out_hasHalfValid_3; // @[IFU.scala 142:46]
  wire  preDecoders_0_io_out_hasHalfValid_4; // @[IFU.scala 142:46]
  wire  preDecoders_0_io_out_hasHalfValid_5; // @[IFU.scala 142:46]
  wire  preDecoders_0_io_out_hasHalfValid_6; // @[IFU.scala 142:46]
  wire  preDecoders_0_io_out_hasHalfValid_7; // @[IFU.scala 142:46]
  wire [31:0] preDecoders_0_io_out_instr_0; // @[IFU.scala 142:46]
  wire [31:0] preDecoders_0_io_out_instr_1; // @[IFU.scala 142:46]
  wire [31:0] preDecoders_0_io_out_instr_2; // @[IFU.scala 142:46]
  wire [31:0] preDecoders_0_io_out_instr_3; // @[IFU.scala 142:46]
  wire [31:0] preDecoders_0_io_out_instr_4; // @[IFU.scala 142:46]
  wire [31:0] preDecoders_0_io_out_instr_5; // @[IFU.scala 142:46]
  wire [31:0] preDecoders_0_io_out_instr_6; // @[IFU.scala 142:46]
  wire [31:0] preDecoders_0_io_out_instr_7; // @[IFU.scala 142:46]
  wire [63:0] preDecoders_0_io_out_jumpOffset_0; // @[IFU.scala 142:46]
  wire [63:0] preDecoders_0_io_out_jumpOffset_1; // @[IFU.scala 142:46]
  wire [63:0] preDecoders_0_io_out_jumpOffset_2; // @[IFU.scala 142:46]
  wire [63:0] preDecoders_0_io_out_jumpOffset_3; // @[IFU.scala 142:46]
  wire [63:0] preDecoders_0_io_out_jumpOffset_4; // @[IFU.scala 142:46]
  wire [63:0] preDecoders_0_io_out_jumpOffset_5; // @[IFU.scala 142:46]
  wire [63:0] preDecoders_0_io_out_jumpOffset_6; // @[IFU.scala 142:46]
  wire [63:0] preDecoders_0_io_out_jumpOffset_7; // @[IFU.scala 142:46]
  wire [15:0] preDecoders_1_io_in_data_0; // @[IFU.scala 142:46]
  wire [15:0] preDecoders_1_io_in_data_1; // @[IFU.scala 142:46]
  wire [15:0] preDecoders_1_io_in_data_2; // @[IFU.scala 142:46]
  wire [15:0] preDecoders_1_io_in_data_3; // @[IFU.scala 142:46]
  wire [15:0] preDecoders_1_io_in_data_4; // @[IFU.scala 142:46]
  wire [15:0] preDecoders_1_io_in_data_5; // @[IFU.scala 142:46]
  wire [15:0] preDecoders_1_io_in_data_6; // @[IFU.scala 142:46]
  wire [15:0] preDecoders_1_io_in_data_7; // @[IFU.scala 142:46]
  wire [15:0] preDecoders_1_io_in_data_8; // @[IFU.scala 142:46]
  wire  preDecoders_1_io_out_pd_0_isRVC; // @[IFU.scala 142:46]
  wire [1:0] preDecoders_1_io_out_pd_0_brType; // @[IFU.scala 142:46]
  wire  preDecoders_1_io_out_pd_0_isCall; // @[IFU.scala 142:46]
  wire  preDecoders_1_io_out_pd_0_isRet; // @[IFU.scala 142:46]
  wire  preDecoders_1_io_out_pd_1_valid; // @[IFU.scala 142:46]
  wire  preDecoders_1_io_out_pd_1_isRVC; // @[IFU.scala 142:46]
  wire [1:0] preDecoders_1_io_out_pd_1_brType; // @[IFU.scala 142:46]
  wire  preDecoders_1_io_out_pd_1_isCall; // @[IFU.scala 142:46]
  wire  preDecoders_1_io_out_pd_1_isRet; // @[IFU.scala 142:46]
  wire  preDecoders_1_io_out_pd_2_valid; // @[IFU.scala 142:46]
  wire  preDecoders_1_io_out_pd_2_isRVC; // @[IFU.scala 142:46]
  wire [1:0] preDecoders_1_io_out_pd_2_brType; // @[IFU.scala 142:46]
  wire  preDecoders_1_io_out_pd_2_isCall; // @[IFU.scala 142:46]
  wire  preDecoders_1_io_out_pd_2_isRet; // @[IFU.scala 142:46]
  wire  preDecoders_1_io_out_pd_3_valid; // @[IFU.scala 142:46]
  wire  preDecoders_1_io_out_pd_3_isRVC; // @[IFU.scala 142:46]
  wire [1:0] preDecoders_1_io_out_pd_3_brType; // @[IFU.scala 142:46]
  wire  preDecoders_1_io_out_pd_3_isCall; // @[IFU.scala 142:46]
  wire  preDecoders_1_io_out_pd_3_isRet; // @[IFU.scala 142:46]
  wire  preDecoders_1_io_out_pd_4_valid; // @[IFU.scala 142:46]
  wire  preDecoders_1_io_out_pd_4_isRVC; // @[IFU.scala 142:46]
  wire [1:0] preDecoders_1_io_out_pd_4_brType; // @[IFU.scala 142:46]
  wire  preDecoders_1_io_out_pd_4_isCall; // @[IFU.scala 142:46]
  wire  preDecoders_1_io_out_pd_4_isRet; // @[IFU.scala 142:46]
  wire  preDecoders_1_io_out_pd_5_valid; // @[IFU.scala 142:46]
  wire  preDecoders_1_io_out_pd_5_isRVC; // @[IFU.scala 142:46]
  wire [1:0] preDecoders_1_io_out_pd_5_brType; // @[IFU.scala 142:46]
  wire  preDecoders_1_io_out_pd_5_isCall; // @[IFU.scala 142:46]
  wire  preDecoders_1_io_out_pd_5_isRet; // @[IFU.scala 142:46]
  wire  preDecoders_1_io_out_pd_6_valid; // @[IFU.scala 142:46]
  wire  preDecoders_1_io_out_pd_6_isRVC; // @[IFU.scala 142:46]
  wire [1:0] preDecoders_1_io_out_pd_6_brType; // @[IFU.scala 142:46]
  wire  preDecoders_1_io_out_pd_6_isCall; // @[IFU.scala 142:46]
  wire  preDecoders_1_io_out_pd_6_isRet; // @[IFU.scala 142:46]
  wire  preDecoders_1_io_out_pd_7_valid; // @[IFU.scala 142:46]
  wire  preDecoders_1_io_out_pd_7_isRVC; // @[IFU.scala 142:46]
  wire [1:0] preDecoders_1_io_out_pd_7_brType; // @[IFU.scala 142:46]
  wire  preDecoders_1_io_out_pd_7_isCall; // @[IFU.scala 142:46]
  wire  preDecoders_1_io_out_pd_7_isRet; // @[IFU.scala 142:46]
  wire  preDecoders_1_io_out_hasHalfValid_2; // @[IFU.scala 142:46]
  wire  preDecoders_1_io_out_hasHalfValid_3; // @[IFU.scala 142:46]
  wire  preDecoders_1_io_out_hasHalfValid_4; // @[IFU.scala 142:46]
  wire  preDecoders_1_io_out_hasHalfValid_5; // @[IFU.scala 142:46]
  wire  preDecoders_1_io_out_hasHalfValid_6; // @[IFU.scala 142:46]
  wire  preDecoders_1_io_out_hasHalfValid_7; // @[IFU.scala 142:46]
  wire [31:0] preDecoders_1_io_out_instr_0; // @[IFU.scala 142:46]
  wire [31:0] preDecoders_1_io_out_instr_1; // @[IFU.scala 142:46]
  wire [31:0] preDecoders_1_io_out_instr_2; // @[IFU.scala 142:46]
  wire [31:0] preDecoders_1_io_out_instr_3; // @[IFU.scala 142:46]
  wire [31:0] preDecoders_1_io_out_instr_4; // @[IFU.scala 142:46]
  wire [31:0] preDecoders_1_io_out_instr_5; // @[IFU.scala 142:46]
  wire [31:0] preDecoders_1_io_out_instr_6; // @[IFU.scala 142:46]
  wire [31:0] preDecoders_1_io_out_instr_7; // @[IFU.scala 142:46]
  wire [63:0] preDecoders_1_io_out_jumpOffset_0; // @[IFU.scala 142:46]
  wire [63:0] preDecoders_1_io_out_jumpOffset_1; // @[IFU.scala 142:46]
  wire [63:0] preDecoders_1_io_out_jumpOffset_2; // @[IFU.scala 142:46]
  wire [63:0] preDecoders_1_io_out_jumpOffset_3; // @[IFU.scala 142:46]
  wire [63:0] preDecoders_1_io_out_jumpOffset_4; // @[IFU.scala 142:46]
  wire [63:0] preDecoders_1_io_out_jumpOffset_5; // @[IFU.scala 142:46]
  wire [63:0] preDecoders_1_io_out_jumpOffset_6; // @[IFU.scala 142:46]
  wire [63:0] preDecoders_1_io_out_jumpOffset_7; // @[IFU.scala 142:46]
  wire [15:0] preDecoders_2_io_in_data_0; // @[IFU.scala 142:46]
  wire [15:0] preDecoders_2_io_in_data_1; // @[IFU.scala 142:46]
  wire [15:0] preDecoders_2_io_in_data_2; // @[IFU.scala 142:46]
  wire [15:0] preDecoders_2_io_in_data_3; // @[IFU.scala 142:46]
  wire [15:0] preDecoders_2_io_in_data_4; // @[IFU.scala 142:46]
  wire [15:0] preDecoders_2_io_in_data_5; // @[IFU.scala 142:46]
  wire [15:0] preDecoders_2_io_in_data_6; // @[IFU.scala 142:46]
  wire [15:0] preDecoders_2_io_in_data_7; // @[IFU.scala 142:46]
  wire [15:0] preDecoders_2_io_in_data_8; // @[IFU.scala 142:46]
  wire  preDecoders_2_io_out_pd_0_isRVC; // @[IFU.scala 142:46]
  wire [1:0] preDecoders_2_io_out_pd_0_brType; // @[IFU.scala 142:46]
  wire  preDecoders_2_io_out_pd_0_isCall; // @[IFU.scala 142:46]
  wire  preDecoders_2_io_out_pd_0_isRet; // @[IFU.scala 142:46]
  wire  preDecoders_2_io_out_pd_1_valid; // @[IFU.scala 142:46]
  wire  preDecoders_2_io_out_pd_1_isRVC; // @[IFU.scala 142:46]
  wire [1:0] preDecoders_2_io_out_pd_1_brType; // @[IFU.scala 142:46]
  wire  preDecoders_2_io_out_pd_1_isCall; // @[IFU.scala 142:46]
  wire  preDecoders_2_io_out_pd_1_isRet; // @[IFU.scala 142:46]
  wire  preDecoders_2_io_out_pd_2_valid; // @[IFU.scala 142:46]
  wire  preDecoders_2_io_out_pd_2_isRVC; // @[IFU.scala 142:46]
  wire [1:0] preDecoders_2_io_out_pd_2_brType; // @[IFU.scala 142:46]
  wire  preDecoders_2_io_out_pd_2_isCall; // @[IFU.scala 142:46]
  wire  preDecoders_2_io_out_pd_2_isRet; // @[IFU.scala 142:46]
  wire  preDecoders_2_io_out_pd_3_valid; // @[IFU.scala 142:46]
  wire  preDecoders_2_io_out_pd_3_isRVC; // @[IFU.scala 142:46]
  wire [1:0] preDecoders_2_io_out_pd_3_brType; // @[IFU.scala 142:46]
  wire  preDecoders_2_io_out_pd_3_isCall; // @[IFU.scala 142:46]
  wire  preDecoders_2_io_out_pd_3_isRet; // @[IFU.scala 142:46]
  wire  preDecoders_2_io_out_pd_4_valid; // @[IFU.scala 142:46]
  wire  preDecoders_2_io_out_pd_4_isRVC; // @[IFU.scala 142:46]
  wire [1:0] preDecoders_2_io_out_pd_4_brType; // @[IFU.scala 142:46]
  wire  preDecoders_2_io_out_pd_4_isCall; // @[IFU.scala 142:46]
  wire  preDecoders_2_io_out_pd_4_isRet; // @[IFU.scala 142:46]
  wire  preDecoders_2_io_out_pd_5_valid; // @[IFU.scala 142:46]
  wire  preDecoders_2_io_out_pd_5_isRVC; // @[IFU.scala 142:46]
  wire [1:0] preDecoders_2_io_out_pd_5_brType; // @[IFU.scala 142:46]
  wire  preDecoders_2_io_out_pd_5_isCall; // @[IFU.scala 142:46]
  wire  preDecoders_2_io_out_pd_5_isRet; // @[IFU.scala 142:46]
  wire  preDecoders_2_io_out_pd_6_valid; // @[IFU.scala 142:46]
  wire  preDecoders_2_io_out_pd_6_isRVC; // @[IFU.scala 142:46]
  wire [1:0] preDecoders_2_io_out_pd_6_brType; // @[IFU.scala 142:46]
  wire  preDecoders_2_io_out_pd_6_isCall; // @[IFU.scala 142:46]
  wire  preDecoders_2_io_out_pd_6_isRet; // @[IFU.scala 142:46]
  wire  preDecoders_2_io_out_pd_7_valid; // @[IFU.scala 142:46]
  wire  preDecoders_2_io_out_pd_7_isRVC; // @[IFU.scala 142:46]
  wire [1:0] preDecoders_2_io_out_pd_7_brType; // @[IFU.scala 142:46]
  wire  preDecoders_2_io_out_pd_7_isCall; // @[IFU.scala 142:46]
  wire  preDecoders_2_io_out_pd_7_isRet; // @[IFU.scala 142:46]
  wire  preDecoders_2_io_out_hasHalfValid_2; // @[IFU.scala 142:46]
  wire  preDecoders_2_io_out_hasHalfValid_3; // @[IFU.scala 142:46]
  wire  preDecoders_2_io_out_hasHalfValid_4; // @[IFU.scala 142:46]
  wire  preDecoders_2_io_out_hasHalfValid_5; // @[IFU.scala 142:46]
  wire  preDecoders_2_io_out_hasHalfValid_6; // @[IFU.scala 142:46]
  wire  preDecoders_2_io_out_hasHalfValid_7; // @[IFU.scala 142:46]
  wire [31:0] preDecoders_2_io_out_instr_0; // @[IFU.scala 142:46]
  wire [31:0] preDecoders_2_io_out_instr_1; // @[IFU.scala 142:46]
  wire [31:0] preDecoders_2_io_out_instr_2; // @[IFU.scala 142:46]
  wire [31:0] preDecoders_2_io_out_instr_3; // @[IFU.scala 142:46]
  wire [31:0] preDecoders_2_io_out_instr_4; // @[IFU.scala 142:46]
  wire [31:0] preDecoders_2_io_out_instr_5; // @[IFU.scala 142:46]
  wire [31:0] preDecoders_2_io_out_instr_6; // @[IFU.scala 142:46]
  wire [31:0] preDecoders_2_io_out_instr_7; // @[IFU.scala 142:46]
  wire [63:0] preDecoders_2_io_out_jumpOffset_0; // @[IFU.scala 142:46]
  wire [63:0] preDecoders_2_io_out_jumpOffset_1; // @[IFU.scala 142:46]
  wire [63:0] preDecoders_2_io_out_jumpOffset_2; // @[IFU.scala 142:46]
  wire [63:0] preDecoders_2_io_out_jumpOffset_3; // @[IFU.scala 142:46]
  wire [63:0] preDecoders_2_io_out_jumpOffset_4; // @[IFU.scala 142:46]
  wire [63:0] preDecoders_2_io_out_jumpOffset_5; // @[IFU.scala 142:46]
  wire [63:0] preDecoders_2_io_out_jumpOffset_6; // @[IFU.scala 142:46]
  wire [63:0] preDecoders_2_io_out_jumpOffset_7; // @[IFU.scala 142:46]
  wire [15:0] preDecoders_3_io_in_data_0; // @[IFU.scala 142:46]
  wire [15:0] preDecoders_3_io_in_data_1; // @[IFU.scala 142:46]
  wire [15:0] preDecoders_3_io_in_data_2; // @[IFU.scala 142:46]
  wire [15:0] preDecoders_3_io_in_data_3; // @[IFU.scala 142:46]
  wire [15:0] preDecoders_3_io_in_data_4; // @[IFU.scala 142:46]
  wire [15:0] preDecoders_3_io_in_data_5; // @[IFU.scala 142:46]
  wire [15:0] preDecoders_3_io_in_data_6; // @[IFU.scala 142:46]
  wire [15:0] preDecoders_3_io_in_data_7; // @[IFU.scala 142:46]
  wire [15:0] preDecoders_3_io_in_data_8; // @[IFU.scala 142:46]
  wire  preDecoders_3_io_out_pd_0_isRVC; // @[IFU.scala 142:46]
  wire [1:0] preDecoders_3_io_out_pd_0_brType; // @[IFU.scala 142:46]
  wire  preDecoders_3_io_out_pd_0_isCall; // @[IFU.scala 142:46]
  wire  preDecoders_3_io_out_pd_0_isRet; // @[IFU.scala 142:46]
  wire  preDecoders_3_io_out_pd_1_valid; // @[IFU.scala 142:46]
  wire  preDecoders_3_io_out_pd_1_isRVC; // @[IFU.scala 142:46]
  wire [1:0] preDecoders_3_io_out_pd_1_brType; // @[IFU.scala 142:46]
  wire  preDecoders_3_io_out_pd_1_isCall; // @[IFU.scala 142:46]
  wire  preDecoders_3_io_out_pd_1_isRet; // @[IFU.scala 142:46]
  wire  preDecoders_3_io_out_pd_2_valid; // @[IFU.scala 142:46]
  wire  preDecoders_3_io_out_pd_2_isRVC; // @[IFU.scala 142:46]
  wire [1:0] preDecoders_3_io_out_pd_2_brType; // @[IFU.scala 142:46]
  wire  preDecoders_3_io_out_pd_2_isCall; // @[IFU.scala 142:46]
  wire  preDecoders_3_io_out_pd_2_isRet; // @[IFU.scala 142:46]
  wire  preDecoders_3_io_out_pd_3_valid; // @[IFU.scala 142:46]
  wire  preDecoders_3_io_out_pd_3_isRVC; // @[IFU.scala 142:46]
  wire [1:0] preDecoders_3_io_out_pd_3_brType; // @[IFU.scala 142:46]
  wire  preDecoders_3_io_out_pd_3_isCall; // @[IFU.scala 142:46]
  wire  preDecoders_3_io_out_pd_3_isRet; // @[IFU.scala 142:46]
  wire  preDecoders_3_io_out_pd_4_valid; // @[IFU.scala 142:46]
  wire  preDecoders_3_io_out_pd_4_isRVC; // @[IFU.scala 142:46]
  wire [1:0] preDecoders_3_io_out_pd_4_brType; // @[IFU.scala 142:46]
  wire  preDecoders_3_io_out_pd_4_isCall; // @[IFU.scala 142:46]
  wire  preDecoders_3_io_out_pd_4_isRet; // @[IFU.scala 142:46]
  wire  preDecoders_3_io_out_pd_5_valid; // @[IFU.scala 142:46]
  wire  preDecoders_3_io_out_pd_5_isRVC; // @[IFU.scala 142:46]
  wire [1:0] preDecoders_3_io_out_pd_5_brType; // @[IFU.scala 142:46]
  wire  preDecoders_3_io_out_pd_5_isCall; // @[IFU.scala 142:46]
  wire  preDecoders_3_io_out_pd_5_isRet; // @[IFU.scala 142:46]
  wire  preDecoders_3_io_out_pd_6_valid; // @[IFU.scala 142:46]
  wire  preDecoders_3_io_out_pd_6_isRVC; // @[IFU.scala 142:46]
  wire [1:0] preDecoders_3_io_out_pd_6_brType; // @[IFU.scala 142:46]
  wire  preDecoders_3_io_out_pd_6_isCall; // @[IFU.scala 142:46]
  wire  preDecoders_3_io_out_pd_6_isRet; // @[IFU.scala 142:46]
  wire  preDecoders_3_io_out_pd_7_valid; // @[IFU.scala 142:46]
  wire  preDecoders_3_io_out_pd_7_isRVC; // @[IFU.scala 142:46]
  wire [1:0] preDecoders_3_io_out_pd_7_brType; // @[IFU.scala 142:46]
  wire  preDecoders_3_io_out_pd_7_isCall; // @[IFU.scala 142:46]
  wire  preDecoders_3_io_out_pd_7_isRet; // @[IFU.scala 142:46]
  wire  preDecoders_3_io_out_hasHalfValid_2; // @[IFU.scala 142:46]
  wire  preDecoders_3_io_out_hasHalfValid_3; // @[IFU.scala 142:46]
  wire  preDecoders_3_io_out_hasHalfValid_4; // @[IFU.scala 142:46]
  wire  preDecoders_3_io_out_hasHalfValid_5; // @[IFU.scala 142:46]
  wire  preDecoders_3_io_out_hasHalfValid_6; // @[IFU.scala 142:46]
  wire  preDecoders_3_io_out_hasHalfValid_7; // @[IFU.scala 142:46]
  wire [31:0] preDecoders_3_io_out_instr_0; // @[IFU.scala 142:46]
  wire [31:0] preDecoders_3_io_out_instr_1; // @[IFU.scala 142:46]
  wire [31:0] preDecoders_3_io_out_instr_2; // @[IFU.scala 142:46]
  wire [31:0] preDecoders_3_io_out_instr_3; // @[IFU.scala 142:46]
  wire [31:0] preDecoders_3_io_out_instr_4; // @[IFU.scala 142:46]
  wire [31:0] preDecoders_3_io_out_instr_5; // @[IFU.scala 142:46]
  wire [31:0] preDecoders_3_io_out_instr_6; // @[IFU.scala 142:46]
  wire [31:0] preDecoders_3_io_out_instr_7; // @[IFU.scala 142:46]
  wire [63:0] preDecoders_3_io_out_jumpOffset_0; // @[IFU.scala 142:46]
  wire [63:0] preDecoders_3_io_out_jumpOffset_1; // @[IFU.scala 142:46]
  wire [63:0] preDecoders_3_io_out_jumpOffset_2; // @[IFU.scala 142:46]
  wire [63:0] preDecoders_3_io_out_jumpOffset_3; // @[IFU.scala 142:46]
  wire [63:0] preDecoders_3_io_out_jumpOffset_4; // @[IFU.scala 142:46]
  wire [63:0] preDecoders_3_io_out_jumpOffset_5; // @[IFU.scala 142:46]
  wire [63:0] preDecoders_3_io_out_jumpOffset_6; // @[IFU.scala 142:46]
  wire [63:0] preDecoders_3_io_out_jumpOffset_7; // @[IFU.scala 142:46]
  wire  predChecker_clock; // @[IFU.scala 144:31]
  wire  predChecker_io_in_ftqOffset_valid; // @[IFU.scala 144:31]
  wire [2:0] predChecker_io_in_ftqOffset_bits; // @[IFU.scala 144:31]
  wire [63:0] predChecker_io_in_jumpOffset_0; // @[IFU.scala 144:31]
  wire [63:0] predChecker_io_in_jumpOffset_1; // @[IFU.scala 144:31]
  wire [63:0] predChecker_io_in_jumpOffset_2; // @[IFU.scala 144:31]
  wire [63:0] predChecker_io_in_jumpOffset_3; // @[IFU.scala 144:31]
  wire [63:0] predChecker_io_in_jumpOffset_4; // @[IFU.scala 144:31]
  wire [63:0] predChecker_io_in_jumpOffset_5; // @[IFU.scala 144:31]
  wire [63:0] predChecker_io_in_jumpOffset_6; // @[IFU.scala 144:31]
  wire [63:0] predChecker_io_in_jumpOffset_7; // @[IFU.scala 144:31]
  wire [38:0] predChecker_io_in_target; // @[IFU.scala 144:31]
  wire  predChecker_io_in_instrRange_0; // @[IFU.scala 144:31]
  wire  predChecker_io_in_instrRange_1; // @[IFU.scala 144:31]
  wire  predChecker_io_in_instrRange_2; // @[IFU.scala 144:31]
  wire  predChecker_io_in_instrRange_3; // @[IFU.scala 144:31]
  wire  predChecker_io_in_instrRange_4; // @[IFU.scala 144:31]
  wire  predChecker_io_in_instrRange_5; // @[IFU.scala 144:31]
  wire  predChecker_io_in_instrRange_6; // @[IFU.scala 144:31]
  wire  predChecker_io_in_instrRange_7; // @[IFU.scala 144:31]
  wire  predChecker_io_in_instrValid_0; // @[IFU.scala 144:31]
  wire  predChecker_io_in_instrValid_1; // @[IFU.scala 144:31]
  wire  predChecker_io_in_instrValid_2; // @[IFU.scala 144:31]
  wire  predChecker_io_in_instrValid_3; // @[IFU.scala 144:31]
  wire  predChecker_io_in_instrValid_4; // @[IFU.scala 144:31]
  wire  predChecker_io_in_instrValid_5; // @[IFU.scala 144:31]
  wire  predChecker_io_in_instrValid_6; // @[IFU.scala 144:31]
  wire  predChecker_io_in_instrValid_7; // @[IFU.scala 144:31]
  wire  predChecker_io_in_pds_0_isRVC; // @[IFU.scala 144:31]
  wire [1:0] predChecker_io_in_pds_0_brType; // @[IFU.scala 144:31]
  wire  predChecker_io_in_pds_0_isRet; // @[IFU.scala 144:31]
  wire  predChecker_io_in_pds_1_isRVC; // @[IFU.scala 144:31]
  wire [1:0] predChecker_io_in_pds_1_brType; // @[IFU.scala 144:31]
  wire  predChecker_io_in_pds_1_isRet; // @[IFU.scala 144:31]
  wire  predChecker_io_in_pds_2_isRVC; // @[IFU.scala 144:31]
  wire [1:0] predChecker_io_in_pds_2_brType; // @[IFU.scala 144:31]
  wire  predChecker_io_in_pds_2_isRet; // @[IFU.scala 144:31]
  wire  predChecker_io_in_pds_3_isRVC; // @[IFU.scala 144:31]
  wire [1:0] predChecker_io_in_pds_3_brType; // @[IFU.scala 144:31]
  wire  predChecker_io_in_pds_3_isRet; // @[IFU.scala 144:31]
  wire  predChecker_io_in_pds_4_isRVC; // @[IFU.scala 144:31]
  wire [1:0] predChecker_io_in_pds_4_brType; // @[IFU.scala 144:31]
  wire  predChecker_io_in_pds_4_isRet; // @[IFU.scala 144:31]
  wire  predChecker_io_in_pds_5_isRVC; // @[IFU.scala 144:31]
  wire [1:0] predChecker_io_in_pds_5_brType; // @[IFU.scala 144:31]
  wire  predChecker_io_in_pds_5_isRet; // @[IFU.scala 144:31]
  wire  predChecker_io_in_pds_6_isRVC; // @[IFU.scala 144:31]
  wire [1:0] predChecker_io_in_pds_6_brType; // @[IFU.scala 144:31]
  wire  predChecker_io_in_pds_6_isRet; // @[IFU.scala 144:31]
  wire  predChecker_io_in_pds_7_isRVC; // @[IFU.scala 144:31]
  wire [1:0] predChecker_io_in_pds_7_brType; // @[IFU.scala 144:31]
  wire  predChecker_io_in_pds_7_isRet; // @[IFU.scala 144:31]
  wire [38:0] predChecker_io_in_pc_0; // @[IFU.scala 144:31]
  wire [38:0] predChecker_io_in_pc_1; // @[IFU.scala 144:31]
  wire [38:0] predChecker_io_in_pc_2; // @[IFU.scala 144:31]
  wire [38:0] predChecker_io_in_pc_3; // @[IFU.scala 144:31]
  wire [38:0] predChecker_io_in_pc_4; // @[IFU.scala 144:31]
  wire [38:0] predChecker_io_in_pc_5; // @[IFU.scala 144:31]
  wire [38:0] predChecker_io_in_pc_6; // @[IFU.scala 144:31]
  wire [38:0] predChecker_io_in_pc_7; // @[IFU.scala 144:31]
  wire  predChecker_io_out_stage1Out_fixedRange_0; // @[IFU.scala 144:31]
  wire  predChecker_io_out_stage1Out_fixedRange_1; // @[IFU.scala 144:31]
  wire  predChecker_io_out_stage1Out_fixedRange_2; // @[IFU.scala 144:31]
  wire  predChecker_io_out_stage1Out_fixedRange_3; // @[IFU.scala 144:31]
  wire  predChecker_io_out_stage1Out_fixedRange_4; // @[IFU.scala 144:31]
  wire  predChecker_io_out_stage1Out_fixedRange_5; // @[IFU.scala 144:31]
  wire  predChecker_io_out_stage1Out_fixedRange_6; // @[IFU.scala 144:31]
  wire  predChecker_io_out_stage1Out_fixedRange_7; // @[IFU.scala 144:31]
  wire  predChecker_io_out_stage1Out_fixedTaken_0; // @[IFU.scala 144:31]
  wire  predChecker_io_out_stage1Out_fixedTaken_1; // @[IFU.scala 144:31]
  wire  predChecker_io_out_stage1Out_fixedTaken_2; // @[IFU.scala 144:31]
  wire  predChecker_io_out_stage1Out_fixedTaken_3; // @[IFU.scala 144:31]
  wire  predChecker_io_out_stage1Out_fixedTaken_4; // @[IFU.scala 144:31]
  wire  predChecker_io_out_stage1Out_fixedTaken_5; // @[IFU.scala 144:31]
  wire  predChecker_io_out_stage1Out_fixedTaken_6; // @[IFU.scala 144:31]
  wire  predChecker_io_out_stage1Out_fixedTaken_7; // @[IFU.scala 144:31]
  wire [38:0] predChecker_io_out_stage2Out_fixedTarget_0; // @[IFU.scala 144:31]
  wire [38:0] predChecker_io_out_stage2Out_fixedTarget_1; // @[IFU.scala 144:31]
  wire [38:0] predChecker_io_out_stage2Out_fixedTarget_2; // @[IFU.scala 144:31]
  wire [38:0] predChecker_io_out_stage2Out_fixedTarget_3; // @[IFU.scala 144:31]
  wire [38:0] predChecker_io_out_stage2Out_fixedTarget_4; // @[IFU.scala 144:31]
  wire [38:0] predChecker_io_out_stage2Out_fixedTarget_5; // @[IFU.scala 144:31]
  wire [38:0] predChecker_io_out_stage2Out_fixedTarget_6; // @[IFU.scala 144:31]
  wire [38:0] predChecker_io_out_stage2Out_fixedTarget_7; // @[IFU.scala 144:31]
  wire  predChecker_io_out_stage2Out_fixedMissPred_0; // @[IFU.scala 144:31]
  wire  predChecker_io_out_stage2Out_fixedMissPred_1; // @[IFU.scala 144:31]
  wire  predChecker_io_out_stage2Out_fixedMissPred_2; // @[IFU.scala 144:31]
  wire  predChecker_io_out_stage2Out_fixedMissPred_3; // @[IFU.scala 144:31]
  wire  predChecker_io_out_stage2Out_fixedMissPred_4; // @[IFU.scala 144:31]
  wire  predChecker_io_out_stage2Out_fixedMissPred_5; // @[IFU.scala 144:31]
  wire  predChecker_io_out_stage2Out_fixedMissPred_6; // @[IFU.scala 144:31]
  wire  predChecker_io_out_stage2Out_fixedMissPred_7; // @[IFU.scala 144:31]
  wire [2:0] predChecker_io_out_stage2Out_faultType_0_value; // @[IFU.scala 144:31]
  wire [2:0] predChecker_io_out_stage2Out_faultType_1_value; // @[IFU.scala 144:31]
  wire [2:0] predChecker_io_out_stage2Out_faultType_2_value; // @[IFU.scala 144:31]
  wire [2:0] predChecker_io_out_stage2Out_faultType_3_value; // @[IFU.scala 144:31]
  wire [2:0] predChecker_io_out_stage2Out_faultType_4_value; // @[IFU.scala 144:31]
  wire [2:0] predChecker_io_out_stage2Out_faultType_5_value; // @[IFU.scala 144:31]
  wire [2:0] predChecker_io_out_stage2Out_faultType_6_value; // @[IFU.scala 144:31]
  wire [2:0] predChecker_io_out_stage2Out_faultType_7_value; // @[IFU.scala 144:31]
  wire  frontendTrigger_clock; // @[IFU.scala 145:31]
  wire  frontendTrigger_reset; // @[IFU.scala 145:31]
  wire  frontendTrigger_io_frontendTrigger_t_valid; // @[IFU.scala 145:31]
  wire [1:0] frontendTrigger_io_frontendTrigger_t_bits_addr; // @[IFU.scala 145:31]
  wire [1:0] frontendTrigger_io_frontendTrigger_t_bits_tdata_matchType; // @[IFU.scala 145:31]
  wire  frontendTrigger_io_frontendTrigger_t_bits_tdata_select; // @[IFU.scala 145:31]
  wire  frontendTrigger_io_frontendTrigger_t_bits_tdata_timing; // @[IFU.scala 145:31]
  wire  frontendTrigger_io_frontendTrigger_t_bits_tdata_chain; // @[IFU.scala 145:31]
  wire [63:0] frontendTrigger_io_frontendTrigger_t_bits_tdata_tdata2; // @[IFU.scala 145:31]
  wire  frontendTrigger_io_csrTriggerEnable_0; // @[IFU.scala 145:31]
  wire  frontendTrigger_io_csrTriggerEnable_1; // @[IFU.scala 145:31]
  wire  frontendTrigger_io_csrTriggerEnable_2; // @[IFU.scala 145:31]
  wire  frontendTrigger_io_csrTriggerEnable_3; // @[IFU.scala 145:31]
  wire  frontendTrigger_io_triggered_0_frontendHit_0; // @[IFU.scala 145:31]
  wire  frontendTrigger_io_triggered_0_frontendHit_1; // @[IFU.scala 145:31]
  wire  frontendTrigger_io_triggered_0_frontendHit_2; // @[IFU.scala 145:31]
  wire  frontendTrigger_io_triggered_0_frontendHit_3; // @[IFU.scala 145:31]
  wire  frontendTrigger_io_triggered_0_backendEn_0; // @[IFU.scala 145:31]
  wire  frontendTrigger_io_triggered_0_backendEn_1; // @[IFU.scala 145:31]
  wire  frontendTrigger_io_triggered_1_frontendHit_0; // @[IFU.scala 145:31]
  wire  frontendTrigger_io_triggered_1_frontendHit_1; // @[IFU.scala 145:31]
  wire  frontendTrigger_io_triggered_1_frontendHit_2; // @[IFU.scala 145:31]
  wire  frontendTrigger_io_triggered_1_frontendHit_3; // @[IFU.scala 145:31]
  wire  frontendTrigger_io_triggered_1_backendEn_0; // @[IFU.scala 145:31]
  wire  frontendTrigger_io_triggered_1_backendEn_1; // @[IFU.scala 145:31]
  wire  frontendTrigger_io_triggered_2_frontendHit_0; // @[IFU.scala 145:31]
  wire  frontendTrigger_io_triggered_2_frontendHit_1; // @[IFU.scala 145:31]
  wire  frontendTrigger_io_triggered_2_frontendHit_2; // @[IFU.scala 145:31]
  wire  frontendTrigger_io_triggered_2_frontendHit_3; // @[IFU.scala 145:31]
  wire  frontendTrigger_io_triggered_2_backendEn_0; // @[IFU.scala 145:31]
  wire  frontendTrigger_io_triggered_2_backendEn_1; // @[IFU.scala 145:31]
  wire  frontendTrigger_io_triggered_3_frontendHit_0; // @[IFU.scala 145:31]
  wire  frontendTrigger_io_triggered_3_frontendHit_1; // @[IFU.scala 145:31]
  wire  frontendTrigger_io_triggered_3_frontendHit_2; // @[IFU.scala 145:31]
  wire  frontendTrigger_io_triggered_3_frontendHit_3; // @[IFU.scala 145:31]
  wire  frontendTrigger_io_triggered_3_backendEn_0; // @[IFU.scala 145:31]
  wire  frontendTrigger_io_triggered_3_backendEn_1; // @[IFU.scala 145:31]
  wire  frontendTrigger_io_triggered_4_frontendHit_0; // @[IFU.scala 145:31]
  wire  frontendTrigger_io_triggered_4_frontendHit_1; // @[IFU.scala 145:31]
  wire  frontendTrigger_io_triggered_4_frontendHit_2; // @[IFU.scala 145:31]
  wire  frontendTrigger_io_triggered_4_frontendHit_3; // @[IFU.scala 145:31]
  wire  frontendTrigger_io_triggered_4_backendEn_0; // @[IFU.scala 145:31]
  wire  frontendTrigger_io_triggered_4_backendEn_1; // @[IFU.scala 145:31]
  wire  frontendTrigger_io_triggered_5_frontendHit_0; // @[IFU.scala 145:31]
  wire  frontendTrigger_io_triggered_5_frontendHit_1; // @[IFU.scala 145:31]
  wire  frontendTrigger_io_triggered_5_frontendHit_2; // @[IFU.scala 145:31]
  wire  frontendTrigger_io_triggered_5_frontendHit_3; // @[IFU.scala 145:31]
  wire  frontendTrigger_io_triggered_5_backendEn_0; // @[IFU.scala 145:31]
  wire  frontendTrigger_io_triggered_5_backendEn_1; // @[IFU.scala 145:31]
  wire  frontendTrigger_io_triggered_6_frontendHit_0; // @[IFU.scala 145:31]
  wire  frontendTrigger_io_triggered_6_frontendHit_1; // @[IFU.scala 145:31]
  wire  frontendTrigger_io_triggered_6_frontendHit_2; // @[IFU.scala 145:31]
  wire  frontendTrigger_io_triggered_6_frontendHit_3; // @[IFU.scala 145:31]
  wire  frontendTrigger_io_triggered_6_backendEn_0; // @[IFU.scala 145:31]
  wire  frontendTrigger_io_triggered_6_backendEn_1; // @[IFU.scala 145:31]
  wire  frontendTrigger_io_triggered_7_frontendHit_0; // @[IFU.scala 145:31]
  wire  frontendTrigger_io_triggered_7_frontendHit_1; // @[IFU.scala 145:31]
  wire  frontendTrigger_io_triggered_7_frontendHit_2; // @[IFU.scala 145:31]
  wire  frontendTrigger_io_triggered_7_frontendHit_3; // @[IFU.scala 145:31]
  wire  frontendTrigger_io_triggered_7_backendEn_0; // @[IFU.scala 145:31]
  wire  frontendTrigger_io_triggered_7_backendEn_1; // @[IFU.scala 145:31]
  wire  frontendTrigger_io_pds_0_isRVC; // @[IFU.scala 145:31]
  wire  frontendTrigger_io_pds_1_isRVC; // @[IFU.scala 145:31]
  wire  frontendTrigger_io_pds_2_isRVC; // @[IFU.scala 145:31]
  wire  frontendTrigger_io_pds_3_isRVC; // @[IFU.scala 145:31]
  wire  frontendTrigger_io_pds_4_isRVC; // @[IFU.scala 145:31]
  wire  frontendTrigger_io_pds_5_isRVC; // @[IFU.scala 145:31]
  wire  frontendTrigger_io_pds_6_isRVC; // @[IFU.scala 145:31]
  wire  frontendTrigger_io_pds_7_isRVC; // @[IFU.scala 145:31]
  wire [38:0] frontendTrigger_io_pc_0; // @[IFU.scala 145:31]
  wire [38:0] frontendTrigger_io_pc_1; // @[IFU.scala 145:31]
  wire [38:0] frontendTrigger_io_pc_2; // @[IFU.scala 145:31]
  wire [38:0] frontendTrigger_io_pc_3; // @[IFU.scala 145:31]
  wire [38:0] frontendTrigger_io_pc_4; // @[IFU.scala 145:31]
  wire [38:0] frontendTrigger_io_pc_5; // @[IFU.scala 145:31]
  wire [38:0] frontendTrigger_io_pc_6; // @[IFU.scala 145:31]
  wire [38:0] frontendTrigger_io_pc_7; // @[IFU.scala 145:31]
  wire [15:0] frontendTrigger_io_data_0; // @[IFU.scala 145:31]
  wire [15:0] frontendTrigger_io_data_1; // @[IFU.scala 145:31]
  wire [15:0] frontendTrigger_io_data_2; // @[IFU.scala 145:31]
  wire [15:0] frontendTrigger_io_data_3; // @[IFU.scala 145:31]
  wire [15:0] frontendTrigger_io_data_4; // @[IFU.scala 145:31]
  wire [15:0] frontendTrigger_io_data_5; // @[IFU.scala 145:31]
  wire [15:0] frontendTrigger_io_data_6; // @[IFU.scala 145:31]
  wire [15:0] frontendTrigger_io_data_7; // @[IFU.scala 145:31]
  wire [15:0] frontendTrigger_io_data_8; // @[IFU.scala 145:31]
  wire [31:0] f3_expd_instr_expander_io_in; // @[IFU.scala 382:32]
  wire [31:0] f3_expd_instr_expander_io_out_bits; // @[IFU.scala 382:32]
  wire [31:0] f3_expd_instr_expander_1_io_in; // @[IFU.scala 382:32]
  wire [31:0] f3_expd_instr_expander_1_io_out_bits; // @[IFU.scala 382:32]
  wire [31:0] f3_expd_instr_expander_2_io_in; // @[IFU.scala 382:32]
  wire [31:0] f3_expd_instr_expander_2_io_out_bits; // @[IFU.scala 382:32]
  wire [31:0] f3_expd_instr_expander_3_io_in; // @[IFU.scala 382:32]
  wire [31:0] f3_expd_instr_expander_3_io_out_bits; // @[IFU.scala 382:32]
  wire [31:0] f3_expd_instr_expander_4_io_in; // @[IFU.scala 382:32]
  wire [31:0] f3_expd_instr_expander_4_io_out_bits; // @[IFU.scala 382:32]
  wire [31:0] f3_expd_instr_expander_5_io_in; // @[IFU.scala 382:32]
  wire [31:0] f3_expd_instr_expander_5_io_out_bits; // @[IFU.scala 382:32]
  wire [31:0] f3_expd_instr_expander_6_io_in; // @[IFU.scala 382:32]
  wire [31:0] f3_expd_instr_expander_6_io_out_bits; // @[IFU.scala 382:32]
  wire [31:0] f3_expd_instr_expander_7_io_in; // @[IFU.scala 382:32]
  wire [31:0] f3_expd_instr_expander_7_io_out_bits; // @[IFU.scala 382:32]
  wire  writer_clock; // @[ChiselDB.scala 132:24]
  wire  writer_reset; // @[ChiselDB.scala 132:24]
  wire  writer_en; // @[ChiselDB.scala 132:24]
  wire [63:0] writer_stamp; // @[ChiselDB.scala 132:24]
  wire [38:0] writer_data_start_addr; // @[ChiselDB.scala 132:24]
  wire [31:0] writer_data_instr_count; // @[ChiselDB.scala 132:24]
  wire  writer_data_exception; // @[ChiselDB.scala 132:24]
  wire  writer_data_is_cache_hit; // @[ChiselDB.scala 132:24]
  wire  writer_1_clock; // @[ChiselDB.scala 132:24]
  wire  writer_1_reset; // @[ChiselDB.scala 132:24]
  wire  writer_1_en; // @[ChiselDB.scala 132:24]
  wire [63:0] writer_1_stamp; // @[ChiselDB.scala 132:24]
  wire [38:0] writer_1_data_start_addr; // @[ChiselDB.scala 132:24]
  wire  writer_1_data_is_miss_pred; // @[ChiselDB.scala 132:24]
  wire [31:0] writer_1_data_miss_pred_offset; // @[ChiselDB.scala 132:24]
  wire  writer_1_data_checkJalFault; // @[ChiselDB.scala 132:24]
  wire  writer_1_data_checkRetFault; // @[ChiselDB.scala 132:24]
  wire  writer_1_data_checkTargetFault; // @[ChiselDB.scala 132:24]
  wire  writer_1_data_checkNotCFIFault; // @[ChiselDB.scala 132:24]
  wire  writer_1_data_checkInvalidTaken; // @[ChiselDB.scala 132:24]
  wire  f0_doubleLine = io_ftqInter_fromFtq_req_bits_startAddr[5]; // @[FrontendBundle.scala 39:34]
  wire  f0_fire = io_ftqInter_fromFtq_req_ready & io_ftqInter_fromFtq_req_valid; // @[Decoupled.scala 50:35]
  wire  from_bpu_f0_flush_differentFlag = io_ftqInter_fromFtq_flushFromBpu_s2_bits_flag ^
    io_ftqInter_fromFtq_req_bits_ftqIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  from_bpu_f0_flush_compare = io_ftqInter_fromFtq_flushFromBpu_s2_bits_value >
    io_ftqInter_fromFtq_req_bits_ftqIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _from_bpu_f0_flush_T = from_bpu_f0_flush_differentFlag ^ from_bpu_f0_flush_compare; // @[CircularQueuePtr.scala 88:19]
  wire  _from_bpu_f0_flush_T_2 = io_ftqInter_fromFtq_flushFromBpu_s2_valid & ~_from_bpu_f0_flush_T; // @[NewFtq.scala 186:17]
  wire  from_bpu_f0_flush_differentFlag_1 = io_ftqInter_fromFtq_flushFromBpu_s3_bits_flag ^
    io_ftqInter_fromFtq_req_bits_ftqIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  from_bpu_f0_flush_compare_1 = io_ftqInter_fromFtq_flushFromBpu_s3_bits_value >
    io_ftqInter_fromFtq_req_bits_ftqIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _from_bpu_f0_flush_T_3 = from_bpu_f0_flush_differentFlag_1 ^ from_bpu_f0_flush_compare_1; // @[CircularQueuePtr.scala 88:19]
  wire  _from_bpu_f0_flush_T_5 = io_ftqInter_fromFtq_flushFromBpu_s3_valid & ~_from_bpu_f0_flush_T_3; // @[NewFtq.scala 186:17]
  wire  from_bpu_f0_flush = _from_bpu_f0_flush_T_2 | _from_bpu_f0_flush_T_5; // @[IFU.scala 167:84]
  reg  wb_ftq_req_ftqIdx_flag; // @[IFU.scala 707:34]
  reg [2:0] wb_ftq_req_ftqIdx_value; // @[IFU.scala 707:34]
  wire [3:0] _f3_wb_not_flush_T = {wb_ftq_req_ftqIdx_flag,wb_ftq_req_ftqIdx_value}; // @[CircularQueuePtr.scala 61:50]
  reg  f3_ftq_req_ftqIdx_flag; // @[Reg.scala 16:16]
  reg [2:0] f3_ftq_req_ftqIdx_value; // @[Reg.scala 16:16]
  wire [3:0] _f3_wb_not_flush_T_1 = {f3_ftq_req_ftqIdx_flag,f3_ftq_req_ftqIdx_value}; // @[CircularQueuePtr.scala 61:70]
  wire  _f3_wb_not_flush_T_2 = _f3_wb_not_flush_T == _f3_wb_not_flush_T_1; // @[CircularQueuePtr.scala 61:52]
  reg  f3_valid; // @[IFU.scala 365:34]
  reg  wb_valid; // @[IFU.scala 706:34]
  wire  f3_wb_not_flush = _f3_wb_not_flush_T_2 & f3_valid & wb_valid; // @[IFU.scala 729:74]
  wire  _checkFlushWb_bits_misOffset_valid_T = predChecker_io_out_stage2Out_fixedMissPred_0 |
    predChecker_io_out_stage2Out_fixedMissPred_1; // @[ParallelMux.scala 36:53]
  wire  _checkFlushWb_bits_misOffset_valid_T_2 = predChecker_io_out_stage2Out_fixedMissPred_0 |
    predChecker_io_out_stage2Out_fixedMissPred_1 | (predChecker_io_out_stage2Out_fixedMissPred_2 |
    predChecker_io_out_stage2Out_fixedMissPred_3); // @[ParallelMux.scala 36:53]
  wire  _checkFlushWb_bits_misOffset_valid_T_3 = predChecker_io_out_stage2Out_fixedMissPred_4 |
    predChecker_io_out_stage2Out_fixedMissPred_5; // @[ParallelMux.scala 36:53]
  wire  _checkFlushWb_bits_misOffset_valid_T_6 = predChecker_io_out_stage2Out_fixedMissPred_0 |
    predChecker_io_out_stage2Out_fixedMissPred_1 | (predChecker_io_out_stage2Out_fixedMissPred_2 |
    predChecker_io_out_stage2Out_fixedMissPred_3) | (predChecker_io_out_stage2Out_fixedMissPred_4 |
    predChecker_io_out_stage2Out_fixedMissPred_5 | (predChecker_io_out_stage2Out_fixedMissPred_6 |
    predChecker_io_out_stage2Out_fixedMissPred_7)); // @[ParallelMux.scala 36:53]
  reg  wb_false_lastHalf_REG; // @[IFU.scala 718:34]
  reg [2:0] wb_lastIdx; // @[IFU.scala 717:34]
  wire  wb_false_lastHalf = wb_false_lastHalf_REG & wb_lastIdx != 3'h7; // @[IFU.scala 718:54]
  wire  checkFlushWb_bits_misOffset_valid = _checkFlushWb_bits_misOffset_valid_T_6 | wb_false_lastHalf; // @[IFU.scala 755:91]
  wire  wb_redirect = checkFlushWb_bits_misOffset_valid & wb_valid; // @[IFU.scala 765:52]
  wire  f3_flush = io_ftqInter_fromFtq_redirect_valid | wb_redirect & ~f3_wb_not_flush; // @[IFU.scala 174:32]
  reg  f3_mmio; // @[Reg.scala 16:16]
  wire  f3_req_is_mmio = f3_mmio & f3_valid; // @[IFU.scala 420:36]
  reg [3:0] mmio_state; // @[IFU.scala 418:27]
  wire  _mmio_redirect_T = mmio_state == 4'h9; // @[IFU.scala 692:50]
  wire  _mmio_redirect_T_1 = f3_req_is_mmio & mmio_state == 4'h9; // @[IFU.scala 692:36]
  reg  mmio_redirect_REG; // @[IFU.scala 692:77]
  reg  f3_mmio_use_seq_pc; // @[IFU.scala 445:35]
  wire  mmio_redirect = f3_req_is_mmio & mmio_state == 4'h9 & mmio_redirect_REG & f3_mmio_use_seq_pc; // @[IFU.scala 692:99]
  wire  f2_flush = io_ftqInter_fromFtq_redirect_valid | mmio_redirect | wb_redirect; // @[IFU.scala 175:49]
  reg  f1_ftq_req_ftqIdx_flag; // @[Reg.scala 16:16]
  wire  from_bpu_f1_flush_differentFlag = io_ftqInter_fromFtq_flushFromBpu_s3_bits_flag ^ f1_ftq_req_ftqIdx_flag; // @[CircularQueuePtr.scala 86:35]
  reg [2:0] f1_ftq_req_ftqIdx_value; // @[Reg.scala 16:16]
  wire  from_bpu_f1_flush_compare = io_ftqInter_fromFtq_flushFromBpu_s3_bits_value > f1_ftq_req_ftqIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _from_bpu_f1_flush_T = from_bpu_f1_flush_differentFlag ^ from_bpu_f1_flush_compare; // @[CircularQueuePtr.scala 88:19]
  wire  _from_bpu_f1_flush_T_2 = io_ftqInter_fromFtq_flushFromBpu_s3_valid & ~_from_bpu_f1_flush_T; // @[NewFtq.scala 186:17]
  reg  f1_valid; // @[IFU.scala 202:30]
  wire  from_bpu_f1_flush = _from_bpu_f1_flush_T_2 & f1_valid; // @[IFU.scala 211:84]
  wire  f1_flush = f2_flush | from_bpu_f1_flush; // @[IFU.scala 176:24]
  wire  f0_flush = f1_flush | from_bpu_f0_flush; // @[IFU.scala 177:24]
  reg  f2_valid; // @[IFU.scala 236:30]
  wire  f3_mmio_req_commit = f3_req_is_mmio & mmio_state == 4'ha; // @[IFU.scala 422:43]
  wire  f3_ready = f3_req_is_mmio ? io_toIbuffer_ready & f3_mmio_req_commit | ~f3_valid : io_toIbuffer_ready | ~f3_valid
    ; // @[IFU.scala 453:18]
  reg  f2_icache_all_resp_reg; // @[IFU.scala 246:46]
  reg [38:0] f2_ftq_req_startAddr; // @[Reg.scala 16:16]
  reg [38:0] f2_ftq_req_nextlineStart; // @[Reg.scala 16:16]
  reg  f2_doubleLine; // @[Reg.scala 16:16]
  wire  f2_icache_all_resp_wire = io_icacheInter_resp_0_valid & io_icacheInter_resp_0_bits_vaddr == f2_ftq_req_startAddr
     & (io_icacheInter_resp_1_valid & io_icacheInter_resp_1_bits_vaddr == f2_ftq_req_nextlineStart | ~f2_doubleLine); // @[IFU.scala 245:116]
  wire  icacheRespAllValid = f2_icache_all_resp_reg | f2_icache_all_resp_wire; // @[IFU.scala 248:48]
  wire  f2_fire = f2_valid & f3_ready & icacheRespAllValid; // @[IFU.scala 241:44]
  wire  f2_ready = f2_fire | ~f2_valid; // @[IFU.scala 243:23]
  wire  f1_fire = f1_valid & f2_ready; // @[IFU.scala 207:32]
  wire  f1_ready = f1_fire | ~f1_valid; // @[IFU.scala 209:23]
  reg [38:0] f1_ftq_req_startAddr; // @[Reg.scala 16:16]
  reg [38:0] f1_ftq_req_nextlineStart; // @[Reg.scala 16:16]
  reg [38:0] f1_ftq_req_nextStartAddr; // @[Reg.scala 16:16]
  reg  f1_ftq_req_ftqOffset_valid; // @[Reg.scala 16:16]
  reg [2:0] f1_ftq_req_ftqOffset_bits; // @[Reg.scala 16:16]
  reg  f1_doubleLine; // @[Reg.scala 16:16]
  wire  _GEN_10 = f1_fire ? 1'h0 : f1_valid; // @[IFU.scala 202:30 216:{35,46}]
  wire  _GEN_11 = f0_fire & ~f0_flush | _GEN_10; // @[IFU.scala 215:{35,46}]
  wire [39:0] _f1_pc_T = {{1'd0}, f1_ftq_req_startAddr}; // @[IFU.scala 218:92]
  wire [38:0] f1_pc_0 = _f1_pc_T[38:0]; // @[IFU.scala 218:92]
  wire [38:0] f1_pc_1 = f1_ftq_req_startAddr + 39'h2; // @[IFU.scala 218:92]
  wire [38:0] f1_pc_2 = f1_ftq_req_startAddr + 39'h4; // @[IFU.scala 218:92]
  wire [38:0] f1_pc_3 = f1_ftq_req_startAddr + 39'h6; // @[IFU.scala 218:92]
  wire [38:0] f1_pc_4 = f1_ftq_req_startAddr + 39'h8; // @[IFU.scala 218:92]
  wire [38:0] f1_pc_5 = f1_ftq_req_startAddr + 39'ha; // @[IFU.scala 218:92]
  wire [38:0] f1_pc_6 = f1_ftq_req_startAddr + 39'hc; // @[IFU.scala 218:92]
  wire [38:0] f1_pc_7 = f1_ftq_req_startAddr + 39'he; // @[IFU.scala 218:92]
  wire [38:0] f1_half_snpc_6 = f1_ftq_req_startAddr + 39'h10; // @[IFU.scala 219:92]
  wire [38:0] f1_half_snpc_7 = f1_ftq_req_startAddr + 39'h12; // @[IFU.scala 219:92]
  wire [5:0] _f1_cut_ptr_T_1 = {1'h0,f1_ftq_req_startAddr[5:1]}; // @[Cat.scala 31:58]
  wire [6:0] _f1_cut_ptr_T_2 = {{1'd0}, _f1_cut_ptr_T_1}; // @[IFU.scala 220:150]
  wire [5:0] f1_cut_ptr_0 = _f1_cut_ptr_T_2[5:0]; // @[IFU.scala 220:150]
  wire [5:0] f1_cut_ptr_1 = _f1_cut_ptr_T_1 + 6'h1; // @[IFU.scala 220:150]
  wire [5:0] f1_cut_ptr_2 = _f1_cut_ptr_T_1 + 6'h2; // @[IFU.scala 220:150]
  wire [5:0] f1_cut_ptr_3 = _f1_cut_ptr_T_1 + 6'h3; // @[IFU.scala 220:150]
  wire [5:0] f1_cut_ptr_4 = _f1_cut_ptr_T_1 + 6'h4; // @[IFU.scala 220:150]
  wire [5:0] f1_cut_ptr_5 = _f1_cut_ptr_T_1 + 6'h5; // @[IFU.scala 220:150]
  wire [5:0] f1_cut_ptr_6 = _f1_cut_ptr_T_1 + 6'h6; // @[IFU.scala 220:150]
  wire [5:0] f1_cut_ptr_7 = _f1_cut_ptr_T_1 + 6'h7; // @[IFU.scala 220:150]
  wire [5:0] f1_cut_ptr_8 = _f1_cut_ptr_T_1 + 6'h8; // @[IFU.scala 220:150]
  reg [38:0] f2_ftq_req_nextStartAddr; // @[Reg.scala 16:16]
  reg  f2_ftq_req_ftqIdx_flag; // @[Reg.scala 16:16]
  reg [2:0] f2_ftq_req_ftqIdx_value; // @[Reg.scala 16:16]
  reg  f2_ftq_req_ftqOffset_valid; // @[Reg.scala 16:16]
  reg [2:0] f2_ftq_req_ftqOffset_bits; // @[Reg.scala 16:16]
  wire  _io_icacheStop_T = ~f3_ready; // @[IFU.scala 250:20]
  wire  _GEN_23 = f2_fire & f2_icache_all_resp_reg ? 1'h0 : f2_icache_all_resp_reg; // @[IFU.scala 246:46 254:{63,87}]
  wire  _GEN_24 = f2_valid & f2_icache_all_resp_wire & _io_icacheStop_T | _GEN_23; // @[IFU.scala 253:{63,87}]
  wire  _GEN_26 = f2_fire ? 1'h0 : f2_valid; // @[IFU.scala 236:30 258:{35,45}]
  wire  _GEN_27 = f1_fire & ~f1_flush | _GEN_26; // @[IFU.scala 257:{35,45}]
  wire  _f2_mmio_T_2 = ~io_icacheInter_resp_0_bits_tlbExcp_pageFault; // @[IFU.scala 269:60]
  wire  f2_mmio = io_icacheInter_resp_0_bits_tlbExcp_mmio & ~io_icacheInter_resp_0_bits_tlbExcp_accessFault &
    _f2_mmio_T_2; // @[IFU.scala 268:100]
  reg [38:0] f2_pc_0; // @[Reg.scala 16:16]
  reg [38:0] f2_pc_1; // @[Reg.scala 16:16]
  reg [38:0] f2_pc_2; // @[Reg.scala 16:16]
  reg [38:0] f2_pc_3; // @[Reg.scala 16:16]
  reg [38:0] f2_pc_4; // @[Reg.scala 16:16]
  reg [38:0] f2_pc_5; // @[Reg.scala 16:16]
  reg [38:0] f2_pc_6; // @[Reg.scala 16:16]
  reg [38:0] f2_pc_7; // @[Reg.scala 16:16]
  reg [38:0] f2_half_snpc_0; // @[Reg.scala 16:16]
  reg [38:0] f2_half_snpc_1; // @[Reg.scala 16:16]
  reg [38:0] f2_half_snpc_2; // @[Reg.scala 16:16]
  reg [38:0] f2_half_snpc_3; // @[Reg.scala 16:16]
  reg [38:0] f2_half_snpc_4; // @[Reg.scala 16:16]
  reg [38:0] f2_half_snpc_5; // @[Reg.scala 16:16]
  reg [38:0] f2_half_snpc_6; // @[Reg.scala 16:16]
  reg [38:0] f2_half_snpc_7; // @[Reg.scala 16:16]
  reg [5:0] f2_cut_ptr_0; // @[Reg.scala 16:16]
  reg [5:0] f2_cut_ptr_1; // @[Reg.scala 16:16]
  reg [5:0] f2_cut_ptr_2; // @[Reg.scala 16:16]
  reg [5:0] f2_cut_ptr_3; // @[Reg.scala 16:16]
  reg [5:0] f2_cut_ptr_4; // @[Reg.scala 16:16]
  reg [5:0] f2_cut_ptr_5; // @[Reg.scala 16:16]
  reg [5:0] f2_cut_ptr_6; // @[Reg.scala 16:16]
  reg [5:0] f2_cut_ptr_7; // @[Reg.scala 16:16]
  reg [5:0] f2_cut_ptr_8; // @[Reg.scala 16:16]
  reg [38:0] f2_resend_vaddr; // @[Reg.scala 16:16]
  wire [39:0] f2_foldpc_value = {2'h0,f2_pc_0[38:1]}; // @[Cat.scala 31:58]
  wire [9:0] _f2_foldpc_T_5 = f2_foldpc_value[9:0] ^ f2_foldpc_value[19:10]; // @[ParallelMux.scala 58:52]
  wire [9:0] _f2_foldpc_T_6 = f2_foldpc_value[29:20] ^ f2_foldpc_value[39:30]; // @[ParallelMux.scala 58:52]
  wire [9:0] f2_foldpc_0 = _f2_foldpc_T_5 ^ _f2_foldpc_T_6; // @[ParallelMux.scala 58:52]
  wire [39:0] f2_foldpc_value_1 = {2'h0,f2_pc_1[38:1]}; // @[Cat.scala 31:58]
  wire [9:0] _f2_foldpc_T_13 = f2_foldpc_value_1[9:0] ^ f2_foldpc_value_1[19:10]; // @[ParallelMux.scala 58:52]
  wire [9:0] _f2_foldpc_T_14 = f2_foldpc_value_1[29:20] ^ f2_foldpc_value_1[39:30]; // @[ParallelMux.scala 58:52]
  wire [9:0] f2_foldpc_1 = _f2_foldpc_T_13 ^ _f2_foldpc_T_14; // @[ParallelMux.scala 58:52]
  wire [39:0] f2_foldpc_value_2 = {2'h0,f2_pc_2[38:1]}; // @[Cat.scala 31:58]
  wire [9:0] _f2_foldpc_T_21 = f2_foldpc_value_2[9:0] ^ f2_foldpc_value_2[19:10]; // @[ParallelMux.scala 58:52]
  wire [9:0] _f2_foldpc_T_22 = f2_foldpc_value_2[29:20] ^ f2_foldpc_value_2[39:30]; // @[ParallelMux.scala 58:52]
  wire [9:0] f2_foldpc_2 = _f2_foldpc_T_21 ^ _f2_foldpc_T_22; // @[ParallelMux.scala 58:52]
  wire [39:0] f2_foldpc_value_3 = {2'h0,f2_pc_3[38:1]}; // @[Cat.scala 31:58]
  wire [9:0] _f2_foldpc_T_29 = f2_foldpc_value_3[9:0] ^ f2_foldpc_value_3[19:10]; // @[ParallelMux.scala 58:52]
  wire [9:0] _f2_foldpc_T_30 = f2_foldpc_value_3[29:20] ^ f2_foldpc_value_3[39:30]; // @[ParallelMux.scala 58:52]
  wire [9:0] f2_foldpc_3 = _f2_foldpc_T_29 ^ _f2_foldpc_T_30; // @[ParallelMux.scala 58:52]
  wire [39:0] f2_foldpc_value_4 = {2'h0,f2_pc_4[38:1]}; // @[Cat.scala 31:58]
  wire [9:0] _f2_foldpc_T_37 = f2_foldpc_value_4[9:0] ^ f2_foldpc_value_4[19:10]; // @[ParallelMux.scala 58:52]
  wire [9:0] _f2_foldpc_T_38 = f2_foldpc_value_4[29:20] ^ f2_foldpc_value_4[39:30]; // @[ParallelMux.scala 58:52]
  wire [9:0] f2_foldpc_4 = _f2_foldpc_T_37 ^ _f2_foldpc_T_38; // @[ParallelMux.scala 58:52]
  wire [39:0] f2_foldpc_value_5 = {2'h0,f2_pc_5[38:1]}; // @[Cat.scala 31:58]
  wire [9:0] _f2_foldpc_T_45 = f2_foldpc_value_5[9:0] ^ f2_foldpc_value_5[19:10]; // @[ParallelMux.scala 58:52]
  wire [9:0] _f2_foldpc_T_46 = f2_foldpc_value_5[29:20] ^ f2_foldpc_value_5[39:30]; // @[ParallelMux.scala 58:52]
  wire [9:0] f2_foldpc_5 = _f2_foldpc_T_45 ^ _f2_foldpc_T_46; // @[ParallelMux.scala 58:52]
  wire [39:0] f2_foldpc_value_6 = {2'h0,f2_pc_6[38:1]}; // @[Cat.scala 31:58]
  wire [9:0] _f2_foldpc_T_53 = f2_foldpc_value_6[9:0] ^ f2_foldpc_value_6[19:10]; // @[ParallelMux.scala 58:52]
  wire [9:0] _f2_foldpc_T_54 = f2_foldpc_value_6[29:20] ^ f2_foldpc_value_6[39:30]; // @[ParallelMux.scala 58:52]
  wire [9:0] f2_foldpc_6 = _f2_foldpc_T_53 ^ _f2_foldpc_T_54; // @[ParallelMux.scala 58:52]
  wire [39:0] f2_foldpc_value_7 = {2'h0,f2_pc_7[38:1]}; // @[Cat.scala 31:58]
  wire [9:0] _f2_foldpc_T_61 = f2_foldpc_value_7[9:0] ^ f2_foldpc_value_7[19:10]; // @[ParallelMux.scala 58:52]
  wire [9:0] _f2_foldpc_T_62 = f2_foldpc_value_7[29:20] ^ f2_foldpc_value_7[39:30]; // @[ParallelMux.scala 58:52]
  wire [9:0] f2_foldpc_7 = _f2_foldpc_T_61 ^ _f2_foldpc_T_62; // @[ParallelMux.scala 58:52]
  wire  _f2_jump_range_T = ~f2_ftq_req_ftqOffset_valid; // @[IFU.scala 286:42]
  wire [7:0] _f2_jump_range_T_2 = _f2_jump_range_T ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [2:0] _f2_jump_range_T_4 = ~f2_ftq_req_ftqOffset_bits; // @[IFU.scala 286:105]
  wire [7:0] _f2_jump_range_T_5 = 8'hff >> _f2_jump_range_T_4; // @[IFU.scala 286:102]
  wire [7:0] f2_jump_range = _f2_jump_range_T_2 | _f2_jump_range_T_5; // @[IFU.scala 286:71]
  wire [7:0] _f2_ftr_range_T_1 = f2_ftq_req_ftqOffset_valid ? 8'hff : 8'h0; // @[Bitwise.scala 74:12]
  wire [38:0] f2_ftr_range_byteOffset = f2_ftq_req_nextStartAddr - f2_ftq_req_startAddr; // @[IFU.scala 42:25]
  wire [38:0] _f2_ftr_range_T_4 = f2_ftr_range_byteOffset - 39'h2; // @[IFU.scala 43:17]
  wire [2:0] _f2_ftr_range_T_6 = ~_f2_ftr_range_T_4[3:1]; // @[IFU.scala 287:105]
  wire [7:0] _f2_ftr_range_T_7 = 8'hff >> _f2_ftr_range_T_6; // @[IFU.scala 287:102]
  wire [7:0] f2_ftr_range = _f2_ftr_range_T_1 | _f2_ftr_range_T_7; // @[IFU.scala 287:71]
  wire [7:0] f2_instr_range = f2_jump_range & f2_ftr_range; // @[IFU.scala 288:38]
  wire  _f2_pf_vec_T_2 = f2_ftq_req_startAddr[6] ^ f2_pc_0[6]; // @[IFU.scala 278:29]
  wire  _f2_pf_vec_T_3 = ~_f2_pf_vec_T_2; // @[IFU.scala 289:60]
  wire  _f2_pf_vec_T_8 = _f2_pf_vec_T_2 & f2_doubleLine; // @[IFU.scala 289:172]
  wire  f2_pf_vec_0 = ~_f2_pf_vec_T_2 & io_icacheInter_resp_0_bits_tlbExcp_pageFault | _f2_pf_vec_T_2 & f2_doubleLine &
    io_icacheInter_resp_1_bits_tlbExcp_pageFault; // @[IFU.scala 289:125]
  wire  _f2_pf_vec_T_13 = f2_ftq_req_startAddr[6] ^ f2_pc_1[6]; // @[IFU.scala 278:29]
  wire  _f2_pf_vec_T_14 = ~_f2_pf_vec_T_13; // @[IFU.scala 289:60]
  wire  _f2_pf_vec_T_19 = _f2_pf_vec_T_13 & f2_doubleLine; // @[IFU.scala 289:172]
  wire  f2_pf_vec_1 = ~_f2_pf_vec_T_13 & io_icacheInter_resp_0_bits_tlbExcp_pageFault | _f2_pf_vec_T_13 & f2_doubleLine
     & io_icacheInter_resp_1_bits_tlbExcp_pageFault; // @[IFU.scala 289:125]
  wire  _f2_pf_vec_T_24 = f2_ftq_req_startAddr[6] ^ f2_pc_2[6]; // @[IFU.scala 278:29]
  wire  _f2_pf_vec_T_25 = ~_f2_pf_vec_T_24; // @[IFU.scala 289:60]
  wire  _f2_pf_vec_T_30 = _f2_pf_vec_T_24 & f2_doubleLine; // @[IFU.scala 289:172]
  wire  f2_pf_vec_2 = ~_f2_pf_vec_T_24 & io_icacheInter_resp_0_bits_tlbExcp_pageFault | _f2_pf_vec_T_24 & f2_doubleLine
     & io_icacheInter_resp_1_bits_tlbExcp_pageFault; // @[IFU.scala 289:125]
  wire  _f2_pf_vec_T_35 = f2_ftq_req_startAddr[6] ^ f2_pc_3[6]; // @[IFU.scala 278:29]
  wire  _f2_pf_vec_T_36 = ~_f2_pf_vec_T_35; // @[IFU.scala 289:60]
  wire  _f2_pf_vec_T_41 = _f2_pf_vec_T_35 & f2_doubleLine; // @[IFU.scala 289:172]
  wire  f2_pf_vec_3 = ~_f2_pf_vec_T_35 & io_icacheInter_resp_0_bits_tlbExcp_pageFault | _f2_pf_vec_T_35 & f2_doubleLine
     & io_icacheInter_resp_1_bits_tlbExcp_pageFault; // @[IFU.scala 289:125]
  wire  _f2_pf_vec_T_46 = f2_ftq_req_startAddr[6] ^ f2_pc_4[6]; // @[IFU.scala 278:29]
  wire  _f2_pf_vec_T_47 = ~_f2_pf_vec_T_46; // @[IFU.scala 289:60]
  wire  _f2_pf_vec_T_52 = _f2_pf_vec_T_46 & f2_doubleLine; // @[IFU.scala 289:172]
  wire  f2_pf_vec_4 = ~_f2_pf_vec_T_46 & io_icacheInter_resp_0_bits_tlbExcp_pageFault | _f2_pf_vec_T_46 & f2_doubleLine
     & io_icacheInter_resp_1_bits_tlbExcp_pageFault; // @[IFU.scala 289:125]
  wire  _f2_pf_vec_T_57 = f2_ftq_req_startAddr[6] ^ f2_pc_5[6]; // @[IFU.scala 278:29]
  wire  _f2_pf_vec_T_58 = ~_f2_pf_vec_T_57; // @[IFU.scala 289:60]
  wire  _f2_pf_vec_T_63 = _f2_pf_vec_T_57 & f2_doubleLine; // @[IFU.scala 289:172]
  wire  f2_pf_vec_5 = ~_f2_pf_vec_T_57 & io_icacheInter_resp_0_bits_tlbExcp_pageFault | _f2_pf_vec_T_57 & f2_doubleLine
     & io_icacheInter_resp_1_bits_tlbExcp_pageFault; // @[IFU.scala 289:125]
  wire  _f2_pf_vec_T_68 = f2_ftq_req_startAddr[6] ^ f2_pc_6[6]; // @[IFU.scala 278:29]
  wire  _f2_pf_vec_T_69 = ~_f2_pf_vec_T_68; // @[IFU.scala 289:60]
  wire  _f2_pf_vec_T_74 = _f2_pf_vec_T_68 & f2_doubleLine; // @[IFU.scala 289:172]
  wire  f2_pf_vec_6 = ~_f2_pf_vec_T_68 & io_icacheInter_resp_0_bits_tlbExcp_pageFault | _f2_pf_vec_T_68 & f2_doubleLine
     & io_icacheInter_resp_1_bits_tlbExcp_pageFault; // @[IFU.scala 289:125]
  wire  _f2_pf_vec_T_79 = f2_ftq_req_startAddr[6] ^ f2_pc_7[6]; // @[IFU.scala 278:29]
  wire  _f2_pf_vec_T_80 = ~_f2_pf_vec_T_79; // @[IFU.scala 289:60]
  wire  _f2_pf_vec_T_85 = _f2_pf_vec_T_79 & f2_doubleLine; // @[IFU.scala 289:172]
  wire  f2_pf_vec_7 = ~_f2_pf_vec_T_79 & io_icacheInter_resp_0_bits_tlbExcp_pageFault | _f2_pf_vec_T_79 & f2_doubleLine
     & io_icacheInter_resp_1_bits_tlbExcp_pageFault; // @[IFU.scala 289:125]
  wire  f2_af_vec_0 = _f2_pf_vec_T_3 & io_icacheInter_resp_0_bits_tlbExcp_accessFault | _f2_pf_vec_T_8 &
    io_icacheInter_resp_1_bits_tlbExcp_accessFault; // @[IFU.scala 290:125]
  wire  f2_af_vec_1 = _f2_pf_vec_T_14 & io_icacheInter_resp_0_bits_tlbExcp_accessFault | _f2_pf_vec_T_19 &
    io_icacheInter_resp_1_bits_tlbExcp_accessFault; // @[IFU.scala 290:125]
  wire  f2_af_vec_2 = _f2_pf_vec_T_25 & io_icacheInter_resp_0_bits_tlbExcp_accessFault | _f2_pf_vec_T_30 &
    io_icacheInter_resp_1_bits_tlbExcp_accessFault; // @[IFU.scala 290:125]
  wire  f2_af_vec_3 = _f2_pf_vec_T_36 & io_icacheInter_resp_0_bits_tlbExcp_accessFault | _f2_pf_vec_T_41 &
    io_icacheInter_resp_1_bits_tlbExcp_accessFault; // @[IFU.scala 290:125]
  wire  f2_af_vec_4 = _f2_pf_vec_T_47 & io_icacheInter_resp_0_bits_tlbExcp_accessFault | _f2_pf_vec_T_52 &
    io_icacheInter_resp_1_bits_tlbExcp_accessFault; // @[IFU.scala 290:125]
  wire  f2_af_vec_5 = _f2_pf_vec_T_58 & io_icacheInter_resp_0_bits_tlbExcp_accessFault | _f2_pf_vec_T_63 &
    io_icacheInter_resp_1_bits_tlbExcp_accessFault; // @[IFU.scala 290:125]
  wire  f2_af_vec_6 = _f2_pf_vec_T_69 & io_icacheInter_resp_0_bits_tlbExcp_accessFault | _f2_pf_vec_T_74 &
    io_icacheInter_resp_1_bits_tlbExcp_accessFault; // @[IFU.scala 290:125]
  wire  f2_af_vec_7 = _f2_pf_vec_T_80 & io_icacheInter_resp_0_bits_tlbExcp_accessFault | _f2_pf_vec_T_85 &
    io_icacheInter_resp_1_bits_tlbExcp_accessFault; // @[IFU.scala 290:125]
  wire [1023:0] f2_data_2_cacheline_0 = {io_icacheInter_resp_1_bits_registerData,io_icacheInter_resp_0_bits_registerData
    }; // @[Cat.scala 31:58]
  wire [1023:0] f2_data_2_cacheline_1 = {io_icacheInter_resp_1_bits_registerData,io_icacheInter_resp_0_bits_sramData}; // @[Cat.scala 31:58]
  wire [1023:0] f2_data_2_cacheline_2 = {io_icacheInter_resp_1_bits_sramData,io_icacheInter_resp_0_bits_registerData}; // @[Cat.scala 31:58]
  wire [1023:0] f2_data_2_cacheline_3 = {io_icacheInter_resp_1_bits_sramData,io_icacheInter_resp_0_bits_sramData}; // @[Cat.scala 31:58]
  wire [767:0] f2_cut_data_partCacheline = f2_data_2_cacheline_0[767:0]; // @[IFU.scala 298:36]
  wire [15:0] f2_cut_data_dataVec__0 = f2_cut_data_partCacheline[15:0]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec__1 = f2_cut_data_partCacheline[31:16]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec__2 = f2_cut_data_partCacheline[47:32]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec__3 = f2_cut_data_partCacheline[63:48]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec__4 = f2_cut_data_partCacheline[79:64]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec__5 = f2_cut_data_partCacheline[95:80]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec__6 = f2_cut_data_partCacheline[111:96]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec__7 = f2_cut_data_partCacheline[127:112]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec__8 = f2_cut_data_partCacheline[143:128]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec__9 = f2_cut_data_partCacheline[159:144]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec__10 = f2_cut_data_partCacheline[175:160]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec__11 = f2_cut_data_partCacheline[191:176]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec__12 = f2_cut_data_partCacheline[207:192]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec__13 = f2_cut_data_partCacheline[223:208]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec__14 = f2_cut_data_partCacheline[239:224]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec__15 = f2_cut_data_partCacheline[255:240]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec__16 = f2_cut_data_partCacheline[271:256]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec__17 = f2_cut_data_partCacheline[287:272]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec__18 = f2_cut_data_partCacheline[303:288]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec__19 = f2_cut_data_partCacheline[319:304]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec__20 = f2_cut_data_partCacheline[335:320]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec__21 = f2_cut_data_partCacheline[351:336]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec__22 = f2_cut_data_partCacheline[367:352]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec__23 = f2_cut_data_partCacheline[383:368]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec__24 = f2_cut_data_partCacheline[399:384]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec__25 = f2_cut_data_partCacheline[415:400]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec__26 = f2_cut_data_partCacheline[431:416]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec__27 = f2_cut_data_partCacheline[447:432]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec__28 = f2_cut_data_partCacheline[463:448]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec__29 = f2_cut_data_partCacheline[479:464]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec__30 = f2_cut_data_partCacheline[495:480]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec__31 = f2_cut_data_partCacheline[511:496]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec__32 = f2_cut_data_partCacheline[527:512]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec__33 = f2_cut_data_partCacheline[543:528]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec__34 = f2_cut_data_partCacheline[559:544]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec__35 = f2_cut_data_partCacheline[575:560]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec__36 = f2_cut_data_partCacheline[591:576]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec__37 = f2_cut_data_partCacheline[607:592]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec__38 = f2_cut_data_partCacheline[623:608]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec__39 = f2_cut_data_partCacheline[639:624]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec__40 = f2_cut_data_partCacheline[655:640]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec__41 = f2_cut_data_partCacheline[671:656]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec__42 = f2_cut_data_partCacheline[687:672]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec__43 = f2_cut_data_partCacheline[703:688]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec__44 = f2_cut_data_partCacheline[719:704]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec__45 = f2_cut_data_partCacheline[735:720]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec__46 = f2_cut_data_partCacheline[751:736]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec__47 = f2_cut_data_partCacheline[767:752]; // @[IFU.scala 300:40]
  wire [15:0] _GEN_56 = 6'h1 == f2_cut_ptr_0 ? f2_cut_data_dataVec__1 : f2_cut_data_dataVec__0; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_57 = 6'h2 == f2_cut_ptr_0 ? f2_cut_data_dataVec__2 : _GEN_56; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_58 = 6'h3 == f2_cut_ptr_0 ? f2_cut_data_dataVec__3 : _GEN_57; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_59 = 6'h4 == f2_cut_ptr_0 ? f2_cut_data_dataVec__4 : _GEN_58; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_60 = 6'h5 == f2_cut_ptr_0 ? f2_cut_data_dataVec__5 : _GEN_59; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_61 = 6'h6 == f2_cut_ptr_0 ? f2_cut_data_dataVec__6 : _GEN_60; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_62 = 6'h7 == f2_cut_ptr_0 ? f2_cut_data_dataVec__7 : _GEN_61; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_63 = 6'h8 == f2_cut_ptr_0 ? f2_cut_data_dataVec__8 : _GEN_62; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_64 = 6'h9 == f2_cut_ptr_0 ? f2_cut_data_dataVec__9 : _GEN_63; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_65 = 6'ha == f2_cut_ptr_0 ? f2_cut_data_dataVec__10 : _GEN_64; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_66 = 6'hb == f2_cut_ptr_0 ? f2_cut_data_dataVec__11 : _GEN_65; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_67 = 6'hc == f2_cut_ptr_0 ? f2_cut_data_dataVec__12 : _GEN_66; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_68 = 6'hd == f2_cut_ptr_0 ? f2_cut_data_dataVec__13 : _GEN_67; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_69 = 6'he == f2_cut_ptr_0 ? f2_cut_data_dataVec__14 : _GEN_68; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_70 = 6'hf == f2_cut_ptr_0 ? f2_cut_data_dataVec__15 : _GEN_69; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_71 = 6'h10 == f2_cut_ptr_0 ? f2_cut_data_dataVec__16 : _GEN_70; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_72 = 6'h11 == f2_cut_ptr_0 ? f2_cut_data_dataVec__17 : _GEN_71; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_73 = 6'h12 == f2_cut_ptr_0 ? f2_cut_data_dataVec__18 : _GEN_72; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_74 = 6'h13 == f2_cut_ptr_0 ? f2_cut_data_dataVec__19 : _GEN_73; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_75 = 6'h14 == f2_cut_ptr_0 ? f2_cut_data_dataVec__20 : _GEN_74; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_76 = 6'h15 == f2_cut_ptr_0 ? f2_cut_data_dataVec__21 : _GEN_75; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_77 = 6'h16 == f2_cut_ptr_0 ? f2_cut_data_dataVec__22 : _GEN_76; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_78 = 6'h17 == f2_cut_ptr_0 ? f2_cut_data_dataVec__23 : _GEN_77; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_79 = 6'h18 == f2_cut_ptr_0 ? f2_cut_data_dataVec__24 : _GEN_78; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_80 = 6'h19 == f2_cut_ptr_0 ? f2_cut_data_dataVec__25 : _GEN_79; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_81 = 6'h1a == f2_cut_ptr_0 ? f2_cut_data_dataVec__26 : _GEN_80; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_82 = 6'h1b == f2_cut_ptr_0 ? f2_cut_data_dataVec__27 : _GEN_81; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_83 = 6'h1c == f2_cut_ptr_0 ? f2_cut_data_dataVec__28 : _GEN_82; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_84 = 6'h1d == f2_cut_ptr_0 ? f2_cut_data_dataVec__29 : _GEN_83; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_85 = 6'h1e == f2_cut_ptr_0 ? f2_cut_data_dataVec__30 : _GEN_84; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_86 = 6'h1f == f2_cut_ptr_0 ? f2_cut_data_dataVec__31 : _GEN_85; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_87 = 6'h20 == f2_cut_ptr_0 ? f2_cut_data_dataVec__32 : _GEN_86; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_88 = 6'h21 == f2_cut_ptr_0 ? f2_cut_data_dataVec__33 : _GEN_87; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_89 = 6'h22 == f2_cut_ptr_0 ? f2_cut_data_dataVec__34 : _GEN_88; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_90 = 6'h23 == f2_cut_ptr_0 ? f2_cut_data_dataVec__35 : _GEN_89; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_91 = 6'h24 == f2_cut_ptr_0 ? f2_cut_data_dataVec__36 : _GEN_90; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_92 = 6'h25 == f2_cut_ptr_0 ? f2_cut_data_dataVec__37 : _GEN_91; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_93 = 6'h26 == f2_cut_ptr_0 ? f2_cut_data_dataVec__38 : _GEN_92; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_94 = 6'h27 == f2_cut_ptr_0 ? f2_cut_data_dataVec__39 : _GEN_93; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_95 = 6'h28 == f2_cut_ptr_0 ? f2_cut_data_dataVec__40 : _GEN_94; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_96 = 6'h29 == f2_cut_ptr_0 ? f2_cut_data_dataVec__41 : _GEN_95; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_97 = 6'h2a == f2_cut_ptr_0 ? f2_cut_data_dataVec__42 : _GEN_96; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_98 = 6'h2b == f2_cut_ptr_0 ? f2_cut_data_dataVec__43 : _GEN_97; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_99 = 6'h2c == f2_cut_ptr_0 ? f2_cut_data_dataVec__44 : _GEN_98; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_100 = 6'h2d == f2_cut_ptr_0 ? f2_cut_data_dataVec__45 : _GEN_99; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_101 = 6'h2e == f2_cut_ptr_0 ? f2_cut_data_dataVec__46 : _GEN_100; // @[IFU.scala 302:{19,19}]
  wire [15:0] f2_cut_data_result__0 = 6'h2f == f2_cut_ptr_0 ? f2_cut_data_dataVec__47 : _GEN_101; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_104 = 6'h1 == f2_cut_ptr_1 ? f2_cut_data_dataVec__1 : f2_cut_data_dataVec__0; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_105 = 6'h2 == f2_cut_ptr_1 ? f2_cut_data_dataVec__2 : _GEN_104; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_106 = 6'h3 == f2_cut_ptr_1 ? f2_cut_data_dataVec__3 : _GEN_105; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_107 = 6'h4 == f2_cut_ptr_1 ? f2_cut_data_dataVec__4 : _GEN_106; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_108 = 6'h5 == f2_cut_ptr_1 ? f2_cut_data_dataVec__5 : _GEN_107; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_109 = 6'h6 == f2_cut_ptr_1 ? f2_cut_data_dataVec__6 : _GEN_108; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_110 = 6'h7 == f2_cut_ptr_1 ? f2_cut_data_dataVec__7 : _GEN_109; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_111 = 6'h8 == f2_cut_ptr_1 ? f2_cut_data_dataVec__8 : _GEN_110; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_112 = 6'h9 == f2_cut_ptr_1 ? f2_cut_data_dataVec__9 : _GEN_111; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_113 = 6'ha == f2_cut_ptr_1 ? f2_cut_data_dataVec__10 : _GEN_112; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_114 = 6'hb == f2_cut_ptr_1 ? f2_cut_data_dataVec__11 : _GEN_113; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_115 = 6'hc == f2_cut_ptr_1 ? f2_cut_data_dataVec__12 : _GEN_114; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_116 = 6'hd == f2_cut_ptr_1 ? f2_cut_data_dataVec__13 : _GEN_115; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_117 = 6'he == f2_cut_ptr_1 ? f2_cut_data_dataVec__14 : _GEN_116; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_118 = 6'hf == f2_cut_ptr_1 ? f2_cut_data_dataVec__15 : _GEN_117; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_119 = 6'h10 == f2_cut_ptr_1 ? f2_cut_data_dataVec__16 : _GEN_118; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_120 = 6'h11 == f2_cut_ptr_1 ? f2_cut_data_dataVec__17 : _GEN_119; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_121 = 6'h12 == f2_cut_ptr_1 ? f2_cut_data_dataVec__18 : _GEN_120; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_122 = 6'h13 == f2_cut_ptr_1 ? f2_cut_data_dataVec__19 : _GEN_121; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_123 = 6'h14 == f2_cut_ptr_1 ? f2_cut_data_dataVec__20 : _GEN_122; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_124 = 6'h15 == f2_cut_ptr_1 ? f2_cut_data_dataVec__21 : _GEN_123; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_125 = 6'h16 == f2_cut_ptr_1 ? f2_cut_data_dataVec__22 : _GEN_124; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_126 = 6'h17 == f2_cut_ptr_1 ? f2_cut_data_dataVec__23 : _GEN_125; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_127 = 6'h18 == f2_cut_ptr_1 ? f2_cut_data_dataVec__24 : _GEN_126; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_128 = 6'h19 == f2_cut_ptr_1 ? f2_cut_data_dataVec__25 : _GEN_127; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_129 = 6'h1a == f2_cut_ptr_1 ? f2_cut_data_dataVec__26 : _GEN_128; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_130 = 6'h1b == f2_cut_ptr_1 ? f2_cut_data_dataVec__27 : _GEN_129; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_131 = 6'h1c == f2_cut_ptr_1 ? f2_cut_data_dataVec__28 : _GEN_130; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_132 = 6'h1d == f2_cut_ptr_1 ? f2_cut_data_dataVec__29 : _GEN_131; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_133 = 6'h1e == f2_cut_ptr_1 ? f2_cut_data_dataVec__30 : _GEN_132; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_134 = 6'h1f == f2_cut_ptr_1 ? f2_cut_data_dataVec__31 : _GEN_133; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_135 = 6'h20 == f2_cut_ptr_1 ? f2_cut_data_dataVec__32 : _GEN_134; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_136 = 6'h21 == f2_cut_ptr_1 ? f2_cut_data_dataVec__33 : _GEN_135; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_137 = 6'h22 == f2_cut_ptr_1 ? f2_cut_data_dataVec__34 : _GEN_136; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_138 = 6'h23 == f2_cut_ptr_1 ? f2_cut_data_dataVec__35 : _GEN_137; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_139 = 6'h24 == f2_cut_ptr_1 ? f2_cut_data_dataVec__36 : _GEN_138; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_140 = 6'h25 == f2_cut_ptr_1 ? f2_cut_data_dataVec__37 : _GEN_139; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_141 = 6'h26 == f2_cut_ptr_1 ? f2_cut_data_dataVec__38 : _GEN_140; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_142 = 6'h27 == f2_cut_ptr_1 ? f2_cut_data_dataVec__39 : _GEN_141; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_143 = 6'h28 == f2_cut_ptr_1 ? f2_cut_data_dataVec__40 : _GEN_142; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_144 = 6'h29 == f2_cut_ptr_1 ? f2_cut_data_dataVec__41 : _GEN_143; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_145 = 6'h2a == f2_cut_ptr_1 ? f2_cut_data_dataVec__42 : _GEN_144; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_146 = 6'h2b == f2_cut_ptr_1 ? f2_cut_data_dataVec__43 : _GEN_145; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_147 = 6'h2c == f2_cut_ptr_1 ? f2_cut_data_dataVec__44 : _GEN_146; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_148 = 6'h2d == f2_cut_ptr_1 ? f2_cut_data_dataVec__45 : _GEN_147; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_149 = 6'h2e == f2_cut_ptr_1 ? f2_cut_data_dataVec__46 : _GEN_148; // @[IFU.scala 302:{19,19}]
  wire [15:0] f2_cut_data_result__1 = 6'h2f == f2_cut_ptr_1 ? f2_cut_data_dataVec__47 : _GEN_149; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_152 = 6'h1 == f2_cut_ptr_2 ? f2_cut_data_dataVec__1 : f2_cut_data_dataVec__0; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_153 = 6'h2 == f2_cut_ptr_2 ? f2_cut_data_dataVec__2 : _GEN_152; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_154 = 6'h3 == f2_cut_ptr_2 ? f2_cut_data_dataVec__3 : _GEN_153; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_155 = 6'h4 == f2_cut_ptr_2 ? f2_cut_data_dataVec__4 : _GEN_154; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_156 = 6'h5 == f2_cut_ptr_2 ? f2_cut_data_dataVec__5 : _GEN_155; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_157 = 6'h6 == f2_cut_ptr_2 ? f2_cut_data_dataVec__6 : _GEN_156; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_158 = 6'h7 == f2_cut_ptr_2 ? f2_cut_data_dataVec__7 : _GEN_157; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_159 = 6'h8 == f2_cut_ptr_2 ? f2_cut_data_dataVec__8 : _GEN_158; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_160 = 6'h9 == f2_cut_ptr_2 ? f2_cut_data_dataVec__9 : _GEN_159; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_161 = 6'ha == f2_cut_ptr_2 ? f2_cut_data_dataVec__10 : _GEN_160; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_162 = 6'hb == f2_cut_ptr_2 ? f2_cut_data_dataVec__11 : _GEN_161; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_163 = 6'hc == f2_cut_ptr_2 ? f2_cut_data_dataVec__12 : _GEN_162; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_164 = 6'hd == f2_cut_ptr_2 ? f2_cut_data_dataVec__13 : _GEN_163; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_165 = 6'he == f2_cut_ptr_2 ? f2_cut_data_dataVec__14 : _GEN_164; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_166 = 6'hf == f2_cut_ptr_2 ? f2_cut_data_dataVec__15 : _GEN_165; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_167 = 6'h10 == f2_cut_ptr_2 ? f2_cut_data_dataVec__16 : _GEN_166; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_168 = 6'h11 == f2_cut_ptr_2 ? f2_cut_data_dataVec__17 : _GEN_167; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_169 = 6'h12 == f2_cut_ptr_2 ? f2_cut_data_dataVec__18 : _GEN_168; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_170 = 6'h13 == f2_cut_ptr_2 ? f2_cut_data_dataVec__19 : _GEN_169; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_171 = 6'h14 == f2_cut_ptr_2 ? f2_cut_data_dataVec__20 : _GEN_170; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_172 = 6'h15 == f2_cut_ptr_2 ? f2_cut_data_dataVec__21 : _GEN_171; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_173 = 6'h16 == f2_cut_ptr_2 ? f2_cut_data_dataVec__22 : _GEN_172; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_174 = 6'h17 == f2_cut_ptr_2 ? f2_cut_data_dataVec__23 : _GEN_173; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_175 = 6'h18 == f2_cut_ptr_2 ? f2_cut_data_dataVec__24 : _GEN_174; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_176 = 6'h19 == f2_cut_ptr_2 ? f2_cut_data_dataVec__25 : _GEN_175; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_177 = 6'h1a == f2_cut_ptr_2 ? f2_cut_data_dataVec__26 : _GEN_176; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_178 = 6'h1b == f2_cut_ptr_2 ? f2_cut_data_dataVec__27 : _GEN_177; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_179 = 6'h1c == f2_cut_ptr_2 ? f2_cut_data_dataVec__28 : _GEN_178; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_180 = 6'h1d == f2_cut_ptr_2 ? f2_cut_data_dataVec__29 : _GEN_179; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_181 = 6'h1e == f2_cut_ptr_2 ? f2_cut_data_dataVec__30 : _GEN_180; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_182 = 6'h1f == f2_cut_ptr_2 ? f2_cut_data_dataVec__31 : _GEN_181; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_183 = 6'h20 == f2_cut_ptr_2 ? f2_cut_data_dataVec__32 : _GEN_182; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_184 = 6'h21 == f2_cut_ptr_2 ? f2_cut_data_dataVec__33 : _GEN_183; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_185 = 6'h22 == f2_cut_ptr_2 ? f2_cut_data_dataVec__34 : _GEN_184; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_186 = 6'h23 == f2_cut_ptr_2 ? f2_cut_data_dataVec__35 : _GEN_185; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_187 = 6'h24 == f2_cut_ptr_2 ? f2_cut_data_dataVec__36 : _GEN_186; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_188 = 6'h25 == f2_cut_ptr_2 ? f2_cut_data_dataVec__37 : _GEN_187; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_189 = 6'h26 == f2_cut_ptr_2 ? f2_cut_data_dataVec__38 : _GEN_188; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_190 = 6'h27 == f2_cut_ptr_2 ? f2_cut_data_dataVec__39 : _GEN_189; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_191 = 6'h28 == f2_cut_ptr_2 ? f2_cut_data_dataVec__40 : _GEN_190; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_192 = 6'h29 == f2_cut_ptr_2 ? f2_cut_data_dataVec__41 : _GEN_191; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_193 = 6'h2a == f2_cut_ptr_2 ? f2_cut_data_dataVec__42 : _GEN_192; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_194 = 6'h2b == f2_cut_ptr_2 ? f2_cut_data_dataVec__43 : _GEN_193; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_195 = 6'h2c == f2_cut_ptr_2 ? f2_cut_data_dataVec__44 : _GEN_194; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_196 = 6'h2d == f2_cut_ptr_2 ? f2_cut_data_dataVec__45 : _GEN_195; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_197 = 6'h2e == f2_cut_ptr_2 ? f2_cut_data_dataVec__46 : _GEN_196; // @[IFU.scala 302:{19,19}]
  wire [15:0] f2_cut_data_result__2 = 6'h2f == f2_cut_ptr_2 ? f2_cut_data_dataVec__47 : _GEN_197; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_200 = 6'h1 == f2_cut_ptr_3 ? f2_cut_data_dataVec__1 : f2_cut_data_dataVec__0; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_201 = 6'h2 == f2_cut_ptr_3 ? f2_cut_data_dataVec__2 : _GEN_200; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_202 = 6'h3 == f2_cut_ptr_3 ? f2_cut_data_dataVec__3 : _GEN_201; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_203 = 6'h4 == f2_cut_ptr_3 ? f2_cut_data_dataVec__4 : _GEN_202; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_204 = 6'h5 == f2_cut_ptr_3 ? f2_cut_data_dataVec__5 : _GEN_203; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_205 = 6'h6 == f2_cut_ptr_3 ? f2_cut_data_dataVec__6 : _GEN_204; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_206 = 6'h7 == f2_cut_ptr_3 ? f2_cut_data_dataVec__7 : _GEN_205; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_207 = 6'h8 == f2_cut_ptr_3 ? f2_cut_data_dataVec__8 : _GEN_206; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_208 = 6'h9 == f2_cut_ptr_3 ? f2_cut_data_dataVec__9 : _GEN_207; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_209 = 6'ha == f2_cut_ptr_3 ? f2_cut_data_dataVec__10 : _GEN_208; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_210 = 6'hb == f2_cut_ptr_3 ? f2_cut_data_dataVec__11 : _GEN_209; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_211 = 6'hc == f2_cut_ptr_3 ? f2_cut_data_dataVec__12 : _GEN_210; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_212 = 6'hd == f2_cut_ptr_3 ? f2_cut_data_dataVec__13 : _GEN_211; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_213 = 6'he == f2_cut_ptr_3 ? f2_cut_data_dataVec__14 : _GEN_212; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_214 = 6'hf == f2_cut_ptr_3 ? f2_cut_data_dataVec__15 : _GEN_213; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_215 = 6'h10 == f2_cut_ptr_3 ? f2_cut_data_dataVec__16 : _GEN_214; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_216 = 6'h11 == f2_cut_ptr_3 ? f2_cut_data_dataVec__17 : _GEN_215; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_217 = 6'h12 == f2_cut_ptr_3 ? f2_cut_data_dataVec__18 : _GEN_216; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_218 = 6'h13 == f2_cut_ptr_3 ? f2_cut_data_dataVec__19 : _GEN_217; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_219 = 6'h14 == f2_cut_ptr_3 ? f2_cut_data_dataVec__20 : _GEN_218; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_220 = 6'h15 == f2_cut_ptr_3 ? f2_cut_data_dataVec__21 : _GEN_219; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_221 = 6'h16 == f2_cut_ptr_3 ? f2_cut_data_dataVec__22 : _GEN_220; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_222 = 6'h17 == f2_cut_ptr_3 ? f2_cut_data_dataVec__23 : _GEN_221; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_223 = 6'h18 == f2_cut_ptr_3 ? f2_cut_data_dataVec__24 : _GEN_222; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_224 = 6'h19 == f2_cut_ptr_3 ? f2_cut_data_dataVec__25 : _GEN_223; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_225 = 6'h1a == f2_cut_ptr_3 ? f2_cut_data_dataVec__26 : _GEN_224; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_226 = 6'h1b == f2_cut_ptr_3 ? f2_cut_data_dataVec__27 : _GEN_225; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_227 = 6'h1c == f2_cut_ptr_3 ? f2_cut_data_dataVec__28 : _GEN_226; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_228 = 6'h1d == f2_cut_ptr_3 ? f2_cut_data_dataVec__29 : _GEN_227; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_229 = 6'h1e == f2_cut_ptr_3 ? f2_cut_data_dataVec__30 : _GEN_228; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_230 = 6'h1f == f2_cut_ptr_3 ? f2_cut_data_dataVec__31 : _GEN_229; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_231 = 6'h20 == f2_cut_ptr_3 ? f2_cut_data_dataVec__32 : _GEN_230; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_232 = 6'h21 == f2_cut_ptr_3 ? f2_cut_data_dataVec__33 : _GEN_231; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_233 = 6'h22 == f2_cut_ptr_3 ? f2_cut_data_dataVec__34 : _GEN_232; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_234 = 6'h23 == f2_cut_ptr_3 ? f2_cut_data_dataVec__35 : _GEN_233; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_235 = 6'h24 == f2_cut_ptr_3 ? f2_cut_data_dataVec__36 : _GEN_234; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_236 = 6'h25 == f2_cut_ptr_3 ? f2_cut_data_dataVec__37 : _GEN_235; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_237 = 6'h26 == f2_cut_ptr_3 ? f2_cut_data_dataVec__38 : _GEN_236; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_238 = 6'h27 == f2_cut_ptr_3 ? f2_cut_data_dataVec__39 : _GEN_237; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_239 = 6'h28 == f2_cut_ptr_3 ? f2_cut_data_dataVec__40 : _GEN_238; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_240 = 6'h29 == f2_cut_ptr_3 ? f2_cut_data_dataVec__41 : _GEN_239; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_241 = 6'h2a == f2_cut_ptr_3 ? f2_cut_data_dataVec__42 : _GEN_240; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_242 = 6'h2b == f2_cut_ptr_3 ? f2_cut_data_dataVec__43 : _GEN_241; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_243 = 6'h2c == f2_cut_ptr_3 ? f2_cut_data_dataVec__44 : _GEN_242; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_244 = 6'h2d == f2_cut_ptr_3 ? f2_cut_data_dataVec__45 : _GEN_243; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_245 = 6'h2e == f2_cut_ptr_3 ? f2_cut_data_dataVec__46 : _GEN_244; // @[IFU.scala 302:{19,19}]
  wire [15:0] f2_cut_data_result__3 = 6'h2f == f2_cut_ptr_3 ? f2_cut_data_dataVec__47 : _GEN_245; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_248 = 6'h1 == f2_cut_ptr_4 ? f2_cut_data_dataVec__1 : f2_cut_data_dataVec__0; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_249 = 6'h2 == f2_cut_ptr_4 ? f2_cut_data_dataVec__2 : _GEN_248; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_250 = 6'h3 == f2_cut_ptr_4 ? f2_cut_data_dataVec__3 : _GEN_249; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_251 = 6'h4 == f2_cut_ptr_4 ? f2_cut_data_dataVec__4 : _GEN_250; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_252 = 6'h5 == f2_cut_ptr_4 ? f2_cut_data_dataVec__5 : _GEN_251; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_253 = 6'h6 == f2_cut_ptr_4 ? f2_cut_data_dataVec__6 : _GEN_252; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_254 = 6'h7 == f2_cut_ptr_4 ? f2_cut_data_dataVec__7 : _GEN_253; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_255 = 6'h8 == f2_cut_ptr_4 ? f2_cut_data_dataVec__8 : _GEN_254; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_256 = 6'h9 == f2_cut_ptr_4 ? f2_cut_data_dataVec__9 : _GEN_255; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_257 = 6'ha == f2_cut_ptr_4 ? f2_cut_data_dataVec__10 : _GEN_256; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_258 = 6'hb == f2_cut_ptr_4 ? f2_cut_data_dataVec__11 : _GEN_257; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_259 = 6'hc == f2_cut_ptr_4 ? f2_cut_data_dataVec__12 : _GEN_258; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_260 = 6'hd == f2_cut_ptr_4 ? f2_cut_data_dataVec__13 : _GEN_259; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_261 = 6'he == f2_cut_ptr_4 ? f2_cut_data_dataVec__14 : _GEN_260; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_262 = 6'hf == f2_cut_ptr_4 ? f2_cut_data_dataVec__15 : _GEN_261; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_263 = 6'h10 == f2_cut_ptr_4 ? f2_cut_data_dataVec__16 : _GEN_262; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_264 = 6'h11 == f2_cut_ptr_4 ? f2_cut_data_dataVec__17 : _GEN_263; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_265 = 6'h12 == f2_cut_ptr_4 ? f2_cut_data_dataVec__18 : _GEN_264; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_266 = 6'h13 == f2_cut_ptr_4 ? f2_cut_data_dataVec__19 : _GEN_265; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_267 = 6'h14 == f2_cut_ptr_4 ? f2_cut_data_dataVec__20 : _GEN_266; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_268 = 6'h15 == f2_cut_ptr_4 ? f2_cut_data_dataVec__21 : _GEN_267; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_269 = 6'h16 == f2_cut_ptr_4 ? f2_cut_data_dataVec__22 : _GEN_268; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_270 = 6'h17 == f2_cut_ptr_4 ? f2_cut_data_dataVec__23 : _GEN_269; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_271 = 6'h18 == f2_cut_ptr_4 ? f2_cut_data_dataVec__24 : _GEN_270; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_272 = 6'h19 == f2_cut_ptr_4 ? f2_cut_data_dataVec__25 : _GEN_271; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_273 = 6'h1a == f2_cut_ptr_4 ? f2_cut_data_dataVec__26 : _GEN_272; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_274 = 6'h1b == f2_cut_ptr_4 ? f2_cut_data_dataVec__27 : _GEN_273; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_275 = 6'h1c == f2_cut_ptr_4 ? f2_cut_data_dataVec__28 : _GEN_274; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_276 = 6'h1d == f2_cut_ptr_4 ? f2_cut_data_dataVec__29 : _GEN_275; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_277 = 6'h1e == f2_cut_ptr_4 ? f2_cut_data_dataVec__30 : _GEN_276; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_278 = 6'h1f == f2_cut_ptr_4 ? f2_cut_data_dataVec__31 : _GEN_277; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_279 = 6'h20 == f2_cut_ptr_4 ? f2_cut_data_dataVec__32 : _GEN_278; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_280 = 6'h21 == f2_cut_ptr_4 ? f2_cut_data_dataVec__33 : _GEN_279; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_281 = 6'h22 == f2_cut_ptr_4 ? f2_cut_data_dataVec__34 : _GEN_280; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_282 = 6'h23 == f2_cut_ptr_4 ? f2_cut_data_dataVec__35 : _GEN_281; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_283 = 6'h24 == f2_cut_ptr_4 ? f2_cut_data_dataVec__36 : _GEN_282; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_284 = 6'h25 == f2_cut_ptr_4 ? f2_cut_data_dataVec__37 : _GEN_283; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_285 = 6'h26 == f2_cut_ptr_4 ? f2_cut_data_dataVec__38 : _GEN_284; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_286 = 6'h27 == f2_cut_ptr_4 ? f2_cut_data_dataVec__39 : _GEN_285; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_287 = 6'h28 == f2_cut_ptr_4 ? f2_cut_data_dataVec__40 : _GEN_286; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_288 = 6'h29 == f2_cut_ptr_4 ? f2_cut_data_dataVec__41 : _GEN_287; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_289 = 6'h2a == f2_cut_ptr_4 ? f2_cut_data_dataVec__42 : _GEN_288; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_290 = 6'h2b == f2_cut_ptr_4 ? f2_cut_data_dataVec__43 : _GEN_289; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_291 = 6'h2c == f2_cut_ptr_4 ? f2_cut_data_dataVec__44 : _GEN_290; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_292 = 6'h2d == f2_cut_ptr_4 ? f2_cut_data_dataVec__45 : _GEN_291; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_293 = 6'h2e == f2_cut_ptr_4 ? f2_cut_data_dataVec__46 : _GEN_292; // @[IFU.scala 302:{19,19}]
  wire [15:0] f2_cut_data_result__4 = 6'h2f == f2_cut_ptr_4 ? f2_cut_data_dataVec__47 : _GEN_293; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_296 = 6'h1 == f2_cut_ptr_5 ? f2_cut_data_dataVec__1 : f2_cut_data_dataVec__0; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_297 = 6'h2 == f2_cut_ptr_5 ? f2_cut_data_dataVec__2 : _GEN_296; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_298 = 6'h3 == f2_cut_ptr_5 ? f2_cut_data_dataVec__3 : _GEN_297; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_299 = 6'h4 == f2_cut_ptr_5 ? f2_cut_data_dataVec__4 : _GEN_298; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_300 = 6'h5 == f2_cut_ptr_5 ? f2_cut_data_dataVec__5 : _GEN_299; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_301 = 6'h6 == f2_cut_ptr_5 ? f2_cut_data_dataVec__6 : _GEN_300; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_302 = 6'h7 == f2_cut_ptr_5 ? f2_cut_data_dataVec__7 : _GEN_301; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_303 = 6'h8 == f2_cut_ptr_5 ? f2_cut_data_dataVec__8 : _GEN_302; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_304 = 6'h9 == f2_cut_ptr_5 ? f2_cut_data_dataVec__9 : _GEN_303; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_305 = 6'ha == f2_cut_ptr_5 ? f2_cut_data_dataVec__10 : _GEN_304; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_306 = 6'hb == f2_cut_ptr_5 ? f2_cut_data_dataVec__11 : _GEN_305; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_307 = 6'hc == f2_cut_ptr_5 ? f2_cut_data_dataVec__12 : _GEN_306; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_308 = 6'hd == f2_cut_ptr_5 ? f2_cut_data_dataVec__13 : _GEN_307; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_309 = 6'he == f2_cut_ptr_5 ? f2_cut_data_dataVec__14 : _GEN_308; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_310 = 6'hf == f2_cut_ptr_5 ? f2_cut_data_dataVec__15 : _GEN_309; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_311 = 6'h10 == f2_cut_ptr_5 ? f2_cut_data_dataVec__16 : _GEN_310; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_312 = 6'h11 == f2_cut_ptr_5 ? f2_cut_data_dataVec__17 : _GEN_311; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_313 = 6'h12 == f2_cut_ptr_5 ? f2_cut_data_dataVec__18 : _GEN_312; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_314 = 6'h13 == f2_cut_ptr_5 ? f2_cut_data_dataVec__19 : _GEN_313; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_315 = 6'h14 == f2_cut_ptr_5 ? f2_cut_data_dataVec__20 : _GEN_314; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_316 = 6'h15 == f2_cut_ptr_5 ? f2_cut_data_dataVec__21 : _GEN_315; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_317 = 6'h16 == f2_cut_ptr_5 ? f2_cut_data_dataVec__22 : _GEN_316; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_318 = 6'h17 == f2_cut_ptr_5 ? f2_cut_data_dataVec__23 : _GEN_317; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_319 = 6'h18 == f2_cut_ptr_5 ? f2_cut_data_dataVec__24 : _GEN_318; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_320 = 6'h19 == f2_cut_ptr_5 ? f2_cut_data_dataVec__25 : _GEN_319; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_321 = 6'h1a == f2_cut_ptr_5 ? f2_cut_data_dataVec__26 : _GEN_320; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_322 = 6'h1b == f2_cut_ptr_5 ? f2_cut_data_dataVec__27 : _GEN_321; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_323 = 6'h1c == f2_cut_ptr_5 ? f2_cut_data_dataVec__28 : _GEN_322; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_324 = 6'h1d == f2_cut_ptr_5 ? f2_cut_data_dataVec__29 : _GEN_323; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_325 = 6'h1e == f2_cut_ptr_5 ? f2_cut_data_dataVec__30 : _GEN_324; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_326 = 6'h1f == f2_cut_ptr_5 ? f2_cut_data_dataVec__31 : _GEN_325; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_327 = 6'h20 == f2_cut_ptr_5 ? f2_cut_data_dataVec__32 : _GEN_326; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_328 = 6'h21 == f2_cut_ptr_5 ? f2_cut_data_dataVec__33 : _GEN_327; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_329 = 6'h22 == f2_cut_ptr_5 ? f2_cut_data_dataVec__34 : _GEN_328; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_330 = 6'h23 == f2_cut_ptr_5 ? f2_cut_data_dataVec__35 : _GEN_329; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_331 = 6'h24 == f2_cut_ptr_5 ? f2_cut_data_dataVec__36 : _GEN_330; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_332 = 6'h25 == f2_cut_ptr_5 ? f2_cut_data_dataVec__37 : _GEN_331; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_333 = 6'h26 == f2_cut_ptr_5 ? f2_cut_data_dataVec__38 : _GEN_332; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_334 = 6'h27 == f2_cut_ptr_5 ? f2_cut_data_dataVec__39 : _GEN_333; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_335 = 6'h28 == f2_cut_ptr_5 ? f2_cut_data_dataVec__40 : _GEN_334; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_336 = 6'h29 == f2_cut_ptr_5 ? f2_cut_data_dataVec__41 : _GEN_335; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_337 = 6'h2a == f2_cut_ptr_5 ? f2_cut_data_dataVec__42 : _GEN_336; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_338 = 6'h2b == f2_cut_ptr_5 ? f2_cut_data_dataVec__43 : _GEN_337; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_339 = 6'h2c == f2_cut_ptr_5 ? f2_cut_data_dataVec__44 : _GEN_338; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_340 = 6'h2d == f2_cut_ptr_5 ? f2_cut_data_dataVec__45 : _GEN_339; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_341 = 6'h2e == f2_cut_ptr_5 ? f2_cut_data_dataVec__46 : _GEN_340; // @[IFU.scala 302:{19,19}]
  wire [15:0] f2_cut_data_result__5 = 6'h2f == f2_cut_ptr_5 ? f2_cut_data_dataVec__47 : _GEN_341; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_344 = 6'h1 == f2_cut_ptr_6 ? f2_cut_data_dataVec__1 : f2_cut_data_dataVec__0; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_345 = 6'h2 == f2_cut_ptr_6 ? f2_cut_data_dataVec__2 : _GEN_344; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_346 = 6'h3 == f2_cut_ptr_6 ? f2_cut_data_dataVec__3 : _GEN_345; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_347 = 6'h4 == f2_cut_ptr_6 ? f2_cut_data_dataVec__4 : _GEN_346; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_348 = 6'h5 == f2_cut_ptr_6 ? f2_cut_data_dataVec__5 : _GEN_347; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_349 = 6'h6 == f2_cut_ptr_6 ? f2_cut_data_dataVec__6 : _GEN_348; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_350 = 6'h7 == f2_cut_ptr_6 ? f2_cut_data_dataVec__7 : _GEN_349; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_351 = 6'h8 == f2_cut_ptr_6 ? f2_cut_data_dataVec__8 : _GEN_350; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_352 = 6'h9 == f2_cut_ptr_6 ? f2_cut_data_dataVec__9 : _GEN_351; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_353 = 6'ha == f2_cut_ptr_6 ? f2_cut_data_dataVec__10 : _GEN_352; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_354 = 6'hb == f2_cut_ptr_6 ? f2_cut_data_dataVec__11 : _GEN_353; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_355 = 6'hc == f2_cut_ptr_6 ? f2_cut_data_dataVec__12 : _GEN_354; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_356 = 6'hd == f2_cut_ptr_6 ? f2_cut_data_dataVec__13 : _GEN_355; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_357 = 6'he == f2_cut_ptr_6 ? f2_cut_data_dataVec__14 : _GEN_356; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_358 = 6'hf == f2_cut_ptr_6 ? f2_cut_data_dataVec__15 : _GEN_357; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_359 = 6'h10 == f2_cut_ptr_6 ? f2_cut_data_dataVec__16 : _GEN_358; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_360 = 6'h11 == f2_cut_ptr_6 ? f2_cut_data_dataVec__17 : _GEN_359; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_361 = 6'h12 == f2_cut_ptr_6 ? f2_cut_data_dataVec__18 : _GEN_360; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_362 = 6'h13 == f2_cut_ptr_6 ? f2_cut_data_dataVec__19 : _GEN_361; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_363 = 6'h14 == f2_cut_ptr_6 ? f2_cut_data_dataVec__20 : _GEN_362; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_364 = 6'h15 == f2_cut_ptr_6 ? f2_cut_data_dataVec__21 : _GEN_363; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_365 = 6'h16 == f2_cut_ptr_6 ? f2_cut_data_dataVec__22 : _GEN_364; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_366 = 6'h17 == f2_cut_ptr_6 ? f2_cut_data_dataVec__23 : _GEN_365; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_367 = 6'h18 == f2_cut_ptr_6 ? f2_cut_data_dataVec__24 : _GEN_366; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_368 = 6'h19 == f2_cut_ptr_6 ? f2_cut_data_dataVec__25 : _GEN_367; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_369 = 6'h1a == f2_cut_ptr_6 ? f2_cut_data_dataVec__26 : _GEN_368; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_370 = 6'h1b == f2_cut_ptr_6 ? f2_cut_data_dataVec__27 : _GEN_369; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_371 = 6'h1c == f2_cut_ptr_6 ? f2_cut_data_dataVec__28 : _GEN_370; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_372 = 6'h1d == f2_cut_ptr_6 ? f2_cut_data_dataVec__29 : _GEN_371; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_373 = 6'h1e == f2_cut_ptr_6 ? f2_cut_data_dataVec__30 : _GEN_372; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_374 = 6'h1f == f2_cut_ptr_6 ? f2_cut_data_dataVec__31 : _GEN_373; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_375 = 6'h20 == f2_cut_ptr_6 ? f2_cut_data_dataVec__32 : _GEN_374; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_376 = 6'h21 == f2_cut_ptr_6 ? f2_cut_data_dataVec__33 : _GEN_375; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_377 = 6'h22 == f2_cut_ptr_6 ? f2_cut_data_dataVec__34 : _GEN_376; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_378 = 6'h23 == f2_cut_ptr_6 ? f2_cut_data_dataVec__35 : _GEN_377; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_379 = 6'h24 == f2_cut_ptr_6 ? f2_cut_data_dataVec__36 : _GEN_378; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_380 = 6'h25 == f2_cut_ptr_6 ? f2_cut_data_dataVec__37 : _GEN_379; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_381 = 6'h26 == f2_cut_ptr_6 ? f2_cut_data_dataVec__38 : _GEN_380; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_382 = 6'h27 == f2_cut_ptr_6 ? f2_cut_data_dataVec__39 : _GEN_381; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_383 = 6'h28 == f2_cut_ptr_6 ? f2_cut_data_dataVec__40 : _GEN_382; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_384 = 6'h29 == f2_cut_ptr_6 ? f2_cut_data_dataVec__41 : _GEN_383; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_385 = 6'h2a == f2_cut_ptr_6 ? f2_cut_data_dataVec__42 : _GEN_384; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_386 = 6'h2b == f2_cut_ptr_6 ? f2_cut_data_dataVec__43 : _GEN_385; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_387 = 6'h2c == f2_cut_ptr_6 ? f2_cut_data_dataVec__44 : _GEN_386; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_388 = 6'h2d == f2_cut_ptr_6 ? f2_cut_data_dataVec__45 : _GEN_387; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_389 = 6'h2e == f2_cut_ptr_6 ? f2_cut_data_dataVec__46 : _GEN_388; // @[IFU.scala 302:{19,19}]
  wire [15:0] f2_cut_data_result__6 = 6'h2f == f2_cut_ptr_6 ? f2_cut_data_dataVec__47 : _GEN_389; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_392 = 6'h1 == f2_cut_ptr_7 ? f2_cut_data_dataVec__1 : f2_cut_data_dataVec__0; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_393 = 6'h2 == f2_cut_ptr_7 ? f2_cut_data_dataVec__2 : _GEN_392; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_394 = 6'h3 == f2_cut_ptr_7 ? f2_cut_data_dataVec__3 : _GEN_393; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_395 = 6'h4 == f2_cut_ptr_7 ? f2_cut_data_dataVec__4 : _GEN_394; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_396 = 6'h5 == f2_cut_ptr_7 ? f2_cut_data_dataVec__5 : _GEN_395; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_397 = 6'h6 == f2_cut_ptr_7 ? f2_cut_data_dataVec__6 : _GEN_396; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_398 = 6'h7 == f2_cut_ptr_7 ? f2_cut_data_dataVec__7 : _GEN_397; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_399 = 6'h8 == f2_cut_ptr_7 ? f2_cut_data_dataVec__8 : _GEN_398; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_400 = 6'h9 == f2_cut_ptr_7 ? f2_cut_data_dataVec__9 : _GEN_399; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_401 = 6'ha == f2_cut_ptr_7 ? f2_cut_data_dataVec__10 : _GEN_400; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_402 = 6'hb == f2_cut_ptr_7 ? f2_cut_data_dataVec__11 : _GEN_401; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_403 = 6'hc == f2_cut_ptr_7 ? f2_cut_data_dataVec__12 : _GEN_402; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_404 = 6'hd == f2_cut_ptr_7 ? f2_cut_data_dataVec__13 : _GEN_403; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_405 = 6'he == f2_cut_ptr_7 ? f2_cut_data_dataVec__14 : _GEN_404; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_406 = 6'hf == f2_cut_ptr_7 ? f2_cut_data_dataVec__15 : _GEN_405; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_407 = 6'h10 == f2_cut_ptr_7 ? f2_cut_data_dataVec__16 : _GEN_406; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_408 = 6'h11 == f2_cut_ptr_7 ? f2_cut_data_dataVec__17 : _GEN_407; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_409 = 6'h12 == f2_cut_ptr_7 ? f2_cut_data_dataVec__18 : _GEN_408; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_410 = 6'h13 == f2_cut_ptr_7 ? f2_cut_data_dataVec__19 : _GEN_409; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_411 = 6'h14 == f2_cut_ptr_7 ? f2_cut_data_dataVec__20 : _GEN_410; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_412 = 6'h15 == f2_cut_ptr_7 ? f2_cut_data_dataVec__21 : _GEN_411; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_413 = 6'h16 == f2_cut_ptr_7 ? f2_cut_data_dataVec__22 : _GEN_412; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_414 = 6'h17 == f2_cut_ptr_7 ? f2_cut_data_dataVec__23 : _GEN_413; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_415 = 6'h18 == f2_cut_ptr_7 ? f2_cut_data_dataVec__24 : _GEN_414; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_416 = 6'h19 == f2_cut_ptr_7 ? f2_cut_data_dataVec__25 : _GEN_415; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_417 = 6'h1a == f2_cut_ptr_7 ? f2_cut_data_dataVec__26 : _GEN_416; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_418 = 6'h1b == f2_cut_ptr_7 ? f2_cut_data_dataVec__27 : _GEN_417; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_419 = 6'h1c == f2_cut_ptr_7 ? f2_cut_data_dataVec__28 : _GEN_418; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_420 = 6'h1d == f2_cut_ptr_7 ? f2_cut_data_dataVec__29 : _GEN_419; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_421 = 6'h1e == f2_cut_ptr_7 ? f2_cut_data_dataVec__30 : _GEN_420; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_422 = 6'h1f == f2_cut_ptr_7 ? f2_cut_data_dataVec__31 : _GEN_421; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_423 = 6'h20 == f2_cut_ptr_7 ? f2_cut_data_dataVec__32 : _GEN_422; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_424 = 6'h21 == f2_cut_ptr_7 ? f2_cut_data_dataVec__33 : _GEN_423; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_425 = 6'h22 == f2_cut_ptr_7 ? f2_cut_data_dataVec__34 : _GEN_424; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_426 = 6'h23 == f2_cut_ptr_7 ? f2_cut_data_dataVec__35 : _GEN_425; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_427 = 6'h24 == f2_cut_ptr_7 ? f2_cut_data_dataVec__36 : _GEN_426; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_428 = 6'h25 == f2_cut_ptr_7 ? f2_cut_data_dataVec__37 : _GEN_427; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_429 = 6'h26 == f2_cut_ptr_7 ? f2_cut_data_dataVec__38 : _GEN_428; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_430 = 6'h27 == f2_cut_ptr_7 ? f2_cut_data_dataVec__39 : _GEN_429; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_431 = 6'h28 == f2_cut_ptr_7 ? f2_cut_data_dataVec__40 : _GEN_430; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_432 = 6'h29 == f2_cut_ptr_7 ? f2_cut_data_dataVec__41 : _GEN_431; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_433 = 6'h2a == f2_cut_ptr_7 ? f2_cut_data_dataVec__42 : _GEN_432; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_434 = 6'h2b == f2_cut_ptr_7 ? f2_cut_data_dataVec__43 : _GEN_433; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_435 = 6'h2c == f2_cut_ptr_7 ? f2_cut_data_dataVec__44 : _GEN_434; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_436 = 6'h2d == f2_cut_ptr_7 ? f2_cut_data_dataVec__45 : _GEN_435; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_437 = 6'h2e == f2_cut_ptr_7 ? f2_cut_data_dataVec__46 : _GEN_436; // @[IFU.scala 302:{19,19}]
  wire [15:0] f2_cut_data_result__7 = 6'h2f == f2_cut_ptr_7 ? f2_cut_data_dataVec__47 : _GEN_437; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_440 = 6'h1 == f2_cut_ptr_8 ? f2_cut_data_dataVec__1 : f2_cut_data_dataVec__0; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_441 = 6'h2 == f2_cut_ptr_8 ? f2_cut_data_dataVec__2 : _GEN_440; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_442 = 6'h3 == f2_cut_ptr_8 ? f2_cut_data_dataVec__3 : _GEN_441; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_443 = 6'h4 == f2_cut_ptr_8 ? f2_cut_data_dataVec__4 : _GEN_442; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_444 = 6'h5 == f2_cut_ptr_8 ? f2_cut_data_dataVec__5 : _GEN_443; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_445 = 6'h6 == f2_cut_ptr_8 ? f2_cut_data_dataVec__6 : _GEN_444; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_446 = 6'h7 == f2_cut_ptr_8 ? f2_cut_data_dataVec__7 : _GEN_445; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_447 = 6'h8 == f2_cut_ptr_8 ? f2_cut_data_dataVec__8 : _GEN_446; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_448 = 6'h9 == f2_cut_ptr_8 ? f2_cut_data_dataVec__9 : _GEN_447; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_449 = 6'ha == f2_cut_ptr_8 ? f2_cut_data_dataVec__10 : _GEN_448; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_450 = 6'hb == f2_cut_ptr_8 ? f2_cut_data_dataVec__11 : _GEN_449; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_451 = 6'hc == f2_cut_ptr_8 ? f2_cut_data_dataVec__12 : _GEN_450; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_452 = 6'hd == f2_cut_ptr_8 ? f2_cut_data_dataVec__13 : _GEN_451; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_453 = 6'he == f2_cut_ptr_8 ? f2_cut_data_dataVec__14 : _GEN_452; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_454 = 6'hf == f2_cut_ptr_8 ? f2_cut_data_dataVec__15 : _GEN_453; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_455 = 6'h10 == f2_cut_ptr_8 ? f2_cut_data_dataVec__16 : _GEN_454; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_456 = 6'h11 == f2_cut_ptr_8 ? f2_cut_data_dataVec__17 : _GEN_455; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_457 = 6'h12 == f2_cut_ptr_8 ? f2_cut_data_dataVec__18 : _GEN_456; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_458 = 6'h13 == f2_cut_ptr_8 ? f2_cut_data_dataVec__19 : _GEN_457; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_459 = 6'h14 == f2_cut_ptr_8 ? f2_cut_data_dataVec__20 : _GEN_458; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_460 = 6'h15 == f2_cut_ptr_8 ? f2_cut_data_dataVec__21 : _GEN_459; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_461 = 6'h16 == f2_cut_ptr_8 ? f2_cut_data_dataVec__22 : _GEN_460; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_462 = 6'h17 == f2_cut_ptr_8 ? f2_cut_data_dataVec__23 : _GEN_461; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_463 = 6'h18 == f2_cut_ptr_8 ? f2_cut_data_dataVec__24 : _GEN_462; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_464 = 6'h19 == f2_cut_ptr_8 ? f2_cut_data_dataVec__25 : _GEN_463; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_465 = 6'h1a == f2_cut_ptr_8 ? f2_cut_data_dataVec__26 : _GEN_464; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_466 = 6'h1b == f2_cut_ptr_8 ? f2_cut_data_dataVec__27 : _GEN_465; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_467 = 6'h1c == f2_cut_ptr_8 ? f2_cut_data_dataVec__28 : _GEN_466; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_468 = 6'h1d == f2_cut_ptr_8 ? f2_cut_data_dataVec__29 : _GEN_467; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_469 = 6'h1e == f2_cut_ptr_8 ? f2_cut_data_dataVec__30 : _GEN_468; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_470 = 6'h1f == f2_cut_ptr_8 ? f2_cut_data_dataVec__31 : _GEN_469; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_471 = 6'h20 == f2_cut_ptr_8 ? f2_cut_data_dataVec__32 : _GEN_470; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_472 = 6'h21 == f2_cut_ptr_8 ? f2_cut_data_dataVec__33 : _GEN_471; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_473 = 6'h22 == f2_cut_ptr_8 ? f2_cut_data_dataVec__34 : _GEN_472; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_474 = 6'h23 == f2_cut_ptr_8 ? f2_cut_data_dataVec__35 : _GEN_473; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_475 = 6'h24 == f2_cut_ptr_8 ? f2_cut_data_dataVec__36 : _GEN_474; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_476 = 6'h25 == f2_cut_ptr_8 ? f2_cut_data_dataVec__37 : _GEN_475; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_477 = 6'h26 == f2_cut_ptr_8 ? f2_cut_data_dataVec__38 : _GEN_476; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_478 = 6'h27 == f2_cut_ptr_8 ? f2_cut_data_dataVec__39 : _GEN_477; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_479 = 6'h28 == f2_cut_ptr_8 ? f2_cut_data_dataVec__40 : _GEN_478; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_480 = 6'h29 == f2_cut_ptr_8 ? f2_cut_data_dataVec__41 : _GEN_479; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_481 = 6'h2a == f2_cut_ptr_8 ? f2_cut_data_dataVec__42 : _GEN_480; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_482 = 6'h2b == f2_cut_ptr_8 ? f2_cut_data_dataVec__43 : _GEN_481; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_483 = 6'h2c == f2_cut_ptr_8 ? f2_cut_data_dataVec__44 : _GEN_482; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_484 = 6'h2d == f2_cut_ptr_8 ? f2_cut_data_dataVec__45 : _GEN_483; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_485 = 6'h2e == f2_cut_ptr_8 ? f2_cut_data_dataVec__46 : _GEN_484; // @[IFU.scala 302:{19,19}]
  wire [15:0] f2_cut_data_result__8 = 6'h2f == f2_cut_ptr_8 ? f2_cut_data_dataVec__47 : _GEN_485; // @[IFU.scala 302:{19,19}]
  wire [767:0] f2_cut_data_partCacheline_1 = f2_data_2_cacheline_1[767:0]; // @[IFU.scala 298:36]
  wire [15:0] f2_cut_data_dataVec_1_0 = f2_cut_data_partCacheline_1[15:0]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_1_1 = f2_cut_data_partCacheline_1[31:16]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_1_2 = f2_cut_data_partCacheline_1[47:32]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_1_3 = f2_cut_data_partCacheline_1[63:48]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_1_4 = f2_cut_data_partCacheline_1[79:64]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_1_5 = f2_cut_data_partCacheline_1[95:80]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_1_6 = f2_cut_data_partCacheline_1[111:96]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_1_7 = f2_cut_data_partCacheline_1[127:112]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_1_8 = f2_cut_data_partCacheline_1[143:128]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_1_9 = f2_cut_data_partCacheline_1[159:144]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_1_10 = f2_cut_data_partCacheline_1[175:160]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_1_11 = f2_cut_data_partCacheline_1[191:176]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_1_12 = f2_cut_data_partCacheline_1[207:192]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_1_13 = f2_cut_data_partCacheline_1[223:208]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_1_14 = f2_cut_data_partCacheline_1[239:224]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_1_15 = f2_cut_data_partCacheline_1[255:240]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_1_16 = f2_cut_data_partCacheline_1[271:256]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_1_17 = f2_cut_data_partCacheline_1[287:272]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_1_18 = f2_cut_data_partCacheline_1[303:288]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_1_19 = f2_cut_data_partCacheline_1[319:304]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_1_20 = f2_cut_data_partCacheline_1[335:320]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_1_21 = f2_cut_data_partCacheline_1[351:336]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_1_22 = f2_cut_data_partCacheline_1[367:352]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_1_23 = f2_cut_data_partCacheline_1[383:368]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_1_24 = f2_cut_data_partCacheline_1[399:384]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_1_25 = f2_cut_data_partCacheline_1[415:400]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_1_26 = f2_cut_data_partCacheline_1[431:416]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_1_27 = f2_cut_data_partCacheline_1[447:432]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_1_28 = f2_cut_data_partCacheline_1[463:448]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_1_29 = f2_cut_data_partCacheline_1[479:464]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_1_30 = f2_cut_data_partCacheline_1[495:480]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_1_31 = f2_cut_data_partCacheline_1[511:496]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_1_32 = f2_cut_data_partCacheline_1[527:512]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_1_33 = f2_cut_data_partCacheline_1[543:528]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_1_34 = f2_cut_data_partCacheline_1[559:544]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_1_35 = f2_cut_data_partCacheline_1[575:560]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_1_36 = f2_cut_data_partCacheline_1[591:576]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_1_37 = f2_cut_data_partCacheline_1[607:592]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_1_38 = f2_cut_data_partCacheline_1[623:608]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_1_39 = f2_cut_data_partCacheline_1[639:624]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_1_40 = f2_cut_data_partCacheline_1[655:640]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_1_41 = f2_cut_data_partCacheline_1[671:656]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_1_42 = f2_cut_data_partCacheline_1[687:672]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_1_43 = f2_cut_data_partCacheline_1[703:688]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_1_44 = f2_cut_data_partCacheline_1[719:704]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_1_45 = f2_cut_data_partCacheline_1[735:720]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_1_46 = f2_cut_data_partCacheline_1[751:736]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_1_47 = f2_cut_data_partCacheline_1[767:752]; // @[IFU.scala 300:40]
  wire [15:0] _GEN_488 = 6'h1 == f2_cut_ptr_0 ? f2_cut_data_dataVec_1_1 : f2_cut_data_dataVec_1_0; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_489 = 6'h2 == f2_cut_ptr_0 ? f2_cut_data_dataVec_1_2 : _GEN_488; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_490 = 6'h3 == f2_cut_ptr_0 ? f2_cut_data_dataVec_1_3 : _GEN_489; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_491 = 6'h4 == f2_cut_ptr_0 ? f2_cut_data_dataVec_1_4 : _GEN_490; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_492 = 6'h5 == f2_cut_ptr_0 ? f2_cut_data_dataVec_1_5 : _GEN_491; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_493 = 6'h6 == f2_cut_ptr_0 ? f2_cut_data_dataVec_1_6 : _GEN_492; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_494 = 6'h7 == f2_cut_ptr_0 ? f2_cut_data_dataVec_1_7 : _GEN_493; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_495 = 6'h8 == f2_cut_ptr_0 ? f2_cut_data_dataVec_1_8 : _GEN_494; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_496 = 6'h9 == f2_cut_ptr_0 ? f2_cut_data_dataVec_1_9 : _GEN_495; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_497 = 6'ha == f2_cut_ptr_0 ? f2_cut_data_dataVec_1_10 : _GEN_496; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_498 = 6'hb == f2_cut_ptr_0 ? f2_cut_data_dataVec_1_11 : _GEN_497; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_499 = 6'hc == f2_cut_ptr_0 ? f2_cut_data_dataVec_1_12 : _GEN_498; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_500 = 6'hd == f2_cut_ptr_0 ? f2_cut_data_dataVec_1_13 : _GEN_499; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_501 = 6'he == f2_cut_ptr_0 ? f2_cut_data_dataVec_1_14 : _GEN_500; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_502 = 6'hf == f2_cut_ptr_0 ? f2_cut_data_dataVec_1_15 : _GEN_501; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_503 = 6'h10 == f2_cut_ptr_0 ? f2_cut_data_dataVec_1_16 : _GEN_502; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_504 = 6'h11 == f2_cut_ptr_0 ? f2_cut_data_dataVec_1_17 : _GEN_503; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_505 = 6'h12 == f2_cut_ptr_0 ? f2_cut_data_dataVec_1_18 : _GEN_504; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_506 = 6'h13 == f2_cut_ptr_0 ? f2_cut_data_dataVec_1_19 : _GEN_505; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_507 = 6'h14 == f2_cut_ptr_0 ? f2_cut_data_dataVec_1_20 : _GEN_506; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_508 = 6'h15 == f2_cut_ptr_0 ? f2_cut_data_dataVec_1_21 : _GEN_507; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_509 = 6'h16 == f2_cut_ptr_0 ? f2_cut_data_dataVec_1_22 : _GEN_508; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_510 = 6'h17 == f2_cut_ptr_0 ? f2_cut_data_dataVec_1_23 : _GEN_509; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_511 = 6'h18 == f2_cut_ptr_0 ? f2_cut_data_dataVec_1_24 : _GEN_510; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_512 = 6'h19 == f2_cut_ptr_0 ? f2_cut_data_dataVec_1_25 : _GEN_511; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_513 = 6'h1a == f2_cut_ptr_0 ? f2_cut_data_dataVec_1_26 : _GEN_512; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_514 = 6'h1b == f2_cut_ptr_0 ? f2_cut_data_dataVec_1_27 : _GEN_513; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_515 = 6'h1c == f2_cut_ptr_0 ? f2_cut_data_dataVec_1_28 : _GEN_514; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_516 = 6'h1d == f2_cut_ptr_0 ? f2_cut_data_dataVec_1_29 : _GEN_515; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_517 = 6'h1e == f2_cut_ptr_0 ? f2_cut_data_dataVec_1_30 : _GEN_516; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_518 = 6'h1f == f2_cut_ptr_0 ? f2_cut_data_dataVec_1_31 : _GEN_517; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_519 = 6'h20 == f2_cut_ptr_0 ? f2_cut_data_dataVec_1_32 : _GEN_518; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_520 = 6'h21 == f2_cut_ptr_0 ? f2_cut_data_dataVec_1_33 : _GEN_519; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_521 = 6'h22 == f2_cut_ptr_0 ? f2_cut_data_dataVec_1_34 : _GEN_520; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_522 = 6'h23 == f2_cut_ptr_0 ? f2_cut_data_dataVec_1_35 : _GEN_521; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_523 = 6'h24 == f2_cut_ptr_0 ? f2_cut_data_dataVec_1_36 : _GEN_522; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_524 = 6'h25 == f2_cut_ptr_0 ? f2_cut_data_dataVec_1_37 : _GEN_523; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_525 = 6'h26 == f2_cut_ptr_0 ? f2_cut_data_dataVec_1_38 : _GEN_524; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_526 = 6'h27 == f2_cut_ptr_0 ? f2_cut_data_dataVec_1_39 : _GEN_525; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_527 = 6'h28 == f2_cut_ptr_0 ? f2_cut_data_dataVec_1_40 : _GEN_526; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_528 = 6'h29 == f2_cut_ptr_0 ? f2_cut_data_dataVec_1_41 : _GEN_527; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_529 = 6'h2a == f2_cut_ptr_0 ? f2_cut_data_dataVec_1_42 : _GEN_528; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_530 = 6'h2b == f2_cut_ptr_0 ? f2_cut_data_dataVec_1_43 : _GEN_529; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_531 = 6'h2c == f2_cut_ptr_0 ? f2_cut_data_dataVec_1_44 : _GEN_530; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_532 = 6'h2d == f2_cut_ptr_0 ? f2_cut_data_dataVec_1_45 : _GEN_531; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_533 = 6'h2e == f2_cut_ptr_0 ? f2_cut_data_dataVec_1_46 : _GEN_532; // @[IFU.scala 302:{19,19}]
  wire [15:0] f2_cut_data_result_1_0 = 6'h2f == f2_cut_ptr_0 ? f2_cut_data_dataVec_1_47 : _GEN_533; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_536 = 6'h1 == f2_cut_ptr_1 ? f2_cut_data_dataVec_1_1 : f2_cut_data_dataVec_1_0; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_537 = 6'h2 == f2_cut_ptr_1 ? f2_cut_data_dataVec_1_2 : _GEN_536; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_538 = 6'h3 == f2_cut_ptr_1 ? f2_cut_data_dataVec_1_3 : _GEN_537; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_539 = 6'h4 == f2_cut_ptr_1 ? f2_cut_data_dataVec_1_4 : _GEN_538; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_540 = 6'h5 == f2_cut_ptr_1 ? f2_cut_data_dataVec_1_5 : _GEN_539; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_541 = 6'h6 == f2_cut_ptr_1 ? f2_cut_data_dataVec_1_6 : _GEN_540; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_542 = 6'h7 == f2_cut_ptr_1 ? f2_cut_data_dataVec_1_7 : _GEN_541; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_543 = 6'h8 == f2_cut_ptr_1 ? f2_cut_data_dataVec_1_8 : _GEN_542; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_544 = 6'h9 == f2_cut_ptr_1 ? f2_cut_data_dataVec_1_9 : _GEN_543; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_545 = 6'ha == f2_cut_ptr_1 ? f2_cut_data_dataVec_1_10 : _GEN_544; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_546 = 6'hb == f2_cut_ptr_1 ? f2_cut_data_dataVec_1_11 : _GEN_545; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_547 = 6'hc == f2_cut_ptr_1 ? f2_cut_data_dataVec_1_12 : _GEN_546; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_548 = 6'hd == f2_cut_ptr_1 ? f2_cut_data_dataVec_1_13 : _GEN_547; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_549 = 6'he == f2_cut_ptr_1 ? f2_cut_data_dataVec_1_14 : _GEN_548; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_550 = 6'hf == f2_cut_ptr_1 ? f2_cut_data_dataVec_1_15 : _GEN_549; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_551 = 6'h10 == f2_cut_ptr_1 ? f2_cut_data_dataVec_1_16 : _GEN_550; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_552 = 6'h11 == f2_cut_ptr_1 ? f2_cut_data_dataVec_1_17 : _GEN_551; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_553 = 6'h12 == f2_cut_ptr_1 ? f2_cut_data_dataVec_1_18 : _GEN_552; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_554 = 6'h13 == f2_cut_ptr_1 ? f2_cut_data_dataVec_1_19 : _GEN_553; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_555 = 6'h14 == f2_cut_ptr_1 ? f2_cut_data_dataVec_1_20 : _GEN_554; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_556 = 6'h15 == f2_cut_ptr_1 ? f2_cut_data_dataVec_1_21 : _GEN_555; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_557 = 6'h16 == f2_cut_ptr_1 ? f2_cut_data_dataVec_1_22 : _GEN_556; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_558 = 6'h17 == f2_cut_ptr_1 ? f2_cut_data_dataVec_1_23 : _GEN_557; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_559 = 6'h18 == f2_cut_ptr_1 ? f2_cut_data_dataVec_1_24 : _GEN_558; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_560 = 6'h19 == f2_cut_ptr_1 ? f2_cut_data_dataVec_1_25 : _GEN_559; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_561 = 6'h1a == f2_cut_ptr_1 ? f2_cut_data_dataVec_1_26 : _GEN_560; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_562 = 6'h1b == f2_cut_ptr_1 ? f2_cut_data_dataVec_1_27 : _GEN_561; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_563 = 6'h1c == f2_cut_ptr_1 ? f2_cut_data_dataVec_1_28 : _GEN_562; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_564 = 6'h1d == f2_cut_ptr_1 ? f2_cut_data_dataVec_1_29 : _GEN_563; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_565 = 6'h1e == f2_cut_ptr_1 ? f2_cut_data_dataVec_1_30 : _GEN_564; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_566 = 6'h1f == f2_cut_ptr_1 ? f2_cut_data_dataVec_1_31 : _GEN_565; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_567 = 6'h20 == f2_cut_ptr_1 ? f2_cut_data_dataVec_1_32 : _GEN_566; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_568 = 6'h21 == f2_cut_ptr_1 ? f2_cut_data_dataVec_1_33 : _GEN_567; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_569 = 6'h22 == f2_cut_ptr_1 ? f2_cut_data_dataVec_1_34 : _GEN_568; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_570 = 6'h23 == f2_cut_ptr_1 ? f2_cut_data_dataVec_1_35 : _GEN_569; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_571 = 6'h24 == f2_cut_ptr_1 ? f2_cut_data_dataVec_1_36 : _GEN_570; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_572 = 6'h25 == f2_cut_ptr_1 ? f2_cut_data_dataVec_1_37 : _GEN_571; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_573 = 6'h26 == f2_cut_ptr_1 ? f2_cut_data_dataVec_1_38 : _GEN_572; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_574 = 6'h27 == f2_cut_ptr_1 ? f2_cut_data_dataVec_1_39 : _GEN_573; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_575 = 6'h28 == f2_cut_ptr_1 ? f2_cut_data_dataVec_1_40 : _GEN_574; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_576 = 6'h29 == f2_cut_ptr_1 ? f2_cut_data_dataVec_1_41 : _GEN_575; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_577 = 6'h2a == f2_cut_ptr_1 ? f2_cut_data_dataVec_1_42 : _GEN_576; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_578 = 6'h2b == f2_cut_ptr_1 ? f2_cut_data_dataVec_1_43 : _GEN_577; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_579 = 6'h2c == f2_cut_ptr_1 ? f2_cut_data_dataVec_1_44 : _GEN_578; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_580 = 6'h2d == f2_cut_ptr_1 ? f2_cut_data_dataVec_1_45 : _GEN_579; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_581 = 6'h2e == f2_cut_ptr_1 ? f2_cut_data_dataVec_1_46 : _GEN_580; // @[IFU.scala 302:{19,19}]
  wire [15:0] f2_cut_data_result_1_1 = 6'h2f == f2_cut_ptr_1 ? f2_cut_data_dataVec_1_47 : _GEN_581; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_584 = 6'h1 == f2_cut_ptr_2 ? f2_cut_data_dataVec_1_1 : f2_cut_data_dataVec_1_0; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_585 = 6'h2 == f2_cut_ptr_2 ? f2_cut_data_dataVec_1_2 : _GEN_584; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_586 = 6'h3 == f2_cut_ptr_2 ? f2_cut_data_dataVec_1_3 : _GEN_585; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_587 = 6'h4 == f2_cut_ptr_2 ? f2_cut_data_dataVec_1_4 : _GEN_586; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_588 = 6'h5 == f2_cut_ptr_2 ? f2_cut_data_dataVec_1_5 : _GEN_587; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_589 = 6'h6 == f2_cut_ptr_2 ? f2_cut_data_dataVec_1_6 : _GEN_588; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_590 = 6'h7 == f2_cut_ptr_2 ? f2_cut_data_dataVec_1_7 : _GEN_589; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_591 = 6'h8 == f2_cut_ptr_2 ? f2_cut_data_dataVec_1_8 : _GEN_590; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_592 = 6'h9 == f2_cut_ptr_2 ? f2_cut_data_dataVec_1_9 : _GEN_591; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_593 = 6'ha == f2_cut_ptr_2 ? f2_cut_data_dataVec_1_10 : _GEN_592; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_594 = 6'hb == f2_cut_ptr_2 ? f2_cut_data_dataVec_1_11 : _GEN_593; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_595 = 6'hc == f2_cut_ptr_2 ? f2_cut_data_dataVec_1_12 : _GEN_594; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_596 = 6'hd == f2_cut_ptr_2 ? f2_cut_data_dataVec_1_13 : _GEN_595; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_597 = 6'he == f2_cut_ptr_2 ? f2_cut_data_dataVec_1_14 : _GEN_596; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_598 = 6'hf == f2_cut_ptr_2 ? f2_cut_data_dataVec_1_15 : _GEN_597; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_599 = 6'h10 == f2_cut_ptr_2 ? f2_cut_data_dataVec_1_16 : _GEN_598; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_600 = 6'h11 == f2_cut_ptr_2 ? f2_cut_data_dataVec_1_17 : _GEN_599; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_601 = 6'h12 == f2_cut_ptr_2 ? f2_cut_data_dataVec_1_18 : _GEN_600; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_602 = 6'h13 == f2_cut_ptr_2 ? f2_cut_data_dataVec_1_19 : _GEN_601; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_603 = 6'h14 == f2_cut_ptr_2 ? f2_cut_data_dataVec_1_20 : _GEN_602; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_604 = 6'h15 == f2_cut_ptr_2 ? f2_cut_data_dataVec_1_21 : _GEN_603; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_605 = 6'h16 == f2_cut_ptr_2 ? f2_cut_data_dataVec_1_22 : _GEN_604; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_606 = 6'h17 == f2_cut_ptr_2 ? f2_cut_data_dataVec_1_23 : _GEN_605; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_607 = 6'h18 == f2_cut_ptr_2 ? f2_cut_data_dataVec_1_24 : _GEN_606; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_608 = 6'h19 == f2_cut_ptr_2 ? f2_cut_data_dataVec_1_25 : _GEN_607; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_609 = 6'h1a == f2_cut_ptr_2 ? f2_cut_data_dataVec_1_26 : _GEN_608; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_610 = 6'h1b == f2_cut_ptr_2 ? f2_cut_data_dataVec_1_27 : _GEN_609; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_611 = 6'h1c == f2_cut_ptr_2 ? f2_cut_data_dataVec_1_28 : _GEN_610; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_612 = 6'h1d == f2_cut_ptr_2 ? f2_cut_data_dataVec_1_29 : _GEN_611; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_613 = 6'h1e == f2_cut_ptr_2 ? f2_cut_data_dataVec_1_30 : _GEN_612; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_614 = 6'h1f == f2_cut_ptr_2 ? f2_cut_data_dataVec_1_31 : _GEN_613; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_615 = 6'h20 == f2_cut_ptr_2 ? f2_cut_data_dataVec_1_32 : _GEN_614; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_616 = 6'h21 == f2_cut_ptr_2 ? f2_cut_data_dataVec_1_33 : _GEN_615; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_617 = 6'h22 == f2_cut_ptr_2 ? f2_cut_data_dataVec_1_34 : _GEN_616; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_618 = 6'h23 == f2_cut_ptr_2 ? f2_cut_data_dataVec_1_35 : _GEN_617; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_619 = 6'h24 == f2_cut_ptr_2 ? f2_cut_data_dataVec_1_36 : _GEN_618; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_620 = 6'h25 == f2_cut_ptr_2 ? f2_cut_data_dataVec_1_37 : _GEN_619; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_621 = 6'h26 == f2_cut_ptr_2 ? f2_cut_data_dataVec_1_38 : _GEN_620; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_622 = 6'h27 == f2_cut_ptr_2 ? f2_cut_data_dataVec_1_39 : _GEN_621; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_623 = 6'h28 == f2_cut_ptr_2 ? f2_cut_data_dataVec_1_40 : _GEN_622; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_624 = 6'h29 == f2_cut_ptr_2 ? f2_cut_data_dataVec_1_41 : _GEN_623; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_625 = 6'h2a == f2_cut_ptr_2 ? f2_cut_data_dataVec_1_42 : _GEN_624; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_626 = 6'h2b == f2_cut_ptr_2 ? f2_cut_data_dataVec_1_43 : _GEN_625; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_627 = 6'h2c == f2_cut_ptr_2 ? f2_cut_data_dataVec_1_44 : _GEN_626; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_628 = 6'h2d == f2_cut_ptr_2 ? f2_cut_data_dataVec_1_45 : _GEN_627; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_629 = 6'h2e == f2_cut_ptr_2 ? f2_cut_data_dataVec_1_46 : _GEN_628; // @[IFU.scala 302:{19,19}]
  wire [15:0] f2_cut_data_result_1_2 = 6'h2f == f2_cut_ptr_2 ? f2_cut_data_dataVec_1_47 : _GEN_629; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_632 = 6'h1 == f2_cut_ptr_3 ? f2_cut_data_dataVec_1_1 : f2_cut_data_dataVec_1_0; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_633 = 6'h2 == f2_cut_ptr_3 ? f2_cut_data_dataVec_1_2 : _GEN_632; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_634 = 6'h3 == f2_cut_ptr_3 ? f2_cut_data_dataVec_1_3 : _GEN_633; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_635 = 6'h4 == f2_cut_ptr_3 ? f2_cut_data_dataVec_1_4 : _GEN_634; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_636 = 6'h5 == f2_cut_ptr_3 ? f2_cut_data_dataVec_1_5 : _GEN_635; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_637 = 6'h6 == f2_cut_ptr_3 ? f2_cut_data_dataVec_1_6 : _GEN_636; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_638 = 6'h7 == f2_cut_ptr_3 ? f2_cut_data_dataVec_1_7 : _GEN_637; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_639 = 6'h8 == f2_cut_ptr_3 ? f2_cut_data_dataVec_1_8 : _GEN_638; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_640 = 6'h9 == f2_cut_ptr_3 ? f2_cut_data_dataVec_1_9 : _GEN_639; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_641 = 6'ha == f2_cut_ptr_3 ? f2_cut_data_dataVec_1_10 : _GEN_640; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_642 = 6'hb == f2_cut_ptr_3 ? f2_cut_data_dataVec_1_11 : _GEN_641; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_643 = 6'hc == f2_cut_ptr_3 ? f2_cut_data_dataVec_1_12 : _GEN_642; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_644 = 6'hd == f2_cut_ptr_3 ? f2_cut_data_dataVec_1_13 : _GEN_643; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_645 = 6'he == f2_cut_ptr_3 ? f2_cut_data_dataVec_1_14 : _GEN_644; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_646 = 6'hf == f2_cut_ptr_3 ? f2_cut_data_dataVec_1_15 : _GEN_645; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_647 = 6'h10 == f2_cut_ptr_3 ? f2_cut_data_dataVec_1_16 : _GEN_646; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_648 = 6'h11 == f2_cut_ptr_3 ? f2_cut_data_dataVec_1_17 : _GEN_647; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_649 = 6'h12 == f2_cut_ptr_3 ? f2_cut_data_dataVec_1_18 : _GEN_648; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_650 = 6'h13 == f2_cut_ptr_3 ? f2_cut_data_dataVec_1_19 : _GEN_649; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_651 = 6'h14 == f2_cut_ptr_3 ? f2_cut_data_dataVec_1_20 : _GEN_650; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_652 = 6'h15 == f2_cut_ptr_3 ? f2_cut_data_dataVec_1_21 : _GEN_651; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_653 = 6'h16 == f2_cut_ptr_3 ? f2_cut_data_dataVec_1_22 : _GEN_652; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_654 = 6'h17 == f2_cut_ptr_3 ? f2_cut_data_dataVec_1_23 : _GEN_653; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_655 = 6'h18 == f2_cut_ptr_3 ? f2_cut_data_dataVec_1_24 : _GEN_654; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_656 = 6'h19 == f2_cut_ptr_3 ? f2_cut_data_dataVec_1_25 : _GEN_655; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_657 = 6'h1a == f2_cut_ptr_3 ? f2_cut_data_dataVec_1_26 : _GEN_656; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_658 = 6'h1b == f2_cut_ptr_3 ? f2_cut_data_dataVec_1_27 : _GEN_657; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_659 = 6'h1c == f2_cut_ptr_3 ? f2_cut_data_dataVec_1_28 : _GEN_658; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_660 = 6'h1d == f2_cut_ptr_3 ? f2_cut_data_dataVec_1_29 : _GEN_659; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_661 = 6'h1e == f2_cut_ptr_3 ? f2_cut_data_dataVec_1_30 : _GEN_660; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_662 = 6'h1f == f2_cut_ptr_3 ? f2_cut_data_dataVec_1_31 : _GEN_661; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_663 = 6'h20 == f2_cut_ptr_3 ? f2_cut_data_dataVec_1_32 : _GEN_662; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_664 = 6'h21 == f2_cut_ptr_3 ? f2_cut_data_dataVec_1_33 : _GEN_663; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_665 = 6'h22 == f2_cut_ptr_3 ? f2_cut_data_dataVec_1_34 : _GEN_664; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_666 = 6'h23 == f2_cut_ptr_3 ? f2_cut_data_dataVec_1_35 : _GEN_665; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_667 = 6'h24 == f2_cut_ptr_3 ? f2_cut_data_dataVec_1_36 : _GEN_666; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_668 = 6'h25 == f2_cut_ptr_3 ? f2_cut_data_dataVec_1_37 : _GEN_667; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_669 = 6'h26 == f2_cut_ptr_3 ? f2_cut_data_dataVec_1_38 : _GEN_668; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_670 = 6'h27 == f2_cut_ptr_3 ? f2_cut_data_dataVec_1_39 : _GEN_669; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_671 = 6'h28 == f2_cut_ptr_3 ? f2_cut_data_dataVec_1_40 : _GEN_670; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_672 = 6'h29 == f2_cut_ptr_3 ? f2_cut_data_dataVec_1_41 : _GEN_671; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_673 = 6'h2a == f2_cut_ptr_3 ? f2_cut_data_dataVec_1_42 : _GEN_672; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_674 = 6'h2b == f2_cut_ptr_3 ? f2_cut_data_dataVec_1_43 : _GEN_673; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_675 = 6'h2c == f2_cut_ptr_3 ? f2_cut_data_dataVec_1_44 : _GEN_674; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_676 = 6'h2d == f2_cut_ptr_3 ? f2_cut_data_dataVec_1_45 : _GEN_675; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_677 = 6'h2e == f2_cut_ptr_3 ? f2_cut_data_dataVec_1_46 : _GEN_676; // @[IFU.scala 302:{19,19}]
  wire [15:0] f2_cut_data_result_1_3 = 6'h2f == f2_cut_ptr_3 ? f2_cut_data_dataVec_1_47 : _GEN_677; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_680 = 6'h1 == f2_cut_ptr_4 ? f2_cut_data_dataVec_1_1 : f2_cut_data_dataVec_1_0; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_681 = 6'h2 == f2_cut_ptr_4 ? f2_cut_data_dataVec_1_2 : _GEN_680; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_682 = 6'h3 == f2_cut_ptr_4 ? f2_cut_data_dataVec_1_3 : _GEN_681; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_683 = 6'h4 == f2_cut_ptr_4 ? f2_cut_data_dataVec_1_4 : _GEN_682; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_684 = 6'h5 == f2_cut_ptr_4 ? f2_cut_data_dataVec_1_5 : _GEN_683; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_685 = 6'h6 == f2_cut_ptr_4 ? f2_cut_data_dataVec_1_6 : _GEN_684; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_686 = 6'h7 == f2_cut_ptr_4 ? f2_cut_data_dataVec_1_7 : _GEN_685; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_687 = 6'h8 == f2_cut_ptr_4 ? f2_cut_data_dataVec_1_8 : _GEN_686; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_688 = 6'h9 == f2_cut_ptr_4 ? f2_cut_data_dataVec_1_9 : _GEN_687; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_689 = 6'ha == f2_cut_ptr_4 ? f2_cut_data_dataVec_1_10 : _GEN_688; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_690 = 6'hb == f2_cut_ptr_4 ? f2_cut_data_dataVec_1_11 : _GEN_689; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_691 = 6'hc == f2_cut_ptr_4 ? f2_cut_data_dataVec_1_12 : _GEN_690; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_692 = 6'hd == f2_cut_ptr_4 ? f2_cut_data_dataVec_1_13 : _GEN_691; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_693 = 6'he == f2_cut_ptr_4 ? f2_cut_data_dataVec_1_14 : _GEN_692; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_694 = 6'hf == f2_cut_ptr_4 ? f2_cut_data_dataVec_1_15 : _GEN_693; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_695 = 6'h10 == f2_cut_ptr_4 ? f2_cut_data_dataVec_1_16 : _GEN_694; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_696 = 6'h11 == f2_cut_ptr_4 ? f2_cut_data_dataVec_1_17 : _GEN_695; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_697 = 6'h12 == f2_cut_ptr_4 ? f2_cut_data_dataVec_1_18 : _GEN_696; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_698 = 6'h13 == f2_cut_ptr_4 ? f2_cut_data_dataVec_1_19 : _GEN_697; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_699 = 6'h14 == f2_cut_ptr_4 ? f2_cut_data_dataVec_1_20 : _GEN_698; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_700 = 6'h15 == f2_cut_ptr_4 ? f2_cut_data_dataVec_1_21 : _GEN_699; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_701 = 6'h16 == f2_cut_ptr_4 ? f2_cut_data_dataVec_1_22 : _GEN_700; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_702 = 6'h17 == f2_cut_ptr_4 ? f2_cut_data_dataVec_1_23 : _GEN_701; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_703 = 6'h18 == f2_cut_ptr_4 ? f2_cut_data_dataVec_1_24 : _GEN_702; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_704 = 6'h19 == f2_cut_ptr_4 ? f2_cut_data_dataVec_1_25 : _GEN_703; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_705 = 6'h1a == f2_cut_ptr_4 ? f2_cut_data_dataVec_1_26 : _GEN_704; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_706 = 6'h1b == f2_cut_ptr_4 ? f2_cut_data_dataVec_1_27 : _GEN_705; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_707 = 6'h1c == f2_cut_ptr_4 ? f2_cut_data_dataVec_1_28 : _GEN_706; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_708 = 6'h1d == f2_cut_ptr_4 ? f2_cut_data_dataVec_1_29 : _GEN_707; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_709 = 6'h1e == f2_cut_ptr_4 ? f2_cut_data_dataVec_1_30 : _GEN_708; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_710 = 6'h1f == f2_cut_ptr_4 ? f2_cut_data_dataVec_1_31 : _GEN_709; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_711 = 6'h20 == f2_cut_ptr_4 ? f2_cut_data_dataVec_1_32 : _GEN_710; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_712 = 6'h21 == f2_cut_ptr_4 ? f2_cut_data_dataVec_1_33 : _GEN_711; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_713 = 6'h22 == f2_cut_ptr_4 ? f2_cut_data_dataVec_1_34 : _GEN_712; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_714 = 6'h23 == f2_cut_ptr_4 ? f2_cut_data_dataVec_1_35 : _GEN_713; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_715 = 6'h24 == f2_cut_ptr_4 ? f2_cut_data_dataVec_1_36 : _GEN_714; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_716 = 6'h25 == f2_cut_ptr_4 ? f2_cut_data_dataVec_1_37 : _GEN_715; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_717 = 6'h26 == f2_cut_ptr_4 ? f2_cut_data_dataVec_1_38 : _GEN_716; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_718 = 6'h27 == f2_cut_ptr_4 ? f2_cut_data_dataVec_1_39 : _GEN_717; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_719 = 6'h28 == f2_cut_ptr_4 ? f2_cut_data_dataVec_1_40 : _GEN_718; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_720 = 6'h29 == f2_cut_ptr_4 ? f2_cut_data_dataVec_1_41 : _GEN_719; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_721 = 6'h2a == f2_cut_ptr_4 ? f2_cut_data_dataVec_1_42 : _GEN_720; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_722 = 6'h2b == f2_cut_ptr_4 ? f2_cut_data_dataVec_1_43 : _GEN_721; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_723 = 6'h2c == f2_cut_ptr_4 ? f2_cut_data_dataVec_1_44 : _GEN_722; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_724 = 6'h2d == f2_cut_ptr_4 ? f2_cut_data_dataVec_1_45 : _GEN_723; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_725 = 6'h2e == f2_cut_ptr_4 ? f2_cut_data_dataVec_1_46 : _GEN_724; // @[IFU.scala 302:{19,19}]
  wire [15:0] f2_cut_data_result_1_4 = 6'h2f == f2_cut_ptr_4 ? f2_cut_data_dataVec_1_47 : _GEN_725; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_728 = 6'h1 == f2_cut_ptr_5 ? f2_cut_data_dataVec_1_1 : f2_cut_data_dataVec_1_0; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_729 = 6'h2 == f2_cut_ptr_5 ? f2_cut_data_dataVec_1_2 : _GEN_728; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_730 = 6'h3 == f2_cut_ptr_5 ? f2_cut_data_dataVec_1_3 : _GEN_729; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_731 = 6'h4 == f2_cut_ptr_5 ? f2_cut_data_dataVec_1_4 : _GEN_730; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_732 = 6'h5 == f2_cut_ptr_5 ? f2_cut_data_dataVec_1_5 : _GEN_731; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_733 = 6'h6 == f2_cut_ptr_5 ? f2_cut_data_dataVec_1_6 : _GEN_732; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_734 = 6'h7 == f2_cut_ptr_5 ? f2_cut_data_dataVec_1_7 : _GEN_733; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_735 = 6'h8 == f2_cut_ptr_5 ? f2_cut_data_dataVec_1_8 : _GEN_734; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_736 = 6'h9 == f2_cut_ptr_5 ? f2_cut_data_dataVec_1_9 : _GEN_735; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_737 = 6'ha == f2_cut_ptr_5 ? f2_cut_data_dataVec_1_10 : _GEN_736; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_738 = 6'hb == f2_cut_ptr_5 ? f2_cut_data_dataVec_1_11 : _GEN_737; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_739 = 6'hc == f2_cut_ptr_5 ? f2_cut_data_dataVec_1_12 : _GEN_738; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_740 = 6'hd == f2_cut_ptr_5 ? f2_cut_data_dataVec_1_13 : _GEN_739; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_741 = 6'he == f2_cut_ptr_5 ? f2_cut_data_dataVec_1_14 : _GEN_740; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_742 = 6'hf == f2_cut_ptr_5 ? f2_cut_data_dataVec_1_15 : _GEN_741; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_743 = 6'h10 == f2_cut_ptr_5 ? f2_cut_data_dataVec_1_16 : _GEN_742; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_744 = 6'h11 == f2_cut_ptr_5 ? f2_cut_data_dataVec_1_17 : _GEN_743; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_745 = 6'h12 == f2_cut_ptr_5 ? f2_cut_data_dataVec_1_18 : _GEN_744; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_746 = 6'h13 == f2_cut_ptr_5 ? f2_cut_data_dataVec_1_19 : _GEN_745; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_747 = 6'h14 == f2_cut_ptr_5 ? f2_cut_data_dataVec_1_20 : _GEN_746; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_748 = 6'h15 == f2_cut_ptr_5 ? f2_cut_data_dataVec_1_21 : _GEN_747; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_749 = 6'h16 == f2_cut_ptr_5 ? f2_cut_data_dataVec_1_22 : _GEN_748; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_750 = 6'h17 == f2_cut_ptr_5 ? f2_cut_data_dataVec_1_23 : _GEN_749; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_751 = 6'h18 == f2_cut_ptr_5 ? f2_cut_data_dataVec_1_24 : _GEN_750; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_752 = 6'h19 == f2_cut_ptr_5 ? f2_cut_data_dataVec_1_25 : _GEN_751; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_753 = 6'h1a == f2_cut_ptr_5 ? f2_cut_data_dataVec_1_26 : _GEN_752; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_754 = 6'h1b == f2_cut_ptr_5 ? f2_cut_data_dataVec_1_27 : _GEN_753; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_755 = 6'h1c == f2_cut_ptr_5 ? f2_cut_data_dataVec_1_28 : _GEN_754; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_756 = 6'h1d == f2_cut_ptr_5 ? f2_cut_data_dataVec_1_29 : _GEN_755; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_757 = 6'h1e == f2_cut_ptr_5 ? f2_cut_data_dataVec_1_30 : _GEN_756; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_758 = 6'h1f == f2_cut_ptr_5 ? f2_cut_data_dataVec_1_31 : _GEN_757; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_759 = 6'h20 == f2_cut_ptr_5 ? f2_cut_data_dataVec_1_32 : _GEN_758; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_760 = 6'h21 == f2_cut_ptr_5 ? f2_cut_data_dataVec_1_33 : _GEN_759; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_761 = 6'h22 == f2_cut_ptr_5 ? f2_cut_data_dataVec_1_34 : _GEN_760; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_762 = 6'h23 == f2_cut_ptr_5 ? f2_cut_data_dataVec_1_35 : _GEN_761; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_763 = 6'h24 == f2_cut_ptr_5 ? f2_cut_data_dataVec_1_36 : _GEN_762; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_764 = 6'h25 == f2_cut_ptr_5 ? f2_cut_data_dataVec_1_37 : _GEN_763; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_765 = 6'h26 == f2_cut_ptr_5 ? f2_cut_data_dataVec_1_38 : _GEN_764; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_766 = 6'h27 == f2_cut_ptr_5 ? f2_cut_data_dataVec_1_39 : _GEN_765; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_767 = 6'h28 == f2_cut_ptr_5 ? f2_cut_data_dataVec_1_40 : _GEN_766; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_768 = 6'h29 == f2_cut_ptr_5 ? f2_cut_data_dataVec_1_41 : _GEN_767; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_769 = 6'h2a == f2_cut_ptr_5 ? f2_cut_data_dataVec_1_42 : _GEN_768; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_770 = 6'h2b == f2_cut_ptr_5 ? f2_cut_data_dataVec_1_43 : _GEN_769; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_771 = 6'h2c == f2_cut_ptr_5 ? f2_cut_data_dataVec_1_44 : _GEN_770; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_772 = 6'h2d == f2_cut_ptr_5 ? f2_cut_data_dataVec_1_45 : _GEN_771; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_773 = 6'h2e == f2_cut_ptr_5 ? f2_cut_data_dataVec_1_46 : _GEN_772; // @[IFU.scala 302:{19,19}]
  wire [15:0] f2_cut_data_result_1_5 = 6'h2f == f2_cut_ptr_5 ? f2_cut_data_dataVec_1_47 : _GEN_773; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_776 = 6'h1 == f2_cut_ptr_6 ? f2_cut_data_dataVec_1_1 : f2_cut_data_dataVec_1_0; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_777 = 6'h2 == f2_cut_ptr_6 ? f2_cut_data_dataVec_1_2 : _GEN_776; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_778 = 6'h3 == f2_cut_ptr_6 ? f2_cut_data_dataVec_1_3 : _GEN_777; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_779 = 6'h4 == f2_cut_ptr_6 ? f2_cut_data_dataVec_1_4 : _GEN_778; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_780 = 6'h5 == f2_cut_ptr_6 ? f2_cut_data_dataVec_1_5 : _GEN_779; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_781 = 6'h6 == f2_cut_ptr_6 ? f2_cut_data_dataVec_1_6 : _GEN_780; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_782 = 6'h7 == f2_cut_ptr_6 ? f2_cut_data_dataVec_1_7 : _GEN_781; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_783 = 6'h8 == f2_cut_ptr_6 ? f2_cut_data_dataVec_1_8 : _GEN_782; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_784 = 6'h9 == f2_cut_ptr_6 ? f2_cut_data_dataVec_1_9 : _GEN_783; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_785 = 6'ha == f2_cut_ptr_6 ? f2_cut_data_dataVec_1_10 : _GEN_784; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_786 = 6'hb == f2_cut_ptr_6 ? f2_cut_data_dataVec_1_11 : _GEN_785; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_787 = 6'hc == f2_cut_ptr_6 ? f2_cut_data_dataVec_1_12 : _GEN_786; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_788 = 6'hd == f2_cut_ptr_6 ? f2_cut_data_dataVec_1_13 : _GEN_787; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_789 = 6'he == f2_cut_ptr_6 ? f2_cut_data_dataVec_1_14 : _GEN_788; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_790 = 6'hf == f2_cut_ptr_6 ? f2_cut_data_dataVec_1_15 : _GEN_789; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_791 = 6'h10 == f2_cut_ptr_6 ? f2_cut_data_dataVec_1_16 : _GEN_790; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_792 = 6'h11 == f2_cut_ptr_6 ? f2_cut_data_dataVec_1_17 : _GEN_791; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_793 = 6'h12 == f2_cut_ptr_6 ? f2_cut_data_dataVec_1_18 : _GEN_792; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_794 = 6'h13 == f2_cut_ptr_6 ? f2_cut_data_dataVec_1_19 : _GEN_793; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_795 = 6'h14 == f2_cut_ptr_6 ? f2_cut_data_dataVec_1_20 : _GEN_794; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_796 = 6'h15 == f2_cut_ptr_6 ? f2_cut_data_dataVec_1_21 : _GEN_795; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_797 = 6'h16 == f2_cut_ptr_6 ? f2_cut_data_dataVec_1_22 : _GEN_796; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_798 = 6'h17 == f2_cut_ptr_6 ? f2_cut_data_dataVec_1_23 : _GEN_797; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_799 = 6'h18 == f2_cut_ptr_6 ? f2_cut_data_dataVec_1_24 : _GEN_798; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_800 = 6'h19 == f2_cut_ptr_6 ? f2_cut_data_dataVec_1_25 : _GEN_799; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_801 = 6'h1a == f2_cut_ptr_6 ? f2_cut_data_dataVec_1_26 : _GEN_800; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_802 = 6'h1b == f2_cut_ptr_6 ? f2_cut_data_dataVec_1_27 : _GEN_801; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_803 = 6'h1c == f2_cut_ptr_6 ? f2_cut_data_dataVec_1_28 : _GEN_802; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_804 = 6'h1d == f2_cut_ptr_6 ? f2_cut_data_dataVec_1_29 : _GEN_803; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_805 = 6'h1e == f2_cut_ptr_6 ? f2_cut_data_dataVec_1_30 : _GEN_804; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_806 = 6'h1f == f2_cut_ptr_6 ? f2_cut_data_dataVec_1_31 : _GEN_805; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_807 = 6'h20 == f2_cut_ptr_6 ? f2_cut_data_dataVec_1_32 : _GEN_806; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_808 = 6'h21 == f2_cut_ptr_6 ? f2_cut_data_dataVec_1_33 : _GEN_807; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_809 = 6'h22 == f2_cut_ptr_6 ? f2_cut_data_dataVec_1_34 : _GEN_808; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_810 = 6'h23 == f2_cut_ptr_6 ? f2_cut_data_dataVec_1_35 : _GEN_809; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_811 = 6'h24 == f2_cut_ptr_6 ? f2_cut_data_dataVec_1_36 : _GEN_810; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_812 = 6'h25 == f2_cut_ptr_6 ? f2_cut_data_dataVec_1_37 : _GEN_811; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_813 = 6'h26 == f2_cut_ptr_6 ? f2_cut_data_dataVec_1_38 : _GEN_812; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_814 = 6'h27 == f2_cut_ptr_6 ? f2_cut_data_dataVec_1_39 : _GEN_813; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_815 = 6'h28 == f2_cut_ptr_6 ? f2_cut_data_dataVec_1_40 : _GEN_814; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_816 = 6'h29 == f2_cut_ptr_6 ? f2_cut_data_dataVec_1_41 : _GEN_815; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_817 = 6'h2a == f2_cut_ptr_6 ? f2_cut_data_dataVec_1_42 : _GEN_816; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_818 = 6'h2b == f2_cut_ptr_6 ? f2_cut_data_dataVec_1_43 : _GEN_817; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_819 = 6'h2c == f2_cut_ptr_6 ? f2_cut_data_dataVec_1_44 : _GEN_818; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_820 = 6'h2d == f2_cut_ptr_6 ? f2_cut_data_dataVec_1_45 : _GEN_819; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_821 = 6'h2e == f2_cut_ptr_6 ? f2_cut_data_dataVec_1_46 : _GEN_820; // @[IFU.scala 302:{19,19}]
  wire [15:0] f2_cut_data_result_1_6 = 6'h2f == f2_cut_ptr_6 ? f2_cut_data_dataVec_1_47 : _GEN_821; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_824 = 6'h1 == f2_cut_ptr_7 ? f2_cut_data_dataVec_1_1 : f2_cut_data_dataVec_1_0; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_825 = 6'h2 == f2_cut_ptr_7 ? f2_cut_data_dataVec_1_2 : _GEN_824; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_826 = 6'h3 == f2_cut_ptr_7 ? f2_cut_data_dataVec_1_3 : _GEN_825; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_827 = 6'h4 == f2_cut_ptr_7 ? f2_cut_data_dataVec_1_4 : _GEN_826; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_828 = 6'h5 == f2_cut_ptr_7 ? f2_cut_data_dataVec_1_5 : _GEN_827; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_829 = 6'h6 == f2_cut_ptr_7 ? f2_cut_data_dataVec_1_6 : _GEN_828; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_830 = 6'h7 == f2_cut_ptr_7 ? f2_cut_data_dataVec_1_7 : _GEN_829; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_831 = 6'h8 == f2_cut_ptr_7 ? f2_cut_data_dataVec_1_8 : _GEN_830; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_832 = 6'h9 == f2_cut_ptr_7 ? f2_cut_data_dataVec_1_9 : _GEN_831; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_833 = 6'ha == f2_cut_ptr_7 ? f2_cut_data_dataVec_1_10 : _GEN_832; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_834 = 6'hb == f2_cut_ptr_7 ? f2_cut_data_dataVec_1_11 : _GEN_833; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_835 = 6'hc == f2_cut_ptr_7 ? f2_cut_data_dataVec_1_12 : _GEN_834; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_836 = 6'hd == f2_cut_ptr_7 ? f2_cut_data_dataVec_1_13 : _GEN_835; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_837 = 6'he == f2_cut_ptr_7 ? f2_cut_data_dataVec_1_14 : _GEN_836; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_838 = 6'hf == f2_cut_ptr_7 ? f2_cut_data_dataVec_1_15 : _GEN_837; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_839 = 6'h10 == f2_cut_ptr_7 ? f2_cut_data_dataVec_1_16 : _GEN_838; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_840 = 6'h11 == f2_cut_ptr_7 ? f2_cut_data_dataVec_1_17 : _GEN_839; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_841 = 6'h12 == f2_cut_ptr_7 ? f2_cut_data_dataVec_1_18 : _GEN_840; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_842 = 6'h13 == f2_cut_ptr_7 ? f2_cut_data_dataVec_1_19 : _GEN_841; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_843 = 6'h14 == f2_cut_ptr_7 ? f2_cut_data_dataVec_1_20 : _GEN_842; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_844 = 6'h15 == f2_cut_ptr_7 ? f2_cut_data_dataVec_1_21 : _GEN_843; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_845 = 6'h16 == f2_cut_ptr_7 ? f2_cut_data_dataVec_1_22 : _GEN_844; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_846 = 6'h17 == f2_cut_ptr_7 ? f2_cut_data_dataVec_1_23 : _GEN_845; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_847 = 6'h18 == f2_cut_ptr_7 ? f2_cut_data_dataVec_1_24 : _GEN_846; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_848 = 6'h19 == f2_cut_ptr_7 ? f2_cut_data_dataVec_1_25 : _GEN_847; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_849 = 6'h1a == f2_cut_ptr_7 ? f2_cut_data_dataVec_1_26 : _GEN_848; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_850 = 6'h1b == f2_cut_ptr_7 ? f2_cut_data_dataVec_1_27 : _GEN_849; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_851 = 6'h1c == f2_cut_ptr_7 ? f2_cut_data_dataVec_1_28 : _GEN_850; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_852 = 6'h1d == f2_cut_ptr_7 ? f2_cut_data_dataVec_1_29 : _GEN_851; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_853 = 6'h1e == f2_cut_ptr_7 ? f2_cut_data_dataVec_1_30 : _GEN_852; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_854 = 6'h1f == f2_cut_ptr_7 ? f2_cut_data_dataVec_1_31 : _GEN_853; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_855 = 6'h20 == f2_cut_ptr_7 ? f2_cut_data_dataVec_1_32 : _GEN_854; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_856 = 6'h21 == f2_cut_ptr_7 ? f2_cut_data_dataVec_1_33 : _GEN_855; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_857 = 6'h22 == f2_cut_ptr_7 ? f2_cut_data_dataVec_1_34 : _GEN_856; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_858 = 6'h23 == f2_cut_ptr_7 ? f2_cut_data_dataVec_1_35 : _GEN_857; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_859 = 6'h24 == f2_cut_ptr_7 ? f2_cut_data_dataVec_1_36 : _GEN_858; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_860 = 6'h25 == f2_cut_ptr_7 ? f2_cut_data_dataVec_1_37 : _GEN_859; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_861 = 6'h26 == f2_cut_ptr_7 ? f2_cut_data_dataVec_1_38 : _GEN_860; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_862 = 6'h27 == f2_cut_ptr_7 ? f2_cut_data_dataVec_1_39 : _GEN_861; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_863 = 6'h28 == f2_cut_ptr_7 ? f2_cut_data_dataVec_1_40 : _GEN_862; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_864 = 6'h29 == f2_cut_ptr_7 ? f2_cut_data_dataVec_1_41 : _GEN_863; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_865 = 6'h2a == f2_cut_ptr_7 ? f2_cut_data_dataVec_1_42 : _GEN_864; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_866 = 6'h2b == f2_cut_ptr_7 ? f2_cut_data_dataVec_1_43 : _GEN_865; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_867 = 6'h2c == f2_cut_ptr_7 ? f2_cut_data_dataVec_1_44 : _GEN_866; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_868 = 6'h2d == f2_cut_ptr_7 ? f2_cut_data_dataVec_1_45 : _GEN_867; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_869 = 6'h2e == f2_cut_ptr_7 ? f2_cut_data_dataVec_1_46 : _GEN_868; // @[IFU.scala 302:{19,19}]
  wire [15:0] f2_cut_data_result_1_7 = 6'h2f == f2_cut_ptr_7 ? f2_cut_data_dataVec_1_47 : _GEN_869; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_872 = 6'h1 == f2_cut_ptr_8 ? f2_cut_data_dataVec_1_1 : f2_cut_data_dataVec_1_0; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_873 = 6'h2 == f2_cut_ptr_8 ? f2_cut_data_dataVec_1_2 : _GEN_872; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_874 = 6'h3 == f2_cut_ptr_8 ? f2_cut_data_dataVec_1_3 : _GEN_873; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_875 = 6'h4 == f2_cut_ptr_8 ? f2_cut_data_dataVec_1_4 : _GEN_874; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_876 = 6'h5 == f2_cut_ptr_8 ? f2_cut_data_dataVec_1_5 : _GEN_875; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_877 = 6'h6 == f2_cut_ptr_8 ? f2_cut_data_dataVec_1_6 : _GEN_876; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_878 = 6'h7 == f2_cut_ptr_8 ? f2_cut_data_dataVec_1_7 : _GEN_877; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_879 = 6'h8 == f2_cut_ptr_8 ? f2_cut_data_dataVec_1_8 : _GEN_878; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_880 = 6'h9 == f2_cut_ptr_8 ? f2_cut_data_dataVec_1_9 : _GEN_879; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_881 = 6'ha == f2_cut_ptr_8 ? f2_cut_data_dataVec_1_10 : _GEN_880; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_882 = 6'hb == f2_cut_ptr_8 ? f2_cut_data_dataVec_1_11 : _GEN_881; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_883 = 6'hc == f2_cut_ptr_8 ? f2_cut_data_dataVec_1_12 : _GEN_882; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_884 = 6'hd == f2_cut_ptr_8 ? f2_cut_data_dataVec_1_13 : _GEN_883; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_885 = 6'he == f2_cut_ptr_8 ? f2_cut_data_dataVec_1_14 : _GEN_884; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_886 = 6'hf == f2_cut_ptr_8 ? f2_cut_data_dataVec_1_15 : _GEN_885; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_887 = 6'h10 == f2_cut_ptr_8 ? f2_cut_data_dataVec_1_16 : _GEN_886; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_888 = 6'h11 == f2_cut_ptr_8 ? f2_cut_data_dataVec_1_17 : _GEN_887; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_889 = 6'h12 == f2_cut_ptr_8 ? f2_cut_data_dataVec_1_18 : _GEN_888; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_890 = 6'h13 == f2_cut_ptr_8 ? f2_cut_data_dataVec_1_19 : _GEN_889; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_891 = 6'h14 == f2_cut_ptr_8 ? f2_cut_data_dataVec_1_20 : _GEN_890; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_892 = 6'h15 == f2_cut_ptr_8 ? f2_cut_data_dataVec_1_21 : _GEN_891; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_893 = 6'h16 == f2_cut_ptr_8 ? f2_cut_data_dataVec_1_22 : _GEN_892; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_894 = 6'h17 == f2_cut_ptr_8 ? f2_cut_data_dataVec_1_23 : _GEN_893; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_895 = 6'h18 == f2_cut_ptr_8 ? f2_cut_data_dataVec_1_24 : _GEN_894; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_896 = 6'h19 == f2_cut_ptr_8 ? f2_cut_data_dataVec_1_25 : _GEN_895; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_897 = 6'h1a == f2_cut_ptr_8 ? f2_cut_data_dataVec_1_26 : _GEN_896; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_898 = 6'h1b == f2_cut_ptr_8 ? f2_cut_data_dataVec_1_27 : _GEN_897; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_899 = 6'h1c == f2_cut_ptr_8 ? f2_cut_data_dataVec_1_28 : _GEN_898; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_900 = 6'h1d == f2_cut_ptr_8 ? f2_cut_data_dataVec_1_29 : _GEN_899; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_901 = 6'h1e == f2_cut_ptr_8 ? f2_cut_data_dataVec_1_30 : _GEN_900; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_902 = 6'h1f == f2_cut_ptr_8 ? f2_cut_data_dataVec_1_31 : _GEN_901; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_903 = 6'h20 == f2_cut_ptr_8 ? f2_cut_data_dataVec_1_32 : _GEN_902; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_904 = 6'h21 == f2_cut_ptr_8 ? f2_cut_data_dataVec_1_33 : _GEN_903; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_905 = 6'h22 == f2_cut_ptr_8 ? f2_cut_data_dataVec_1_34 : _GEN_904; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_906 = 6'h23 == f2_cut_ptr_8 ? f2_cut_data_dataVec_1_35 : _GEN_905; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_907 = 6'h24 == f2_cut_ptr_8 ? f2_cut_data_dataVec_1_36 : _GEN_906; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_908 = 6'h25 == f2_cut_ptr_8 ? f2_cut_data_dataVec_1_37 : _GEN_907; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_909 = 6'h26 == f2_cut_ptr_8 ? f2_cut_data_dataVec_1_38 : _GEN_908; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_910 = 6'h27 == f2_cut_ptr_8 ? f2_cut_data_dataVec_1_39 : _GEN_909; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_911 = 6'h28 == f2_cut_ptr_8 ? f2_cut_data_dataVec_1_40 : _GEN_910; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_912 = 6'h29 == f2_cut_ptr_8 ? f2_cut_data_dataVec_1_41 : _GEN_911; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_913 = 6'h2a == f2_cut_ptr_8 ? f2_cut_data_dataVec_1_42 : _GEN_912; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_914 = 6'h2b == f2_cut_ptr_8 ? f2_cut_data_dataVec_1_43 : _GEN_913; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_915 = 6'h2c == f2_cut_ptr_8 ? f2_cut_data_dataVec_1_44 : _GEN_914; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_916 = 6'h2d == f2_cut_ptr_8 ? f2_cut_data_dataVec_1_45 : _GEN_915; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_917 = 6'h2e == f2_cut_ptr_8 ? f2_cut_data_dataVec_1_46 : _GEN_916; // @[IFU.scala 302:{19,19}]
  wire [15:0] f2_cut_data_result_1_8 = 6'h2f == f2_cut_ptr_8 ? f2_cut_data_dataVec_1_47 : _GEN_917; // @[IFU.scala 302:{19,19}]
  wire [767:0] f2_cut_data_partCacheline_2 = f2_data_2_cacheline_2[767:0]; // @[IFU.scala 298:36]
  wire [15:0] f2_cut_data_dataVec_2_0 = f2_cut_data_partCacheline_2[15:0]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_2_1 = f2_cut_data_partCacheline_2[31:16]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_2_2 = f2_cut_data_partCacheline_2[47:32]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_2_3 = f2_cut_data_partCacheline_2[63:48]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_2_4 = f2_cut_data_partCacheline_2[79:64]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_2_5 = f2_cut_data_partCacheline_2[95:80]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_2_6 = f2_cut_data_partCacheline_2[111:96]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_2_7 = f2_cut_data_partCacheline_2[127:112]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_2_8 = f2_cut_data_partCacheline_2[143:128]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_2_9 = f2_cut_data_partCacheline_2[159:144]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_2_10 = f2_cut_data_partCacheline_2[175:160]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_2_11 = f2_cut_data_partCacheline_2[191:176]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_2_12 = f2_cut_data_partCacheline_2[207:192]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_2_13 = f2_cut_data_partCacheline_2[223:208]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_2_14 = f2_cut_data_partCacheline_2[239:224]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_2_15 = f2_cut_data_partCacheline_2[255:240]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_2_16 = f2_cut_data_partCacheline_2[271:256]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_2_17 = f2_cut_data_partCacheline_2[287:272]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_2_18 = f2_cut_data_partCacheline_2[303:288]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_2_19 = f2_cut_data_partCacheline_2[319:304]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_2_20 = f2_cut_data_partCacheline_2[335:320]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_2_21 = f2_cut_data_partCacheline_2[351:336]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_2_22 = f2_cut_data_partCacheline_2[367:352]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_2_23 = f2_cut_data_partCacheline_2[383:368]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_2_24 = f2_cut_data_partCacheline_2[399:384]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_2_25 = f2_cut_data_partCacheline_2[415:400]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_2_26 = f2_cut_data_partCacheline_2[431:416]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_2_27 = f2_cut_data_partCacheline_2[447:432]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_2_28 = f2_cut_data_partCacheline_2[463:448]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_2_29 = f2_cut_data_partCacheline_2[479:464]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_2_30 = f2_cut_data_partCacheline_2[495:480]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_2_31 = f2_cut_data_partCacheline_2[511:496]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_2_32 = f2_cut_data_partCacheline_2[527:512]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_2_33 = f2_cut_data_partCacheline_2[543:528]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_2_34 = f2_cut_data_partCacheline_2[559:544]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_2_35 = f2_cut_data_partCacheline_2[575:560]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_2_36 = f2_cut_data_partCacheline_2[591:576]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_2_37 = f2_cut_data_partCacheline_2[607:592]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_2_38 = f2_cut_data_partCacheline_2[623:608]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_2_39 = f2_cut_data_partCacheline_2[639:624]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_2_40 = f2_cut_data_partCacheline_2[655:640]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_2_41 = f2_cut_data_partCacheline_2[671:656]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_2_42 = f2_cut_data_partCacheline_2[687:672]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_2_43 = f2_cut_data_partCacheline_2[703:688]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_2_44 = f2_cut_data_partCacheline_2[719:704]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_2_45 = f2_cut_data_partCacheline_2[735:720]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_2_46 = f2_cut_data_partCacheline_2[751:736]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_2_47 = f2_cut_data_partCacheline_2[767:752]; // @[IFU.scala 300:40]
  wire [15:0] _GEN_920 = 6'h1 == f2_cut_ptr_0 ? f2_cut_data_dataVec_2_1 : f2_cut_data_dataVec_2_0; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_921 = 6'h2 == f2_cut_ptr_0 ? f2_cut_data_dataVec_2_2 : _GEN_920; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_922 = 6'h3 == f2_cut_ptr_0 ? f2_cut_data_dataVec_2_3 : _GEN_921; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_923 = 6'h4 == f2_cut_ptr_0 ? f2_cut_data_dataVec_2_4 : _GEN_922; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_924 = 6'h5 == f2_cut_ptr_0 ? f2_cut_data_dataVec_2_5 : _GEN_923; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_925 = 6'h6 == f2_cut_ptr_0 ? f2_cut_data_dataVec_2_6 : _GEN_924; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_926 = 6'h7 == f2_cut_ptr_0 ? f2_cut_data_dataVec_2_7 : _GEN_925; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_927 = 6'h8 == f2_cut_ptr_0 ? f2_cut_data_dataVec_2_8 : _GEN_926; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_928 = 6'h9 == f2_cut_ptr_0 ? f2_cut_data_dataVec_2_9 : _GEN_927; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_929 = 6'ha == f2_cut_ptr_0 ? f2_cut_data_dataVec_2_10 : _GEN_928; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_930 = 6'hb == f2_cut_ptr_0 ? f2_cut_data_dataVec_2_11 : _GEN_929; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_931 = 6'hc == f2_cut_ptr_0 ? f2_cut_data_dataVec_2_12 : _GEN_930; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_932 = 6'hd == f2_cut_ptr_0 ? f2_cut_data_dataVec_2_13 : _GEN_931; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_933 = 6'he == f2_cut_ptr_0 ? f2_cut_data_dataVec_2_14 : _GEN_932; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_934 = 6'hf == f2_cut_ptr_0 ? f2_cut_data_dataVec_2_15 : _GEN_933; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_935 = 6'h10 == f2_cut_ptr_0 ? f2_cut_data_dataVec_2_16 : _GEN_934; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_936 = 6'h11 == f2_cut_ptr_0 ? f2_cut_data_dataVec_2_17 : _GEN_935; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_937 = 6'h12 == f2_cut_ptr_0 ? f2_cut_data_dataVec_2_18 : _GEN_936; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_938 = 6'h13 == f2_cut_ptr_0 ? f2_cut_data_dataVec_2_19 : _GEN_937; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_939 = 6'h14 == f2_cut_ptr_0 ? f2_cut_data_dataVec_2_20 : _GEN_938; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_940 = 6'h15 == f2_cut_ptr_0 ? f2_cut_data_dataVec_2_21 : _GEN_939; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_941 = 6'h16 == f2_cut_ptr_0 ? f2_cut_data_dataVec_2_22 : _GEN_940; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_942 = 6'h17 == f2_cut_ptr_0 ? f2_cut_data_dataVec_2_23 : _GEN_941; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_943 = 6'h18 == f2_cut_ptr_0 ? f2_cut_data_dataVec_2_24 : _GEN_942; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_944 = 6'h19 == f2_cut_ptr_0 ? f2_cut_data_dataVec_2_25 : _GEN_943; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_945 = 6'h1a == f2_cut_ptr_0 ? f2_cut_data_dataVec_2_26 : _GEN_944; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_946 = 6'h1b == f2_cut_ptr_0 ? f2_cut_data_dataVec_2_27 : _GEN_945; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_947 = 6'h1c == f2_cut_ptr_0 ? f2_cut_data_dataVec_2_28 : _GEN_946; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_948 = 6'h1d == f2_cut_ptr_0 ? f2_cut_data_dataVec_2_29 : _GEN_947; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_949 = 6'h1e == f2_cut_ptr_0 ? f2_cut_data_dataVec_2_30 : _GEN_948; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_950 = 6'h1f == f2_cut_ptr_0 ? f2_cut_data_dataVec_2_31 : _GEN_949; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_951 = 6'h20 == f2_cut_ptr_0 ? f2_cut_data_dataVec_2_32 : _GEN_950; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_952 = 6'h21 == f2_cut_ptr_0 ? f2_cut_data_dataVec_2_33 : _GEN_951; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_953 = 6'h22 == f2_cut_ptr_0 ? f2_cut_data_dataVec_2_34 : _GEN_952; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_954 = 6'h23 == f2_cut_ptr_0 ? f2_cut_data_dataVec_2_35 : _GEN_953; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_955 = 6'h24 == f2_cut_ptr_0 ? f2_cut_data_dataVec_2_36 : _GEN_954; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_956 = 6'h25 == f2_cut_ptr_0 ? f2_cut_data_dataVec_2_37 : _GEN_955; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_957 = 6'h26 == f2_cut_ptr_0 ? f2_cut_data_dataVec_2_38 : _GEN_956; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_958 = 6'h27 == f2_cut_ptr_0 ? f2_cut_data_dataVec_2_39 : _GEN_957; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_959 = 6'h28 == f2_cut_ptr_0 ? f2_cut_data_dataVec_2_40 : _GEN_958; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_960 = 6'h29 == f2_cut_ptr_0 ? f2_cut_data_dataVec_2_41 : _GEN_959; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_961 = 6'h2a == f2_cut_ptr_0 ? f2_cut_data_dataVec_2_42 : _GEN_960; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_962 = 6'h2b == f2_cut_ptr_0 ? f2_cut_data_dataVec_2_43 : _GEN_961; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_963 = 6'h2c == f2_cut_ptr_0 ? f2_cut_data_dataVec_2_44 : _GEN_962; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_964 = 6'h2d == f2_cut_ptr_0 ? f2_cut_data_dataVec_2_45 : _GEN_963; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_965 = 6'h2e == f2_cut_ptr_0 ? f2_cut_data_dataVec_2_46 : _GEN_964; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_968 = 6'h1 == f2_cut_ptr_1 ? f2_cut_data_dataVec_2_1 : f2_cut_data_dataVec_2_0; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_969 = 6'h2 == f2_cut_ptr_1 ? f2_cut_data_dataVec_2_2 : _GEN_968; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_970 = 6'h3 == f2_cut_ptr_1 ? f2_cut_data_dataVec_2_3 : _GEN_969; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_971 = 6'h4 == f2_cut_ptr_1 ? f2_cut_data_dataVec_2_4 : _GEN_970; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_972 = 6'h5 == f2_cut_ptr_1 ? f2_cut_data_dataVec_2_5 : _GEN_971; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_973 = 6'h6 == f2_cut_ptr_1 ? f2_cut_data_dataVec_2_6 : _GEN_972; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_974 = 6'h7 == f2_cut_ptr_1 ? f2_cut_data_dataVec_2_7 : _GEN_973; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_975 = 6'h8 == f2_cut_ptr_1 ? f2_cut_data_dataVec_2_8 : _GEN_974; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_976 = 6'h9 == f2_cut_ptr_1 ? f2_cut_data_dataVec_2_9 : _GEN_975; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_977 = 6'ha == f2_cut_ptr_1 ? f2_cut_data_dataVec_2_10 : _GEN_976; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_978 = 6'hb == f2_cut_ptr_1 ? f2_cut_data_dataVec_2_11 : _GEN_977; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_979 = 6'hc == f2_cut_ptr_1 ? f2_cut_data_dataVec_2_12 : _GEN_978; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_980 = 6'hd == f2_cut_ptr_1 ? f2_cut_data_dataVec_2_13 : _GEN_979; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_981 = 6'he == f2_cut_ptr_1 ? f2_cut_data_dataVec_2_14 : _GEN_980; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_982 = 6'hf == f2_cut_ptr_1 ? f2_cut_data_dataVec_2_15 : _GEN_981; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_983 = 6'h10 == f2_cut_ptr_1 ? f2_cut_data_dataVec_2_16 : _GEN_982; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_984 = 6'h11 == f2_cut_ptr_1 ? f2_cut_data_dataVec_2_17 : _GEN_983; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_985 = 6'h12 == f2_cut_ptr_1 ? f2_cut_data_dataVec_2_18 : _GEN_984; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_986 = 6'h13 == f2_cut_ptr_1 ? f2_cut_data_dataVec_2_19 : _GEN_985; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_987 = 6'h14 == f2_cut_ptr_1 ? f2_cut_data_dataVec_2_20 : _GEN_986; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_988 = 6'h15 == f2_cut_ptr_1 ? f2_cut_data_dataVec_2_21 : _GEN_987; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_989 = 6'h16 == f2_cut_ptr_1 ? f2_cut_data_dataVec_2_22 : _GEN_988; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_990 = 6'h17 == f2_cut_ptr_1 ? f2_cut_data_dataVec_2_23 : _GEN_989; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_991 = 6'h18 == f2_cut_ptr_1 ? f2_cut_data_dataVec_2_24 : _GEN_990; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_992 = 6'h19 == f2_cut_ptr_1 ? f2_cut_data_dataVec_2_25 : _GEN_991; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_993 = 6'h1a == f2_cut_ptr_1 ? f2_cut_data_dataVec_2_26 : _GEN_992; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_994 = 6'h1b == f2_cut_ptr_1 ? f2_cut_data_dataVec_2_27 : _GEN_993; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_995 = 6'h1c == f2_cut_ptr_1 ? f2_cut_data_dataVec_2_28 : _GEN_994; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_996 = 6'h1d == f2_cut_ptr_1 ? f2_cut_data_dataVec_2_29 : _GEN_995; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_997 = 6'h1e == f2_cut_ptr_1 ? f2_cut_data_dataVec_2_30 : _GEN_996; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_998 = 6'h1f == f2_cut_ptr_1 ? f2_cut_data_dataVec_2_31 : _GEN_997; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_999 = 6'h20 == f2_cut_ptr_1 ? f2_cut_data_dataVec_2_32 : _GEN_998; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1000 = 6'h21 == f2_cut_ptr_1 ? f2_cut_data_dataVec_2_33 : _GEN_999; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1001 = 6'h22 == f2_cut_ptr_1 ? f2_cut_data_dataVec_2_34 : _GEN_1000; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1002 = 6'h23 == f2_cut_ptr_1 ? f2_cut_data_dataVec_2_35 : _GEN_1001; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1003 = 6'h24 == f2_cut_ptr_1 ? f2_cut_data_dataVec_2_36 : _GEN_1002; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1004 = 6'h25 == f2_cut_ptr_1 ? f2_cut_data_dataVec_2_37 : _GEN_1003; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1005 = 6'h26 == f2_cut_ptr_1 ? f2_cut_data_dataVec_2_38 : _GEN_1004; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1006 = 6'h27 == f2_cut_ptr_1 ? f2_cut_data_dataVec_2_39 : _GEN_1005; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1007 = 6'h28 == f2_cut_ptr_1 ? f2_cut_data_dataVec_2_40 : _GEN_1006; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1008 = 6'h29 == f2_cut_ptr_1 ? f2_cut_data_dataVec_2_41 : _GEN_1007; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1009 = 6'h2a == f2_cut_ptr_1 ? f2_cut_data_dataVec_2_42 : _GEN_1008; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1010 = 6'h2b == f2_cut_ptr_1 ? f2_cut_data_dataVec_2_43 : _GEN_1009; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1011 = 6'h2c == f2_cut_ptr_1 ? f2_cut_data_dataVec_2_44 : _GEN_1010; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1012 = 6'h2d == f2_cut_ptr_1 ? f2_cut_data_dataVec_2_45 : _GEN_1011; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1013 = 6'h2e == f2_cut_ptr_1 ? f2_cut_data_dataVec_2_46 : _GEN_1012; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1016 = 6'h1 == f2_cut_ptr_2 ? f2_cut_data_dataVec_2_1 : f2_cut_data_dataVec_2_0; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1017 = 6'h2 == f2_cut_ptr_2 ? f2_cut_data_dataVec_2_2 : _GEN_1016; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1018 = 6'h3 == f2_cut_ptr_2 ? f2_cut_data_dataVec_2_3 : _GEN_1017; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1019 = 6'h4 == f2_cut_ptr_2 ? f2_cut_data_dataVec_2_4 : _GEN_1018; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1020 = 6'h5 == f2_cut_ptr_2 ? f2_cut_data_dataVec_2_5 : _GEN_1019; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1021 = 6'h6 == f2_cut_ptr_2 ? f2_cut_data_dataVec_2_6 : _GEN_1020; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1022 = 6'h7 == f2_cut_ptr_2 ? f2_cut_data_dataVec_2_7 : _GEN_1021; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1023 = 6'h8 == f2_cut_ptr_2 ? f2_cut_data_dataVec_2_8 : _GEN_1022; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1024 = 6'h9 == f2_cut_ptr_2 ? f2_cut_data_dataVec_2_9 : _GEN_1023; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1025 = 6'ha == f2_cut_ptr_2 ? f2_cut_data_dataVec_2_10 : _GEN_1024; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1026 = 6'hb == f2_cut_ptr_2 ? f2_cut_data_dataVec_2_11 : _GEN_1025; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1027 = 6'hc == f2_cut_ptr_2 ? f2_cut_data_dataVec_2_12 : _GEN_1026; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1028 = 6'hd == f2_cut_ptr_2 ? f2_cut_data_dataVec_2_13 : _GEN_1027; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1029 = 6'he == f2_cut_ptr_2 ? f2_cut_data_dataVec_2_14 : _GEN_1028; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1030 = 6'hf == f2_cut_ptr_2 ? f2_cut_data_dataVec_2_15 : _GEN_1029; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1031 = 6'h10 == f2_cut_ptr_2 ? f2_cut_data_dataVec_2_16 : _GEN_1030; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1032 = 6'h11 == f2_cut_ptr_2 ? f2_cut_data_dataVec_2_17 : _GEN_1031; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1033 = 6'h12 == f2_cut_ptr_2 ? f2_cut_data_dataVec_2_18 : _GEN_1032; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1034 = 6'h13 == f2_cut_ptr_2 ? f2_cut_data_dataVec_2_19 : _GEN_1033; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1035 = 6'h14 == f2_cut_ptr_2 ? f2_cut_data_dataVec_2_20 : _GEN_1034; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1036 = 6'h15 == f2_cut_ptr_2 ? f2_cut_data_dataVec_2_21 : _GEN_1035; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1037 = 6'h16 == f2_cut_ptr_2 ? f2_cut_data_dataVec_2_22 : _GEN_1036; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1038 = 6'h17 == f2_cut_ptr_2 ? f2_cut_data_dataVec_2_23 : _GEN_1037; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1039 = 6'h18 == f2_cut_ptr_2 ? f2_cut_data_dataVec_2_24 : _GEN_1038; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1040 = 6'h19 == f2_cut_ptr_2 ? f2_cut_data_dataVec_2_25 : _GEN_1039; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1041 = 6'h1a == f2_cut_ptr_2 ? f2_cut_data_dataVec_2_26 : _GEN_1040; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1042 = 6'h1b == f2_cut_ptr_2 ? f2_cut_data_dataVec_2_27 : _GEN_1041; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1043 = 6'h1c == f2_cut_ptr_2 ? f2_cut_data_dataVec_2_28 : _GEN_1042; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1044 = 6'h1d == f2_cut_ptr_2 ? f2_cut_data_dataVec_2_29 : _GEN_1043; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1045 = 6'h1e == f2_cut_ptr_2 ? f2_cut_data_dataVec_2_30 : _GEN_1044; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1046 = 6'h1f == f2_cut_ptr_2 ? f2_cut_data_dataVec_2_31 : _GEN_1045; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1047 = 6'h20 == f2_cut_ptr_2 ? f2_cut_data_dataVec_2_32 : _GEN_1046; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1048 = 6'h21 == f2_cut_ptr_2 ? f2_cut_data_dataVec_2_33 : _GEN_1047; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1049 = 6'h22 == f2_cut_ptr_2 ? f2_cut_data_dataVec_2_34 : _GEN_1048; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1050 = 6'h23 == f2_cut_ptr_2 ? f2_cut_data_dataVec_2_35 : _GEN_1049; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1051 = 6'h24 == f2_cut_ptr_2 ? f2_cut_data_dataVec_2_36 : _GEN_1050; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1052 = 6'h25 == f2_cut_ptr_2 ? f2_cut_data_dataVec_2_37 : _GEN_1051; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1053 = 6'h26 == f2_cut_ptr_2 ? f2_cut_data_dataVec_2_38 : _GEN_1052; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1054 = 6'h27 == f2_cut_ptr_2 ? f2_cut_data_dataVec_2_39 : _GEN_1053; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1055 = 6'h28 == f2_cut_ptr_2 ? f2_cut_data_dataVec_2_40 : _GEN_1054; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1056 = 6'h29 == f2_cut_ptr_2 ? f2_cut_data_dataVec_2_41 : _GEN_1055; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1057 = 6'h2a == f2_cut_ptr_2 ? f2_cut_data_dataVec_2_42 : _GEN_1056; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1058 = 6'h2b == f2_cut_ptr_2 ? f2_cut_data_dataVec_2_43 : _GEN_1057; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1059 = 6'h2c == f2_cut_ptr_2 ? f2_cut_data_dataVec_2_44 : _GEN_1058; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1060 = 6'h2d == f2_cut_ptr_2 ? f2_cut_data_dataVec_2_45 : _GEN_1059; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1061 = 6'h2e == f2_cut_ptr_2 ? f2_cut_data_dataVec_2_46 : _GEN_1060; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1064 = 6'h1 == f2_cut_ptr_3 ? f2_cut_data_dataVec_2_1 : f2_cut_data_dataVec_2_0; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1065 = 6'h2 == f2_cut_ptr_3 ? f2_cut_data_dataVec_2_2 : _GEN_1064; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1066 = 6'h3 == f2_cut_ptr_3 ? f2_cut_data_dataVec_2_3 : _GEN_1065; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1067 = 6'h4 == f2_cut_ptr_3 ? f2_cut_data_dataVec_2_4 : _GEN_1066; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1068 = 6'h5 == f2_cut_ptr_3 ? f2_cut_data_dataVec_2_5 : _GEN_1067; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1069 = 6'h6 == f2_cut_ptr_3 ? f2_cut_data_dataVec_2_6 : _GEN_1068; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1070 = 6'h7 == f2_cut_ptr_3 ? f2_cut_data_dataVec_2_7 : _GEN_1069; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1071 = 6'h8 == f2_cut_ptr_3 ? f2_cut_data_dataVec_2_8 : _GEN_1070; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1072 = 6'h9 == f2_cut_ptr_3 ? f2_cut_data_dataVec_2_9 : _GEN_1071; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1073 = 6'ha == f2_cut_ptr_3 ? f2_cut_data_dataVec_2_10 : _GEN_1072; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1074 = 6'hb == f2_cut_ptr_3 ? f2_cut_data_dataVec_2_11 : _GEN_1073; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1075 = 6'hc == f2_cut_ptr_3 ? f2_cut_data_dataVec_2_12 : _GEN_1074; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1076 = 6'hd == f2_cut_ptr_3 ? f2_cut_data_dataVec_2_13 : _GEN_1075; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1077 = 6'he == f2_cut_ptr_3 ? f2_cut_data_dataVec_2_14 : _GEN_1076; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1078 = 6'hf == f2_cut_ptr_3 ? f2_cut_data_dataVec_2_15 : _GEN_1077; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1079 = 6'h10 == f2_cut_ptr_3 ? f2_cut_data_dataVec_2_16 : _GEN_1078; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1080 = 6'h11 == f2_cut_ptr_3 ? f2_cut_data_dataVec_2_17 : _GEN_1079; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1081 = 6'h12 == f2_cut_ptr_3 ? f2_cut_data_dataVec_2_18 : _GEN_1080; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1082 = 6'h13 == f2_cut_ptr_3 ? f2_cut_data_dataVec_2_19 : _GEN_1081; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1083 = 6'h14 == f2_cut_ptr_3 ? f2_cut_data_dataVec_2_20 : _GEN_1082; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1084 = 6'h15 == f2_cut_ptr_3 ? f2_cut_data_dataVec_2_21 : _GEN_1083; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1085 = 6'h16 == f2_cut_ptr_3 ? f2_cut_data_dataVec_2_22 : _GEN_1084; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1086 = 6'h17 == f2_cut_ptr_3 ? f2_cut_data_dataVec_2_23 : _GEN_1085; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1087 = 6'h18 == f2_cut_ptr_3 ? f2_cut_data_dataVec_2_24 : _GEN_1086; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1088 = 6'h19 == f2_cut_ptr_3 ? f2_cut_data_dataVec_2_25 : _GEN_1087; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1089 = 6'h1a == f2_cut_ptr_3 ? f2_cut_data_dataVec_2_26 : _GEN_1088; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1090 = 6'h1b == f2_cut_ptr_3 ? f2_cut_data_dataVec_2_27 : _GEN_1089; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1091 = 6'h1c == f2_cut_ptr_3 ? f2_cut_data_dataVec_2_28 : _GEN_1090; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1092 = 6'h1d == f2_cut_ptr_3 ? f2_cut_data_dataVec_2_29 : _GEN_1091; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1093 = 6'h1e == f2_cut_ptr_3 ? f2_cut_data_dataVec_2_30 : _GEN_1092; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1094 = 6'h1f == f2_cut_ptr_3 ? f2_cut_data_dataVec_2_31 : _GEN_1093; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1095 = 6'h20 == f2_cut_ptr_3 ? f2_cut_data_dataVec_2_32 : _GEN_1094; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1096 = 6'h21 == f2_cut_ptr_3 ? f2_cut_data_dataVec_2_33 : _GEN_1095; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1097 = 6'h22 == f2_cut_ptr_3 ? f2_cut_data_dataVec_2_34 : _GEN_1096; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1098 = 6'h23 == f2_cut_ptr_3 ? f2_cut_data_dataVec_2_35 : _GEN_1097; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1099 = 6'h24 == f2_cut_ptr_3 ? f2_cut_data_dataVec_2_36 : _GEN_1098; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1100 = 6'h25 == f2_cut_ptr_3 ? f2_cut_data_dataVec_2_37 : _GEN_1099; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1101 = 6'h26 == f2_cut_ptr_3 ? f2_cut_data_dataVec_2_38 : _GEN_1100; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1102 = 6'h27 == f2_cut_ptr_3 ? f2_cut_data_dataVec_2_39 : _GEN_1101; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1103 = 6'h28 == f2_cut_ptr_3 ? f2_cut_data_dataVec_2_40 : _GEN_1102; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1104 = 6'h29 == f2_cut_ptr_3 ? f2_cut_data_dataVec_2_41 : _GEN_1103; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1105 = 6'h2a == f2_cut_ptr_3 ? f2_cut_data_dataVec_2_42 : _GEN_1104; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1106 = 6'h2b == f2_cut_ptr_3 ? f2_cut_data_dataVec_2_43 : _GEN_1105; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1107 = 6'h2c == f2_cut_ptr_3 ? f2_cut_data_dataVec_2_44 : _GEN_1106; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1108 = 6'h2d == f2_cut_ptr_3 ? f2_cut_data_dataVec_2_45 : _GEN_1107; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1109 = 6'h2e == f2_cut_ptr_3 ? f2_cut_data_dataVec_2_46 : _GEN_1108; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1112 = 6'h1 == f2_cut_ptr_4 ? f2_cut_data_dataVec_2_1 : f2_cut_data_dataVec_2_0; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1113 = 6'h2 == f2_cut_ptr_4 ? f2_cut_data_dataVec_2_2 : _GEN_1112; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1114 = 6'h3 == f2_cut_ptr_4 ? f2_cut_data_dataVec_2_3 : _GEN_1113; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1115 = 6'h4 == f2_cut_ptr_4 ? f2_cut_data_dataVec_2_4 : _GEN_1114; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1116 = 6'h5 == f2_cut_ptr_4 ? f2_cut_data_dataVec_2_5 : _GEN_1115; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1117 = 6'h6 == f2_cut_ptr_4 ? f2_cut_data_dataVec_2_6 : _GEN_1116; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1118 = 6'h7 == f2_cut_ptr_4 ? f2_cut_data_dataVec_2_7 : _GEN_1117; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1119 = 6'h8 == f2_cut_ptr_4 ? f2_cut_data_dataVec_2_8 : _GEN_1118; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1120 = 6'h9 == f2_cut_ptr_4 ? f2_cut_data_dataVec_2_9 : _GEN_1119; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1121 = 6'ha == f2_cut_ptr_4 ? f2_cut_data_dataVec_2_10 : _GEN_1120; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1122 = 6'hb == f2_cut_ptr_4 ? f2_cut_data_dataVec_2_11 : _GEN_1121; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1123 = 6'hc == f2_cut_ptr_4 ? f2_cut_data_dataVec_2_12 : _GEN_1122; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1124 = 6'hd == f2_cut_ptr_4 ? f2_cut_data_dataVec_2_13 : _GEN_1123; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1125 = 6'he == f2_cut_ptr_4 ? f2_cut_data_dataVec_2_14 : _GEN_1124; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1126 = 6'hf == f2_cut_ptr_4 ? f2_cut_data_dataVec_2_15 : _GEN_1125; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1127 = 6'h10 == f2_cut_ptr_4 ? f2_cut_data_dataVec_2_16 : _GEN_1126; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1128 = 6'h11 == f2_cut_ptr_4 ? f2_cut_data_dataVec_2_17 : _GEN_1127; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1129 = 6'h12 == f2_cut_ptr_4 ? f2_cut_data_dataVec_2_18 : _GEN_1128; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1130 = 6'h13 == f2_cut_ptr_4 ? f2_cut_data_dataVec_2_19 : _GEN_1129; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1131 = 6'h14 == f2_cut_ptr_4 ? f2_cut_data_dataVec_2_20 : _GEN_1130; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1132 = 6'h15 == f2_cut_ptr_4 ? f2_cut_data_dataVec_2_21 : _GEN_1131; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1133 = 6'h16 == f2_cut_ptr_4 ? f2_cut_data_dataVec_2_22 : _GEN_1132; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1134 = 6'h17 == f2_cut_ptr_4 ? f2_cut_data_dataVec_2_23 : _GEN_1133; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1135 = 6'h18 == f2_cut_ptr_4 ? f2_cut_data_dataVec_2_24 : _GEN_1134; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1136 = 6'h19 == f2_cut_ptr_4 ? f2_cut_data_dataVec_2_25 : _GEN_1135; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1137 = 6'h1a == f2_cut_ptr_4 ? f2_cut_data_dataVec_2_26 : _GEN_1136; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1138 = 6'h1b == f2_cut_ptr_4 ? f2_cut_data_dataVec_2_27 : _GEN_1137; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1139 = 6'h1c == f2_cut_ptr_4 ? f2_cut_data_dataVec_2_28 : _GEN_1138; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1140 = 6'h1d == f2_cut_ptr_4 ? f2_cut_data_dataVec_2_29 : _GEN_1139; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1141 = 6'h1e == f2_cut_ptr_4 ? f2_cut_data_dataVec_2_30 : _GEN_1140; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1142 = 6'h1f == f2_cut_ptr_4 ? f2_cut_data_dataVec_2_31 : _GEN_1141; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1143 = 6'h20 == f2_cut_ptr_4 ? f2_cut_data_dataVec_2_32 : _GEN_1142; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1144 = 6'h21 == f2_cut_ptr_4 ? f2_cut_data_dataVec_2_33 : _GEN_1143; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1145 = 6'h22 == f2_cut_ptr_4 ? f2_cut_data_dataVec_2_34 : _GEN_1144; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1146 = 6'h23 == f2_cut_ptr_4 ? f2_cut_data_dataVec_2_35 : _GEN_1145; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1147 = 6'h24 == f2_cut_ptr_4 ? f2_cut_data_dataVec_2_36 : _GEN_1146; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1148 = 6'h25 == f2_cut_ptr_4 ? f2_cut_data_dataVec_2_37 : _GEN_1147; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1149 = 6'h26 == f2_cut_ptr_4 ? f2_cut_data_dataVec_2_38 : _GEN_1148; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1150 = 6'h27 == f2_cut_ptr_4 ? f2_cut_data_dataVec_2_39 : _GEN_1149; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1151 = 6'h28 == f2_cut_ptr_4 ? f2_cut_data_dataVec_2_40 : _GEN_1150; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1152 = 6'h29 == f2_cut_ptr_4 ? f2_cut_data_dataVec_2_41 : _GEN_1151; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1153 = 6'h2a == f2_cut_ptr_4 ? f2_cut_data_dataVec_2_42 : _GEN_1152; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1154 = 6'h2b == f2_cut_ptr_4 ? f2_cut_data_dataVec_2_43 : _GEN_1153; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1155 = 6'h2c == f2_cut_ptr_4 ? f2_cut_data_dataVec_2_44 : _GEN_1154; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1156 = 6'h2d == f2_cut_ptr_4 ? f2_cut_data_dataVec_2_45 : _GEN_1155; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1157 = 6'h2e == f2_cut_ptr_4 ? f2_cut_data_dataVec_2_46 : _GEN_1156; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1160 = 6'h1 == f2_cut_ptr_5 ? f2_cut_data_dataVec_2_1 : f2_cut_data_dataVec_2_0; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1161 = 6'h2 == f2_cut_ptr_5 ? f2_cut_data_dataVec_2_2 : _GEN_1160; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1162 = 6'h3 == f2_cut_ptr_5 ? f2_cut_data_dataVec_2_3 : _GEN_1161; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1163 = 6'h4 == f2_cut_ptr_5 ? f2_cut_data_dataVec_2_4 : _GEN_1162; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1164 = 6'h5 == f2_cut_ptr_5 ? f2_cut_data_dataVec_2_5 : _GEN_1163; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1165 = 6'h6 == f2_cut_ptr_5 ? f2_cut_data_dataVec_2_6 : _GEN_1164; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1166 = 6'h7 == f2_cut_ptr_5 ? f2_cut_data_dataVec_2_7 : _GEN_1165; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1167 = 6'h8 == f2_cut_ptr_5 ? f2_cut_data_dataVec_2_8 : _GEN_1166; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1168 = 6'h9 == f2_cut_ptr_5 ? f2_cut_data_dataVec_2_9 : _GEN_1167; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1169 = 6'ha == f2_cut_ptr_5 ? f2_cut_data_dataVec_2_10 : _GEN_1168; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1170 = 6'hb == f2_cut_ptr_5 ? f2_cut_data_dataVec_2_11 : _GEN_1169; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1171 = 6'hc == f2_cut_ptr_5 ? f2_cut_data_dataVec_2_12 : _GEN_1170; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1172 = 6'hd == f2_cut_ptr_5 ? f2_cut_data_dataVec_2_13 : _GEN_1171; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1173 = 6'he == f2_cut_ptr_5 ? f2_cut_data_dataVec_2_14 : _GEN_1172; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1174 = 6'hf == f2_cut_ptr_5 ? f2_cut_data_dataVec_2_15 : _GEN_1173; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1175 = 6'h10 == f2_cut_ptr_5 ? f2_cut_data_dataVec_2_16 : _GEN_1174; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1176 = 6'h11 == f2_cut_ptr_5 ? f2_cut_data_dataVec_2_17 : _GEN_1175; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1177 = 6'h12 == f2_cut_ptr_5 ? f2_cut_data_dataVec_2_18 : _GEN_1176; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1178 = 6'h13 == f2_cut_ptr_5 ? f2_cut_data_dataVec_2_19 : _GEN_1177; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1179 = 6'h14 == f2_cut_ptr_5 ? f2_cut_data_dataVec_2_20 : _GEN_1178; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1180 = 6'h15 == f2_cut_ptr_5 ? f2_cut_data_dataVec_2_21 : _GEN_1179; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1181 = 6'h16 == f2_cut_ptr_5 ? f2_cut_data_dataVec_2_22 : _GEN_1180; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1182 = 6'h17 == f2_cut_ptr_5 ? f2_cut_data_dataVec_2_23 : _GEN_1181; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1183 = 6'h18 == f2_cut_ptr_5 ? f2_cut_data_dataVec_2_24 : _GEN_1182; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1184 = 6'h19 == f2_cut_ptr_5 ? f2_cut_data_dataVec_2_25 : _GEN_1183; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1185 = 6'h1a == f2_cut_ptr_5 ? f2_cut_data_dataVec_2_26 : _GEN_1184; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1186 = 6'h1b == f2_cut_ptr_5 ? f2_cut_data_dataVec_2_27 : _GEN_1185; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1187 = 6'h1c == f2_cut_ptr_5 ? f2_cut_data_dataVec_2_28 : _GEN_1186; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1188 = 6'h1d == f2_cut_ptr_5 ? f2_cut_data_dataVec_2_29 : _GEN_1187; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1189 = 6'h1e == f2_cut_ptr_5 ? f2_cut_data_dataVec_2_30 : _GEN_1188; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1190 = 6'h1f == f2_cut_ptr_5 ? f2_cut_data_dataVec_2_31 : _GEN_1189; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1191 = 6'h20 == f2_cut_ptr_5 ? f2_cut_data_dataVec_2_32 : _GEN_1190; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1192 = 6'h21 == f2_cut_ptr_5 ? f2_cut_data_dataVec_2_33 : _GEN_1191; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1193 = 6'h22 == f2_cut_ptr_5 ? f2_cut_data_dataVec_2_34 : _GEN_1192; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1194 = 6'h23 == f2_cut_ptr_5 ? f2_cut_data_dataVec_2_35 : _GEN_1193; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1195 = 6'h24 == f2_cut_ptr_5 ? f2_cut_data_dataVec_2_36 : _GEN_1194; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1196 = 6'h25 == f2_cut_ptr_5 ? f2_cut_data_dataVec_2_37 : _GEN_1195; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1197 = 6'h26 == f2_cut_ptr_5 ? f2_cut_data_dataVec_2_38 : _GEN_1196; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1198 = 6'h27 == f2_cut_ptr_5 ? f2_cut_data_dataVec_2_39 : _GEN_1197; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1199 = 6'h28 == f2_cut_ptr_5 ? f2_cut_data_dataVec_2_40 : _GEN_1198; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1200 = 6'h29 == f2_cut_ptr_5 ? f2_cut_data_dataVec_2_41 : _GEN_1199; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1201 = 6'h2a == f2_cut_ptr_5 ? f2_cut_data_dataVec_2_42 : _GEN_1200; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1202 = 6'h2b == f2_cut_ptr_5 ? f2_cut_data_dataVec_2_43 : _GEN_1201; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1203 = 6'h2c == f2_cut_ptr_5 ? f2_cut_data_dataVec_2_44 : _GEN_1202; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1204 = 6'h2d == f2_cut_ptr_5 ? f2_cut_data_dataVec_2_45 : _GEN_1203; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1205 = 6'h2e == f2_cut_ptr_5 ? f2_cut_data_dataVec_2_46 : _GEN_1204; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1208 = 6'h1 == f2_cut_ptr_6 ? f2_cut_data_dataVec_2_1 : f2_cut_data_dataVec_2_0; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1209 = 6'h2 == f2_cut_ptr_6 ? f2_cut_data_dataVec_2_2 : _GEN_1208; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1210 = 6'h3 == f2_cut_ptr_6 ? f2_cut_data_dataVec_2_3 : _GEN_1209; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1211 = 6'h4 == f2_cut_ptr_6 ? f2_cut_data_dataVec_2_4 : _GEN_1210; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1212 = 6'h5 == f2_cut_ptr_6 ? f2_cut_data_dataVec_2_5 : _GEN_1211; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1213 = 6'h6 == f2_cut_ptr_6 ? f2_cut_data_dataVec_2_6 : _GEN_1212; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1214 = 6'h7 == f2_cut_ptr_6 ? f2_cut_data_dataVec_2_7 : _GEN_1213; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1215 = 6'h8 == f2_cut_ptr_6 ? f2_cut_data_dataVec_2_8 : _GEN_1214; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1216 = 6'h9 == f2_cut_ptr_6 ? f2_cut_data_dataVec_2_9 : _GEN_1215; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1217 = 6'ha == f2_cut_ptr_6 ? f2_cut_data_dataVec_2_10 : _GEN_1216; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1218 = 6'hb == f2_cut_ptr_6 ? f2_cut_data_dataVec_2_11 : _GEN_1217; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1219 = 6'hc == f2_cut_ptr_6 ? f2_cut_data_dataVec_2_12 : _GEN_1218; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1220 = 6'hd == f2_cut_ptr_6 ? f2_cut_data_dataVec_2_13 : _GEN_1219; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1221 = 6'he == f2_cut_ptr_6 ? f2_cut_data_dataVec_2_14 : _GEN_1220; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1222 = 6'hf == f2_cut_ptr_6 ? f2_cut_data_dataVec_2_15 : _GEN_1221; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1223 = 6'h10 == f2_cut_ptr_6 ? f2_cut_data_dataVec_2_16 : _GEN_1222; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1224 = 6'h11 == f2_cut_ptr_6 ? f2_cut_data_dataVec_2_17 : _GEN_1223; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1225 = 6'h12 == f2_cut_ptr_6 ? f2_cut_data_dataVec_2_18 : _GEN_1224; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1226 = 6'h13 == f2_cut_ptr_6 ? f2_cut_data_dataVec_2_19 : _GEN_1225; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1227 = 6'h14 == f2_cut_ptr_6 ? f2_cut_data_dataVec_2_20 : _GEN_1226; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1228 = 6'h15 == f2_cut_ptr_6 ? f2_cut_data_dataVec_2_21 : _GEN_1227; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1229 = 6'h16 == f2_cut_ptr_6 ? f2_cut_data_dataVec_2_22 : _GEN_1228; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1230 = 6'h17 == f2_cut_ptr_6 ? f2_cut_data_dataVec_2_23 : _GEN_1229; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1231 = 6'h18 == f2_cut_ptr_6 ? f2_cut_data_dataVec_2_24 : _GEN_1230; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1232 = 6'h19 == f2_cut_ptr_6 ? f2_cut_data_dataVec_2_25 : _GEN_1231; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1233 = 6'h1a == f2_cut_ptr_6 ? f2_cut_data_dataVec_2_26 : _GEN_1232; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1234 = 6'h1b == f2_cut_ptr_6 ? f2_cut_data_dataVec_2_27 : _GEN_1233; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1235 = 6'h1c == f2_cut_ptr_6 ? f2_cut_data_dataVec_2_28 : _GEN_1234; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1236 = 6'h1d == f2_cut_ptr_6 ? f2_cut_data_dataVec_2_29 : _GEN_1235; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1237 = 6'h1e == f2_cut_ptr_6 ? f2_cut_data_dataVec_2_30 : _GEN_1236; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1238 = 6'h1f == f2_cut_ptr_6 ? f2_cut_data_dataVec_2_31 : _GEN_1237; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1239 = 6'h20 == f2_cut_ptr_6 ? f2_cut_data_dataVec_2_32 : _GEN_1238; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1240 = 6'h21 == f2_cut_ptr_6 ? f2_cut_data_dataVec_2_33 : _GEN_1239; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1241 = 6'h22 == f2_cut_ptr_6 ? f2_cut_data_dataVec_2_34 : _GEN_1240; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1242 = 6'h23 == f2_cut_ptr_6 ? f2_cut_data_dataVec_2_35 : _GEN_1241; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1243 = 6'h24 == f2_cut_ptr_6 ? f2_cut_data_dataVec_2_36 : _GEN_1242; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1244 = 6'h25 == f2_cut_ptr_6 ? f2_cut_data_dataVec_2_37 : _GEN_1243; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1245 = 6'h26 == f2_cut_ptr_6 ? f2_cut_data_dataVec_2_38 : _GEN_1244; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1246 = 6'h27 == f2_cut_ptr_6 ? f2_cut_data_dataVec_2_39 : _GEN_1245; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1247 = 6'h28 == f2_cut_ptr_6 ? f2_cut_data_dataVec_2_40 : _GEN_1246; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1248 = 6'h29 == f2_cut_ptr_6 ? f2_cut_data_dataVec_2_41 : _GEN_1247; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1249 = 6'h2a == f2_cut_ptr_6 ? f2_cut_data_dataVec_2_42 : _GEN_1248; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1250 = 6'h2b == f2_cut_ptr_6 ? f2_cut_data_dataVec_2_43 : _GEN_1249; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1251 = 6'h2c == f2_cut_ptr_6 ? f2_cut_data_dataVec_2_44 : _GEN_1250; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1252 = 6'h2d == f2_cut_ptr_6 ? f2_cut_data_dataVec_2_45 : _GEN_1251; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1253 = 6'h2e == f2_cut_ptr_6 ? f2_cut_data_dataVec_2_46 : _GEN_1252; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1256 = 6'h1 == f2_cut_ptr_7 ? f2_cut_data_dataVec_2_1 : f2_cut_data_dataVec_2_0; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1257 = 6'h2 == f2_cut_ptr_7 ? f2_cut_data_dataVec_2_2 : _GEN_1256; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1258 = 6'h3 == f2_cut_ptr_7 ? f2_cut_data_dataVec_2_3 : _GEN_1257; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1259 = 6'h4 == f2_cut_ptr_7 ? f2_cut_data_dataVec_2_4 : _GEN_1258; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1260 = 6'h5 == f2_cut_ptr_7 ? f2_cut_data_dataVec_2_5 : _GEN_1259; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1261 = 6'h6 == f2_cut_ptr_7 ? f2_cut_data_dataVec_2_6 : _GEN_1260; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1262 = 6'h7 == f2_cut_ptr_7 ? f2_cut_data_dataVec_2_7 : _GEN_1261; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1263 = 6'h8 == f2_cut_ptr_7 ? f2_cut_data_dataVec_2_8 : _GEN_1262; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1264 = 6'h9 == f2_cut_ptr_7 ? f2_cut_data_dataVec_2_9 : _GEN_1263; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1265 = 6'ha == f2_cut_ptr_7 ? f2_cut_data_dataVec_2_10 : _GEN_1264; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1266 = 6'hb == f2_cut_ptr_7 ? f2_cut_data_dataVec_2_11 : _GEN_1265; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1267 = 6'hc == f2_cut_ptr_7 ? f2_cut_data_dataVec_2_12 : _GEN_1266; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1268 = 6'hd == f2_cut_ptr_7 ? f2_cut_data_dataVec_2_13 : _GEN_1267; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1269 = 6'he == f2_cut_ptr_7 ? f2_cut_data_dataVec_2_14 : _GEN_1268; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1270 = 6'hf == f2_cut_ptr_7 ? f2_cut_data_dataVec_2_15 : _GEN_1269; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1271 = 6'h10 == f2_cut_ptr_7 ? f2_cut_data_dataVec_2_16 : _GEN_1270; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1272 = 6'h11 == f2_cut_ptr_7 ? f2_cut_data_dataVec_2_17 : _GEN_1271; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1273 = 6'h12 == f2_cut_ptr_7 ? f2_cut_data_dataVec_2_18 : _GEN_1272; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1274 = 6'h13 == f2_cut_ptr_7 ? f2_cut_data_dataVec_2_19 : _GEN_1273; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1275 = 6'h14 == f2_cut_ptr_7 ? f2_cut_data_dataVec_2_20 : _GEN_1274; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1276 = 6'h15 == f2_cut_ptr_7 ? f2_cut_data_dataVec_2_21 : _GEN_1275; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1277 = 6'h16 == f2_cut_ptr_7 ? f2_cut_data_dataVec_2_22 : _GEN_1276; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1278 = 6'h17 == f2_cut_ptr_7 ? f2_cut_data_dataVec_2_23 : _GEN_1277; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1279 = 6'h18 == f2_cut_ptr_7 ? f2_cut_data_dataVec_2_24 : _GEN_1278; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1280 = 6'h19 == f2_cut_ptr_7 ? f2_cut_data_dataVec_2_25 : _GEN_1279; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1281 = 6'h1a == f2_cut_ptr_7 ? f2_cut_data_dataVec_2_26 : _GEN_1280; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1282 = 6'h1b == f2_cut_ptr_7 ? f2_cut_data_dataVec_2_27 : _GEN_1281; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1283 = 6'h1c == f2_cut_ptr_7 ? f2_cut_data_dataVec_2_28 : _GEN_1282; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1284 = 6'h1d == f2_cut_ptr_7 ? f2_cut_data_dataVec_2_29 : _GEN_1283; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1285 = 6'h1e == f2_cut_ptr_7 ? f2_cut_data_dataVec_2_30 : _GEN_1284; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1286 = 6'h1f == f2_cut_ptr_7 ? f2_cut_data_dataVec_2_31 : _GEN_1285; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1287 = 6'h20 == f2_cut_ptr_7 ? f2_cut_data_dataVec_2_32 : _GEN_1286; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1288 = 6'h21 == f2_cut_ptr_7 ? f2_cut_data_dataVec_2_33 : _GEN_1287; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1289 = 6'h22 == f2_cut_ptr_7 ? f2_cut_data_dataVec_2_34 : _GEN_1288; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1290 = 6'h23 == f2_cut_ptr_7 ? f2_cut_data_dataVec_2_35 : _GEN_1289; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1291 = 6'h24 == f2_cut_ptr_7 ? f2_cut_data_dataVec_2_36 : _GEN_1290; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1292 = 6'h25 == f2_cut_ptr_7 ? f2_cut_data_dataVec_2_37 : _GEN_1291; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1293 = 6'h26 == f2_cut_ptr_7 ? f2_cut_data_dataVec_2_38 : _GEN_1292; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1294 = 6'h27 == f2_cut_ptr_7 ? f2_cut_data_dataVec_2_39 : _GEN_1293; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1295 = 6'h28 == f2_cut_ptr_7 ? f2_cut_data_dataVec_2_40 : _GEN_1294; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1296 = 6'h29 == f2_cut_ptr_7 ? f2_cut_data_dataVec_2_41 : _GEN_1295; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1297 = 6'h2a == f2_cut_ptr_7 ? f2_cut_data_dataVec_2_42 : _GEN_1296; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1298 = 6'h2b == f2_cut_ptr_7 ? f2_cut_data_dataVec_2_43 : _GEN_1297; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1299 = 6'h2c == f2_cut_ptr_7 ? f2_cut_data_dataVec_2_44 : _GEN_1298; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1300 = 6'h2d == f2_cut_ptr_7 ? f2_cut_data_dataVec_2_45 : _GEN_1299; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1301 = 6'h2e == f2_cut_ptr_7 ? f2_cut_data_dataVec_2_46 : _GEN_1300; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1304 = 6'h1 == f2_cut_ptr_8 ? f2_cut_data_dataVec_2_1 : f2_cut_data_dataVec_2_0; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1305 = 6'h2 == f2_cut_ptr_8 ? f2_cut_data_dataVec_2_2 : _GEN_1304; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1306 = 6'h3 == f2_cut_ptr_8 ? f2_cut_data_dataVec_2_3 : _GEN_1305; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1307 = 6'h4 == f2_cut_ptr_8 ? f2_cut_data_dataVec_2_4 : _GEN_1306; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1308 = 6'h5 == f2_cut_ptr_8 ? f2_cut_data_dataVec_2_5 : _GEN_1307; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1309 = 6'h6 == f2_cut_ptr_8 ? f2_cut_data_dataVec_2_6 : _GEN_1308; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1310 = 6'h7 == f2_cut_ptr_8 ? f2_cut_data_dataVec_2_7 : _GEN_1309; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1311 = 6'h8 == f2_cut_ptr_8 ? f2_cut_data_dataVec_2_8 : _GEN_1310; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1312 = 6'h9 == f2_cut_ptr_8 ? f2_cut_data_dataVec_2_9 : _GEN_1311; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1313 = 6'ha == f2_cut_ptr_8 ? f2_cut_data_dataVec_2_10 : _GEN_1312; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1314 = 6'hb == f2_cut_ptr_8 ? f2_cut_data_dataVec_2_11 : _GEN_1313; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1315 = 6'hc == f2_cut_ptr_8 ? f2_cut_data_dataVec_2_12 : _GEN_1314; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1316 = 6'hd == f2_cut_ptr_8 ? f2_cut_data_dataVec_2_13 : _GEN_1315; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1317 = 6'he == f2_cut_ptr_8 ? f2_cut_data_dataVec_2_14 : _GEN_1316; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1318 = 6'hf == f2_cut_ptr_8 ? f2_cut_data_dataVec_2_15 : _GEN_1317; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1319 = 6'h10 == f2_cut_ptr_8 ? f2_cut_data_dataVec_2_16 : _GEN_1318; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1320 = 6'h11 == f2_cut_ptr_8 ? f2_cut_data_dataVec_2_17 : _GEN_1319; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1321 = 6'h12 == f2_cut_ptr_8 ? f2_cut_data_dataVec_2_18 : _GEN_1320; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1322 = 6'h13 == f2_cut_ptr_8 ? f2_cut_data_dataVec_2_19 : _GEN_1321; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1323 = 6'h14 == f2_cut_ptr_8 ? f2_cut_data_dataVec_2_20 : _GEN_1322; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1324 = 6'h15 == f2_cut_ptr_8 ? f2_cut_data_dataVec_2_21 : _GEN_1323; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1325 = 6'h16 == f2_cut_ptr_8 ? f2_cut_data_dataVec_2_22 : _GEN_1324; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1326 = 6'h17 == f2_cut_ptr_8 ? f2_cut_data_dataVec_2_23 : _GEN_1325; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1327 = 6'h18 == f2_cut_ptr_8 ? f2_cut_data_dataVec_2_24 : _GEN_1326; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1328 = 6'h19 == f2_cut_ptr_8 ? f2_cut_data_dataVec_2_25 : _GEN_1327; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1329 = 6'h1a == f2_cut_ptr_8 ? f2_cut_data_dataVec_2_26 : _GEN_1328; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1330 = 6'h1b == f2_cut_ptr_8 ? f2_cut_data_dataVec_2_27 : _GEN_1329; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1331 = 6'h1c == f2_cut_ptr_8 ? f2_cut_data_dataVec_2_28 : _GEN_1330; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1332 = 6'h1d == f2_cut_ptr_8 ? f2_cut_data_dataVec_2_29 : _GEN_1331; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1333 = 6'h1e == f2_cut_ptr_8 ? f2_cut_data_dataVec_2_30 : _GEN_1332; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1334 = 6'h1f == f2_cut_ptr_8 ? f2_cut_data_dataVec_2_31 : _GEN_1333; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1335 = 6'h20 == f2_cut_ptr_8 ? f2_cut_data_dataVec_2_32 : _GEN_1334; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1336 = 6'h21 == f2_cut_ptr_8 ? f2_cut_data_dataVec_2_33 : _GEN_1335; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1337 = 6'h22 == f2_cut_ptr_8 ? f2_cut_data_dataVec_2_34 : _GEN_1336; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1338 = 6'h23 == f2_cut_ptr_8 ? f2_cut_data_dataVec_2_35 : _GEN_1337; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1339 = 6'h24 == f2_cut_ptr_8 ? f2_cut_data_dataVec_2_36 : _GEN_1338; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1340 = 6'h25 == f2_cut_ptr_8 ? f2_cut_data_dataVec_2_37 : _GEN_1339; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1341 = 6'h26 == f2_cut_ptr_8 ? f2_cut_data_dataVec_2_38 : _GEN_1340; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1342 = 6'h27 == f2_cut_ptr_8 ? f2_cut_data_dataVec_2_39 : _GEN_1341; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1343 = 6'h28 == f2_cut_ptr_8 ? f2_cut_data_dataVec_2_40 : _GEN_1342; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1344 = 6'h29 == f2_cut_ptr_8 ? f2_cut_data_dataVec_2_41 : _GEN_1343; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1345 = 6'h2a == f2_cut_ptr_8 ? f2_cut_data_dataVec_2_42 : _GEN_1344; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1346 = 6'h2b == f2_cut_ptr_8 ? f2_cut_data_dataVec_2_43 : _GEN_1345; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1347 = 6'h2c == f2_cut_ptr_8 ? f2_cut_data_dataVec_2_44 : _GEN_1346; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1348 = 6'h2d == f2_cut_ptr_8 ? f2_cut_data_dataVec_2_45 : _GEN_1347; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1349 = 6'h2e == f2_cut_ptr_8 ? f2_cut_data_dataVec_2_46 : _GEN_1348; // @[IFU.scala 302:{19,19}]
  wire [767:0] f2_cut_data_partCacheline_3 = f2_data_2_cacheline_3[767:0]; // @[IFU.scala 298:36]
  wire [15:0] f2_cut_data_dataVec_3_0 = f2_cut_data_partCacheline_3[15:0]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_3_1 = f2_cut_data_partCacheline_3[31:16]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_3_2 = f2_cut_data_partCacheline_3[47:32]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_3_3 = f2_cut_data_partCacheline_3[63:48]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_3_4 = f2_cut_data_partCacheline_3[79:64]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_3_5 = f2_cut_data_partCacheline_3[95:80]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_3_6 = f2_cut_data_partCacheline_3[111:96]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_3_7 = f2_cut_data_partCacheline_3[127:112]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_3_8 = f2_cut_data_partCacheline_3[143:128]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_3_9 = f2_cut_data_partCacheline_3[159:144]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_3_10 = f2_cut_data_partCacheline_3[175:160]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_3_11 = f2_cut_data_partCacheline_3[191:176]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_3_12 = f2_cut_data_partCacheline_3[207:192]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_3_13 = f2_cut_data_partCacheline_3[223:208]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_3_14 = f2_cut_data_partCacheline_3[239:224]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_3_15 = f2_cut_data_partCacheline_3[255:240]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_3_16 = f2_cut_data_partCacheline_3[271:256]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_3_17 = f2_cut_data_partCacheline_3[287:272]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_3_18 = f2_cut_data_partCacheline_3[303:288]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_3_19 = f2_cut_data_partCacheline_3[319:304]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_3_20 = f2_cut_data_partCacheline_3[335:320]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_3_21 = f2_cut_data_partCacheline_3[351:336]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_3_22 = f2_cut_data_partCacheline_3[367:352]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_3_23 = f2_cut_data_partCacheline_3[383:368]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_3_24 = f2_cut_data_partCacheline_3[399:384]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_3_25 = f2_cut_data_partCacheline_3[415:400]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_3_26 = f2_cut_data_partCacheline_3[431:416]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_3_27 = f2_cut_data_partCacheline_3[447:432]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_3_28 = f2_cut_data_partCacheline_3[463:448]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_3_29 = f2_cut_data_partCacheline_3[479:464]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_3_30 = f2_cut_data_partCacheline_3[495:480]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_3_31 = f2_cut_data_partCacheline_3[511:496]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_3_32 = f2_cut_data_partCacheline_3[527:512]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_3_33 = f2_cut_data_partCacheline_3[543:528]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_3_34 = f2_cut_data_partCacheline_3[559:544]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_3_35 = f2_cut_data_partCacheline_3[575:560]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_3_36 = f2_cut_data_partCacheline_3[591:576]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_3_37 = f2_cut_data_partCacheline_3[607:592]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_3_38 = f2_cut_data_partCacheline_3[623:608]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_3_39 = f2_cut_data_partCacheline_3[639:624]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_3_40 = f2_cut_data_partCacheline_3[655:640]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_3_41 = f2_cut_data_partCacheline_3[671:656]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_3_42 = f2_cut_data_partCacheline_3[687:672]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_3_43 = f2_cut_data_partCacheline_3[703:688]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_3_44 = f2_cut_data_partCacheline_3[719:704]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_3_45 = f2_cut_data_partCacheline_3[735:720]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_3_46 = f2_cut_data_partCacheline_3[751:736]; // @[IFU.scala 300:40]
  wire [15:0] f2_cut_data_dataVec_3_47 = f2_cut_data_partCacheline_3[767:752]; // @[IFU.scala 300:40]
  wire [15:0] _GEN_1352 = 6'h1 == f2_cut_ptr_0 ? f2_cut_data_dataVec_3_1 : f2_cut_data_dataVec_3_0; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1353 = 6'h2 == f2_cut_ptr_0 ? f2_cut_data_dataVec_3_2 : _GEN_1352; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1354 = 6'h3 == f2_cut_ptr_0 ? f2_cut_data_dataVec_3_3 : _GEN_1353; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1355 = 6'h4 == f2_cut_ptr_0 ? f2_cut_data_dataVec_3_4 : _GEN_1354; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1356 = 6'h5 == f2_cut_ptr_0 ? f2_cut_data_dataVec_3_5 : _GEN_1355; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1357 = 6'h6 == f2_cut_ptr_0 ? f2_cut_data_dataVec_3_6 : _GEN_1356; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1358 = 6'h7 == f2_cut_ptr_0 ? f2_cut_data_dataVec_3_7 : _GEN_1357; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1359 = 6'h8 == f2_cut_ptr_0 ? f2_cut_data_dataVec_3_8 : _GEN_1358; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1360 = 6'h9 == f2_cut_ptr_0 ? f2_cut_data_dataVec_3_9 : _GEN_1359; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1361 = 6'ha == f2_cut_ptr_0 ? f2_cut_data_dataVec_3_10 : _GEN_1360; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1362 = 6'hb == f2_cut_ptr_0 ? f2_cut_data_dataVec_3_11 : _GEN_1361; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1363 = 6'hc == f2_cut_ptr_0 ? f2_cut_data_dataVec_3_12 : _GEN_1362; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1364 = 6'hd == f2_cut_ptr_0 ? f2_cut_data_dataVec_3_13 : _GEN_1363; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1365 = 6'he == f2_cut_ptr_0 ? f2_cut_data_dataVec_3_14 : _GEN_1364; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1366 = 6'hf == f2_cut_ptr_0 ? f2_cut_data_dataVec_3_15 : _GEN_1365; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1367 = 6'h10 == f2_cut_ptr_0 ? f2_cut_data_dataVec_3_16 : _GEN_1366; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1368 = 6'h11 == f2_cut_ptr_0 ? f2_cut_data_dataVec_3_17 : _GEN_1367; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1369 = 6'h12 == f2_cut_ptr_0 ? f2_cut_data_dataVec_3_18 : _GEN_1368; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1370 = 6'h13 == f2_cut_ptr_0 ? f2_cut_data_dataVec_3_19 : _GEN_1369; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1371 = 6'h14 == f2_cut_ptr_0 ? f2_cut_data_dataVec_3_20 : _GEN_1370; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1372 = 6'h15 == f2_cut_ptr_0 ? f2_cut_data_dataVec_3_21 : _GEN_1371; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1373 = 6'h16 == f2_cut_ptr_0 ? f2_cut_data_dataVec_3_22 : _GEN_1372; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1374 = 6'h17 == f2_cut_ptr_0 ? f2_cut_data_dataVec_3_23 : _GEN_1373; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1375 = 6'h18 == f2_cut_ptr_0 ? f2_cut_data_dataVec_3_24 : _GEN_1374; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1376 = 6'h19 == f2_cut_ptr_0 ? f2_cut_data_dataVec_3_25 : _GEN_1375; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1377 = 6'h1a == f2_cut_ptr_0 ? f2_cut_data_dataVec_3_26 : _GEN_1376; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1378 = 6'h1b == f2_cut_ptr_0 ? f2_cut_data_dataVec_3_27 : _GEN_1377; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1379 = 6'h1c == f2_cut_ptr_0 ? f2_cut_data_dataVec_3_28 : _GEN_1378; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1380 = 6'h1d == f2_cut_ptr_0 ? f2_cut_data_dataVec_3_29 : _GEN_1379; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1381 = 6'h1e == f2_cut_ptr_0 ? f2_cut_data_dataVec_3_30 : _GEN_1380; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1382 = 6'h1f == f2_cut_ptr_0 ? f2_cut_data_dataVec_3_31 : _GEN_1381; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1383 = 6'h20 == f2_cut_ptr_0 ? f2_cut_data_dataVec_3_32 : _GEN_1382; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1384 = 6'h21 == f2_cut_ptr_0 ? f2_cut_data_dataVec_3_33 : _GEN_1383; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1385 = 6'h22 == f2_cut_ptr_0 ? f2_cut_data_dataVec_3_34 : _GEN_1384; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1386 = 6'h23 == f2_cut_ptr_0 ? f2_cut_data_dataVec_3_35 : _GEN_1385; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1387 = 6'h24 == f2_cut_ptr_0 ? f2_cut_data_dataVec_3_36 : _GEN_1386; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1388 = 6'h25 == f2_cut_ptr_0 ? f2_cut_data_dataVec_3_37 : _GEN_1387; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1389 = 6'h26 == f2_cut_ptr_0 ? f2_cut_data_dataVec_3_38 : _GEN_1388; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1390 = 6'h27 == f2_cut_ptr_0 ? f2_cut_data_dataVec_3_39 : _GEN_1389; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1391 = 6'h28 == f2_cut_ptr_0 ? f2_cut_data_dataVec_3_40 : _GEN_1390; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1392 = 6'h29 == f2_cut_ptr_0 ? f2_cut_data_dataVec_3_41 : _GEN_1391; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1393 = 6'h2a == f2_cut_ptr_0 ? f2_cut_data_dataVec_3_42 : _GEN_1392; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1394 = 6'h2b == f2_cut_ptr_0 ? f2_cut_data_dataVec_3_43 : _GEN_1393; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1395 = 6'h2c == f2_cut_ptr_0 ? f2_cut_data_dataVec_3_44 : _GEN_1394; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1396 = 6'h2d == f2_cut_ptr_0 ? f2_cut_data_dataVec_3_45 : _GEN_1395; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1397 = 6'h2e == f2_cut_ptr_0 ? f2_cut_data_dataVec_3_46 : _GEN_1396; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1400 = 6'h1 == f2_cut_ptr_1 ? f2_cut_data_dataVec_3_1 : f2_cut_data_dataVec_3_0; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1401 = 6'h2 == f2_cut_ptr_1 ? f2_cut_data_dataVec_3_2 : _GEN_1400; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1402 = 6'h3 == f2_cut_ptr_1 ? f2_cut_data_dataVec_3_3 : _GEN_1401; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1403 = 6'h4 == f2_cut_ptr_1 ? f2_cut_data_dataVec_3_4 : _GEN_1402; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1404 = 6'h5 == f2_cut_ptr_1 ? f2_cut_data_dataVec_3_5 : _GEN_1403; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1405 = 6'h6 == f2_cut_ptr_1 ? f2_cut_data_dataVec_3_6 : _GEN_1404; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1406 = 6'h7 == f2_cut_ptr_1 ? f2_cut_data_dataVec_3_7 : _GEN_1405; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1407 = 6'h8 == f2_cut_ptr_1 ? f2_cut_data_dataVec_3_8 : _GEN_1406; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1408 = 6'h9 == f2_cut_ptr_1 ? f2_cut_data_dataVec_3_9 : _GEN_1407; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1409 = 6'ha == f2_cut_ptr_1 ? f2_cut_data_dataVec_3_10 : _GEN_1408; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1410 = 6'hb == f2_cut_ptr_1 ? f2_cut_data_dataVec_3_11 : _GEN_1409; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1411 = 6'hc == f2_cut_ptr_1 ? f2_cut_data_dataVec_3_12 : _GEN_1410; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1412 = 6'hd == f2_cut_ptr_1 ? f2_cut_data_dataVec_3_13 : _GEN_1411; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1413 = 6'he == f2_cut_ptr_1 ? f2_cut_data_dataVec_3_14 : _GEN_1412; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1414 = 6'hf == f2_cut_ptr_1 ? f2_cut_data_dataVec_3_15 : _GEN_1413; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1415 = 6'h10 == f2_cut_ptr_1 ? f2_cut_data_dataVec_3_16 : _GEN_1414; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1416 = 6'h11 == f2_cut_ptr_1 ? f2_cut_data_dataVec_3_17 : _GEN_1415; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1417 = 6'h12 == f2_cut_ptr_1 ? f2_cut_data_dataVec_3_18 : _GEN_1416; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1418 = 6'h13 == f2_cut_ptr_1 ? f2_cut_data_dataVec_3_19 : _GEN_1417; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1419 = 6'h14 == f2_cut_ptr_1 ? f2_cut_data_dataVec_3_20 : _GEN_1418; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1420 = 6'h15 == f2_cut_ptr_1 ? f2_cut_data_dataVec_3_21 : _GEN_1419; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1421 = 6'h16 == f2_cut_ptr_1 ? f2_cut_data_dataVec_3_22 : _GEN_1420; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1422 = 6'h17 == f2_cut_ptr_1 ? f2_cut_data_dataVec_3_23 : _GEN_1421; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1423 = 6'h18 == f2_cut_ptr_1 ? f2_cut_data_dataVec_3_24 : _GEN_1422; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1424 = 6'h19 == f2_cut_ptr_1 ? f2_cut_data_dataVec_3_25 : _GEN_1423; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1425 = 6'h1a == f2_cut_ptr_1 ? f2_cut_data_dataVec_3_26 : _GEN_1424; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1426 = 6'h1b == f2_cut_ptr_1 ? f2_cut_data_dataVec_3_27 : _GEN_1425; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1427 = 6'h1c == f2_cut_ptr_1 ? f2_cut_data_dataVec_3_28 : _GEN_1426; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1428 = 6'h1d == f2_cut_ptr_1 ? f2_cut_data_dataVec_3_29 : _GEN_1427; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1429 = 6'h1e == f2_cut_ptr_1 ? f2_cut_data_dataVec_3_30 : _GEN_1428; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1430 = 6'h1f == f2_cut_ptr_1 ? f2_cut_data_dataVec_3_31 : _GEN_1429; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1431 = 6'h20 == f2_cut_ptr_1 ? f2_cut_data_dataVec_3_32 : _GEN_1430; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1432 = 6'h21 == f2_cut_ptr_1 ? f2_cut_data_dataVec_3_33 : _GEN_1431; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1433 = 6'h22 == f2_cut_ptr_1 ? f2_cut_data_dataVec_3_34 : _GEN_1432; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1434 = 6'h23 == f2_cut_ptr_1 ? f2_cut_data_dataVec_3_35 : _GEN_1433; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1435 = 6'h24 == f2_cut_ptr_1 ? f2_cut_data_dataVec_3_36 : _GEN_1434; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1436 = 6'h25 == f2_cut_ptr_1 ? f2_cut_data_dataVec_3_37 : _GEN_1435; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1437 = 6'h26 == f2_cut_ptr_1 ? f2_cut_data_dataVec_3_38 : _GEN_1436; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1438 = 6'h27 == f2_cut_ptr_1 ? f2_cut_data_dataVec_3_39 : _GEN_1437; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1439 = 6'h28 == f2_cut_ptr_1 ? f2_cut_data_dataVec_3_40 : _GEN_1438; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1440 = 6'h29 == f2_cut_ptr_1 ? f2_cut_data_dataVec_3_41 : _GEN_1439; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1441 = 6'h2a == f2_cut_ptr_1 ? f2_cut_data_dataVec_3_42 : _GEN_1440; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1442 = 6'h2b == f2_cut_ptr_1 ? f2_cut_data_dataVec_3_43 : _GEN_1441; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1443 = 6'h2c == f2_cut_ptr_1 ? f2_cut_data_dataVec_3_44 : _GEN_1442; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1444 = 6'h2d == f2_cut_ptr_1 ? f2_cut_data_dataVec_3_45 : _GEN_1443; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1445 = 6'h2e == f2_cut_ptr_1 ? f2_cut_data_dataVec_3_46 : _GEN_1444; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1448 = 6'h1 == f2_cut_ptr_2 ? f2_cut_data_dataVec_3_1 : f2_cut_data_dataVec_3_0; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1449 = 6'h2 == f2_cut_ptr_2 ? f2_cut_data_dataVec_3_2 : _GEN_1448; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1450 = 6'h3 == f2_cut_ptr_2 ? f2_cut_data_dataVec_3_3 : _GEN_1449; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1451 = 6'h4 == f2_cut_ptr_2 ? f2_cut_data_dataVec_3_4 : _GEN_1450; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1452 = 6'h5 == f2_cut_ptr_2 ? f2_cut_data_dataVec_3_5 : _GEN_1451; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1453 = 6'h6 == f2_cut_ptr_2 ? f2_cut_data_dataVec_3_6 : _GEN_1452; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1454 = 6'h7 == f2_cut_ptr_2 ? f2_cut_data_dataVec_3_7 : _GEN_1453; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1455 = 6'h8 == f2_cut_ptr_2 ? f2_cut_data_dataVec_3_8 : _GEN_1454; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1456 = 6'h9 == f2_cut_ptr_2 ? f2_cut_data_dataVec_3_9 : _GEN_1455; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1457 = 6'ha == f2_cut_ptr_2 ? f2_cut_data_dataVec_3_10 : _GEN_1456; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1458 = 6'hb == f2_cut_ptr_2 ? f2_cut_data_dataVec_3_11 : _GEN_1457; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1459 = 6'hc == f2_cut_ptr_2 ? f2_cut_data_dataVec_3_12 : _GEN_1458; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1460 = 6'hd == f2_cut_ptr_2 ? f2_cut_data_dataVec_3_13 : _GEN_1459; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1461 = 6'he == f2_cut_ptr_2 ? f2_cut_data_dataVec_3_14 : _GEN_1460; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1462 = 6'hf == f2_cut_ptr_2 ? f2_cut_data_dataVec_3_15 : _GEN_1461; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1463 = 6'h10 == f2_cut_ptr_2 ? f2_cut_data_dataVec_3_16 : _GEN_1462; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1464 = 6'h11 == f2_cut_ptr_2 ? f2_cut_data_dataVec_3_17 : _GEN_1463; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1465 = 6'h12 == f2_cut_ptr_2 ? f2_cut_data_dataVec_3_18 : _GEN_1464; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1466 = 6'h13 == f2_cut_ptr_2 ? f2_cut_data_dataVec_3_19 : _GEN_1465; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1467 = 6'h14 == f2_cut_ptr_2 ? f2_cut_data_dataVec_3_20 : _GEN_1466; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1468 = 6'h15 == f2_cut_ptr_2 ? f2_cut_data_dataVec_3_21 : _GEN_1467; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1469 = 6'h16 == f2_cut_ptr_2 ? f2_cut_data_dataVec_3_22 : _GEN_1468; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1470 = 6'h17 == f2_cut_ptr_2 ? f2_cut_data_dataVec_3_23 : _GEN_1469; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1471 = 6'h18 == f2_cut_ptr_2 ? f2_cut_data_dataVec_3_24 : _GEN_1470; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1472 = 6'h19 == f2_cut_ptr_2 ? f2_cut_data_dataVec_3_25 : _GEN_1471; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1473 = 6'h1a == f2_cut_ptr_2 ? f2_cut_data_dataVec_3_26 : _GEN_1472; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1474 = 6'h1b == f2_cut_ptr_2 ? f2_cut_data_dataVec_3_27 : _GEN_1473; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1475 = 6'h1c == f2_cut_ptr_2 ? f2_cut_data_dataVec_3_28 : _GEN_1474; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1476 = 6'h1d == f2_cut_ptr_2 ? f2_cut_data_dataVec_3_29 : _GEN_1475; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1477 = 6'h1e == f2_cut_ptr_2 ? f2_cut_data_dataVec_3_30 : _GEN_1476; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1478 = 6'h1f == f2_cut_ptr_2 ? f2_cut_data_dataVec_3_31 : _GEN_1477; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1479 = 6'h20 == f2_cut_ptr_2 ? f2_cut_data_dataVec_3_32 : _GEN_1478; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1480 = 6'h21 == f2_cut_ptr_2 ? f2_cut_data_dataVec_3_33 : _GEN_1479; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1481 = 6'h22 == f2_cut_ptr_2 ? f2_cut_data_dataVec_3_34 : _GEN_1480; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1482 = 6'h23 == f2_cut_ptr_2 ? f2_cut_data_dataVec_3_35 : _GEN_1481; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1483 = 6'h24 == f2_cut_ptr_2 ? f2_cut_data_dataVec_3_36 : _GEN_1482; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1484 = 6'h25 == f2_cut_ptr_2 ? f2_cut_data_dataVec_3_37 : _GEN_1483; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1485 = 6'h26 == f2_cut_ptr_2 ? f2_cut_data_dataVec_3_38 : _GEN_1484; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1486 = 6'h27 == f2_cut_ptr_2 ? f2_cut_data_dataVec_3_39 : _GEN_1485; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1487 = 6'h28 == f2_cut_ptr_2 ? f2_cut_data_dataVec_3_40 : _GEN_1486; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1488 = 6'h29 == f2_cut_ptr_2 ? f2_cut_data_dataVec_3_41 : _GEN_1487; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1489 = 6'h2a == f2_cut_ptr_2 ? f2_cut_data_dataVec_3_42 : _GEN_1488; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1490 = 6'h2b == f2_cut_ptr_2 ? f2_cut_data_dataVec_3_43 : _GEN_1489; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1491 = 6'h2c == f2_cut_ptr_2 ? f2_cut_data_dataVec_3_44 : _GEN_1490; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1492 = 6'h2d == f2_cut_ptr_2 ? f2_cut_data_dataVec_3_45 : _GEN_1491; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1493 = 6'h2e == f2_cut_ptr_2 ? f2_cut_data_dataVec_3_46 : _GEN_1492; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1496 = 6'h1 == f2_cut_ptr_3 ? f2_cut_data_dataVec_3_1 : f2_cut_data_dataVec_3_0; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1497 = 6'h2 == f2_cut_ptr_3 ? f2_cut_data_dataVec_3_2 : _GEN_1496; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1498 = 6'h3 == f2_cut_ptr_3 ? f2_cut_data_dataVec_3_3 : _GEN_1497; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1499 = 6'h4 == f2_cut_ptr_3 ? f2_cut_data_dataVec_3_4 : _GEN_1498; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1500 = 6'h5 == f2_cut_ptr_3 ? f2_cut_data_dataVec_3_5 : _GEN_1499; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1501 = 6'h6 == f2_cut_ptr_3 ? f2_cut_data_dataVec_3_6 : _GEN_1500; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1502 = 6'h7 == f2_cut_ptr_3 ? f2_cut_data_dataVec_3_7 : _GEN_1501; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1503 = 6'h8 == f2_cut_ptr_3 ? f2_cut_data_dataVec_3_8 : _GEN_1502; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1504 = 6'h9 == f2_cut_ptr_3 ? f2_cut_data_dataVec_3_9 : _GEN_1503; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1505 = 6'ha == f2_cut_ptr_3 ? f2_cut_data_dataVec_3_10 : _GEN_1504; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1506 = 6'hb == f2_cut_ptr_3 ? f2_cut_data_dataVec_3_11 : _GEN_1505; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1507 = 6'hc == f2_cut_ptr_3 ? f2_cut_data_dataVec_3_12 : _GEN_1506; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1508 = 6'hd == f2_cut_ptr_3 ? f2_cut_data_dataVec_3_13 : _GEN_1507; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1509 = 6'he == f2_cut_ptr_3 ? f2_cut_data_dataVec_3_14 : _GEN_1508; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1510 = 6'hf == f2_cut_ptr_3 ? f2_cut_data_dataVec_3_15 : _GEN_1509; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1511 = 6'h10 == f2_cut_ptr_3 ? f2_cut_data_dataVec_3_16 : _GEN_1510; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1512 = 6'h11 == f2_cut_ptr_3 ? f2_cut_data_dataVec_3_17 : _GEN_1511; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1513 = 6'h12 == f2_cut_ptr_3 ? f2_cut_data_dataVec_3_18 : _GEN_1512; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1514 = 6'h13 == f2_cut_ptr_3 ? f2_cut_data_dataVec_3_19 : _GEN_1513; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1515 = 6'h14 == f2_cut_ptr_3 ? f2_cut_data_dataVec_3_20 : _GEN_1514; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1516 = 6'h15 == f2_cut_ptr_3 ? f2_cut_data_dataVec_3_21 : _GEN_1515; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1517 = 6'h16 == f2_cut_ptr_3 ? f2_cut_data_dataVec_3_22 : _GEN_1516; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1518 = 6'h17 == f2_cut_ptr_3 ? f2_cut_data_dataVec_3_23 : _GEN_1517; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1519 = 6'h18 == f2_cut_ptr_3 ? f2_cut_data_dataVec_3_24 : _GEN_1518; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1520 = 6'h19 == f2_cut_ptr_3 ? f2_cut_data_dataVec_3_25 : _GEN_1519; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1521 = 6'h1a == f2_cut_ptr_3 ? f2_cut_data_dataVec_3_26 : _GEN_1520; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1522 = 6'h1b == f2_cut_ptr_3 ? f2_cut_data_dataVec_3_27 : _GEN_1521; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1523 = 6'h1c == f2_cut_ptr_3 ? f2_cut_data_dataVec_3_28 : _GEN_1522; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1524 = 6'h1d == f2_cut_ptr_3 ? f2_cut_data_dataVec_3_29 : _GEN_1523; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1525 = 6'h1e == f2_cut_ptr_3 ? f2_cut_data_dataVec_3_30 : _GEN_1524; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1526 = 6'h1f == f2_cut_ptr_3 ? f2_cut_data_dataVec_3_31 : _GEN_1525; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1527 = 6'h20 == f2_cut_ptr_3 ? f2_cut_data_dataVec_3_32 : _GEN_1526; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1528 = 6'h21 == f2_cut_ptr_3 ? f2_cut_data_dataVec_3_33 : _GEN_1527; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1529 = 6'h22 == f2_cut_ptr_3 ? f2_cut_data_dataVec_3_34 : _GEN_1528; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1530 = 6'h23 == f2_cut_ptr_3 ? f2_cut_data_dataVec_3_35 : _GEN_1529; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1531 = 6'h24 == f2_cut_ptr_3 ? f2_cut_data_dataVec_3_36 : _GEN_1530; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1532 = 6'h25 == f2_cut_ptr_3 ? f2_cut_data_dataVec_3_37 : _GEN_1531; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1533 = 6'h26 == f2_cut_ptr_3 ? f2_cut_data_dataVec_3_38 : _GEN_1532; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1534 = 6'h27 == f2_cut_ptr_3 ? f2_cut_data_dataVec_3_39 : _GEN_1533; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1535 = 6'h28 == f2_cut_ptr_3 ? f2_cut_data_dataVec_3_40 : _GEN_1534; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1536 = 6'h29 == f2_cut_ptr_3 ? f2_cut_data_dataVec_3_41 : _GEN_1535; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1537 = 6'h2a == f2_cut_ptr_3 ? f2_cut_data_dataVec_3_42 : _GEN_1536; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1538 = 6'h2b == f2_cut_ptr_3 ? f2_cut_data_dataVec_3_43 : _GEN_1537; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1539 = 6'h2c == f2_cut_ptr_3 ? f2_cut_data_dataVec_3_44 : _GEN_1538; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1540 = 6'h2d == f2_cut_ptr_3 ? f2_cut_data_dataVec_3_45 : _GEN_1539; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1541 = 6'h2e == f2_cut_ptr_3 ? f2_cut_data_dataVec_3_46 : _GEN_1540; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1544 = 6'h1 == f2_cut_ptr_4 ? f2_cut_data_dataVec_3_1 : f2_cut_data_dataVec_3_0; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1545 = 6'h2 == f2_cut_ptr_4 ? f2_cut_data_dataVec_3_2 : _GEN_1544; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1546 = 6'h3 == f2_cut_ptr_4 ? f2_cut_data_dataVec_3_3 : _GEN_1545; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1547 = 6'h4 == f2_cut_ptr_4 ? f2_cut_data_dataVec_3_4 : _GEN_1546; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1548 = 6'h5 == f2_cut_ptr_4 ? f2_cut_data_dataVec_3_5 : _GEN_1547; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1549 = 6'h6 == f2_cut_ptr_4 ? f2_cut_data_dataVec_3_6 : _GEN_1548; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1550 = 6'h7 == f2_cut_ptr_4 ? f2_cut_data_dataVec_3_7 : _GEN_1549; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1551 = 6'h8 == f2_cut_ptr_4 ? f2_cut_data_dataVec_3_8 : _GEN_1550; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1552 = 6'h9 == f2_cut_ptr_4 ? f2_cut_data_dataVec_3_9 : _GEN_1551; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1553 = 6'ha == f2_cut_ptr_4 ? f2_cut_data_dataVec_3_10 : _GEN_1552; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1554 = 6'hb == f2_cut_ptr_4 ? f2_cut_data_dataVec_3_11 : _GEN_1553; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1555 = 6'hc == f2_cut_ptr_4 ? f2_cut_data_dataVec_3_12 : _GEN_1554; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1556 = 6'hd == f2_cut_ptr_4 ? f2_cut_data_dataVec_3_13 : _GEN_1555; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1557 = 6'he == f2_cut_ptr_4 ? f2_cut_data_dataVec_3_14 : _GEN_1556; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1558 = 6'hf == f2_cut_ptr_4 ? f2_cut_data_dataVec_3_15 : _GEN_1557; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1559 = 6'h10 == f2_cut_ptr_4 ? f2_cut_data_dataVec_3_16 : _GEN_1558; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1560 = 6'h11 == f2_cut_ptr_4 ? f2_cut_data_dataVec_3_17 : _GEN_1559; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1561 = 6'h12 == f2_cut_ptr_4 ? f2_cut_data_dataVec_3_18 : _GEN_1560; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1562 = 6'h13 == f2_cut_ptr_4 ? f2_cut_data_dataVec_3_19 : _GEN_1561; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1563 = 6'h14 == f2_cut_ptr_4 ? f2_cut_data_dataVec_3_20 : _GEN_1562; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1564 = 6'h15 == f2_cut_ptr_4 ? f2_cut_data_dataVec_3_21 : _GEN_1563; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1565 = 6'h16 == f2_cut_ptr_4 ? f2_cut_data_dataVec_3_22 : _GEN_1564; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1566 = 6'h17 == f2_cut_ptr_4 ? f2_cut_data_dataVec_3_23 : _GEN_1565; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1567 = 6'h18 == f2_cut_ptr_4 ? f2_cut_data_dataVec_3_24 : _GEN_1566; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1568 = 6'h19 == f2_cut_ptr_4 ? f2_cut_data_dataVec_3_25 : _GEN_1567; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1569 = 6'h1a == f2_cut_ptr_4 ? f2_cut_data_dataVec_3_26 : _GEN_1568; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1570 = 6'h1b == f2_cut_ptr_4 ? f2_cut_data_dataVec_3_27 : _GEN_1569; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1571 = 6'h1c == f2_cut_ptr_4 ? f2_cut_data_dataVec_3_28 : _GEN_1570; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1572 = 6'h1d == f2_cut_ptr_4 ? f2_cut_data_dataVec_3_29 : _GEN_1571; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1573 = 6'h1e == f2_cut_ptr_4 ? f2_cut_data_dataVec_3_30 : _GEN_1572; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1574 = 6'h1f == f2_cut_ptr_4 ? f2_cut_data_dataVec_3_31 : _GEN_1573; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1575 = 6'h20 == f2_cut_ptr_4 ? f2_cut_data_dataVec_3_32 : _GEN_1574; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1576 = 6'h21 == f2_cut_ptr_4 ? f2_cut_data_dataVec_3_33 : _GEN_1575; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1577 = 6'h22 == f2_cut_ptr_4 ? f2_cut_data_dataVec_3_34 : _GEN_1576; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1578 = 6'h23 == f2_cut_ptr_4 ? f2_cut_data_dataVec_3_35 : _GEN_1577; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1579 = 6'h24 == f2_cut_ptr_4 ? f2_cut_data_dataVec_3_36 : _GEN_1578; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1580 = 6'h25 == f2_cut_ptr_4 ? f2_cut_data_dataVec_3_37 : _GEN_1579; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1581 = 6'h26 == f2_cut_ptr_4 ? f2_cut_data_dataVec_3_38 : _GEN_1580; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1582 = 6'h27 == f2_cut_ptr_4 ? f2_cut_data_dataVec_3_39 : _GEN_1581; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1583 = 6'h28 == f2_cut_ptr_4 ? f2_cut_data_dataVec_3_40 : _GEN_1582; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1584 = 6'h29 == f2_cut_ptr_4 ? f2_cut_data_dataVec_3_41 : _GEN_1583; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1585 = 6'h2a == f2_cut_ptr_4 ? f2_cut_data_dataVec_3_42 : _GEN_1584; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1586 = 6'h2b == f2_cut_ptr_4 ? f2_cut_data_dataVec_3_43 : _GEN_1585; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1587 = 6'h2c == f2_cut_ptr_4 ? f2_cut_data_dataVec_3_44 : _GEN_1586; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1588 = 6'h2d == f2_cut_ptr_4 ? f2_cut_data_dataVec_3_45 : _GEN_1587; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1589 = 6'h2e == f2_cut_ptr_4 ? f2_cut_data_dataVec_3_46 : _GEN_1588; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1592 = 6'h1 == f2_cut_ptr_5 ? f2_cut_data_dataVec_3_1 : f2_cut_data_dataVec_3_0; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1593 = 6'h2 == f2_cut_ptr_5 ? f2_cut_data_dataVec_3_2 : _GEN_1592; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1594 = 6'h3 == f2_cut_ptr_5 ? f2_cut_data_dataVec_3_3 : _GEN_1593; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1595 = 6'h4 == f2_cut_ptr_5 ? f2_cut_data_dataVec_3_4 : _GEN_1594; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1596 = 6'h5 == f2_cut_ptr_5 ? f2_cut_data_dataVec_3_5 : _GEN_1595; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1597 = 6'h6 == f2_cut_ptr_5 ? f2_cut_data_dataVec_3_6 : _GEN_1596; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1598 = 6'h7 == f2_cut_ptr_5 ? f2_cut_data_dataVec_3_7 : _GEN_1597; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1599 = 6'h8 == f2_cut_ptr_5 ? f2_cut_data_dataVec_3_8 : _GEN_1598; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1600 = 6'h9 == f2_cut_ptr_5 ? f2_cut_data_dataVec_3_9 : _GEN_1599; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1601 = 6'ha == f2_cut_ptr_5 ? f2_cut_data_dataVec_3_10 : _GEN_1600; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1602 = 6'hb == f2_cut_ptr_5 ? f2_cut_data_dataVec_3_11 : _GEN_1601; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1603 = 6'hc == f2_cut_ptr_5 ? f2_cut_data_dataVec_3_12 : _GEN_1602; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1604 = 6'hd == f2_cut_ptr_5 ? f2_cut_data_dataVec_3_13 : _GEN_1603; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1605 = 6'he == f2_cut_ptr_5 ? f2_cut_data_dataVec_3_14 : _GEN_1604; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1606 = 6'hf == f2_cut_ptr_5 ? f2_cut_data_dataVec_3_15 : _GEN_1605; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1607 = 6'h10 == f2_cut_ptr_5 ? f2_cut_data_dataVec_3_16 : _GEN_1606; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1608 = 6'h11 == f2_cut_ptr_5 ? f2_cut_data_dataVec_3_17 : _GEN_1607; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1609 = 6'h12 == f2_cut_ptr_5 ? f2_cut_data_dataVec_3_18 : _GEN_1608; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1610 = 6'h13 == f2_cut_ptr_5 ? f2_cut_data_dataVec_3_19 : _GEN_1609; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1611 = 6'h14 == f2_cut_ptr_5 ? f2_cut_data_dataVec_3_20 : _GEN_1610; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1612 = 6'h15 == f2_cut_ptr_5 ? f2_cut_data_dataVec_3_21 : _GEN_1611; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1613 = 6'h16 == f2_cut_ptr_5 ? f2_cut_data_dataVec_3_22 : _GEN_1612; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1614 = 6'h17 == f2_cut_ptr_5 ? f2_cut_data_dataVec_3_23 : _GEN_1613; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1615 = 6'h18 == f2_cut_ptr_5 ? f2_cut_data_dataVec_3_24 : _GEN_1614; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1616 = 6'h19 == f2_cut_ptr_5 ? f2_cut_data_dataVec_3_25 : _GEN_1615; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1617 = 6'h1a == f2_cut_ptr_5 ? f2_cut_data_dataVec_3_26 : _GEN_1616; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1618 = 6'h1b == f2_cut_ptr_5 ? f2_cut_data_dataVec_3_27 : _GEN_1617; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1619 = 6'h1c == f2_cut_ptr_5 ? f2_cut_data_dataVec_3_28 : _GEN_1618; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1620 = 6'h1d == f2_cut_ptr_5 ? f2_cut_data_dataVec_3_29 : _GEN_1619; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1621 = 6'h1e == f2_cut_ptr_5 ? f2_cut_data_dataVec_3_30 : _GEN_1620; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1622 = 6'h1f == f2_cut_ptr_5 ? f2_cut_data_dataVec_3_31 : _GEN_1621; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1623 = 6'h20 == f2_cut_ptr_5 ? f2_cut_data_dataVec_3_32 : _GEN_1622; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1624 = 6'h21 == f2_cut_ptr_5 ? f2_cut_data_dataVec_3_33 : _GEN_1623; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1625 = 6'h22 == f2_cut_ptr_5 ? f2_cut_data_dataVec_3_34 : _GEN_1624; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1626 = 6'h23 == f2_cut_ptr_5 ? f2_cut_data_dataVec_3_35 : _GEN_1625; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1627 = 6'h24 == f2_cut_ptr_5 ? f2_cut_data_dataVec_3_36 : _GEN_1626; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1628 = 6'h25 == f2_cut_ptr_5 ? f2_cut_data_dataVec_3_37 : _GEN_1627; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1629 = 6'h26 == f2_cut_ptr_5 ? f2_cut_data_dataVec_3_38 : _GEN_1628; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1630 = 6'h27 == f2_cut_ptr_5 ? f2_cut_data_dataVec_3_39 : _GEN_1629; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1631 = 6'h28 == f2_cut_ptr_5 ? f2_cut_data_dataVec_3_40 : _GEN_1630; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1632 = 6'h29 == f2_cut_ptr_5 ? f2_cut_data_dataVec_3_41 : _GEN_1631; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1633 = 6'h2a == f2_cut_ptr_5 ? f2_cut_data_dataVec_3_42 : _GEN_1632; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1634 = 6'h2b == f2_cut_ptr_5 ? f2_cut_data_dataVec_3_43 : _GEN_1633; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1635 = 6'h2c == f2_cut_ptr_5 ? f2_cut_data_dataVec_3_44 : _GEN_1634; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1636 = 6'h2d == f2_cut_ptr_5 ? f2_cut_data_dataVec_3_45 : _GEN_1635; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1637 = 6'h2e == f2_cut_ptr_5 ? f2_cut_data_dataVec_3_46 : _GEN_1636; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1640 = 6'h1 == f2_cut_ptr_6 ? f2_cut_data_dataVec_3_1 : f2_cut_data_dataVec_3_0; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1641 = 6'h2 == f2_cut_ptr_6 ? f2_cut_data_dataVec_3_2 : _GEN_1640; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1642 = 6'h3 == f2_cut_ptr_6 ? f2_cut_data_dataVec_3_3 : _GEN_1641; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1643 = 6'h4 == f2_cut_ptr_6 ? f2_cut_data_dataVec_3_4 : _GEN_1642; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1644 = 6'h5 == f2_cut_ptr_6 ? f2_cut_data_dataVec_3_5 : _GEN_1643; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1645 = 6'h6 == f2_cut_ptr_6 ? f2_cut_data_dataVec_3_6 : _GEN_1644; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1646 = 6'h7 == f2_cut_ptr_6 ? f2_cut_data_dataVec_3_7 : _GEN_1645; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1647 = 6'h8 == f2_cut_ptr_6 ? f2_cut_data_dataVec_3_8 : _GEN_1646; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1648 = 6'h9 == f2_cut_ptr_6 ? f2_cut_data_dataVec_3_9 : _GEN_1647; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1649 = 6'ha == f2_cut_ptr_6 ? f2_cut_data_dataVec_3_10 : _GEN_1648; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1650 = 6'hb == f2_cut_ptr_6 ? f2_cut_data_dataVec_3_11 : _GEN_1649; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1651 = 6'hc == f2_cut_ptr_6 ? f2_cut_data_dataVec_3_12 : _GEN_1650; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1652 = 6'hd == f2_cut_ptr_6 ? f2_cut_data_dataVec_3_13 : _GEN_1651; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1653 = 6'he == f2_cut_ptr_6 ? f2_cut_data_dataVec_3_14 : _GEN_1652; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1654 = 6'hf == f2_cut_ptr_6 ? f2_cut_data_dataVec_3_15 : _GEN_1653; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1655 = 6'h10 == f2_cut_ptr_6 ? f2_cut_data_dataVec_3_16 : _GEN_1654; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1656 = 6'h11 == f2_cut_ptr_6 ? f2_cut_data_dataVec_3_17 : _GEN_1655; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1657 = 6'h12 == f2_cut_ptr_6 ? f2_cut_data_dataVec_3_18 : _GEN_1656; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1658 = 6'h13 == f2_cut_ptr_6 ? f2_cut_data_dataVec_3_19 : _GEN_1657; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1659 = 6'h14 == f2_cut_ptr_6 ? f2_cut_data_dataVec_3_20 : _GEN_1658; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1660 = 6'h15 == f2_cut_ptr_6 ? f2_cut_data_dataVec_3_21 : _GEN_1659; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1661 = 6'h16 == f2_cut_ptr_6 ? f2_cut_data_dataVec_3_22 : _GEN_1660; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1662 = 6'h17 == f2_cut_ptr_6 ? f2_cut_data_dataVec_3_23 : _GEN_1661; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1663 = 6'h18 == f2_cut_ptr_6 ? f2_cut_data_dataVec_3_24 : _GEN_1662; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1664 = 6'h19 == f2_cut_ptr_6 ? f2_cut_data_dataVec_3_25 : _GEN_1663; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1665 = 6'h1a == f2_cut_ptr_6 ? f2_cut_data_dataVec_3_26 : _GEN_1664; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1666 = 6'h1b == f2_cut_ptr_6 ? f2_cut_data_dataVec_3_27 : _GEN_1665; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1667 = 6'h1c == f2_cut_ptr_6 ? f2_cut_data_dataVec_3_28 : _GEN_1666; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1668 = 6'h1d == f2_cut_ptr_6 ? f2_cut_data_dataVec_3_29 : _GEN_1667; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1669 = 6'h1e == f2_cut_ptr_6 ? f2_cut_data_dataVec_3_30 : _GEN_1668; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1670 = 6'h1f == f2_cut_ptr_6 ? f2_cut_data_dataVec_3_31 : _GEN_1669; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1671 = 6'h20 == f2_cut_ptr_6 ? f2_cut_data_dataVec_3_32 : _GEN_1670; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1672 = 6'h21 == f2_cut_ptr_6 ? f2_cut_data_dataVec_3_33 : _GEN_1671; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1673 = 6'h22 == f2_cut_ptr_6 ? f2_cut_data_dataVec_3_34 : _GEN_1672; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1674 = 6'h23 == f2_cut_ptr_6 ? f2_cut_data_dataVec_3_35 : _GEN_1673; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1675 = 6'h24 == f2_cut_ptr_6 ? f2_cut_data_dataVec_3_36 : _GEN_1674; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1676 = 6'h25 == f2_cut_ptr_6 ? f2_cut_data_dataVec_3_37 : _GEN_1675; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1677 = 6'h26 == f2_cut_ptr_6 ? f2_cut_data_dataVec_3_38 : _GEN_1676; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1678 = 6'h27 == f2_cut_ptr_6 ? f2_cut_data_dataVec_3_39 : _GEN_1677; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1679 = 6'h28 == f2_cut_ptr_6 ? f2_cut_data_dataVec_3_40 : _GEN_1678; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1680 = 6'h29 == f2_cut_ptr_6 ? f2_cut_data_dataVec_3_41 : _GEN_1679; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1681 = 6'h2a == f2_cut_ptr_6 ? f2_cut_data_dataVec_3_42 : _GEN_1680; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1682 = 6'h2b == f2_cut_ptr_6 ? f2_cut_data_dataVec_3_43 : _GEN_1681; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1683 = 6'h2c == f2_cut_ptr_6 ? f2_cut_data_dataVec_3_44 : _GEN_1682; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1684 = 6'h2d == f2_cut_ptr_6 ? f2_cut_data_dataVec_3_45 : _GEN_1683; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1685 = 6'h2e == f2_cut_ptr_6 ? f2_cut_data_dataVec_3_46 : _GEN_1684; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1688 = 6'h1 == f2_cut_ptr_7 ? f2_cut_data_dataVec_3_1 : f2_cut_data_dataVec_3_0; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1689 = 6'h2 == f2_cut_ptr_7 ? f2_cut_data_dataVec_3_2 : _GEN_1688; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1690 = 6'h3 == f2_cut_ptr_7 ? f2_cut_data_dataVec_3_3 : _GEN_1689; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1691 = 6'h4 == f2_cut_ptr_7 ? f2_cut_data_dataVec_3_4 : _GEN_1690; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1692 = 6'h5 == f2_cut_ptr_7 ? f2_cut_data_dataVec_3_5 : _GEN_1691; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1693 = 6'h6 == f2_cut_ptr_7 ? f2_cut_data_dataVec_3_6 : _GEN_1692; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1694 = 6'h7 == f2_cut_ptr_7 ? f2_cut_data_dataVec_3_7 : _GEN_1693; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1695 = 6'h8 == f2_cut_ptr_7 ? f2_cut_data_dataVec_3_8 : _GEN_1694; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1696 = 6'h9 == f2_cut_ptr_7 ? f2_cut_data_dataVec_3_9 : _GEN_1695; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1697 = 6'ha == f2_cut_ptr_7 ? f2_cut_data_dataVec_3_10 : _GEN_1696; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1698 = 6'hb == f2_cut_ptr_7 ? f2_cut_data_dataVec_3_11 : _GEN_1697; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1699 = 6'hc == f2_cut_ptr_7 ? f2_cut_data_dataVec_3_12 : _GEN_1698; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1700 = 6'hd == f2_cut_ptr_7 ? f2_cut_data_dataVec_3_13 : _GEN_1699; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1701 = 6'he == f2_cut_ptr_7 ? f2_cut_data_dataVec_3_14 : _GEN_1700; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1702 = 6'hf == f2_cut_ptr_7 ? f2_cut_data_dataVec_3_15 : _GEN_1701; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1703 = 6'h10 == f2_cut_ptr_7 ? f2_cut_data_dataVec_3_16 : _GEN_1702; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1704 = 6'h11 == f2_cut_ptr_7 ? f2_cut_data_dataVec_3_17 : _GEN_1703; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1705 = 6'h12 == f2_cut_ptr_7 ? f2_cut_data_dataVec_3_18 : _GEN_1704; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1706 = 6'h13 == f2_cut_ptr_7 ? f2_cut_data_dataVec_3_19 : _GEN_1705; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1707 = 6'h14 == f2_cut_ptr_7 ? f2_cut_data_dataVec_3_20 : _GEN_1706; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1708 = 6'h15 == f2_cut_ptr_7 ? f2_cut_data_dataVec_3_21 : _GEN_1707; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1709 = 6'h16 == f2_cut_ptr_7 ? f2_cut_data_dataVec_3_22 : _GEN_1708; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1710 = 6'h17 == f2_cut_ptr_7 ? f2_cut_data_dataVec_3_23 : _GEN_1709; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1711 = 6'h18 == f2_cut_ptr_7 ? f2_cut_data_dataVec_3_24 : _GEN_1710; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1712 = 6'h19 == f2_cut_ptr_7 ? f2_cut_data_dataVec_3_25 : _GEN_1711; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1713 = 6'h1a == f2_cut_ptr_7 ? f2_cut_data_dataVec_3_26 : _GEN_1712; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1714 = 6'h1b == f2_cut_ptr_7 ? f2_cut_data_dataVec_3_27 : _GEN_1713; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1715 = 6'h1c == f2_cut_ptr_7 ? f2_cut_data_dataVec_3_28 : _GEN_1714; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1716 = 6'h1d == f2_cut_ptr_7 ? f2_cut_data_dataVec_3_29 : _GEN_1715; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1717 = 6'h1e == f2_cut_ptr_7 ? f2_cut_data_dataVec_3_30 : _GEN_1716; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1718 = 6'h1f == f2_cut_ptr_7 ? f2_cut_data_dataVec_3_31 : _GEN_1717; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1719 = 6'h20 == f2_cut_ptr_7 ? f2_cut_data_dataVec_3_32 : _GEN_1718; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1720 = 6'h21 == f2_cut_ptr_7 ? f2_cut_data_dataVec_3_33 : _GEN_1719; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1721 = 6'h22 == f2_cut_ptr_7 ? f2_cut_data_dataVec_3_34 : _GEN_1720; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1722 = 6'h23 == f2_cut_ptr_7 ? f2_cut_data_dataVec_3_35 : _GEN_1721; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1723 = 6'h24 == f2_cut_ptr_7 ? f2_cut_data_dataVec_3_36 : _GEN_1722; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1724 = 6'h25 == f2_cut_ptr_7 ? f2_cut_data_dataVec_3_37 : _GEN_1723; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1725 = 6'h26 == f2_cut_ptr_7 ? f2_cut_data_dataVec_3_38 : _GEN_1724; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1726 = 6'h27 == f2_cut_ptr_7 ? f2_cut_data_dataVec_3_39 : _GEN_1725; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1727 = 6'h28 == f2_cut_ptr_7 ? f2_cut_data_dataVec_3_40 : _GEN_1726; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1728 = 6'h29 == f2_cut_ptr_7 ? f2_cut_data_dataVec_3_41 : _GEN_1727; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1729 = 6'h2a == f2_cut_ptr_7 ? f2_cut_data_dataVec_3_42 : _GEN_1728; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1730 = 6'h2b == f2_cut_ptr_7 ? f2_cut_data_dataVec_3_43 : _GEN_1729; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1731 = 6'h2c == f2_cut_ptr_7 ? f2_cut_data_dataVec_3_44 : _GEN_1730; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1732 = 6'h2d == f2_cut_ptr_7 ? f2_cut_data_dataVec_3_45 : _GEN_1731; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1733 = 6'h2e == f2_cut_ptr_7 ? f2_cut_data_dataVec_3_46 : _GEN_1732; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1736 = 6'h1 == f2_cut_ptr_8 ? f2_cut_data_dataVec_3_1 : f2_cut_data_dataVec_3_0; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1737 = 6'h2 == f2_cut_ptr_8 ? f2_cut_data_dataVec_3_2 : _GEN_1736; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1738 = 6'h3 == f2_cut_ptr_8 ? f2_cut_data_dataVec_3_3 : _GEN_1737; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1739 = 6'h4 == f2_cut_ptr_8 ? f2_cut_data_dataVec_3_4 : _GEN_1738; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1740 = 6'h5 == f2_cut_ptr_8 ? f2_cut_data_dataVec_3_5 : _GEN_1739; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1741 = 6'h6 == f2_cut_ptr_8 ? f2_cut_data_dataVec_3_6 : _GEN_1740; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1742 = 6'h7 == f2_cut_ptr_8 ? f2_cut_data_dataVec_3_7 : _GEN_1741; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1743 = 6'h8 == f2_cut_ptr_8 ? f2_cut_data_dataVec_3_8 : _GEN_1742; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1744 = 6'h9 == f2_cut_ptr_8 ? f2_cut_data_dataVec_3_9 : _GEN_1743; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1745 = 6'ha == f2_cut_ptr_8 ? f2_cut_data_dataVec_3_10 : _GEN_1744; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1746 = 6'hb == f2_cut_ptr_8 ? f2_cut_data_dataVec_3_11 : _GEN_1745; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1747 = 6'hc == f2_cut_ptr_8 ? f2_cut_data_dataVec_3_12 : _GEN_1746; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1748 = 6'hd == f2_cut_ptr_8 ? f2_cut_data_dataVec_3_13 : _GEN_1747; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1749 = 6'he == f2_cut_ptr_8 ? f2_cut_data_dataVec_3_14 : _GEN_1748; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1750 = 6'hf == f2_cut_ptr_8 ? f2_cut_data_dataVec_3_15 : _GEN_1749; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1751 = 6'h10 == f2_cut_ptr_8 ? f2_cut_data_dataVec_3_16 : _GEN_1750; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1752 = 6'h11 == f2_cut_ptr_8 ? f2_cut_data_dataVec_3_17 : _GEN_1751; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1753 = 6'h12 == f2_cut_ptr_8 ? f2_cut_data_dataVec_3_18 : _GEN_1752; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1754 = 6'h13 == f2_cut_ptr_8 ? f2_cut_data_dataVec_3_19 : _GEN_1753; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1755 = 6'h14 == f2_cut_ptr_8 ? f2_cut_data_dataVec_3_20 : _GEN_1754; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1756 = 6'h15 == f2_cut_ptr_8 ? f2_cut_data_dataVec_3_21 : _GEN_1755; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1757 = 6'h16 == f2_cut_ptr_8 ? f2_cut_data_dataVec_3_22 : _GEN_1756; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1758 = 6'h17 == f2_cut_ptr_8 ? f2_cut_data_dataVec_3_23 : _GEN_1757; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1759 = 6'h18 == f2_cut_ptr_8 ? f2_cut_data_dataVec_3_24 : _GEN_1758; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1760 = 6'h19 == f2_cut_ptr_8 ? f2_cut_data_dataVec_3_25 : _GEN_1759; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1761 = 6'h1a == f2_cut_ptr_8 ? f2_cut_data_dataVec_3_26 : _GEN_1760; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1762 = 6'h1b == f2_cut_ptr_8 ? f2_cut_data_dataVec_3_27 : _GEN_1761; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1763 = 6'h1c == f2_cut_ptr_8 ? f2_cut_data_dataVec_3_28 : _GEN_1762; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1764 = 6'h1d == f2_cut_ptr_8 ? f2_cut_data_dataVec_3_29 : _GEN_1763; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1765 = 6'h1e == f2_cut_ptr_8 ? f2_cut_data_dataVec_3_30 : _GEN_1764; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1766 = 6'h1f == f2_cut_ptr_8 ? f2_cut_data_dataVec_3_31 : _GEN_1765; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1767 = 6'h20 == f2_cut_ptr_8 ? f2_cut_data_dataVec_3_32 : _GEN_1766; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1768 = 6'h21 == f2_cut_ptr_8 ? f2_cut_data_dataVec_3_33 : _GEN_1767; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1769 = 6'h22 == f2_cut_ptr_8 ? f2_cut_data_dataVec_3_34 : _GEN_1768; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1770 = 6'h23 == f2_cut_ptr_8 ? f2_cut_data_dataVec_3_35 : _GEN_1769; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1771 = 6'h24 == f2_cut_ptr_8 ? f2_cut_data_dataVec_3_36 : _GEN_1770; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1772 = 6'h25 == f2_cut_ptr_8 ? f2_cut_data_dataVec_3_37 : _GEN_1771; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1773 = 6'h26 == f2_cut_ptr_8 ? f2_cut_data_dataVec_3_38 : _GEN_1772; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1774 = 6'h27 == f2_cut_ptr_8 ? f2_cut_data_dataVec_3_39 : _GEN_1773; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1775 = 6'h28 == f2_cut_ptr_8 ? f2_cut_data_dataVec_3_40 : _GEN_1774; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1776 = 6'h29 == f2_cut_ptr_8 ? f2_cut_data_dataVec_3_41 : _GEN_1775; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1777 = 6'h2a == f2_cut_ptr_8 ? f2_cut_data_dataVec_3_42 : _GEN_1776; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1778 = 6'h2b == f2_cut_ptr_8 ? f2_cut_data_dataVec_3_43 : _GEN_1777; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1779 = 6'h2c == f2_cut_ptr_8 ? f2_cut_data_dataVec_3_44 : _GEN_1778; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1780 = 6'h2d == f2_cut_ptr_8 ? f2_cut_data_dataVec_3_45 : _GEN_1779; // @[IFU.scala 302:{19,19}]
  wire [15:0] _GEN_1781 = 6'h2e == f2_cut_ptr_8 ? f2_cut_data_dataVec_3_46 : _GEN_1780; // @[IFU.scala 302:{19,19}]
  wire [1:0] f2_predecod_ptr = {io_icacheInter_resp_1_bits_select,io_icacheInter_resp_0_bits_select}; // @[Cat.scala 31:58]
  wire [3:0] _preDecoderOut_T = 4'h1 << f2_predecod_ptr; // @[OneHot.scala 57:35]
  wire [63:0] _preDecoderOut_T_677 = _preDecoderOut_T[0] ? preDecoders_0_io_out_jumpOffset_0 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _preDecoderOut_T_678 = _preDecoderOut_T[1] ? preDecoders_1_io_out_jumpOffset_0 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _preDecoderOut_T_679 = _preDecoderOut_T[2] ? preDecoders_2_io_out_jumpOffset_0 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _preDecoderOut_T_680 = _preDecoderOut_T[3] ? preDecoders_3_io_out_jumpOffset_0 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _preDecoderOut_T_681 = _preDecoderOut_T_677 | _preDecoderOut_T_678; // @[Mux.scala 27:73]
  wire [63:0] _preDecoderOut_T_682 = _preDecoderOut_T_681 | _preDecoderOut_T_679; // @[Mux.scala 27:73]
  wire [63:0] preDecoderOut_jumpOffset_0 = _preDecoderOut_T_682 | _preDecoderOut_T_680; // @[Mux.scala 27:73]
  wire [63:0] _preDecoderOut_T_684 = _preDecoderOut_T[0] ? preDecoders_0_io_out_jumpOffset_1 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _preDecoderOut_T_685 = _preDecoderOut_T[1] ? preDecoders_1_io_out_jumpOffset_1 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _preDecoderOut_T_686 = _preDecoderOut_T[2] ? preDecoders_2_io_out_jumpOffset_1 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _preDecoderOut_T_687 = _preDecoderOut_T[3] ? preDecoders_3_io_out_jumpOffset_1 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _preDecoderOut_T_688 = _preDecoderOut_T_684 | _preDecoderOut_T_685; // @[Mux.scala 27:73]
  wire [63:0] _preDecoderOut_T_689 = _preDecoderOut_T_688 | _preDecoderOut_T_686; // @[Mux.scala 27:73]
  wire [63:0] preDecoderOut_jumpOffset_1 = _preDecoderOut_T_689 | _preDecoderOut_T_687; // @[Mux.scala 27:73]
  wire [63:0] _preDecoderOut_T_691 = _preDecoderOut_T[0] ? preDecoders_0_io_out_jumpOffset_2 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _preDecoderOut_T_692 = _preDecoderOut_T[1] ? preDecoders_1_io_out_jumpOffset_2 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _preDecoderOut_T_693 = _preDecoderOut_T[2] ? preDecoders_2_io_out_jumpOffset_2 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _preDecoderOut_T_694 = _preDecoderOut_T[3] ? preDecoders_3_io_out_jumpOffset_2 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _preDecoderOut_T_695 = _preDecoderOut_T_691 | _preDecoderOut_T_692; // @[Mux.scala 27:73]
  wire [63:0] _preDecoderOut_T_696 = _preDecoderOut_T_695 | _preDecoderOut_T_693; // @[Mux.scala 27:73]
  wire [63:0] preDecoderOut_jumpOffset_2 = _preDecoderOut_T_696 | _preDecoderOut_T_694; // @[Mux.scala 27:73]
  wire [63:0] _preDecoderOut_T_698 = _preDecoderOut_T[0] ? preDecoders_0_io_out_jumpOffset_3 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _preDecoderOut_T_699 = _preDecoderOut_T[1] ? preDecoders_1_io_out_jumpOffset_3 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _preDecoderOut_T_700 = _preDecoderOut_T[2] ? preDecoders_2_io_out_jumpOffset_3 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _preDecoderOut_T_701 = _preDecoderOut_T[3] ? preDecoders_3_io_out_jumpOffset_3 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _preDecoderOut_T_702 = _preDecoderOut_T_698 | _preDecoderOut_T_699; // @[Mux.scala 27:73]
  wire [63:0] _preDecoderOut_T_703 = _preDecoderOut_T_702 | _preDecoderOut_T_700; // @[Mux.scala 27:73]
  wire [63:0] preDecoderOut_jumpOffset_3 = _preDecoderOut_T_703 | _preDecoderOut_T_701; // @[Mux.scala 27:73]
  wire [63:0] _preDecoderOut_T_705 = _preDecoderOut_T[0] ? preDecoders_0_io_out_jumpOffset_4 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _preDecoderOut_T_706 = _preDecoderOut_T[1] ? preDecoders_1_io_out_jumpOffset_4 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _preDecoderOut_T_707 = _preDecoderOut_T[2] ? preDecoders_2_io_out_jumpOffset_4 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _preDecoderOut_T_708 = _preDecoderOut_T[3] ? preDecoders_3_io_out_jumpOffset_4 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _preDecoderOut_T_709 = _preDecoderOut_T_705 | _preDecoderOut_T_706; // @[Mux.scala 27:73]
  wire [63:0] _preDecoderOut_T_710 = _preDecoderOut_T_709 | _preDecoderOut_T_707; // @[Mux.scala 27:73]
  wire [63:0] preDecoderOut_jumpOffset_4 = _preDecoderOut_T_710 | _preDecoderOut_T_708; // @[Mux.scala 27:73]
  wire [63:0] _preDecoderOut_T_712 = _preDecoderOut_T[0] ? preDecoders_0_io_out_jumpOffset_5 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _preDecoderOut_T_713 = _preDecoderOut_T[1] ? preDecoders_1_io_out_jumpOffset_5 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _preDecoderOut_T_714 = _preDecoderOut_T[2] ? preDecoders_2_io_out_jumpOffset_5 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _preDecoderOut_T_715 = _preDecoderOut_T[3] ? preDecoders_3_io_out_jumpOffset_5 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _preDecoderOut_T_716 = _preDecoderOut_T_712 | _preDecoderOut_T_713; // @[Mux.scala 27:73]
  wire [63:0] _preDecoderOut_T_717 = _preDecoderOut_T_716 | _preDecoderOut_T_714; // @[Mux.scala 27:73]
  wire [63:0] preDecoderOut_jumpOffset_5 = _preDecoderOut_T_717 | _preDecoderOut_T_715; // @[Mux.scala 27:73]
  wire [63:0] _preDecoderOut_T_719 = _preDecoderOut_T[0] ? preDecoders_0_io_out_jumpOffset_6 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _preDecoderOut_T_720 = _preDecoderOut_T[1] ? preDecoders_1_io_out_jumpOffset_6 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _preDecoderOut_T_721 = _preDecoderOut_T[2] ? preDecoders_2_io_out_jumpOffset_6 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _preDecoderOut_T_722 = _preDecoderOut_T[3] ? preDecoders_3_io_out_jumpOffset_6 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _preDecoderOut_T_723 = _preDecoderOut_T_719 | _preDecoderOut_T_720; // @[Mux.scala 27:73]
  wire [63:0] _preDecoderOut_T_724 = _preDecoderOut_T_723 | _preDecoderOut_T_721; // @[Mux.scala 27:73]
  wire [63:0] preDecoderOut_jumpOffset_6 = _preDecoderOut_T_724 | _preDecoderOut_T_722; // @[Mux.scala 27:73]
  wire [63:0] _preDecoderOut_T_726 = _preDecoderOut_T[0] ? preDecoders_0_io_out_jumpOffset_7 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _preDecoderOut_T_727 = _preDecoderOut_T[1] ? preDecoders_1_io_out_jumpOffset_7 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _preDecoderOut_T_728 = _preDecoderOut_T[2] ? preDecoders_2_io_out_jumpOffset_7 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _preDecoderOut_T_729 = _preDecoderOut_T[3] ? preDecoders_3_io_out_jumpOffset_7 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _preDecoderOut_T_730 = _preDecoderOut_T_726 | _preDecoderOut_T_727; // @[Mux.scala 27:73]
  wire [63:0] _preDecoderOut_T_731 = _preDecoderOut_T_730 | _preDecoderOut_T_728; // @[Mux.scala 27:73]
  wire [63:0] preDecoderOut_jumpOffset_7 = _preDecoderOut_T_731 | _preDecoderOut_T_729; // @[Mux.scala 27:73]
  wire [31:0] _preDecoderOut_T_733 = _preDecoderOut_T[0] ? preDecoders_0_io_out_instr_0 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _preDecoderOut_T_734 = _preDecoderOut_T[1] ? preDecoders_1_io_out_instr_0 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _preDecoderOut_T_735 = _preDecoderOut_T[2] ? preDecoders_2_io_out_instr_0 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _preDecoderOut_T_736 = _preDecoderOut_T[3] ? preDecoders_3_io_out_instr_0 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _preDecoderOut_T_737 = _preDecoderOut_T_733 | _preDecoderOut_T_734; // @[Mux.scala 27:73]
  wire [31:0] _preDecoderOut_T_738 = _preDecoderOut_T_737 | _preDecoderOut_T_735; // @[Mux.scala 27:73]
  wire [31:0] preDecoderOut_instr_0 = _preDecoderOut_T_738 | _preDecoderOut_T_736; // @[Mux.scala 27:73]
  wire [31:0] _preDecoderOut_T_740 = _preDecoderOut_T[0] ? preDecoders_0_io_out_instr_1 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _preDecoderOut_T_741 = _preDecoderOut_T[1] ? preDecoders_1_io_out_instr_1 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _preDecoderOut_T_742 = _preDecoderOut_T[2] ? preDecoders_2_io_out_instr_1 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _preDecoderOut_T_743 = _preDecoderOut_T[3] ? preDecoders_3_io_out_instr_1 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _preDecoderOut_T_744 = _preDecoderOut_T_740 | _preDecoderOut_T_741; // @[Mux.scala 27:73]
  wire [31:0] _preDecoderOut_T_745 = _preDecoderOut_T_744 | _preDecoderOut_T_742; // @[Mux.scala 27:73]
  wire [31:0] preDecoderOut_instr_1 = _preDecoderOut_T_745 | _preDecoderOut_T_743; // @[Mux.scala 27:73]
  wire [31:0] _preDecoderOut_T_747 = _preDecoderOut_T[0] ? preDecoders_0_io_out_instr_2 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _preDecoderOut_T_748 = _preDecoderOut_T[1] ? preDecoders_1_io_out_instr_2 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _preDecoderOut_T_749 = _preDecoderOut_T[2] ? preDecoders_2_io_out_instr_2 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _preDecoderOut_T_750 = _preDecoderOut_T[3] ? preDecoders_3_io_out_instr_2 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _preDecoderOut_T_751 = _preDecoderOut_T_747 | _preDecoderOut_T_748; // @[Mux.scala 27:73]
  wire [31:0] _preDecoderOut_T_752 = _preDecoderOut_T_751 | _preDecoderOut_T_749; // @[Mux.scala 27:73]
  wire [31:0] preDecoderOut_instr_2 = _preDecoderOut_T_752 | _preDecoderOut_T_750; // @[Mux.scala 27:73]
  wire [31:0] _preDecoderOut_T_754 = _preDecoderOut_T[0] ? preDecoders_0_io_out_instr_3 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _preDecoderOut_T_755 = _preDecoderOut_T[1] ? preDecoders_1_io_out_instr_3 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _preDecoderOut_T_756 = _preDecoderOut_T[2] ? preDecoders_2_io_out_instr_3 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _preDecoderOut_T_757 = _preDecoderOut_T[3] ? preDecoders_3_io_out_instr_3 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _preDecoderOut_T_758 = _preDecoderOut_T_754 | _preDecoderOut_T_755; // @[Mux.scala 27:73]
  wire [31:0] _preDecoderOut_T_759 = _preDecoderOut_T_758 | _preDecoderOut_T_756; // @[Mux.scala 27:73]
  wire [31:0] preDecoderOut_instr_3 = _preDecoderOut_T_759 | _preDecoderOut_T_757; // @[Mux.scala 27:73]
  wire [31:0] _preDecoderOut_T_761 = _preDecoderOut_T[0] ? preDecoders_0_io_out_instr_4 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _preDecoderOut_T_762 = _preDecoderOut_T[1] ? preDecoders_1_io_out_instr_4 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _preDecoderOut_T_763 = _preDecoderOut_T[2] ? preDecoders_2_io_out_instr_4 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _preDecoderOut_T_764 = _preDecoderOut_T[3] ? preDecoders_3_io_out_instr_4 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _preDecoderOut_T_765 = _preDecoderOut_T_761 | _preDecoderOut_T_762; // @[Mux.scala 27:73]
  wire [31:0] _preDecoderOut_T_766 = _preDecoderOut_T_765 | _preDecoderOut_T_763; // @[Mux.scala 27:73]
  wire [31:0] preDecoderOut_instr_4 = _preDecoderOut_T_766 | _preDecoderOut_T_764; // @[Mux.scala 27:73]
  wire [31:0] _preDecoderOut_T_768 = _preDecoderOut_T[0] ? preDecoders_0_io_out_instr_5 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _preDecoderOut_T_769 = _preDecoderOut_T[1] ? preDecoders_1_io_out_instr_5 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _preDecoderOut_T_770 = _preDecoderOut_T[2] ? preDecoders_2_io_out_instr_5 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _preDecoderOut_T_771 = _preDecoderOut_T[3] ? preDecoders_3_io_out_instr_5 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _preDecoderOut_T_772 = _preDecoderOut_T_768 | _preDecoderOut_T_769; // @[Mux.scala 27:73]
  wire [31:0] _preDecoderOut_T_773 = _preDecoderOut_T_772 | _preDecoderOut_T_770; // @[Mux.scala 27:73]
  wire [31:0] preDecoderOut_instr_5 = _preDecoderOut_T_773 | _preDecoderOut_T_771; // @[Mux.scala 27:73]
  wire [31:0] _preDecoderOut_T_775 = _preDecoderOut_T[0] ? preDecoders_0_io_out_instr_6 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _preDecoderOut_T_776 = _preDecoderOut_T[1] ? preDecoders_1_io_out_instr_6 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _preDecoderOut_T_777 = _preDecoderOut_T[2] ? preDecoders_2_io_out_instr_6 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _preDecoderOut_T_778 = _preDecoderOut_T[3] ? preDecoders_3_io_out_instr_6 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _preDecoderOut_T_779 = _preDecoderOut_T_775 | _preDecoderOut_T_776; // @[Mux.scala 27:73]
  wire [31:0] _preDecoderOut_T_780 = _preDecoderOut_T_779 | _preDecoderOut_T_777; // @[Mux.scala 27:73]
  wire [31:0] preDecoderOut_instr_6 = _preDecoderOut_T_780 | _preDecoderOut_T_778; // @[Mux.scala 27:73]
  wire [31:0] _preDecoderOut_T_782 = _preDecoderOut_T[0] ? preDecoders_0_io_out_instr_7 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _preDecoderOut_T_783 = _preDecoderOut_T[1] ? preDecoders_1_io_out_instr_7 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _preDecoderOut_T_784 = _preDecoderOut_T[2] ? preDecoders_2_io_out_instr_7 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _preDecoderOut_T_785 = _preDecoderOut_T[3] ? preDecoders_3_io_out_instr_7 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _preDecoderOut_T_786 = _preDecoderOut_T_782 | _preDecoderOut_T_783; // @[Mux.scala 27:73]
  wire [31:0] _preDecoderOut_T_787 = _preDecoderOut_T_786 | _preDecoderOut_T_784; // @[Mux.scala 27:73]
  wire [31:0] preDecoderOut_instr_7 = _preDecoderOut_T_787 | _preDecoderOut_T_785; // @[Mux.scala 27:73]
  wire  preDecoderOut_hasHalfValid_1 = _preDecoderOut_T[0] | _preDecoderOut_T[1] | _preDecoderOut_T[2] |
    _preDecoderOut_T[3]; // @[Mux.scala 27:73]
  wire  preDecoderOut_hasHalfValid_2 = _preDecoderOut_T[0] & preDecoders_0_io_out_hasHalfValid_2 | _preDecoderOut_T[1]
     & preDecoders_1_io_out_hasHalfValid_2 | _preDecoderOut_T[2] & preDecoders_2_io_out_hasHalfValid_2 |
    _preDecoderOut_T[3] & preDecoders_3_io_out_hasHalfValid_2; // @[Mux.scala 27:73]
  wire  preDecoderOut_hasHalfValid_3 = _preDecoderOut_T[0] & preDecoders_0_io_out_hasHalfValid_3 | _preDecoderOut_T[1]
     & preDecoders_1_io_out_hasHalfValid_3 | _preDecoderOut_T[2] & preDecoders_2_io_out_hasHalfValid_3 |
    _preDecoderOut_T[3] & preDecoders_3_io_out_hasHalfValid_3; // @[Mux.scala 27:73]
  wire  preDecoderOut_hasHalfValid_4 = _preDecoderOut_T[0] & preDecoders_0_io_out_hasHalfValid_4 | _preDecoderOut_T[1]
     & preDecoders_1_io_out_hasHalfValid_4 | _preDecoderOut_T[2] & preDecoders_2_io_out_hasHalfValid_4 |
    _preDecoderOut_T[3] & preDecoders_3_io_out_hasHalfValid_4; // @[Mux.scala 27:73]
  wire  preDecoderOut_hasHalfValid_5 = _preDecoderOut_T[0] & preDecoders_0_io_out_hasHalfValid_5 | _preDecoderOut_T[1]
     & preDecoders_1_io_out_hasHalfValid_5 | _preDecoderOut_T[2] & preDecoders_2_io_out_hasHalfValid_5 |
    _preDecoderOut_T[3] & preDecoders_3_io_out_hasHalfValid_5; // @[Mux.scala 27:73]
  wire  preDecoderOut_hasHalfValid_6 = _preDecoderOut_T[0] & preDecoders_0_io_out_hasHalfValid_6 | _preDecoderOut_T[1]
     & preDecoders_1_io_out_hasHalfValid_6 | _preDecoderOut_T[2] & preDecoders_2_io_out_hasHalfValid_6 |
    _preDecoderOut_T[3] & preDecoders_3_io_out_hasHalfValid_6; // @[Mux.scala 27:73]
  wire  preDecoderOut_hasHalfValid_7 = _preDecoderOut_T[0] & preDecoders_0_io_out_hasHalfValid_7 | _preDecoderOut_T[1]
     & preDecoders_1_io_out_hasHalfValid_7 | _preDecoderOut_T[2] & preDecoders_2_io_out_hasHalfValid_7 |
    _preDecoderOut_T[3] & preDecoders_3_io_out_hasHalfValid_7; // @[Mux.scala 27:73]
  wire  preDecoderOut_pd_0_isRet = _preDecoderOut_T[0] & preDecoders_0_io_out_pd_0_isRet | _preDecoderOut_T[1] &
    preDecoders_1_io_out_pd_0_isRet | _preDecoderOut_T[2] & preDecoders_2_io_out_pd_0_isRet | _preDecoderOut_T[3] &
    preDecoders_3_io_out_pd_0_isRet; // @[Mux.scala 27:73]
  wire  preDecoderOut_pd_0_isCall = _preDecoderOut_T[0] & preDecoders_0_io_out_pd_0_isCall | _preDecoderOut_T[1] &
    preDecoders_1_io_out_pd_0_isCall | _preDecoderOut_T[2] & preDecoders_2_io_out_pd_0_isCall | _preDecoderOut_T[3] &
    preDecoders_3_io_out_pd_0_isCall; // @[Mux.scala 27:73]
  wire [1:0] _preDecoderOut_T_859 = _preDecoderOut_T[0] ? preDecoders_0_io_out_pd_0_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _preDecoderOut_T_860 = _preDecoderOut_T[1] ? preDecoders_1_io_out_pd_0_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _preDecoderOut_T_861 = _preDecoderOut_T[2] ? preDecoders_2_io_out_pd_0_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _preDecoderOut_T_862 = _preDecoderOut_T[3] ? preDecoders_3_io_out_pd_0_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _preDecoderOut_T_863 = _preDecoderOut_T_859 | _preDecoderOut_T_860; // @[Mux.scala 27:73]
  wire [1:0] _preDecoderOut_T_864 = _preDecoderOut_T_863 | _preDecoderOut_T_861; // @[Mux.scala 27:73]
  wire [1:0] preDecoderOut_pd_0_brType = _preDecoderOut_T_864 | _preDecoderOut_T_862; // @[Mux.scala 27:73]
  wire  preDecoderOut_pd_0_isRVC = _preDecoderOut_T[0] & preDecoders_0_io_out_pd_0_isRVC | _preDecoderOut_T[1] &
    preDecoders_1_io_out_pd_0_isRVC | _preDecoderOut_T[2] & preDecoders_2_io_out_pd_0_isRVC | _preDecoderOut_T[3] &
    preDecoders_3_io_out_pd_0_isRVC; // @[Mux.scala 27:73]
  wire  preDecoderOut_pd_1_isRet = _preDecoderOut_T[0] & preDecoders_0_io_out_pd_1_isRet | _preDecoderOut_T[1] &
    preDecoders_1_io_out_pd_1_isRet | _preDecoderOut_T[2] & preDecoders_2_io_out_pd_1_isRet | _preDecoderOut_T[3] &
    preDecoders_3_io_out_pd_1_isRet; // @[Mux.scala 27:73]
  wire  preDecoderOut_pd_1_isCall = _preDecoderOut_T[0] & preDecoders_0_io_out_pd_1_isCall | _preDecoderOut_T[1] &
    preDecoders_1_io_out_pd_1_isCall | _preDecoderOut_T[2] & preDecoders_2_io_out_pd_1_isCall | _preDecoderOut_T[3] &
    preDecoders_3_io_out_pd_1_isCall; // @[Mux.scala 27:73]
  wire [1:0] _preDecoderOut_T_894 = _preDecoderOut_T[0] ? preDecoders_0_io_out_pd_1_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _preDecoderOut_T_895 = _preDecoderOut_T[1] ? preDecoders_1_io_out_pd_1_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _preDecoderOut_T_896 = _preDecoderOut_T[2] ? preDecoders_2_io_out_pd_1_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _preDecoderOut_T_897 = _preDecoderOut_T[3] ? preDecoders_3_io_out_pd_1_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _preDecoderOut_T_898 = _preDecoderOut_T_894 | _preDecoderOut_T_895; // @[Mux.scala 27:73]
  wire [1:0] _preDecoderOut_T_899 = _preDecoderOut_T_898 | _preDecoderOut_T_896; // @[Mux.scala 27:73]
  wire [1:0] preDecoderOut_pd_1_brType = _preDecoderOut_T_899 | _preDecoderOut_T_897; // @[Mux.scala 27:73]
  wire  preDecoderOut_pd_1_isRVC = _preDecoderOut_T[0] & preDecoders_0_io_out_pd_1_isRVC | _preDecoderOut_T[1] &
    preDecoders_1_io_out_pd_1_isRVC | _preDecoderOut_T[2] & preDecoders_2_io_out_pd_1_isRVC | _preDecoderOut_T[3] &
    preDecoders_3_io_out_pd_1_isRVC; // @[Mux.scala 27:73]
  wire  preDecoderOut_pd_1_valid = _preDecoderOut_T[0] & preDecoders_0_io_out_pd_1_valid | _preDecoderOut_T[1] &
    preDecoders_1_io_out_pd_1_valid | _preDecoderOut_T[2] & preDecoders_2_io_out_pd_1_valid | _preDecoderOut_T[3] &
    preDecoders_3_io_out_pd_1_valid; // @[Mux.scala 27:73]
  wire  preDecoderOut_pd_2_isRet = _preDecoderOut_T[0] & preDecoders_0_io_out_pd_2_isRet | _preDecoderOut_T[1] &
    preDecoders_1_io_out_pd_2_isRet | _preDecoderOut_T[2] & preDecoders_2_io_out_pd_2_isRet | _preDecoderOut_T[3] &
    preDecoders_3_io_out_pd_2_isRet; // @[Mux.scala 27:73]
  wire  preDecoderOut_pd_2_isCall = _preDecoderOut_T[0] & preDecoders_0_io_out_pd_2_isCall | _preDecoderOut_T[1] &
    preDecoders_1_io_out_pd_2_isCall | _preDecoderOut_T[2] & preDecoders_2_io_out_pd_2_isCall | _preDecoderOut_T[3] &
    preDecoders_3_io_out_pd_2_isCall; // @[Mux.scala 27:73]
  wire [1:0] _preDecoderOut_T_929 = _preDecoderOut_T[0] ? preDecoders_0_io_out_pd_2_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _preDecoderOut_T_930 = _preDecoderOut_T[1] ? preDecoders_1_io_out_pd_2_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _preDecoderOut_T_931 = _preDecoderOut_T[2] ? preDecoders_2_io_out_pd_2_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _preDecoderOut_T_932 = _preDecoderOut_T[3] ? preDecoders_3_io_out_pd_2_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _preDecoderOut_T_933 = _preDecoderOut_T_929 | _preDecoderOut_T_930; // @[Mux.scala 27:73]
  wire [1:0] _preDecoderOut_T_934 = _preDecoderOut_T_933 | _preDecoderOut_T_931; // @[Mux.scala 27:73]
  wire [1:0] preDecoderOut_pd_2_brType = _preDecoderOut_T_934 | _preDecoderOut_T_932; // @[Mux.scala 27:73]
  wire  preDecoderOut_pd_2_isRVC = _preDecoderOut_T[0] & preDecoders_0_io_out_pd_2_isRVC | _preDecoderOut_T[1] &
    preDecoders_1_io_out_pd_2_isRVC | _preDecoderOut_T[2] & preDecoders_2_io_out_pd_2_isRVC | _preDecoderOut_T[3] &
    preDecoders_3_io_out_pd_2_isRVC; // @[Mux.scala 27:73]
  wire  preDecoderOut_pd_2_valid = _preDecoderOut_T[0] & preDecoders_0_io_out_pd_2_valid | _preDecoderOut_T[1] &
    preDecoders_1_io_out_pd_2_valid | _preDecoderOut_T[2] & preDecoders_2_io_out_pd_2_valid | _preDecoderOut_T[3] &
    preDecoders_3_io_out_pd_2_valid; // @[Mux.scala 27:73]
  wire  preDecoderOut_pd_3_isRet = _preDecoderOut_T[0] & preDecoders_0_io_out_pd_3_isRet | _preDecoderOut_T[1] &
    preDecoders_1_io_out_pd_3_isRet | _preDecoderOut_T[2] & preDecoders_2_io_out_pd_3_isRet | _preDecoderOut_T[3] &
    preDecoders_3_io_out_pd_3_isRet; // @[Mux.scala 27:73]
  wire  preDecoderOut_pd_3_isCall = _preDecoderOut_T[0] & preDecoders_0_io_out_pd_3_isCall | _preDecoderOut_T[1] &
    preDecoders_1_io_out_pd_3_isCall | _preDecoderOut_T[2] & preDecoders_2_io_out_pd_3_isCall | _preDecoderOut_T[3] &
    preDecoders_3_io_out_pd_3_isCall; // @[Mux.scala 27:73]
  wire [1:0] _preDecoderOut_T_964 = _preDecoderOut_T[0] ? preDecoders_0_io_out_pd_3_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _preDecoderOut_T_965 = _preDecoderOut_T[1] ? preDecoders_1_io_out_pd_3_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _preDecoderOut_T_966 = _preDecoderOut_T[2] ? preDecoders_2_io_out_pd_3_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _preDecoderOut_T_967 = _preDecoderOut_T[3] ? preDecoders_3_io_out_pd_3_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _preDecoderOut_T_968 = _preDecoderOut_T_964 | _preDecoderOut_T_965; // @[Mux.scala 27:73]
  wire [1:0] _preDecoderOut_T_969 = _preDecoderOut_T_968 | _preDecoderOut_T_966; // @[Mux.scala 27:73]
  wire [1:0] preDecoderOut_pd_3_brType = _preDecoderOut_T_969 | _preDecoderOut_T_967; // @[Mux.scala 27:73]
  wire  preDecoderOut_pd_3_isRVC = _preDecoderOut_T[0] & preDecoders_0_io_out_pd_3_isRVC | _preDecoderOut_T[1] &
    preDecoders_1_io_out_pd_3_isRVC | _preDecoderOut_T[2] & preDecoders_2_io_out_pd_3_isRVC | _preDecoderOut_T[3] &
    preDecoders_3_io_out_pd_3_isRVC; // @[Mux.scala 27:73]
  wire  preDecoderOut_pd_3_valid = _preDecoderOut_T[0] & preDecoders_0_io_out_pd_3_valid | _preDecoderOut_T[1] &
    preDecoders_1_io_out_pd_3_valid | _preDecoderOut_T[2] & preDecoders_2_io_out_pd_3_valid | _preDecoderOut_T[3] &
    preDecoders_3_io_out_pd_3_valid; // @[Mux.scala 27:73]
  wire  preDecoderOut_pd_4_isRet = _preDecoderOut_T[0] & preDecoders_0_io_out_pd_4_isRet | _preDecoderOut_T[1] &
    preDecoders_1_io_out_pd_4_isRet | _preDecoderOut_T[2] & preDecoders_2_io_out_pd_4_isRet | _preDecoderOut_T[3] &
    preDecoders_3_io_out_pd_4_isRet; // @[Mux.scala 27:73]
  wire  preDecoderOut_pd_4_isCall = _preDecoderOut_T[0] & preDecoders_0_io_out_pd_4_isCall | _preDecoderOut_T[1] &
    preDecoders_1_io_out_pd_4_isCall | _preDecoderOut_T[2] & preDecoders_2_io_out_pd_4_isCall | _preDecoderOut_T[3] &
    preDecoders_3_io_out_pd_4_isCall; // @[Mux.scala 27:73]
  wire [1:0] _preDecoderOut_T_999 = _preDecoderOut_T[0] ? preDecoders_0_io_out_pd_4_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _preDecoderOut_T_1000 = _preDecoderOut_T[1] ? preDecoders_1_io_out_pd_4_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _preDecoderOut_T_1001 = _preDecoderOut_T[2] ? preDecoders_2_io_out_pd_4_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _preDecoderOut_T_1002 = _preDecoderOut_T[3] ? preDecoders_3_io_out_pd_4_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _preDecoderOut_T_1003 = _preDecoderOut_T_999 | _preDecoderOut_T_1000; // @[Mux.scala 27:73]
  wire [1:0] _preDecoderOut_T_1004 = _preDecoderOut_T_1003 | _preDecoderOut_T_1001; // @[Mux.scala 27:73]
  wire [1:0] preDecoderOut_pd_4_brType = _preDecoderOut_T_1004 | _preDecoderOut_T_1002; // @[Mux.scala 27:73]
  wire  preDecoderOut_pd_4_isRVC = _preDecoderOut_T[0] & preDecoders_0_io_out_pd_4_isRVC | _preDecoderOut_T[1] &
    preDecoders_1_io_out_pd_4_isRVC | _preDecoderOut_T[2] & preDecoders_2_io_out_pd_4_isRVC | _preDecoderOut_T[3] &
    preDecoders_3_io_out_pd_4_isRVC; // @[Mux.scala 27:73]
  wire  preDecoderOut_pd_4_valid = _preDecoderOut_T[0] & preDecoders_0_io_out_pd_4_valid | _preDecoderOut_T[1] &
    preDecoders_1_io_out_pd_4_valid | _preDecoderOut_T[2] & preDecoders_2_io_out_pd_4_valid | _preDecoderOut_T[3] &
    preDecoders_3_io_out_pd_4_valid; // @[Mux.scala 27:73]
  wire  preDecoderOut_pd_5_isRet = _preDecoderOut_T[0] & preDecoders_0_io_out_pd_5_isRet | _preDecoderOut_T[1] &
    preDecoders_1_io_out_pd_5_isRet | _preDecoderOut_T[2] & preDecoders_2_io_out_pd_5_isRet | _preDecoderOut_T[3] &
    preDecoders_3_io_out_pd_5_isRet; // @[Mux.scala 27:73]
  wire  preDecoderOut_pd_5_isCall = _preDecoderOut_T[0] & preDecoders_0_io_out_pd_5_isCall | _preDecoderOut_T[1] &
    preDecoders_1_io_out_pd_5_isCall | _preDecoderOut_T[2] & preDecoders_2_io_out_pd_5_isCall | _preDecoderOut_T[3] &
    preDecoders_3_io_out_pd_5_isCall; // @[Mux.scala 27:73]
  wire [1:0] _preDecoderOut_T_1034 = _preDecoderOut_T[0] ? preDecoders_0_io_out_pd_5_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _preDecoderOut_T_1035 = _preDecoderOut_T[1] ? preDecoders_1_io_out_pd_5_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _preDecoderOut_T_1036 = _preDecoderOut_T[2] ? preDecoders_2_io_out_pd_5_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _preDecoderOut_T_1037 = _preDecoderOut_T[3] ? preDecoders_3_io_out_pd_5_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _preDecoderOut_T_1038 = _preDecoderOut_T_1034 | _preDecoderOut_T_1035; // @[Mux.scala 27:73]
  wire [1:0] _preDecoderOut_T_1039 = _preDecoderOut_T_1038 | _preDecoderOut_T_1036; // @[Mux.scala 27:73]
  wire [1:0] preDecoderOut_pd_5_brType = _preDecoderOut_T_1039 | _preDecoderOut_T_1037; // @[Mux.scala 27:73]
  wire  preDecoderOut_pd_5_isRVC = _preDecoderOut_T[0] & preDecoders_0_io_out_pd_5_isRVC | _preDecoderOut_T[1] &
    preDecoders_1_io_out_pd_5_isRVC | _preDecoderOut_T[2] & preDecoders_2_io_out_pd_5_isRVC | _preDecoderOut_T[3] &
    preDecoders_3_io_out_pd_5_isRVC; // @[Mux.scala 27:73]
  wire  preDecoderOut_pd_5_valid = _preDecoderOut_T[0] & preDecoders_0_io_out_pd_5_valid | _preDecoderOut_T[1] &
    preDecoders_1_io_out_pd_5_valid | _preDecoderOut_T[2] & preDecoders_2_io_out_pd_5_valid | _preDecoderOut_T[3] &
    preDecoders_3_io_out_pd_5_valid; // @[Mux.scala 27:73]
  wire  preDecoderOut_pd_6_isRet = _preDecoderOut_T[0] & preDecoders_0_io_out_pd_6_isRet | _preDecoderOut_T[1] &
    preDecoders_1_io_out_pd_6_isRet | _preDecoderOut_T[2] & preDecoders_2_io_out_pd_6_isRet | _preDecoderOut_T[3] &
    preDecoders_3_io_out_pd_6_isRet; // @[Mux.scala 27:73]
  wire  preDecoderOut_pd_6_isCall = _preDecoderOut_T[0] & preDecoders_0_io_out_pd_6_isCall | _preDecoderOut_T[1] &
    preDecoders_1_io_out_pd_6_isCall | _preDecoderOut_T[2] & preDecoders_2_io_out_pd_6_isCall | _preDecoderOut_T[3] &
    preDecoders_3_io_out_pd_6_isCall; // @[Mux.scala 27:73]
  wire [1:0] _preDecoderOut_T_1069 = _preDecoderOut_T[0] ? preDecoders_0_io_out_pd_6_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _preDecoderOut_T_1070 = _preDecoderOut_T[1] ? preDecoders_1_io_out_pd_6_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _preDecoderOut_T_1071 = _preDecoderOut_T[2] ? preDecoders_2_io_out_pd_6_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _preDecoderOut_T_1072 = _preDecoderOut_T[3] ? preDecoders_3_io_out_pd_6_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _preDecoderOut_T_1073 = _preDecoderOut_T_1069 | _preDecoderOut_T_1070; // @[Mux.scala 27:73]
  wire [1:0] _preDecoderOut_T_1074 = _preDecoderOut_T_1073 | _preDecoderOut_T_1071; // @[Mux.scala 27:73]
  wire [1:0] preDecoderOut_pd_6_brType = _preDecoderOut_T_1074 | _preDecoderOut_T_1072; // @[Mux.scala 27:73]
  wire  preDecoderOut_pd_6_isRVC = _preDecoderOut_T[0] & preDecoders_0_io_out_pd_6_isRVC | _preDecoderOut_T[1] &
    preDecoders_1_io_out_pd_6_isRVC | _preDecoderOut_T[2] & preDecoders_2_io_out_pd_6_isRVC | _preDecoderOut_T[3] &
    preDecoders_3_io_out_pd_6_isRVC; // @[Mux.scala 27:73]
  wire  preDecoderOut_pd_6_valid = _preDecoderOut_T[0] & preDecoders_0_io_out_pd_6_valid | _preDecoderOut_T[1] &
    preDecoders_1_io_out_pd_6_valid | _preDecoderOut_T[2] & preDecoders_2_io_out_pd_6_valid | _preDecoderOut_T[3] &
    preDecoders_3_io_out_pd_6_valid; // @[Mux.scala 27:73]
  wire  preDecoderOut_pd_7_isRet = _preDecoderOut_T[0] & preDecoders_0_io_out_pd_7_isRet | _preDecoderOut_T[1] &
    preDecoders_1_io_out_pd_7_isRet | _preDecoderOut_T[2] & preDecoders_2_io_out_pd_7_isRet | _preDecoderOut_T[3] &
    preDecoders_3_io_out_pd_7_isRet; // @[Mux.scala 27:73]
  wire  preDecoderOut_pd_7_isCall = _preDecoderOut_T[0] & preDecoders_0_io_out_pd_7_isCall | _preDecoderOut_T[1] &
    preDecoders_1_io_out_pd_7_isCall | _preDecoderOut_T[2] & preDecoders_2_io_out_pd_7_isCall | _preDecoderOut_T[3] &
    preDecoders_3_io_out_pd_7_isCall; // @[Mux.scala 27:73]
  wire [1:0] _preDecoderOut_T_1104 = _preDecoderOut_T[0] ? preDecoders_0_io_out_pd_7_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _preDecoderOut_T_1105 = _preDecoderOut_T[1] ? preDecoders_1_io_out_pd_7_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _preDecoderOut_T_1106 = _preDecoderOut_T[2] ? preDecoders_2_io_out_pd_7_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _preDecoderOut_T_1107 = _preDecoderOut_T[3] ? preDecoders_3_io_out_pd_7_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _preDecoderOut_T_1108 = _preDecoderOut_T_1104 | _preDecoderOut_T_1105; // @[Mux.scala 27:73]
  wire [1:0] _preDecoderOut_T_1109 = _preDecoderOut_T_1108 | _preDecoderOut_T_1106; // @[Mux.scala 27:73]
  wire [1:0] preDecoderOut_pd_7_brType = _preDecoderOut_T_1109 | _preDecoderOut_T_1107; // @[Mux.scala 27:73]
  wire  preDecoderOut_pd_7_isRVC = _preDecoderOut_T[0] & preDecoders_0_io_out_pd_7_isRVC | _preDecoderOut_T[1] &
    preDecoders_1_io_out_pd_7_isRVC | _preDecoderOut_T[2] & preDecoders_2_io_out_pd_7_isRVC | _preDecoderOut_T[3] &
    preDecoders_3_io_out_pd_7_isRVC; // @[Mux.scala 27:73]
  wire  preDecoderOut_pd_7_valid = _preDecoderOut_T[0] & preDecoders_0_io_out_pd_7_valid | _preDecoderOut_T[1] &
    preDecoders_1_io_out_pd_7_valid | _preDecoderOut_T[2] & preDecoders_2_io_out_pd_7_valid | _preDecoderOut_T[3] &
    preDecoders_3_io_out_pd_7_valid; // @[Mux.scala 27:73]
  wire  _f2_crossPageFault_T_1 = f2_pc_0[5:0] == 6'h3e; // @[IFU.scala 282:29]
  wire  f2_crossPageFault_0 = _f2_crossPageFault_T_1 & _f2_mmio_T_2 & f2_doubleLine &
    io_icacheInter_resp_1_bits_tlbExcp_pageFault & ~preDecoderOut_pd_0_isRVC; // @[IFU.scala 346:147]
  wire  _f2_crossPageFault_T_9 = f2_pc_1[5:0] == 6'h3e; // @[IFU.scala 282:29]
  wire  f2_crossPageFault_1 = _f2_crossPageFault_T_9 & _f2_mmio_T_2 & f2_doubleLine &
    io_icacheInter_resp_1_bits_tlbExcp_pageFault & ~preDecoderOut_pd_1_isRVC; // @[IFU.scala 346:147]
  wire  _f2_crossPageFault_T_17 = f2_pc_2[5:0] == 6'h3e; // @[IFU.scala 282:29]
  wire  f2_crossPageFault_2 = _f2_crossPageFault_T_17 & _f2_mmio_T_2 & f2_doubleLine &
    io_icacheInter_resp_1_bits_tlbExcp_pageFault & ~preDecoderOut_pd_2_isRVC; // @[IFU.scala 346:147]
  wire  _f2_crossPageFault_T_25 = f2_pc_3[5:0] == 6'h3e; // @[IFU.scala 282:29]
  wire  f2_crossPageFault_3 = _f2_crossPageFault_T_25 & _f2_mmio_T_2 & f2_doubleLine &
    io_icacheInter_resp_1_bits_tlbExcp_pageFault & ~preDecoderOut_pd_3_isRVC; // @[IFU.scala 346:147]
  wire  _f2_crossPageFault_T_33 = f2_pc_4[5:0] == 6'h3e; // @[IFU.scala 282:29]
  wire  f2_crossPageFault_4 = _f2_crossPageFault_T_33 & _f2_mmio_T_2 & f2_doubleLine &
    io_icacheInter_resp_1_bits_tlbExcp_pageFault & ~preDecoderOut_pd_4_isRVC; // @[IFU.scala 346:147]
  wire  _f2_crossPageFault_T_41 = f2_pc_5[5:0] == 6'h3e; // @[IFU.scala 282:29]
  wire  f2_crossPageFault_5 = _f2_crossPageFault_T_41 & _f2_mmio_T_2 & f2_doubleLine &
    io_icacheInter_resp_1_bits_tlbExcp_pageFault & ~preDecoderOut_pd_5_isRVC; // @[IFU.scala 346:147]
  wire  _f2_crossPageFault_T_49 = f2_pc_6[5:0] == 6'h3e; // @[IFU.scala 282:29]
  wire  f2_crossPageFault_6 = _f2_crossPageFault_T_49 & _f2_mmio_T_2 & f2_doubleLine &
    io_icacheInter_resp_1_bits_tlbExcp_pageFault & ~preDecoderOut_pd_6_isRVC; // @[IFU.scala 346:147]
  wire  _f2_crossPageFault_T_57 = f2_pc_7[5:0] == 6'h3e; // @[IFU.scala 282:29]
  wire  f2_crossPageFault_7 = _f2_crossPageFault_T_57 & _f2_mmio_T_2 & f2_doubleLine &
    io_icacheInter_resp_1_bits_tlbExcp_pageFault & ~preDecoderOut_pd_7_isRVC; // @[IFU.scala 346:147]
  reg [38:0] f3_ftq_req_startAddr; // @[Reg.scala 16:16]
  reg [38:0] f3_ftq_req_nextStartAddr; // @[Reg.scala 16:16]
  reg  f3_ftq_req_ftqOffset_valid; // @[Reg.scala 16:16]
  reg [2:0] f3_ftq_req_ftqOffset_bits; // @[Reg.scala 16:16]
  reg  f3_doubleLine; // @[Reg.scala 16:16]
  wire  f3_fire = io_toIbuffer_ready & io_toIbuffer_valid; // @[Decoupled.scala 50:35]
  reg [15:0] f3_cut_data_0; // @[Reg.scala 16:16]
  reg [15:0] f3_cut_data_1; // @[Reg.scala 16:16]
  reg [15:0] f3_cut_data_2; // @[Reg.scala 16:16]
  reg [15:0] f3_cut_data_3; // @[Reg.scala 16:16]
  reg [15:0] f3_cut_data_4; // @[Reg.scala 16:16]
  reg [15:0] f3_cut_data_5; // @[Reg.scala 16:16]
  reg [15:0] f3_cut_data_6; // @[Reg.scala 16:16]
  reg [15:0] f3_cut_data_7; // @[Reg.scala 16:16]
  reg [15:0] f3_cut_data_8; // @[Reg.scala 16:16]
  reg [31:0] f3_instr_0; // @[Reg.scala 16:16]
  reg [31:0] f3_instr_1; // @[Reg.scala 16:16]
  reg [31:0] f3_instr_2; // @[Reg.scala 16:16]
  reg [31:0] f3_instr_3; // @[Reg.scala 16:16]
  reg [31:0] f3_instr_4; // @[Reg.scala 16:16]
  reg [31:0] f3_instr_5; // @[Reg.scala 16:16]
  reg [31:0] f3_instr_6; // @[Reg.scala 16:16]
  reg [31:0] f3_instr_7; // @[Reg.scala 16:16]
  reg  f3_pd_0_valid; // @[Reg.scala 16:16]
  reg  f3_pd_0_isRVC; // @[Reg.scala 16:16]
  reg [1:0] f3_pd_0_brType; // @[Reg.scala 16:16]
  reg  f3_pd_0_isCall; // @[Reg.scala 16:16]
  reg  f3_pd_0_isRet; // @[Reg.scala 16:16]
  reg  f3_pd_1_valid; // @[Reg.scala 16:16]
  reg  f3_pd_1_isRVC; // @[Reg.scala 16:16]
  reg [1:0] f3_pd_1_brType; // @[Reg.scala 16:16]
  reg  f3_pd_1_isCall; // @[Reg.scala 16:16]
  reg  f3_pd_1_isRet; // @[Reg.scala 16:16]
  reg  f3_pd_2_valid; // @[Reg.scala 16:16]
  reg  f3_pd_2_isRVC; // @[Reg.scala 16:16]
  reg [1:0] f3_pd_2_brType; // @[Reg.scala 16:16]
  reg  f3_pd_2_isCall; // @[Reg.scala 16:16]
  reg  f3_pd_2_isRet; // @[Reg.scala 16:16]
  reg  f3_pd_3_valid; // @[Reg.scala 16:16]
  reg  f3_pd_3_isRVC; // @[Reg.scala 16:16]
  reg [1:0] f3_pd_3_brType; // @[Reg.scala 16:16]
  reg  f3_pd_3_isCall; // @[Reg.scala 16:16]
  reg  f3_pd_3_isRet; // @[Reg.scala 16:16]
  reg  f3_pd_4_valid; // @[Reg.scala 16:16]
  reg  f3_pd_4_isRVC; // @[Reg.scala 16:16]
  reg [1:0] f3_pd_4_brType; // @[Reg.scala 16:16]
  reg  f3_pd_4_isCall; // @[Reg.scala 16:16]
  reg  f3_pd_4_isRet; // @[Reg.scala 16:16]
  reg  f3_pd_5_valid; // @[Reg.scala 16:16]
  reg  f3_pd_5_isRVC; // @[Reg.scala 16:16]
  reg [1:0] f3_pd_5_brType; // @[Reg.scala 16:16]
  reg  f3_pd_5_isCall; // @[Reg.scala 16:16]
  reg  f3_pd_5_isRet; // @[Reg.scala 16:16]
  reg  f3_pd_6_valid; // @[Reg.scala 16:16]
  reg  f3_pd_6_isRVC; // @[Reg.scala 16:16]
  reg [1:0] f3_pd_6_brType; // @[Reg.scala 16:16]
  reg  f3_pd_6_isCall; // @[Reg.scala 16:16]
  reg  f3_pd_6_isRet; // @[Reg.scala 16:16]
  reg  f3_pd_7_valid; // @[Reg.scala 16:16]
  reg  f3_pd_7_isRVC; // @[Reg.scala 16:16]
  reg [1:0] f3_pd_7_brType; // @[Reg.scala 16:16]
  reg  f3_pd_7_isCall; // @[Reg.scala 16:16]
  reg  f3_pd_7_isRet; // @[Reg.scala 16:16]
  reg [63:0] f3_jump_offset_0; // @[Reg.scala 16:16]
  reg [63:0] f3_jump_offset_1; // @[Reg.scala 16:16]
  reg [63:0] f3_jump_offset_2; // @[Reg.scala 16:16]
  reg [63:0] f3_jump_offset_3; // @[Reg.scala 16:16]
  reg [63:0] f3_jump_offset_4; // @[Reg.scala 16:16]
  reg [63:0] f3_jump_offset_5; // @[Reg.scala 16:16]
  reg [63:0] f3_jump_offset_6; // @[Reg.scala 16:16]
  reg [63:0] f3_jump_offset_7; // @[Reg.scala 16:16]
  reg  f3_af_vec_0; // @[Reg.scala 16:16]
  reg  f3_af_vec_1; // @[Reg.scala 16:16]
  reg  f3_af_vec_2; // @[Reg.scala 16:16]
  reg  f3_af_vec_3; // @[Reg.scala 16:16]
  reg  f3_af_vec_4; // @[Reg.scala 16:16]
  reg  f3_af_vec_5; // @[Reg.scala 16:16]
  reg  f3_af_vec_6; // @[Reg.scala 16:16]
  reg  f3_af_vec_7; // @[Reg.scala 16:16]
  reg  f3_pf_vec_0; // @[Reg.scala 16:16]
  reg  f3_pf_vec_1; // @[Reg.scala 16:16]
  reg  f3_pf_vec_2; // @[Reg.scala 16:16]
  reg  f3_pf_vec_3; // @[Reg.scala 16:16]
  reg  f3_pf_vec_4; // @[Reg.scala 16:16]
  reg  f3_pf_vec_5; // @[Reg.scala 16:16]
  reg  f3_pf_vec_6; // @[Reg.scala 16:16]
  reg  f3_pf_vec_7; // @[Reg.scala 16:16]
  reg [38:0] f3_pc_0; // @[Reg.scala 16:16]
  reg [38:0] f3_pc_1; // @[Reg.scala 16:16]
  reg [38:0] f3_pc_2; // @[Reg.scala 16:16]
  reg [38:0] f3_pc_3; // @[Reg.scala 16:16]
  reg [38:0] f3_pc_4; // @[Reg.scala 16:16]
  reg [38:0] f3_pc_5; // @[Reg.scala 16:16]
  reg [38:0] f3_pc_6; // @[Reg.scala 16:16]
  reg [38:0] f3_pc_7; // @[Reg.scala 16:16]
  reg [38:0] f3_half_snpc_0; // @[Reg.scala 16:16]
  reg [38:0] f3_half_snpc_1; // @[Reg.scala 16:16]
  reg [38:0] f3_half_snpc_2; // @[Reg.scala 16:16]
  reg [38:0] f3_half_snpc_3; // @[Reg.scala 16:16]
  reg [38:0] f3_half_snpc_4; // @[Reg.scala 16:16]
  reg [38:0] f3_half_snpc_5; // @[Reg.scala 16:16]
  reg [38:0] f3_half_snpc_6; // @[Reg.scala 16:16]
  reg [38:0] f3_half_snpc_7; // @[Reg.scala 16:16]
  reg [7:0] f3_instr_range; // @[Reg.scala 16:16]
  reg [9:0] f3_foldpc_0; // @[Reg.scala 16:16]
  reg [9:0] f3_foldpc_1; // @[Reg.scala 16:16]
  reg [9:0] f3_foldpc_2; // @[Reg.scala 16:16]
  reg [9:0] f3_foldpc_3; // @[Reg.scala 16:16]
  reg [9:0] f3_foldpc_4; // @[Reg.scala 16:16]
  reg [9:0] f3_foldpc_5; // @[Reg.scala 16:16]
  reg [9:0] f3_foldpc_6; // @[Reg.scala 16:16]
  reg [9:0] f3_foldpc_7; // @[Reg.scala 16:16]
  reg  f3_crossPageFault_0; // @[Reg.scala 16:16]
  reg  f3_crossPageFault_1; // @[Reg.scala 16:16]
  reg  f3_crossPageFault_2; // @[Reg.scala 16:16]
  reg  f3_crossPageFault_3; // @[Reg.scala 16:16]
  reg  f3_crossPageFault_4; // @[Reg.scala 16:16]
  reg  f3_crossPageFault_5; // @[Reg.scala 16:16]
  reg  f3_crossPageFault_6; // @[Reg.scala 16:16]
  reg  f3_crossPageFault_7; // @[Reg.scala 16:16]
  reg  f3_hasHalfValid_1; // @[Reg.scala 16:16]
  reg  f3_hasHalfValid_2; // @[Reg.scala 16:16]
  reg  f3_hasHalfValid_3; // @[Reg.scala 16:16]
  reg  f3_hasHalfValid_4; // @[Reg.scala 16:16]
  reg  f3_hasHalfValid_5; // @[Reg.scala 16:16]
  reg  f3_hasHalfValid_6; // @[Reg.scala 16:16]
  reg  f3_hasHalfValid_7; // @[Reg.scala 16:16]
  reg [35:0] f3_pAddrs_0; // @[Reg.scala 16:16]
  reg [38:0] f3_resend_vaddr; // @[Reg.scala 16:16]
  reg [15:0] f3_mmio_data_0; // @[IFU.scala 407:28]
  reg [15:0] f3_mmio_data_1; // @[IFU.scala 407:28]
  reg  mmio_is_RVC; // @[IFU.scala 408:32]
  reg [35:0] mmio_resend_addr; // @[IFU.scala 409:32]
  reg  mmio_resend_af; // @[IFU.scala 410:32]
  reg  mmio_resend_pf; // @[IFU.scala 411:32]
  reg  is_first_instr; // @[IFU.scala 414:31]
  wire [3:0] _io_mmioCommitRead_mmioFtqPtr_new_ptr_T_2 = _f3_wb_not_flush_T_1 + 4'h1; // @[CircularQueuePtr.scala 39:46]
  reg  io_mmioCommitRead_mmioFtqPtr_REG_flag; // @[IFU.scala 415:42]
  reg [2:0] io_mmioCommitRead_mmioFtqPtr_REG_value; // @[IFU.scala 415:42]
  wire [3:0] _mmio_commit_T = {io_rob_commits_0_bits_ftqIdx_flag,io_rob_commits_0_bits_ftqIdx_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _mmio_commit_T_2 = _mmio_commit_T == _f3_wb_not_flush_T_1; // @[CircularQueuePtr.scala 61:52]
  wire  _mmio_commit_T_5 = io_rob_commits_0_valid & _mmio_commit_T_2 & io_rob_commits_0_bits_ftqOffset == 3'h0; // @[IFU.scala 421:115]
  wire [3:0] _mmio_commit_T_6 = {io_rob_commits_1_bits_ftqIdx_flag,io_rob_commits_1_bits_ftqIdx_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _mmio_commit_T_8 = _mmio_commit_T_6 == _f3_wb_not_flush_T_1; // @[CircularQueuePtr.scala 61:52]
  wire  _mmio_commit_T_11 = io_rob_commits_1_valid & _mmio_commit_T_8 & io_rob_commits_1_bits_ftqOffset == 3'h0; // @[IFU.scala 421:115]
  wire [1:0] _mmio_commit_T_12 = {_mmio_commit_T_11,_mmio_commit_T_5}; // @[IFU.scala 421:151]
  wire  mmio_commit = |_mmio_commit_T_12; // @[IFU.scala 421:158]
  reg  f3_mmio_to_commit_next; // @[IFU.scala 425:39]
  wire  f3_mmio_can_go = _mmio_redirect_T_1 & ~f3_mmio_to_commit_next; // @[IFU.scala 426:47]
  reg  fromFtqRedirectReg_valid; // @[IFU.scala 428:38]
  reg  fromFtqRedirectReg_bits_ftqIdx_flag; // @[IFU.scala 428:38]
  reg [2:0] fromFtqRedirectReg_bits_ftqIdx_value; // @[IFU.scala 428:38]
  reg [2:0] fromFtqRedirectReg_bits_ftqOffset; // @[IFU.scala 428:38]
  reg  fromFtqRedirectReg_bits_level; // @[IFU.scala 428:38]
  reg  mmioF3Flush; // @[IFU.scala 429:38]
  wire  f3_ftq_flush_self = fromFtqRedirectReg_valid & fromFtqRedirectReg_bits_level; // @[IFU.scala 430:56]
  wire  f3_ftq_flush_by_older_differentFlag = fromFtqRedirectReg_bits_ftqIdx_flag ^ f3_ftq_req_ftqIdx_flag; // @[CircularQueuePtr.scala 92:35]
  wire  f3_ftq_flush_by_older_compare = fromFtqRedirectReg_bits_ftqIdx_value < f3_ftq_req_ftqIdx_value; // @[CircularQueuePtr.scala 93:30]
  wire  _f3_ftq_flush_by_older_T = f3_ftq_flush_by_older_differentFlag ^ f3_ftq_flush_by_older_compare; // @[CircularQueuePtr.scala 94:19]
  wire  f3_ftq_flush_by_older = fromFtqRedirectReg_valid & _f3_ftq_flush_by_older_T; // @[IFU.scala 431:56]
  wire  f3_need_not_flush = f3_req_is_mmio & fromFtqRedirectReg_valid & ~f3_ftq_flush_self & ~f3_ftq_flush_by_older; // @[IFU.scala 433:92]
  wire  _T_21 = ~f3_req_is_mmio; // @[IFU.scala 439:20]
  wire  _T_26 = ~f2_flush; // @[IFU.scala 441:24]
  wire  _GEN_1958 = f3_req_is_mmio & f3_mmio_req_commit ? 1'h0 : f3_valid; // @[IFU.scala 365:34 443:{85,95}]
  wire  _GEN_1959 = f3_fire & _T_21 ? 1'h0 : _GEN_1958; // @[IFU.scala 442:{85,95}]
  wire  _GEN_1960 = f2_fire & ~f2_flush | _GEN_1959; // @[IFU.scala 441:{85,95}]
  wire [3:0] _redirect_mmio_req_T = {fromFtqRedirectReg_bits_ftqIdx_flag,fromFtqRedirectReg_bits_ftqIdx_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _redirect_mmio_req_T_2 = _redirect_mmio_req_T == _f3_wb_not_flush_T_1; // @[CircularQueuePtr.scala 61:52]
  wire  redirect_mmio_req = fromFtqRedirectReg_valid & _redirect_mmio_req_T_2 & fromFtqRedirectReg_bits_ftqOffset == 3'h0
    ; // @[IFU.scala 448:93]
  reg  REG; // @[IFU.scala 450:15]
  wire  _GEN_1963 = redirect_mmio_req ? 1'h0 : f3_mmio_use_seq_pc; // @[IFU.scala 445:35 451:{64,85}]
  wire [3:0] _mmio_state_T = io_mmioCommitRead_mmioLastCommit ? 4'h2 : 4'h1; // @[IFU.scala 467:26]
  wire  _mmio_state_T_1 = io_uncacheInter_toUncache_ready & io_uncacheInter_toUncache_valid; // @[Decoupled.scala 50:35]
  wire [3:0] _mmio_state_T_2 = _mmio_state_T_1 ? 4'h3 : 4'h2; // @[IFU.scala 472:25]
  wire  _T_39 = io_uncacheInter_fromUncache_ready & io_uncacheInter_fromUncache_valid; // @[Decoupled.scala 50:35]
  wire  isRVC = io_uncacheInter_fromUncache_bits_data[1:0] != 2'h3; // @[IFU.scala 477:51]
  wire  needResend = ~isRVC & f3_pAddrs_0[2:1] == 2'h3; // @[IFU.scala 478:35]
  wire [3:0] _mmio_state_T_3 = needResend ? 4'h4 : 4'h9; // @[IFU.scala 479:29]
  wire [3:0] _GEN_1967 = _T_39 ? _mmio_state_T_3 : mmio_state; // @[IFU.scala 476:31 479:22 418:27]
  wire  _GEN_1968 = _T_39 ? isRVC : mmio_is_RVC; // @[IFU.scala 476:31 481:23 408:32]
  wire [15:0] _GEN_1969 = _T_39 ? io_uncacheInter_fromUncache_bits_data[15:0] : f3_mmio_data_0; // @[IFU.scala 407:28 476:31 482:29]
  wire [15:0] _GEN_1970 = _T_39 ? io_uncacheInter_fromUncache_bits_data[31:16] : f3_mmio_data_1; // @[IFU.scala 407:28 476:31 483:29]
  wire [3:0] _GEN_1971 = io_iTLBInter_req_valid & ~io_iTLBInter_resp_bits_miss ? 4'h5 : mmio_state; // @[IFU.scala 488:69 489:20 418:27]
  wire  tlbExept = io_iTLBInter_resp_bits_excp_0_pf_instr | io_iTLBInter_resp_bits_excp_0_af_instr; // @[IFU.scala 494:62]
  wire [3:0] _mmio_state_T_4 = tlbExept ? 4'h9 : 4'h6; // @[IFU.scala 496:25]
  wire  pmpExcpAF = io_pmp_resp_instr | ~io_pmp_resp_mmio; // @[IFU.scala 503:41]
  wire [3:0] _mmio_state_T_5 = pmpExcpAF ? 4'h9 : 4'h7; // @[IFU.scala 504:25]
  wire [3:0] _mmio_state_T_7 = _mmio_state_T_1 ? 4'h8 : 4'h7; // @[IFU.scala 509:25]
  wire [3:0] _GEN_1972 = _T_39 ? 4'h9 : mmio_state; // @[IFU.scala 513:31 514:22 418:27]
  wire [15:0] _GEN_1973 = _T_39 ? io_uncacheInter_fromUncache_bits_data[15:0] : f3_mmio_data_1; // @[IFU.scala 407:28 513:31 515:29]
  wire [3:0] _GEN_1974 = mmio_commit ? 4'ha : mmio_state; // @[IFU.scala 520:24 521:23 418:27]
  wire [3:0] _GEN_1975 = 4'ha == mmio_state ? 4'h0 : mmio_state; // @[IFU.scala 456:21 527:18 418:27]
  wire  _GEN_1976 = 4'ha == mmio_state ? 1'h0 : mmio_is_RVC; // @[IFU.scala 456:21 528:19 408:32]
  wire [35:0] _GEN_1977 = 4'ha == mmio_state ? 36'h0 : mmio_resend_addr; // @[IFU.scala 456:21 529:24 409:32]
  wire [3:0] _GEN_1978 = 4'h9 == mmio_state ? _GEN_1974 : _GEN_1975; // @[IFU.scala 456:21]
  wire  _GEN_1979 = 4'h9 == mmio_state ? mmio_is_RVC : _GEN_1976; // @[IFU.scala 456:21 408:32]
  wire [35:0] _GEN_1980 = 4'h9 == mmio_state ? mmio_resend_addr : _GEN_1977; // @[IFU.scala 456:21 409:32]
  wire [3:0] _GEN_1981 = 4'h8 == mmio_state ? _GEN_1972 : _GEN_1978; // @[IFU.scala 456:21]
  wire [15:0] _GEN_1982 = 4'h8 == mmio_state ? _GEN_1973 : f3_mmio_data_1; // @[IFU.scala 456:21 407:28]
  wire  _GEN_1983 = 4'h8 == mmio_state ? mmio_is_RVC : _GEN_1979; // @[IFU.scala 456:21 408:32]
  wire [35:0] _GEN_1984 = 4'h8 == mmio_state ? mmio_resend_addr : _GEN_1980; // @[IFU.scala 456:21 409:32]
  wire [3:0] _GEN_1985 = 4'h7 == mmio_state ? _mmio_state_T_7 : _GEN_1981; // @[IFU.scala 456:21 509:18]
  wire [15:0] _GEN_1986 = 4'h7 == mmio_state ? f3_mmio_data_1 : _GEN_1982; // @[IFU.scala 456:21 407:28]
  wire  _GEN_1987 = 4'h7 == mmio_state ? mmio_is_RVC : _GEN_1983; // @[IFU.scala 456:21 408:32]
  wire [35:0] _GEN_1988 = 4'h7 == mmio_state ? mmio_resend_addr : _GEN_1984; // @[IFU.scala 456:21 409:32]
  wire [3:0] _GEN_1989 = 4'h6 == mmio_state ? _mmio_state_T_5 : _GEN_1985; // @[IFU.scala 456:21 504:18]
  wire  _GEN_1990 = 4'h6 == mmio_state ? pmpExcpAF : mmio_resend_af; // @[IFU.scala 456:21 505:22 410:32]
  wire [15:0] _GEN_1991 = 4'h6 == mmio_state ? f3_mmio_data_1 : _GEN_1986; // @[IFU.scala 456:21 407:28]
  wire  _GEN_1992 = 4'h6 == mmio_state ? mmio_is_RVC : _GEN_1987; // @[IFU.scala 456:21 408:32]
  wire [35:0] _GEN_1993 = 4'h6 == mmio_state ? mmio_resend_addr : _GEN_1988; // @[IFU.scala 456:21 409:32]
  wire [3:0] _GEN_1994 = 4'h5 == mmio_state ? _mmio_state_T_4 : _GEN_1989; // @[IFU.scala 456:21 496:18]
  wire [35:0] _GEN_1995 = 4'h5 == mmio_state ? io_iTLBInter_resp_bits_paddr_0 : _GEN_1993; // @[IFU.scala 456:21 497:24]
  wire  _GEN_1996 = 4'h5 == mmio_state ? mmio_resend_af | io_iTLBInter_resp_bits_excp_0_af_instr : _GEN_1990; // @[IFU.scala 456:21 498:22]
  wire  _GEN_1997 = 4'h5 == mmio_state ? mmio_resend_pf | io_iTLBInter_resp_bits_excp_0_pf_instr : mmio_resend_pf; // @[IFU.scala 456:21 499:22 411:32]
  wire [15:0] _GEN_1998 = 4'h5 == mmio_state ? f3_mmio_data_1 : _GEN_1991; // @[IFU.scala 456:21 407:28]
  wire  _GEN_1999 = 4'h5 == mmio_state ? mmio_is_RVC : _GEN_1992; // @[IFU.scala 456:21 408:32]
  wire [3:0] _GEN_2000 = 4'h4 == mmio_state ? _GEN_1971 : _GEN_1994; // @[IFU.scala 456:21]
  wire [35:0] _GEN_2001 = 4'h4 == mmio_state ? mmio_resend_addr : _GEN_1995; // @[IFU.scala 456:21 409:32]
  wire  _GEN_2002 = 4'h4 == mmio_state ? mmio_resend_af : _GEN_1996; // @[IFU.scala 456:21 410:32]
  wire  _GEN_2003 = 4'h4 == mmio_state ? mmio_resend_pf : _GEN_1997; // @[IFU.scala 456:21 411:32]
  wire [15:0] _GEN_2004 = 4'h4 == mmio_state ? f3_mmio_data_1 : _GEN_1998; // @[IFU.scala 456:21 407:28]
  wire  _GEN_2005 = 4'h4 == mmio_state ? mmio_is_RVC : _GEN_1999; // @[IFU.scala 456:21 408:32]
  wire [3:0] _GEN_2006 = 4'h3 == mmio_state ? _GEN_1967 : _GEN_2000; // @[IFU.scala 456:21]
  wire  _GEN_2007 = 4'h3 == mmio_state ? _GEN_1968 : _GEN_2005; // @[IFU.scala 456:21]
  wire [15:0] _GEN_2008 = 4'h3 == mmio_state ? _GEN_1969 : f3_mmio_data_0; // @[IFU.scala 456:21 407:28]
  wire [15:0] _GEN_2009 = 4'h3 == mmio_state ? _GEN_1970 : _GEN_2004; // @[IFU.scala 456:21]
  wire [35:0] _GEN_2010 = 4'h3 == mmio_state ? mmio_resend_addr : _GEN_2001; // @[IFU.scala 456:21 409:32]
  wire  _GEN_2011 = 4'h3 == mmio_state ? mmio_resend_af : _GEN_2002; // @[IFU.scala 456:21 410:32]
  wire  _io_uncacheInter_toUncache_valid_T_1 = mmio_state == 4'h7; // @[IFU.scala 542:70]
  reg  f3_lastHalf_valid; // @[IFU.scala 563:34]
  wire  f3_instr_valid_1 = f3_lastHalf_valid ? f3_hasHalfValid_1 : f3_pd_1_valid; // @[IFU.scala 605:24]
  wire  f3_instr_valid_0 = f3_lastHalf_valid ? 1'h0 : f3_pd_0_valid; // @[IFU.scala 605:24]
  wire  f3_instr_valid_3 = f3_lastHalf_valid ? f3_hasHalfValid_3 : f3_pd_3_valid; // @[IFU.scala 605:24]
  wire  f3_instr_valid_2 = f3_lastHalf_valid ? f3_hasHalfValid_2 : f3_pd_2_valid; // @[IFU.scala 605:24]
  wire  f3_instr_valid_5 = f3_lastHalf_valid ? f3_hasHalfValid_5 : f3_pd_5_valid; // @[IFU.scala 605:24]
  wire  f3_instr_valid_4 = f3_lastHalf_valid ? f3_hasHalfValid_4 : f3_pd_4_valid; // @[IFU.scala 605:24]
  wire  f3_instr_valid_7 = f3_lastHalf_valid ? f3_hasHalfValid_7 : f3_pd_7_valid; // @[IFU.scala 605:24]
  wire  f3_instr_valid_6 = f3_lastHalf_valid ? f3_hasHalfValid_6 : f3_pd_6_valid; // @[IFU.scala 605:24]
  wire [7:0] _T_59 = {f3_instr_valid_7,f3_instr_valid_6,f3_instr_valid_5,f3_instr_valid_4,f3_instr_valid_3,
    f3_instr_valid_2,f3_instr_valid_1,f3_instr_valid_0}; // @[IFU.scala 574:51]
  wire  _f3_last_validIdx_T_1 = predChecker_io_out_stage1Out_fixedRange_7 ? 1'h0 : 1'h1; // @[ParallelMux.scala 90:77]
  wire [1:0] _f3_last_validIdx_T_3 = predChecker_io_out_stage1Out_fixedRange_5 ? 2'h2 : 2'h3; // @[ParallelMux.scala 90:77]
  wire [1:0] _f3_last_validIdx_T_5 = predChecker_io_out_stage1Out_fixedRange_7 |
    predChecker_io_out_stage1Out_fixedRange_6 ? {{1'd0}, _f3_last_validIdx_T_1} : _f3_last_validIdx_T_3; // @[ParallelMux.scala 90:77]
  wire [2:0] _f3_last_validIdx_T_7 = predChecker_io_out_stage1Out_fixedRange_3 ? 3'h4 : 3'h5; // @[ParallelMux.scala 90:77]
  wire [2:0] _f3_last_validIdx_T_9 = predChecker_io_out_stage1Out_fixedRange_1 ? 3'h6 : 3'h7; // @[ParallelMux.scala 90:77]
  wire [2:0] _f3_last_validIdx_T_11 = predChecker_io_out_stage1Out_fixedRange_3 |
    predChecker_io_out_stage1Out_fixedRange_2 ? _f3_last_validIdx_T_7 : _f3_last_validIdx_T_9; // @[ParallelMux.scala 90:77]
  wire [2:0] _f3_last_validIdx_T_13 = predChecker_io_out_stage1Out_fixedRange_7 |
    predChecker_io_out_stage1Out_fixedRange_6 | (predChecker_io_out_stage1Out_fixedRange_5 |
    predChecker_io_out_stage1Out_fixedRange_4) ? {{1'd0}, _f3_last_validIdx_T_5} : _f3_last_validIdx_T_11; // @[ParallelMux.scala 90:77]
  wire [2:0] f3_last_validIdx = ~_f3_last_validIdx_T_13; // @[IFU.scala 585:38]
  wire  f3_hasLastHalf = ~f3_pd_7_isRVC & predChecker_io_out_stage1Out_fixedRange_7 & f3_instr_valid_7 & ~
    predChecker_io_out_stage1Out_fixedTaken_7 & _T_21; // @[IFU.scala 582:119]
  wire  _GEN_2041 = 3'h1 == f3_last_validIdx ? f3_pd_1_isRVC : f3_pd_0_isRVC; // @[IFU.scala 582:{5,5}]
  wire  _GEN_2042 = 3'h2 == f3_last_validIdx ? f3_pd_2_isRVC : _GEN_2041; // @[IFU.scala 582:{5,5}]
  wire  _GEN_2043 = 3'h3 == f3_last_validIdx ? f3_pd_3_isRVC : _GEN_2042; // @[IFU.scala 582:{5,5}]
  wire  _GEN_2044 = 3'h4 == f3_last_validIdx ? f3_pd_4_isRVC : _GEN_2043; // @[IFU.scala 582:{5,5}]
  wire  _GEN_2045 = 3'h5 == f3_last_validIdx ? f3_pd_5_isRVC : _GEN_2044; // @[IFU.scala 582:{5,5}]
  wire  _GEN_2046 = 3'h6 == f3_last_validIdx ? f3_pd_6_isRVC : _GEN_2045; // @[IFU.scala 582:{5,5}]
  wire  _GEN_2047 = 3'h7 == f3_last_validIdx ? f3_pd_7_isRVC : _GEN_2046; // @[IFU.scala 582:{5,5}]
  wire  _GEN_2049 = 3'h1 == f3_last_validIdx ? predChecker_io_out_stage1Out_fixedRange_1 :
    predChecker_io_out_stage1Out_fixedRange_0; // @[IFU.scala 582:{23,23}]
  wire  _GEN_2050 = 3'h2 == f3_last_validIdx ? predChecker_io_out_stage1Out_fixedRange_2 : _GEN_2049; // @[IFU.scala 582:{23,23}]
  wire  _GEN_2051 = 3'h3 == f3_last_validIdx ? predChecker_io_out_stage1Out_fixedRange_3 : _GEN_2050; // @[IFU.scala 582:{23,23}]
  wire  _GEN_2052 = 3'h4 == f3_last_validIdx ? predChecker_io_out_stage1Out_fixedRange_4 : _GEN_2051; // @[IFU.scala 582:{23,23}]
  wire  _GEN_2053 = 3'h5 == f3_last_validIdx ? predChecker_io_out_stage1Out_fixedRange_5 : _GEN_2052; // @[IFU.scala 582:{23,23}]
  wire  _GEN_2054 = 3'h6 == f3_last_validIdx ? predChecker_io_out_stage1Out_fixedRange_6 : _GEN_2053; // @[IFU.scala 582:{23,23}]
  wire  _GEN_2055 = 3'h7 == f3_last_validIdx ? predChecker_io_out_stage1Out_fixedRange_7 : _GEN_2054; // @[IFU.scala 582:{23,23}]
  wire  _GEN_2057 = 3'h1 == f3_last_validIdx ? f3_instr_valid_1 : f3_instr_valid_0; // @[IFU.scala 582:{59,59}]
  wire  _GEN_2058 = 3'h2 == f3_last_validIdx ? f3_instr_valid_2 : _GEN_2057; // @[IFU.scala 582:{59,59}]
  wire  _GEN_2059 = 3'h3 == f3_last_validIdx ? f3_instr_valid_3 : _GEN_2058; // @[IFU.scala 582:{59,59}]
  wire  _GEN_2060 = 3'h4 == f3_last_validIdx ? f3_instr_valid_4 : _GEN_2059; // @[IFU.scala 582:{59,59}]
  wire  _GEN_2061 = 3'h5 == f3_last_validIdx ? f3_instr_valid_5 : _GEN_2060; // @[IFU.scala 582:{59,59}]
  wire  _GEN_2062 = 3'h6 == f3_last_validIdx ? f3_instr_valid_6 : _GEN_2061; // @[IFU.scala 582:{59,59}]
  wire  _GEN_2063 = 3'h7 == f3_last_validIdx ? f3_instr_valid_7 : _GEN_2062; // @[IFU.scala 582:{59,59}]
  wire  _GEN_2065 = 3'h1 == f3_last_validIdx ? predChecker_io_out_stage1Out_fixedTaken_1 :
    predChecker_io_out_stage1Out_fixedTaken_0; // @[IFU.scala 582:{85,85}]
  wire  _GEN_2066 = 3'h2 == f3_last_validIdx ? predChecker_io_out_stage1Out_fixedTaken_2 : _GEN_2065; // @[IFU.scala 582:{85,85}]
  wire  _GEN_2067 = 3'h3 == f3_last_validIdx ? predChecker_io_out_stage1Out_fixedTaken_3 : _GEN_2066; // @[IFU.scala 582:{85,85}]
  wire  _GEN_2068 = 3'h4 == f3_last_validIdx ? predChecker_io_out_stage1Out_fixedTaken_4 : _GEN_2067; // @[IFU.scala 582:{85,85}]
  wire  _GEN_2069 = 3'h5 == f3_last_validIdx ? predChecker_io_out_stage1Out_fixedTaken_5 : _GEN_2068; // @[IFU.scala 582:{85,85}]
  wire  _GEN_2070 = 3'h6 == f3_last_validIdx ? predChecker_io_out_stage1Out_fixedTaken_6 : _GEN_2069; // @[IFU.scala 582:{85,85}]
  wire  _GEN_2071 = 3'h7 == f3_last_validIdx ? predChecker_io_out_stage1Out_fixedTaken_7 : _GEN_2070; // @[IFU.scala 582:{85,85}]
  reg  f3_lastHalf_disable; // @[IFU.scala 592:36]
  wire  _GEN_2072 = f3_flush | f3_fire & f3_lastHalf_disable ? 1'h0 : f3_lastHalf_disable; // @[IFU.scala 594:53 595:25 592:36]
  wire  _io_toIbuffer_valid_T_3 = ~f3_flush; // @[IFU.scala 619:87]
  wire [7:0] _io_toIbuffer_bits_enqEnable_T = {predChecker_io_out_stage1Out_fixedRange_7,
    predChecker_io_out_stage1Out_fixedRange_6,predChecker_io_out_stage1Out_fixedRange_5,
    predChecker_io_out_stage1Out_fixedRange_4,predChecker_io_out_stage1Out_fixedRange_3,
    predChecker_io_out_stage1Out_fixedRange_2,predChecker_io_out_stage1Out_fixedRange_1,
    predChecker_io_out_stage1Out_fixedRange_0}; // @[IFU.scala 622:64]
  wire [7:0] _io_toIbuffer_bits_enqEnable_T_2 = _io_toIbuffer_bits_enqEnable_T & _T_59; // @[IFU.scala 622:71]
  wire [7:0] _io_toIbuffer_bits_enqEnable_T_6 = _io_toIbuffer_bits_enqEnable_T_2 & 8'hfe; // @[IFU.scala 634:95]
  wire [7:0] _io_toIbuffer_bits_valid_T_2 = 8'hfe & _T_59; // @[IFU.scala 635:53]
  wire [7:0] _GEN_2077 = f3_lastHalf_valid ? _io_toIbuffer_bits_enqEnable_T_6 : _io_toIbuffer_bits_enqEnable_T_2; // @[IFU.scala 633:26 622:33 634:33]
  reg  mmioFlushWb_valid_REG; // @[IFU.scala 649:91]
  wire  mmioFlushWb_valid = _mmio_redirect_T_1 & mmioFlushWb_valid_REG & f3_mmio_use_seq_pc; // @[IFU.scala 649:113]
  wire [38:0] _mmioFlushWb_bits_target_T_1 = f3_ftq_req_startAddr + 39'h2; // @[IFU.scala 657:72]
  wire [38:0] _mmioFlushWb_bits_target_T_3 = f3_ftq_req_startAddr + 39'h4; // @[IFU.scala 657:101]
  wire [38:0] mmioFlushWb_bits_target = mmio_is_RVC ? _mmioFlushWb_bits_target_T_1 : _mmioFlushWb_bits_target_T_3; // @[IFU.scala 657:37]
  wire [31:0] inst = {f3_mmio_data_1,f3_mmio_data_0}; // @[Cat.scala 31:58]
  wire  currentIsRVC = inst[1:0] != 2'h3; // @[PreDecode.scala 30:38]
  wire [31:0] _brType_T = inst & 32'he003; // @[Lookup.scala 31:38]
  wire  _brType_T_1 = 32'ha001 == _brType_T; // @[Lookup.scala 31:38]
  wire [31:0] _brType_T_2 = inst & 32'he07f; // @[Lookup.scala 31:38]
  wire  _brType_T_3 = 32'h8002 == _brType_T_2; // @[Lookup.scala 31:38]
  wire [31:0] _brType_T_4 = inst & 32'hc003; // @[Lookup.scala 31:38]
  wire  _brType_T_5 = 32'hc001 == _brType_T_4; // @[Lookup.scala 31:38]
  wire [31:0] _brType_T_6 = inst & 32'h7f; // @[Lookup.scala 31:38]
  wire  _brType_T_7 = 32'h6f == _brType_T_6; // @[Lookup.scala 31:38]
  wire [31:0] _brType_T_8 = inst & 32'h707f; // @[Lookup.scala 31:38]
  wire  _brType_T_9 = 32'h67 == _brType_T_8; // @[Lookup.scala 31:38]
  wire  _brType_T_11 = 32'h63 == _brType_T_6; // @[Lookup.scala 31:38]
  wire [1:0] _brType_T_13 = _brType_T_9 ? 2'h3 : {{1'd0}, _brType_T_11}; // @[Lookup.scala 34:39]
  wire [1:0] _brType_T_14 = _brType_T_7 ? 2'h2 : _brType_T_13; // @[Lookup.scala 34:39]
  wire [1:0] _brType_T_15 = _brType_T_5 ? 2'h1 : _brType_T_14; // @[Lookup.scala 34:39]
  wire [1:0] _brType_T_16 = _brType_T_3 ? 2'h3 : _brType_T_15; // @[Lookup.scala 34:39]
  wire [1:0] brType = _brType_T_1 ? 2'h2 : _brType_T_16; // @[Lookup.scala 34:39]
  wire [4:0] rd = currentIsRVC ? {{4'd0}, inst[12]} : inst[11:7]; // @[PreDecode.scala 34:17]
  wire  _rs_T_2 = brType == 2'h2; // @[PreDecode.scala 35:43]
  wire [4:0] _rs_T_4 = brType == 2'h2 ? 5'h0 : inst[11:7]; // @[PreDecode.scala 35:35]
  wire [4:0] rs = currentIsRVC ? _rs_T_4 : inst[19:15]; // @[PreDecode.scala 35:17]
  wire  _isCall_T_5 = brType == 2'h3; // @[PreDecode.scala 36:68]
  wire  _isCall_T_9 = rd == 5'h1 | rd == 5'h5; // @[PreDecode.scala 31:38]
  wire  isCall = (_rs_T_2 & ~currentIsRVC | brType == 2'h3) & _isCall_T_9; // @[PreDecode.scala 36:85]
  wire  _isRet_T_3 = rs == 5'h1 | rs == 5'h5; // @[PreDecode.scala 31:38]
  wire  isRet = _isCall_T_5 & _isRet_T_3 & ~isCall; // @[PreDecode.scala 37:54]
  wire [2:0] brOffset_rvc_offset_hi_hi = {inst[12],inst[6:5]}; // @[Cat.scala 31:58]
  wire [6:0] io_toIbuffer_bits_instrs_0_s_opc = |inst[12:5] ? 7'h13 : 7'h1f; // @[RVC.scala 53:20]
  wire [29:0] _io_toIbuffer_bits_instrs_0_s_T_7 = {inst[10:7],inst[12:11],inst[5],inst[6],2'h0,5'h2,3'h0,2'h1,inst[4:2],
    io_toIbuffer_bits_instrs_0_s_opc}; // @[Cat.scala 31:58]
  wire [7:0] _io_toIbuffer_bits_instrs_0_s_T_15 = {inst[6:5],inst[12:10],3'h0}; // @[Cat.scala 31:58]
  wire [27:0] _io_toIbuffer_bits_instrs_0_s_T_20 = {inst[6:5],inst[12:10],3'h0,2'h1,inst[9:7],3'h3,2'h1,inst[4:2],7'h7}; // @[Cat.scala 31:58]
  wire [6:0] _io_toIbuffer_bits_instrs_0_s_T_31 = {inst[5],inst[12:10],inst[6],2'h0}; // @[Cat.scala 31:58]
  wire [26:0] _io_toIbuffer_bits_instrs_0_s_T_36 = {inst[5],inst[12:10],inst[6],2'h0,2'h1,inst[9:7],3'h2,2'h1,inst[4:2],7'h3
    }; // @[Cat.scala 31:58]
  wire [27:0] _io_toIbuffer_bits_instrs_0_s_T_51 = {inst[6:5],inst[12:10],3'h0,2'h1,inst[9:7],3'h3,2'h1,inst[4:2],7'h3}; // @[Cat.scala 31:58]
  wire [26:0] _io_toIbuffer_bits_instrs_0_s_T_73 = {_io_toIbuffer_bits_instrs_0_s_T_31[6:5],2'h1,inst[4:2],2'h1,inst[9:7
    ],3'h2,_io_toIbuffer_bits_instrs_0_s_T_31[4:0],7'h3f}; // @[Cat.scala 31:58]
  wire [27:0] _io_toIbuffer_bits_instrs_0_s_T_93 = {_io_toIbuffer_bits_instrs_0_s_T_15[7:5],2'h1,inst[4:2],2'h1,inst[9:7
    ],3'h3,_io_toIbuffer_bits_instrs_0_s_T_15[4:0],7'h27}; // @[Cat.scala 31:58]
  wire [26:0] _io_toIbuffer_bits_instrs_0_s_T_115 = {_io_toIbuffer_bits_instrs_0_s_T_31[6:5],2'h1,inst[4:2],2'h1,inst[9:
    7],3'h2,_io_toIbuffer_bits_instrs_0_s_T_31[4:0],7'h23}; // @[Cat.scala 31:58]
  wire [27:0] _io_toIbuffer_bits_instrs_0_s_T_135 = {_io_toIbuffer_bits_instrs_0_s_T_15[7:5],2'h1,inst[4:2],2'h1,inst[9:
    7],3'h3,_io_toIbuffer_bits_instrs_0_s_T_15[4:0],7'h23}; // @[Cat.scala 31:58]
  wire [6:0] _io_toIbuffer_bits_instrs_0_s_T_145 = inst[12] ? 7'h7f : 7'h0; // @[Bitwise.scala 74:12]
  wire [11:0] _io_toIbuffer_bits_instrs_0_s_T_147 = {_io_toIbuffer_bits_instrs_0_s_T_145,inst[6:2]}; // @[Cat.scala 31:58]
  wire [31:0] io_toIbuffer_bits_instrs_0_s_8_bits = {_io_toIbuffer_bits_instrs_0_s_T_145,inst[6:2],inst[11:7],3'h0,inst[
    11:7],7'h13}; // @[Cat.scala 31:58]
  wire  _io_toIbuffer_bits_instrs_0_s_opc_T_3 = |inst[11:7]; // @[RVC.scala 77:24]
  wire [6:0] io_toIbuffer_bits_instrs_0_s_opc_1 = |inst[11:7] ? 7'h1b : 7'h1f; // @[RVC.scala 77:20]
  wire [31:0] io_toIbuffer_bits_instrs_0_s_9_bits = {_io_toIbuffer_bits_instrs_0_s_T_145,inst[6:2],inst[11:7],3'h0,inst[
    11:7],io_toIbuffer_bits_instrs_0_s_opc_1}; // @[Cat.scala 31:58]
  wire [31:0] io_toIbuffer_bits_instrs_0_s_10_bits = {_io_toIbuffer_bits_instrs_0_s_T_145,inst[6:2],5'h0,3'h0,inst[11:7]
    ,7'h13}; // @[Cat.scala 31:58]
  wire  _io_toIbuffer_bits_instrs_0_s_opc_T_9 = |_io_toIbuffer_bits_instrs_0_s_T_147; // @[RVC.scala 90:29]
  wire [6:0] io_toIbuffer_bits_instrs_0_s_opc_2 = |_io_toIbuffer_bits_instrs_0_s_T_147 ? 7'h37 : 7'h3f; // @[RVC.scala 90:20]
  wire [14:0] _io_toIbuffer_bits_instrs_0_s_me_T_2 = inst[12] ? 15'h7fff : 15'h0; // @[Bitwise.scala 74:12]
  wire [31:0] _io_toIbuffer_bits_instrs_0_s_me_T_4 = {_io_toIbuffer_bits_instrs_0_s_me_T_2,inst[6:2],12'h0}; // @[Cat.scala 31:58]
  wire [31:0] io_toIbuffer_bits_instrs_0_s_me_bits = {_io_toIbuffer_bits_instrs_0_s_me_T_4[31:12],inst[11:7],
    io_toIbuffer_bits_instrs_0_s_opc_2}; // @[Cat.scala 31:58]
  wire [6:0] io_toIbuffer_bits_instrs_0_s_opc_3 = _io_toIbuffer_bits_instrs_0_s_opc_T_9 ? 7'h13 : 7'h1f; // @[RVC.scala 86:20]
  wire [2:0] _io_toIbuffer_bits_instrs_0_s_T_187 = inst[12] ? 3'h7 : 3'h0; // @[Bitwise.scala 74:12]
  wire [31:0] io_toIbuffer_bits_instrs_0_s_res_bits = {_io_toIbuffer_bits_instrs_0_s_T_187,inst[4:3],inst[5],inst[2],
    inst[6],4'h0,inst[11:7],3'h0,inst[11:7],io_toIbuffer_bits_instrs_0_s_opc_3}; // @[Cat.scala 31:58]
  wire [31:0] io_toIbuffer_bits_instrs_0_s_11_bits = inst[11:7] == 5'h0 | inst[11:7] == 5'h2 ?
    io_toIbuffer_bits_instrs_0_s_res_bits : io_toIbuffer_bits_instrs_0_s_me_bits; // @[RVC.scala 92:10]
  wire [25:0] _io_toIbuffer_bits_instrs_0_s_T_208 = {inst[12],inst[6:2],2'h1,inst[9:7],3'h5,2'h1,inst[9:7],7'h13}; // @[Cat.scala 31:58]
  wire [30:0] _GEN_2128 = {{5'd0}, _io_toIbuffer_bits_instrs_0_s_T_208}; // @[RVC.scala 99:23]
  wire [30:0] _io_toIbuffer_bits_instrs_0_s_T_217 = _GEN_2128 | 31'h40000000; // @[RVC.scala 99:23]
  wire [31:0] _io_toIbuffer_bits_instrs_0_s_T_227 = {_io_toIbuffer_bits_instrs_0_s_T_145,inst[6:2],2'h1,inst[9:7],3'h7,2'h1
    ,inst[9:7],7'h13}; // @[Cat.scala 31:58]
  wire [2:0] _io_toIbuffer_bits_instrs_0_s_funct_T_4 = brOffset_rvc_offset_hi_hi == 3'h1 ? 3'h4 : 3'h0; // @[package.scala 32:76]
  wire [2:0] _io_toIbuffer_bits_instrs_0_s_funct_T_6 = brOffset_rvc_offset_hi_hi == 3'h2 ? 3'h6 :
    _io_toIbuffer_bits_instrs_0_s_funct_T_4; // @[package.scala 32:76]
  wire [2:0] _io_toIbuffer_bits_instrs_0_s_funct_T_8 = brOffset_rvc_offset_hi_hi == 3'h3 ? 3'h7 :
    _io_toIbuffer_bits_instrs_0_s_funct_T_6; // @[package.scala 32:76]
  wire [2:0] _io_toIbuffer_bits_instrs_0_s_funct_T_10 = brOffset_rvc_offset_hi_hi == 3'h4 ? 3'h0 :
    _io_toIbuffer_bits_instrs_0_s_funct_T_8; // @[package.scala 32:76]
  wire [2:0] _io_toIbuffer_bits_instrs_0_s_funct_T_12 = brOffset_rvc_offset_hi_hi == 3'h5 ? 3'h0 :
    _io_toIbuffer_bits_instrs_0_s_funct_T_10; // @[package.scala 32:76]
  wire [2:0] _io_toIbuffer_bits_instrs_0_s_funct_T_14 = brOffset_rvc_offset_hi_hi == 3'h6 ? 3'h2 :
    _io_toIbuffer_bits_instrs_0_s_funct_T_12; // @[package.scala 32:76]
  wire [2:0] io_toIbuffer_bits_instrs_0_s_funct = brOffset_rvc_offset_hi_hi == 3'h7 ? 3'h3 :
    _io_toIbuffer_bits_instrs_0_s_funct_T_14; // @[package.scala 32:76]
  wire [30:0] io_toIbuffer_bits_instrs_0_s_sub = inst[6:5] == 2'h0 ? 31'h40000000 : 31'h0; // @[RVC.scala 103:22]
  wire [6:0] io_toIbuffer_bits_instrs_0_s_opc_4 = inst[12] ? 7'h3b : 7'h33; // @[RVC.scala 104:22]
  wire [24:0] _io_toIbuffer_bits_instrs_0_s_T_234 = {2'h1,inst[4:2],2'h1,inst[9:7],io_toIbuffer_bits_instrs_0_s_funct,2'h1
    ,inst[9:7],io_toIbuffer_bits_instrs_0_s_opc_4}; // @[Cat.scala 31:58]
  wire [30:0] _GEN_2129 = {{6'd0}, _io_toIbuffer_bits_instrs_0_s_T_234}; // @[RVC.scala 105:43]
  wire [30:0] _io_toIbuffer_bits_instrs_0_s_T_235 = _GEN_2129 | io_toIbuffer_bits_instrs_0_s_sub; // @[RVC.scala 105:43]
  wire [30:0] _io_toIbuffer_bits_instrs_0_s_T_238 = inst[11:10] == 2'h1 ? _io_toIbuffer_bits_instrs_0_s_T_217 : {{5
    'd0}, _io_toIbuffer_bits_instrs_0_s_T_208}; // @[package.scala 32:76]
  wire [31:0] _io_toIbuffer_bits_instrs_0_s_T_240 = inst[11:10] == 2'h2 ? _io_toIbuffer_bits_instrs_0_s_T_227 : {{1
    'd0}, _io_toIbuffer_bits_instrs_0_s_T_238}; // @[package.scala 32:76]
  wire [31:0] io_toIbuffer_bits_instrs_0_s_12_bits = inst[11:10] == 2'h3 ? {{1'd0}, _io_toIbuffer_bits_instrs_0_s_T_235}
     : _io_toIbuffer_bits_instrs_0_s_T_240; // @[package.scala 32:76]
  wire [9:0] _io_toIbuffer_bits_instrs_0_s_T_252 = inst[12] ? 10'h3ff : 10'h0; // @[Bitwise.scala 74:12]
  wire [20:0] _io_toIbuffer_bits_instrs_0_s_T_260 = {_io_toIbuffer_bits_instrs_0_s_T_252,inst[8],inst[10:9],inst[6],inst
    [7],inst[2],inst[11],inst[5:3],1'h0}; // @[Cat.scala 31:58]
  wire [31:0] io_toIbuffer_bits_instrs_0_s_13_bits = {_io_toIbuffer_bits_instrs_0_s_T_260[20],
    _io_toIbuffer_bits_instrs_0_s_T_260[10:1],_io_toIbuffer_bits_instrs_0_s_T_260[11],
    _io_toIbuffer_bits_instrs_0_s_T_260[19:12],5'h0,7'h6f}; // @[Cat.scala 31:58]
  wire [4:0] _io_toIbuffer_bits_instrs_0_s_T_306 = inst[12] ? 5'h1f : 5'h0; // @[Bitwise.scala 74:12]
  wire [12:0] _io_toIbuffer_bits_instrs_0_s_T_311 = {_io_toIbuffer_bits_instrs_0_s_T_306,inst[6:5],inst[2],inst[11:10],
    inst[4:3],1'h0}; // @[Cat.scala 31:58]
  wire [31:0] io_toIbuffer_bits_instrs_0_s_14_bits = {_io_toIbuffer_bits_instrs_0_s_T_311[12],
    _io_toIbuffer_bits_instrs_0_s_T_311[10:5],5'h0,2'h1,inst[9:7],3'h0,_io_toIbuffer_bits_instrs_0_s_T_311[4:1],
    _io_toIbuffer_bits_instrs_0_s_T_311[11],7'h63}; // @[Cat.scala 31:58]
  wire [31:0] io_toIbuffer_bits_instrs_0_s_15_bits = {_io_toIbuffer_bits_instrs_0_s_T_311[12],
    _io_toIbuffer_bits_instrs_0_s_T_311[10:5],5'h0,2'h1,inst[9:7],3'h1,_io_toIbuffer_bits_instrs_0_s_T_311[4:1],
    _io_toIbuffer_bits_instrs_0_s_T_311[11],7'h63}; // @[Cat.scala 31:58]
  wire [6:0] io_toIbuffer_bits_instrs_0_s_load_opc = _io_toIbuffer_bits_instrs_0_s_opc_T_3 ? 7'h3 : 7'h1f; // @[RVC.scala 113:23]
  wire [25:0] _io_toIbuffer_bits_instrs_0_s_T_395 = {inst[12],inst[6:2],inst[11:7],3'h1,inst[11:7],7'h13}; // @[Cat.scala 31:58]
  wire [28:0] _io_toIbuffer_bits_instrs_0_s_T_405 = {inst[4:2],inst[12],inst[6:5],3'h0,5'h2,3'h3,inst[11:7],7'h7}; // @[Cat.scala 31:58]
  wire [27:0] _io_toIbuffer_bits_instrs_0_s_T_414 = {inst[3:2],inst[12],inst[6:4],2'h0,5'h2,3'h2,inst[11:7],
    io_toIbuffer_bits_instrs_0_s_load_opc}; // @[Cat.scala 31:58]
  wire [28:0] _io_toIbuffer_bits_instrs_0_s_T_423 = {inst[4:2],inst[12],inst[6:5],3'h0,5'h2,3'h3,inst[11:7],
    io_toIbuffer_bits_instrs_0_s_load_opc}; // @[Cat.scala 31:58]
  wire [19:0] _io_toIbuffer_bits_instrs_0_s_mv_T_2 = {inst[6:2],3'h0,inst[11:7],7'h13}; // @[Cat.scala 31:58]
  wire [24:0] _io_toIbuffer_bits_instrs_0_s_add_T_3 = {inst[6:2],inst[11:7],3'h0,inst[11:7],7'h33}; // @[Cat.scala 31:58]
  wire [24:0] io_toIbuffer_bits_instrs_0_s_jr = {inst[6:2],inst[11:7],3'h0,12'h67}; // @[Cat.scala 31:58]
  wire [24:0] io_toIbuffer_bits_instrs_0_s_reserved = {io_toIbuffer_bits_instrs_0_s_jr[24:7],7'h1f}; // @[Cat.scala 31:58]
  wire [24:0] _io_toIbuffer_bits_instrs_0_s_jr_reserved_T_2 = _io_toIbuffer_bits_instrs_0_s_opc_T_3 ?
    io_toIbuffer_bits_instrs_0_s_jr : io_toIbuffer_bits_instrs_0_s_reserved; // @[RVC.scala 134:33]
  wire  _io_toIbuffer_bits_instrs_0_s_jr_mv_T_1 = |inst[6:2]; // @[RVC.scala 135:27]
  wire [31:0] io_toIbuffer_bits_instrs_0_s_mv_bits = {{12'd0}, _io_toIbuffer_bits_instrs_0_s_mv_T_2}; // @[RVC.scala 21:19 22:14]
  wire [31:0] io_toIbuffer_bits_instrs_0_s_jr_reserved_bits = {{7'd0}, _io_toIbuffer_bits_instrs_0_s_jr_reserved_T_2}; // @[RVC.scala 21:19 22:14]
  wire [31:0] io_toIbuffer_bits_instrs_0_s_jr_mv_bits = |inst[6:2] ? io_toIbuffer_bits_instrs_0_s_mv_bits :
    io_toIbuffer_bits_instrs_0_s_jr_reserved_bits; // @[RVC.scala 135:22]
  wire [24:0] io_toIbuffer_bits_instrs_0_s_jalr = {inst[6:2],inst[11:7],3'h0,12'he7}; // @[Cat.scala 31:58]
  wire [24:0] _io_toIbuffer_bits_instrs_0_s_ebreak_T_1 = {io_toIbuffer_bits_instrs_0_s_jr[24:7],7'h73}; // @[Cat.scala 31:58]
  wire [24:0] io_toIbuffer_bits_instrs_0_s_ebreak = _io_toIbuffer_bits_instrs_0_s_ebreak_T_1 | 25'h100000; // @[RVC.scala 137:46]
  wire [24:0] _io_toIbuffer_bits_instrs_0_s_jalr_ebreak_T_2 = _io_toIbuffer_bits_instrs_0_s_opc_T_3 ?
    io_toIbuffer_bits_instrs_0_s_jalr : io_toIbuffer_bits_instrs_0_s_ebreak; // @[RVC.scala 138:33]
  wire [31:0] io_toIbuffer_bits_instrs_0_s_add_bits = {{7'd0}, _io_toIbuffer_bits_instrs_0_s_add_T_3}; // @[RVC.scala 21:19 22:14]
  wire [31:0] io_toIbuffer_bits_instrs_0_s_jalr_ebreak_bits = {{7'd0}, _io_toIbuffer_bits_instrs_0_s_jalr_ebreak_T_2}; // @[RVC.scala 21:19 22:14]
  wire [31:0] io_toIbuffer_bits_instrs_0_s_jalr_add_bits = _io_toIbuffer_bits_instrs_0_s_jr_mv_T_1 ?
    io_toIbuffer_bits_instrs_0_s_add_bits : io_toIbuffer_bits_instrs_0_s_jalr_ebreak_bits; // @[RVC.scala 139:25]
  wire [31:0] io_toIbuffer_bits_instrs_0_s_20_bits = inst[12] ? io_toIbuffer_bits_instrs_0_s_jalr_add_bits :
    io_toIbuffer_bits_instrs_0_s_jr_mv_bits; // @[RVC.scala 140:10]
  wire [8:0] _io_toIbuffer_bits_instrs_0_s_T_430 = {inst[9:7],inst[12:10],3'h0}; // @[Cat.scala 31:58]
  wire [28:0] _io_toIbuffer_bits_instrs_0_s_T_437 = {_io_toIbuffer_bits_instrs_0_s_T_430[8:5],inst[6:2],5'h2,3'h3,
    _io_toIbuffer_bits_instrs_0_s_T_430[4:0],7'h27}; // @[Cat.scala 31:58]
  wire [7:0] _io_toIbuffer_bits_instrs_0_s_T_443 = {inst[8:7],inst[12:9],2'h0}; // @[Cat.scala 31:58]
  wire [27:0] _io_toIbuffer_bits_instrs_0_s_T_450 = {_io_toIbuffer_bits_instrs_0_s_T_443[7:5],inst[6:2],5'h2,3'h2,
    _io_toIbuffer_bits_instrs_0_s_T_443[4:0],7'h23}; // @[Cat.scala 31:58]
  wire [28:0] _io_toIbuffer_bits_instrs_0_s_T_463 = {_io_toIbuffer_bits_instrs_0_s_T_430[8:5],inst[6:2],5'h2,3'h3,
    _io_toIbuffer_bits_instrs_0_s_T_430[4:0],7'h23}; // @[Cat.scala 31:58]
  wire [4:0] _io_toIbuffer_bits_instrs_0_T_2 = {inst[1:0],inst[15:13]}; // @[Cat.scala 31:58]
  wire [31:0] io_toIbuffer_bits_instrs_0_s_1_bits = {{4'd0}, _io_toIbuffer_bits_instrs_0_s_T_20}; // @[RVC.scala 21:19 22:14]
  wire [31:0] io_toIbuffer_bits_instrs_0_s_0_bits = {{2'd0}, _io_toIbuffer_bits_instrs_0_s_T_7}; // @[RVC.scala 21:19 22:14]
  wire [31:0] _io_toIbuffer_bits_instrs_0_T_4_bits = _io_toIbuffer_bits_instrs_0_T_2 == 5'h1 ?
    io_toIbuffer_bits_instrs_0_s_1_bits : io_toIbuffer_bits_instrs_0_s_0_bits; // @[package.scala 32:76]
  wire [31:0] io_toIbuffer_bits_instrs_0_s_2_bits = {{5'd0}, _io_toIbuffer_bits_instrs_0_s_T_36}; // @[RVC.scala 21:19 22:14]
  wire [31:0] _io_toIbuffer_bits_instrs_0_T_6_bits = _io_toIbuffer_bits_instrs_0_T_2 == 5'h2 ?
    io_toIbuffer_bits_instrs_0_s_2_bits : _io_toIbuffer_bits_instrs_0_T_4_bits; // @[package.scala 32:76]
  wire [31:0] io_toIbuffer_bits_instrs_0_s_3_bits = {{4'd0}, _io_toIbuffer_bits_instrs_0_s_T_51}; // @[RVC.scala 21:19 22:14]
  wire [31:0] _io_toIbuffer_bits_instrs_0_T_8_bits = _io_toIbuffer_bits_instrs_0_T_2 == 5'h3 ?
    io_toIbuffer_bits_instrs_0_s_3_bits : _io_toIbuffer_bits_instrs_0_T_6_bits; // @[package.scala 32:76]
  wire [31:0] io_toIbuffer_bits_instrs_0_s_4_bits = {{5'd0}, _io_toIbuffer_bits_instrs_0_s_T_73}; // @[RVC.scala 21:19 22:14]
  wire [31:0] _io_toIbuffer_bits_instrs_0_T_10_bits = _io_toIbuffer_bits_instrs_0_T_2 == 5'h4 ?
    io_toIbuffer_bits_instrs_0_s_4_bits : _io_toIbuffer_bits_instrs_0_T_8_bits; // @[package.scala 32:76]
  wire [31:0] io_toIbuffer_bits_instrs_0_s_5_bits = {{4'd0}, _io_toIbuffer_bits_instrs_0_s_T_93}; // @[RVC.scala 21:19 22:14]
  wire [31:0] _io_toIbuffer_bits_instrs_0_T_12_bits = _io_toIbuffer_bits_instrs_0_T_2 == 5'h5 ?
    io_toIbuffer_bits_instrs_0_s_5_bits : _io_toIbuffer_bits_instrs_0_T_10_bits; // @[package.scala 32:76]
  wire [31:0] io_toIbuffer_bits_instrs_0_s_6_bits = {{5'd0}, _io_toIbuffer_bits_instrs_0_s_T_115}; // @[RVC.scala 21:19 22:14]
  wire [31:0] _io_toIbuffer_bits_instrs_0_T_14_bits = _io_toIbuffer_bits_instrs_0_T_2 == 5'h6 ?
    io_toIbuffer_bits_instrs_0_s_6_bits : _io_toIbuffer_bits_instrs_0_T_12_bits; // @[package.scala 32:76]
  wire [31:0] io_toIbuffer_bits_instrs_0_s_7_bits = {{4'd0}, _io_toIbuffer_bits_instrs_0_s_T_135}; // @[RVC.scala 21:19 22:14]
  wire [31:0] _io_toIbuffer_bits_instrs_0_T_16_bits = _io_toIbuffer_bits_instrs_0_T_2 == 5'h7 ?
    io_toIbuffer_bits_instrs_0_s_7_bits : _io_toIbuffer_bits_instrs_0_T_14_bits; // @[package.scala 32:76]
  wire [31:0] _io_toIbuffer_bits_instrs_0_T_18_bits = _io_toIbuffer_bits_instrs_0_T_2 == 5'h8 ?
    io_toIbuffer_bits_instrs_0_s_8_bits : _io_toIbuffer_bits_instrs_0_T_16_bits; // @[package.scala 32:76]
  wire [31:0] _io_toIbuffer_bits_instrs_0_T_20_bits = _io_toIbuffer_bits_instrs_0_T_2 == 5'h9 ?
    io_toIbuffer_bits_instrs_0_s_9_bits : _io_toIbuffer_bits_instrs_0_T_18_bits; // @[package.scala 32:76]
  wire [31:0] _io_toIbuffer_bits_instrs_0_T_22_bits = _io_toIbuffer_bits_instrs_0_T_2 == 5'ha ?
    io_toIbuffer_bits_instrs_0_s_10_bits : _io_toIbuffer_bits_instrs_0_T_20_bits; // @[package.scala 32:76]
  wire [31:0] _io_toIbuffer_bits_instrs_0_T_24_bits = _io_toIbuffer_bits_instrs_0_T_2 == 5'hb ?
    io_toIbuffer_bits_instrs_0_s_11_bits : _io_toIbuffer_bits_instrs_0_T_22_bits; // @[package.scala 32:76]
  wire [31:0] _io_toIbuffer_bits_instrs_0_T_26_bits = _io_toIbuffer_bits_instrs_0_T_2 == 5'hc ?
    io_toIbuffer_bits_instrs_0_s_12_bits : _io_toIbuffer_bits_instrs_0_T_24_bits; // @[package.scala 32:76]
  wire [31:0] _io_toIbuffer_bits_instrs_0_T_28_bits = _io_toIbuffer_bits_instrs_0_T_2 == 5'hd ?
    io_toIbuffer_bits_instrs_0_s_13_bits : _io_toIbuffer_bits_instrs_0_T_26_bits; // @[package.scala 32:76]
  wire [31:0] _io_toIbuffer_bits_instrs_0_T_30_bits = _io_toIbuffer_bits_instrs_0_T_2 == 5'he ?
    io_toIbuffer_bits_instrs_0_s_14_bits : _io_toIbuffer_bits_instrs_0_T_28_bits; // @[package.scala 32:76]
  wire [31:0] _io_toIbuffer_bits_instrs_0_T_32_bits = _io_toIbuffer_bits_instrs_0_T_2 == 5'hf ?
    io_toIbuffer_bits_instrs_0_s_15_bits : _io_toIbuffer_bits_instrs_0_T_30_bits; // @[package.scala 32:76]
  wire [31:0] io_toIbuffer_bits_instrs_0_s_16_bits = {{6'd0}, _io_toIbuffer_bits_instrs_0_s_T_395}; // @[RVC.scala 21:19 22:14]
  wire [31:0] _io_toIbuffer_bits_instrs_0_T_34_bits = _io_toIbuffer_bits_instrs_0_T_2 == 5'h10 ?
    io_toIbuffer_bits_instrs_0_s_16_bits : _io_toIbuffer_bits_instrs_0_T_32_bits; // @[package.scala 32:76]
  wire [31:0] io_toIbuffer_bits_instrs_0_s_17_bits = {{3'd0}, _io_toIbuffer_bits_instrs_0_s_T_405}; // @[RVC.scala 21:19 22:14]
  wire [31:0] _io_toIbuffer_bits_instrs_0_T_36_bits = _io_toIbuffer_bits_instrs_0_T_2 == 5'h11 ?
    io_toIbuffer_bits_instrs_0_s_17_bits : _io_toIbuffer_bits_instrs_0_T_34_bits; // @[package.scala 32:76]
  wire [31:0] io_toIbuffer_bits_instrs_0_s_18_bits = {{4'd0}, _io_toIbuffer_bits_instrs_0_s_T_414}; // @[RVC.scala 21:19 22:14]
  wire [31:0] _io_toIbuffer_bits_instrs_0_T_38_bits = _io_toIbuffer_bits_instrs_0_T_2 == 5'h12 ?
    io_toIbuffer_bits_instrs_0_s_18_bits : _io_toIbuffer_bits_instrs_0_T_36_bits; // @[package.scala 32:76]
  wire [31:0] io_toIbuffer_bits_instrs_0_s_19_bits = {{3'd0}, _io_toIbuffer_bits_instrs_0_s_T_423}; // @[RVC.scala 21:19 22:14]
  wire [31:0] _io_toIbuffer_bits_instrs_0_T_40_bits = _io_toIbuffer_bits_instrs_0_T_2 == 5'h13 ?
    io_toIbuffer_bits_instrs_0_s_19_bits : _io_toIbuffer_bits_instrs_0_T_38_bits; // @[package.scala 32:76]
  wire [31:0] _io_toIbuffer_bits_instrs_0_T_42_bits = _io_toIbuffer_bits_instrs_0_T_2 == 5'h14 ?
    io_toIbuffer_bits_instrs_0_s_20_bits : _io_toIbuffer_bits_instrs_0_T_40_bits; // @[package.scala 32:76]
  wire [31:0] io_toIbuffer_bits_instrs_0_s_21_bits = {{3'd0}, _io_toIbuffer_bits_instrs_0_s_T_437}; // @[RVC.scala 21:19 22:14]
  wire [31:0] _io_toIbuffer_bits_instrs_0_T_44_bits = _io_toIbuffer_bits_instrs_0_T_2 == 5'h15 ?
    io_toIbuffer_bits_instrs_0_s_21_bits : _io_toIbuffer_bits_instrs_0_T_42_bits; // @[package.scala 32:76]
  wire [31:0] io_toIbuffer_bits_instrs_0_s_22_bits = {{4'd0}, _io_toIbuffer_bits_instrs_0_s_T_450}; // @[RVC.scala 21:19 22:14]
  wire [31:0] _io_toIbuffer_bits_instrs_0_T_46_bits = _io_toIbuffer_bits_instrs_0_T_2 == 5'h16 ?
    io_toIbuffer_bits_instrs_0_s_22_bits : _io_toIbuffer_bits_instrs_0_T_44_bits; // @[package.scala 32:76]
  wire [31:0] io_toIbuffer_bits_instrs_0_s_23_bits = {{3'd0}, _io_toIbuffer_bits_instrs_0_s_T_463}; // @[RVC.scala 21:19 22:14]
  wire [31:0] _io_toIbuffer_bits_instrs_0_T_48_bits = _io_toIbuffer_bits_instrs_0_T_2 == 5'h17 ?
    io_toIbuffer_bits_instrs_0_s_23_bits : _io_toIbuffer_bits_instrs_0_T_46_bits; // @[package.scala 32:76]
  wire [31:0] _io_toIbuffer_bits_instrs_0_T_50_bits = _io_toIbuffer_bits_instrs_0_T_2 == 5'h18 ? inst :
    _io_toIbuffer_bits_instrs_0_T_48_bits; // @[package.scala 32:76]
  wire [31:0] _io_toIbuffer_bits_instrs_0_T_52_bits = _io_toIbuffer_bits_instrs_0_T_2 == 5'h19 ? inst :
    _io_toIbuffer_bits_instrs_0_T_50_bits; // @[package.scala 32:76]
  wire [31:0] _io_toIbuffer_bits_instrs_0_T_54_bits = _io_toIbuffer_bits_instrs_0_T_2 == 5'h1a ? inst :
    _io_toIbuffer_bits_instrs_0_T_52_bits; // @[package.scala 32:76]
  wire [31:0] _io_toIbuffer_bits_instrs_0_T_56_bits = _io_toIbuffer_bits_instrs_0_T_2 == 5'h1b ? inst :
    _io_toIbuffer_bits_instrs_0_T_54_bits; // @[package.scala 32:76]
  wire [31:0] _io_toIbuffer_bits_instrs_0_T_58_bits = _io_toIbuffer_bits_instrs_0_T_2 == 5'h1c ? inst :
    _io_toIbuffer_bits_instrs_0_T_56_bits; // @[package.scala 32:76]
  wire [31:0] _io_toIbuffer_bits_instrs_0_T_60_bits = _io_toIbuffer_bits_instrs_0_T_2 == 5'h1d ? inst :
    _io_toIbuffer_bits_instrs_0_T_58_bits; // @[package.scala 32:76]
  wire [31:0] _io_toIbuffer_bits_instrs_0_T_62_bits = _io_toIbuffer_bits_instrs_0_T_2 == 5'h1e ? inst :
    _io_toIbuffer_bits_instrs_0_T_60_bits; // @[package.scala 32:76]
  wire [31:0] _io_toIbuffer_bits_instrs_0_T_64_bits = _io_toIbuffer_bits_instrs_0_T_2 == 5'h1f ? inst :
    _io_toIbuffer_bits_instrs_0_T_62_bits; // @[package.scala 32:76]
  wire [31:0] f3_expd_instr_0 = f3_expd_instr_expander_io_out_bits; // @[IFU.scala 381:{34,34}]
  wire  mmioFlushWb_bits_pd_0_isRVC = f3_req_is_mmio ? currentIsRVC : f3_pd_0_isRVC; // @[IFU.scala 662:23 623:33 674:37]
  wire [1:0] mmioFlushWb_bits_pd_0_brType = f3_req_is_mmio ? brType : f3_pd_0_brType; // @[IFU.scala 662:23 623:33 675:37]
  wire  mmioFlushWb_bits_pd_0_isCall = f3_req_is_mmio ? isCall : f3_pd_0_isCall; // @[IFU.scala 662:23 623:33 676:37]
  wire  mmioFlushWb_bits_pd_0_isRet = f3_req_is_mmio ? isRet : f3_pd_0_isRet; // @[IFU.scala 662:23 623:33 677:37]
  reg  wb_valid_REG; // @[IFU.scala 706:42]
  reg [38:0] wb_ftq_req_startAddr; // @[IFU.scala 707:34]
  reg  wb_check_result_stage1_fixedTaken_0; // @[IFU.scala 709:41]
  reg  wb_check_result_stage1_fixedTaken_1; // @[IFU.scala 709:41]
  reg  wb_check_result_stage1_fixedTaken_2; // @[IFU.scala 709:41]
  reg  wb_check_result_stage1_fixedTaken_3; // @[IFU.scala 709:41]
  reg  wb_check_result_stage1_fixedTaken_4; // @[IFU.scala 709:41]
  reg  wb_check_result_stage1_fixedTaken_5; // @[IFU.scala 709:41]
  reg  wb_check_result_stage1_fixedTaken_6; // @[IFU.scala 709:41]
  reg  wb_check_result_stage1_fixedTaken_7; // @[IFU.scala 709:41]
  reg [7:0] wb_instr_range; // @[IFU.scala 711:34]
  reg [38:0] wb_pc_0; // @[IFU.scala 712:34]
  reg [38:0] wb_pc_1; // @[IFU.scala 712:34]
  reg [38:0] wb_pc_2; // @[IFU.scala 712:34]
  reg [38:0] wb_pc_3; // @[IFU.scala 712:34]
  reg [38:0] wb_pc_4; // @[IFU.scala 712:34]
  reg [38:0] wb_pc_5; // @[IFU.scala 712:34]
  reg [38:0] wb_pc_6; // @[IFU.scala 712:34]
  reg [38:0] wb_pc_7; // @[IFU.scala 712:34]
  reg  wb_pd_0_isRVC; // @[IFU.scala 713:34]
  reg [1:0] wb_pd_0_brType; // @[IFU.scala 713:34]
  reg  wb_pd_0_isCall; // @[IFU.scala 713:34]
  reg  wb_pd_0_isRet; // @[IFU.scala 713:34]
  reg  wb_pd_1_isRVC; // @[IFU.scala 713:34]
  reg [1:0] wb_pd_1_brType; // @[IFU.scala 713:34]
  reg  wb_pd_1_isCall; // @[IFU.scala 713:34]
  reg  wb_pd_1_isRet; // @[IFU.scala 713:34]
  reg  wb_pd_2_isRVC; // @[IFU.scala 713:34]
  reg [1:0] wb_pd_2_brType; // @[IFU.scala 713:34]
  reg  wb_pd_2_isCall; // @[IFU.scala 713:34]
  reg  wb_pd_2_isRet; // @[IFU.scala 713:34]
  reg  wb_pd_3_isRVC; // @[IFU.scala 713:34]
  reg [1:0] wb_pd_3_brType; // @[IFU.scala 713:34]
  reg  wb_pd_3_isCall; // @[IFU.scala 713:34]
  reg  wb_pd_3_isRet; // @[IFU.scala 713:34]
  reg  wb_pd_4_isRVC; // @[IFU.scala 713:34]
  reg [1:0] wb_pd_4_brType; // @[IFU.scala 713:34]
  reg  wb_pd_4_isCall; // @[IFU.scala 713:34]
  reg  wb_pd_4_isRet; // @[IFU.scala 713:34]
  reg  wb_pd_5_isRVC; // @[IFU.scala 713:34]
  reg [1:0] wb_pd_5_brType; // @[IFU.scala 713:34]
  reg  wb_pd_5_isCall; // @[IFU.scala 713:34]
  reg  wb_pd_5_isRet; // @[IFU.scala 713:34]
  reg  wb_pd_6_isRVC; // @[IFU.scala 713:34]
  reg [1:0] wb_pd_6_brType; // @[IFU.scala 713:34]
  reg  wb_pd_6_isCall; // @[IFU.scala 713:34]
  reg  wb_pd_6_isRet; // @[IFU.scala 713:34]
  reg  wb_pd_7_isRVC; // @[IFU.scala 713:34]
  reg [1:0] wb_pd_7_brType; // @[IFU.scala 713:34]
  reg  wb_pd_7_isCall; // @[IFU.scala 713:34]
  reg  wb_pd_7_isRet; // @[IFU.scala 713:34]
  reg  wb_instr_valid_0; // @[IFU.scala 714:34]
  reg  wb_instr_valid_1; // @[IFU.scala 714:34]
  reg  wb_instr_valid_2; // @[IFU.scala 714:34]
  reg  wb_instr_valid_3; // @[IFU.scala 714:34]
  reg  wb_instr_valid_4; // @[IFU.scala 714:34]
  reg  wb_instr_valid_5; // @[IFU.scala 714:34]
  reg  wb_instr_valid_6; // @[IFU.scala 714:34]
  reg  wb_instr_valid_7; // @[IFU.scala 714:34]
  reg [38:0] wb_false_target; // @[IFU.scala 719:34]
  wire [38:0] _GEN_2091 = 3'h1 == f3_last_validIdx ? f3_half_snpc_1 : f3_half_snpc_0; // @[IFU.scala 719:{34,34}]
  wire [38:0] _GEN_2092 = 3'h2 == f3_last_validIdx ? f3_half_snpc_2 : _GEN_2091; // @[IFU.scala 719:{34,34}]
  wire [38:0] _GEN_2093 = 3'h3 == f3_last_validIdx ? f3_half_snpc_3 : _GEN_2092; // @[IFU.scala 719:{34,34}]
  reg  REG_1; // @[IFU.scala 735:27]
  wire  _T_81 = wb_valid & REG_1; // @[IFU.scala 735:17]
  reg  REG_2; // @[IFU.scala 736:91]
  wire  _T_88 = _T_81 & predChecker_io_out_stage2Out_fixedMissPred_7 & ~f3_fire & ~REG_2 & _io_toIbuffer_valid_T_3; // @[IFU.scala 736:116]
  reg  REG_3; // @[IFU.scala 742:27]
  wire  _T_89 = wb_valid & REG_3; // @[IFU.scala 742:17]
  wire  _T_91 = _T_89 & predChecker_io_out_stage2Out_fixedMissPred_7 & f3_fire; // @[IFU.scala 743:67]
  wire  _checkFlushWb_bits_misOffset_bits_T_1 = predChecker_io_out_stage2Out_fixedMissPred_0 ? 1'h0 : 1'h1; // @[ParallelMux.scala 90:77]
  wire [1:0] _checkFlushWb_bits_misOffset_bits_T_3 = predChecker_io_out_stage2Out_fixedMissPred_2 ? 2'h2 : 2'h3; // @[ParallelMux.scala 90:77]
  wire [1:0] _checkFlushWb_bits_misOffset_bits_T_5 = _checkFlushWb_bits_misOffset_valid_T ? {{1'd0},
    _checkFlushWb_bits_misOffset_bits_T_1} : _checkFlushWb_bits_misOffset_bits_T_3; // @[ParallelMux.scala 90:77]
  wire [2:0] _checkFlushWb_bits_misOffset_bits_T_7 = predChecker_io_out_stage2Out_fixedMissPred_4 ? 3'h4 : 3'h5; // @[ParallelMux.scala 90:77]
  wire [2:0] _checkFlushWb_bits_misOffset_bits_T_9 = predChecker_io_out_stage2Out_fixedMissPred_6 ? 3'h6 : 3'h7; // @[ParallelMux.scala 90:77]
  wire [2:0] _checkFlushWb_bits_misOffset_bits_T_11 = _checkFlushWb_bits_misOffset_valid_T_3 ?
    _checkFlushWb_bits_misOffset_bits_T_7 : _checkFlushWb_bits_misOffset_bits_T_9; // @[ParallelMux.scala 90:77]
  wire [2:0] _checkFlushWb_bits_misOffset_bits_T_13 = _checkFlushWb_bits_misOffset_valid_T_2 ? {{1'd0},
    _checkFlushWb_bits_misOffset_bits_T_5} : _checkFlushWb_bits_misOffset_bits_T_11; // @[ParallelMux.scala 90:77]
  wire [2:0] checkFlushWb_bits_misOffset_bits = wb_false_lastHalf ? wb_lastIdx : _checkFlushWb_bits_misOffset_bits_T_13; // @[IFU.scala 756:45]
  wire  checkFlushWb_bits_cfiOffset_valid = wb_check_result_stage1_fixedTaken_0 | wb_check_result_stage1_fixedTaken_1 |
    (wb_check_result_stage1_fixedTaken_2 | wb_check_result_stage1_fixedTaken_3) | (wb_check_result_stage1_fixedTaken_4
     | wb_check_result_stage1_fixedTaken_5 | (wb_check_result_stage1_fixedTaken_6 | wb_check_result_stage1_fixedTaken_7)
    ); // @[ParallelMux.scala 36:53]
  wire [38:0] _GEN_2100 = predChecker_io_out_stage2Out_fixedTarget_0; // @[IFU.scala 759:{45,45}]
  wire [38:0] _GEN_2101 = 3'h1 == _checkFlushWb_bits_misOffset_bits_T_13 ? predChecker_io_out_stage2Out_fixedTarget_1 :
    _GEN_2100; // @[IFU.scala 759:{45,45}]
  wire [38:0] _GEN_2102 = 3'h2 == _checkFlushWb_bits_misOffset_bits_T_13 ? predChecker_io_out_stage2Out_fixedTarget_2 :
    _GEN_2101; // @[IFU.scala 759:{45,45}]
  wire [38:0] _GEN_2103 = 3'h3 == _checkFlushWb_bits_misOffset_bits_T_13 ? predChecker_io_out_stage2Out_fixedTarget_3 :
    _GEN_2102; // @[IFU.scala 759:{45,45}]
  wire [38:0] _GEN_2104 = 3'h4 == _checkFlushWb_bits_misOffset_bits_T_13 ? predChecker_io_out_stage2Out_fixedTarget_4 :
    _GEN_2103; // @[IFU.scala 759:{45,45}]
  wire [38:0] _GEN_2105 = 3'h5 == _checkFlushWb_bits_misOffset_bits_T_13 ? predChecker_io_out_stage2Out_fixedTarget_5 :
    _GEN_2104; // @[IFU.scala 759:{45,45}]
  wire [38:0] _GEN_2106 = 3'h6 == _checkFlushWb_bits_misOffset_bits_T_13 ? predChecker_io_out_stage2Out_fixedTarget_6 :
    _GEN_2105; // @[IFU.scala 759:{45,45}]
  wire [38:0] _GEN_2107 = 3'h7 == _checkFlushWb_bits_misOffset_bits_T_13 ? predChecker_io_out_stage2Out_fixedTarget_7 :
    _GEN_2106; // @[IFU.scala 759:{45,45}]
  wire [38:0] checkFlushWb_bits_target = wb_false_lastHalf ? wb_false_target : _GEN_2107; // @[IFU.scala 759:45]
  wire  _checkFlushWb_bits_jalTarget_T = wb_pd_0_brType == 2'h2; // @[PreDecode.scala 77:24]
  wire  _checkFlushWb_bits_jalTarget_T_1 = wb_instr_valid_0 & _checkFlushWb_bits_jalTarget_T; // @[IFU.scala 760:157]
  wire  _checkFlushWb_bits_jalTarget_T_2 = wb_pd_1_brType == 2'h2; // @[PreDecode.scala 77:24]
  wire  _checkFlushWb_bits_jalTarget_T_3 = wb_instr_valid_1 & _checkFlushWb_bits_jalTarget_T_2; // @[IFU.scala 760:157]
  wire  _checkFlushWb_bits_jalTarget_T_4 = wb_pd_2_brType == 2'h2; // @[PreDecode.scala 77:24]
  wire  _checkFlushWb_bits_jalTarget_T_5 = wb_instr_valid_2 & _checkFlushWb_bits_jalTarget_T_4; // @[IFU.scala 760:157]
  wire  _checkFlushWb_bits_jalTarget_T_6 = wb_pd_3_brType == 2'h2; // @[PreDecode.scala 77:24]
  wire  _checkFlushWb_bits_jalTarget_T_7 = wb_instr_valid_3 & _checkFlushWb_bits_jalTarget_T_6; // @[IFU.scala 760:157]
  wire  _checkFlushWb_bits_jalTarget_T_8 = wb_pd_4_brType == 2'h2; // @[PreDecode.scala 77:24]
  wire  _checkFlushWb_bits_jalTarget_T_9 = wb_instr_valid_4 & _checkFlushWb_bits_jalTarget_T_8; // @[IFU.scala 760:157]
  wire  _checkFlushWb_bits_jalTarget_T_10 = wb_pd_5_brType == 2'h2; // @[PreDecode.scala 77:24]
  wire  _checkFlushWb_bits_jalTarget_T_11 = wb_instr_valid_5 & _checkFlushWb_bits_jalTarget_T_10; // @[IFU.scala 760:157]
  wire  _checkFlushWb_bits_jalTarget_T_12 = wb_pd_6_brType == 2'h2; // @[PreDecode.scala 77:24]
  wire  _checkFlushWb_bits_jalTarget_T_13 = wb_instr_valid_6 & _checkFlushWb_bits_jalTarget_T_12; // @[IFU.scala 760:157]
  wire  _checkFlushWb_bits_jalTarget_T_17 = _checkFlushWb_bits_jalTarget_T_1 ? 1'h0 : 1'h1; // @[ParallelMux.scala 90:77]
  wire [1:0] _checkFlushWb_bits_jalTarget_T_19 = _checkFlushWb_bits_jalTarget_T_5 ? 2'h2 : 2'h3; // @[ParallelMux.scala 90:77]
  wire [1:0] _checkFlushWb_bits_jalTarget_T_21 = _checkFlushWb_bits_jalTarget_T_1 | _checkFlushWb_bits_jalTarget_T_3 ?
    {{1'd0}, _checkFlushWb_bits_jalTarget_T_17} : _checkFlushWb_bits_jalTarget_T_19; // @[ParallelMux.scala 90:77]
  wire [2:0] _checkFlushWb_bits_jalTarget_T_23 = _checkFlushWb_bits_jalTarget_T_9 ? 3'h4 : 3'h5; // @[ParallelMux.scala 90:77]
  wire [2:0] _checkFlushWb_bits_jalTarget_T_25 = _checkFlushWb_bits_jalTarget_T_13 ? 3'h6 : 3'h7; // @[ParallelMux.scala 90:77]
  wire [2:0] _checkFlushWb_bits_jalTarget_T_27 = _checkFlushWb_bits_jalTarget_T_9 | _checkFlushWb_bits_jalTarget_T_11 ?
    _checkFlushWb_bits_jalTarget_T_23 : _checkFlushWb_bits_jalTarget_T_25; // @[ParallelMux.scala 90:77]
  wire [2:0] _checkFlushWb_bits_jalTarget_T_29 = _checkFlushWb_bits_jalTarget_T_1 | _checkFlushWb_bits_jalTarget_T_3 | (
    _checkFlushWb_bits_jalTarget_T_5 | _checkFlushWb_bits_jalTarget_T_7) ? {{1'd0}, _checkFlushWb_bits_jalTarget_T_21}
     : _checkFlushWb_bits_jalTarget_T_27; // @[ParallelMux.scala 90:77]
  wire [38:0] _GEN_2109 = 3'h1 == _checkFlushWb_bits_jalTarget_T_29 ? predChecker_io_out_stage2Out_fixedTarget_1 :
    _GEN_2100; // @[IFU.scala 760:{39,39}]
  wire [38:0] _GEN_2110 = 3'h2 == _checkFlushWb_bits_jalTarget_T_29 ? predChecker_io_out_stage2Out_fixedTarget_2 :
    _GEN_2109; // @[IFU.scala 760:{39,39}]
  wire [38:0] _GEN_2111 = 3'h3 == _checkFlushWb_bits_jalTarget_T_29 ? predChecker_io_out_stage2Out_fixedTarget_3 :
    _GEN_2110; // @[IFU.scala 760:{39,39}]
  wire [38:0] _GEN_2112 = 3'h4 == _checkFlushWb_bits_jalTarget_T_29 ? predChecker_io_out_stage2Out_fixedTarget_4 :
    _GEN_2111; // @[IFU.scala 760:{39,39}]
  wire [38:0] _GEN_2113 = 3'h5 == _checkFlushWb_bits_jalTarget_T_29 ? predChecker_io_out_stage2Out_fixedTarget_5 :
    _GEN_2112; // @[IFU.scala 760:{39,39}]
  wire [38:0] _GEN_2114 = 3'h6 == _checkFlushWb_bits_jalTarget_T_29 ? predChecker_io_out_stage2Out_fixedTarget_6 :
    _GEN_2113; // @[IFU.scala 760:{39,39}]
  wire [38:0] checkFlushWb_bits_jalTarget = 3'h7 == _checkFlushWb_bits_jalTarget_T_29 ?
    predChecker_io_out_stage2Out_fixedTarget_7 : _GEN_2114; // @[IFU.scala 760:{39,39}]
  wire  _checkJalFault_T = predChecker_io_out_stage2Out_faultType_0_value == 3'h1; // @[PreDecode.scala 190:31]
  wire  _checkJalFault_T_1 = predChecker_io_out_stage2Out_faultType_1_value == 3'h1; // @[PreDecode.scala 190:31]
  wire  _checkJalFault_T_2 = predChecker_io_out_stage2Out_faultType_2_value == 3'h1; // @[PreDecode.scala 190:31]
  wire  _checkJalFault_T_3 = predChecker_io_out_stage2Out_faultType_3_value == 3'h1; // @[PreDecode.scala 190:31]
  wire  _checkJalFault_T_4 = predChecker_io_out_stage2Out_faultType_4_value == 3'h1; // @[PreDecode.scala 190:31]
  wire  _checkJalFault_T_5 = predChecker_io_out_stage2Out_faultType_5_value == 3'h1; // @[PreDecode.scala 190:31]
  wire  _checkJalFault_T_6 = predChecker_io_out_stage2Out_faultType_6_value == 3'h1; // @[PreDecode.scala 190:31]
  wire  _checkJalFault_T_7 = predChecker_io_out_stage2Out_faultType_7_value == 3'h1; // @[PreDecode.scala 190:31]
  wire  _checkRetFault_T = predChecker_io_out_stage2Out_faultType_0_value == 3'h2; // @[PreDecode.scala 191:31]
  wire  _checkRetFault_T_1 = predChecker_io_out_stage2Out_faultType_1_value == 3'h2; // @[PreDecode.scala 191:31]
  wire  _checkRetFault_T_2 = predChecker_io_out_stage2Out_faultType_2_value == 3'h2; // @[PreDecode.scala 191:31]
  wire  _checkRetFault_T_3 = predChecker_io_out_stage2Out_faultType_3_value == 3'h2; // @[PreDecode.scala 191:31]
  wire  _checkRetFault_T_4 = predChecker_io_out_stage2Out_faultType_4_value == 3'h2; // @[PreDecode.scala 191:31]
  wire  _checkRetFault_T_5 = predChecker_io_out_stage2Out_faultType_5_value == 3'h2; // @[PreDecode.scala 191:31]
  wire  _checkRetFault_T_6 = predChecker_io_out_stage2Out_faultType_6_value == 3'h2; // @[PreDecode.scala 191:31]
  wire  _checkRetFault_T_7 = predChecker_io_out_stage2Out_faultType_7_value == 3'h2; // @[PreDecode.scala 191:31]
  wire  _checkTargetFault_T = predChecker_io_out_stage2Out_faultType_0_value == 3'h3; // @[PreDecode.scala 192:31]
  wire  _checkTargetFault_T_1 = predChecker_io_out_stage2Out_faultType_1_value == 3'h3; // @[PreDecode.scala 192:31]
  wire  _checkTargetFault_T_2 = predChecker_io_out_stage2Out_faultType_2_value == 3'h3; // @[PreDecode.scala 192:31]
  wire  _checkTargetFault_T_3 = predChecker_io_out_stage2Out_faultType_3_value == 3'h3; // @[PreDecode.scala 192:31]
  wire  _checkTargetFault_T_4 = predChecker_io_out_stage2Out_faultType_4_value == 3'h3; // @[PreDecode.scala 192:31]
  wire  _checkTargetFault_T_5 = predChecker_io_out_stage2Out_faultType_5_value == 3'h3; // @[PreDecode.scala 192:31]
  wire  _checkTargetFault_T_6 = predChecker_io_out_stage2Out_faultType_6_value == 3'h3; // @[PreDecode.scala 192:31]
  wire  _checkTargetFault_T_7 = predChecker_io_out_stage2Out_faultType_7_value == 3'h3; // @[PreDecode.scala 192:31]
  wire  _checkNotCFIFault_T = predChecker_io_out_stage2Out_faultType_0_value == 3'h4; // @[PreDecode.scala 194:36]
  wire  _checkNotCFIFault_T_1 = predChecker_io_out_stage2Out_faultType_1_value == 3'h4; // @[PreDecode.scala 194:36]
  wire  _checkNotCFIFault_T_2 = predChecker_io_out_stage2Out_faultType_2_value == 3'h4; // @[PreDecode.scala 194:36]
  wire  _checkNotCFIFault_T_3 = predChecker_io_out_stage2Out_faultType_3_value == 3'h4; // @[PreDecode.scala 194:36]
  wire  _checkNotCFIFault_T_4 = predChecker_io_out_stage2Out_faultType_4_value == 3'h4; // @[PreDecode.scala 194:36]
  wire  _checkNotCFIFault_T_5 = predChecker_io_out_stage2Out_faultType_5_value == 3'h4; // @[PreDecode.scala 194:36]
  wire  _checkNotCFIFault_T_6 = predChecker_io_out_stage2Out_faultType_6_value == 3'h4; // @[PreDecode.scala 194:36]
  wire  _checkNotCFIFault_T_7 = predChecker_io_out_stage2Out_faultType_7_value == 3'h4; // @[PreDecode.scala 194:36]
  wire  _checkInvalidTaken_T = predChecker_io_out_stage2Out_faultType_0_value == 3'h5; // @[PreDecode.scala 193:36]
  wire  _checkInvalidTaken_T_1 = predChecker_io_out_stage2Out_faultType_1_value == 3'h5; // @[PreDecode.scala 193:36]
  wire  _checkInvalidTaken_T_2 = predChecker_io_out_stage2Out_faultType_2_value == 3'h5; // @[PreDecode.scala 193:36]
  wire  _checkInvalidTaken_T_3 = predChecker_io_out_stage2Out_faultType_3_value == 3'h5; // @[PreDecode.scala 193:36]
  wire  _checkInvalidTaken_T_4 = predChecker_io_out_stage2Out_faultType_4_value == 3'h5; // @[PreDecode.scala 193:36]
  wire  _checkInvalidTaken_T_5 = predChecker_io_out_stage2Out_faultType_5_value == 3'h5; // @[PreDecode.scala 193:36]
  wire  _checkInvalidTaken_T_6 = predChecker_io_out_stage2Out_faultType_6_value == 3'h5; // @[PreDecode.scala 193:36]
  wire  _checkInvalidTaken_T_7 = predChecker_io_out_stage2Out_faultType_7_value == 3'h5; // @[PreDecode.scala 193:36]
  reg  f3_perf_info_only_0_hit; // @[Reg.scala 16:16]
  reg  f3_perf_info_only_0_miss; // @[Reg.scala 16:16]
  reg  f3_perf_info_hit_0_hit_1; // @[Reg.scala 16:16]
  reg  f3_perf_info_hit_0_miss_1; // @[Reg.scala 16:16]
  reg  f3_perf_info_miss_0_hit_1; // @[Reg.scala 16:16]
  reg  f3_perf_info_miss_0_miss_1; // @[Reg.scala 16:16]
  reg  f3_perf_info_hit_0_except_1; // @[Reg.scala 16:16]
  reg  f3_perf_info_miss_0_except_1; // @[Reg.scala 16:16]
  reg  f3_perf_info_except_0; // @[Reg.scala 16:16]
  reg  f3_perf_info_bank_hit_1; // @[Reg.scala 16:16]
  reg  f3_perf_info_hit; // @[Reg.scala 16:16]
  wire  f3_req_1 = f3_fire & f3_doubleLine; // @[IFU.scala 791:41]
  reg  io_perf_0_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg  io_perf_0_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg  io_perf_1_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg  io_perf_1_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg  io_perf_2_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg  io_perf_2_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg  io_perf_3_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg  io_perf_3_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg  io_perf_4_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg  io_perf_4_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg  io_perf_5_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg  io_perf_5_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg  io_perf_6_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg  io_perf_6_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg  io_perf_7_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg  io_perf_7_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg  io_perf_8_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg  io_perf_8_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg  io_perf_9_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg  io_perf_9_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg  io_perf_10_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg  io_perf_10_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg  io_perf_11_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg  io_perf_11_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg  io_perf_12_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg  io_perf_12_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  wire  _T_133 = f3_perf_info_hit_0_except_1 & f3_fire; // @[IFU.scala 825:68]
  wire  _T_135 = f3_perf_info_miss_0_except_1 & f3_fire; // @[IFU.scala 826:70]
  wire  _T_137 = f3_perf_info_except_0 & f3_fire; // @[IFU.scala 827:56]
  wire [1:0] _fetchIBufferDumpData_instr_count_T_8 = io_toIbuffer_bits_enqEnable[0] + io_toIbuffer_bits_enqEnable[1]; // @[Bitwise.scala 48:55]
  wire [1:0] _fetchIBufferDumpData_instr_count_T_10 = io_toIbuffer_bits_enqEnable[2] + io_toIbuffer_bits_enqEnable[3]; // @[Bitwise.scala 48:55]
  wire [2:0] _fetchIBufferDumpData_instr_count_T_12 = _fetchIBufferDumpData_instr_count_T_8 +
    _fetchIBufferDumpData_instr_count_T_10; // @[Bitwise.scala 48:55]
  wire [1:0] _fetchIBufferDumpData_instr_count_T_14 = io_toIbuffer_bits_enqEnable[4] + io_toIbuffer_bits_enqEnable[5]; // @[Bitwise.scala 48:55]
  wire [1:0] _fetchIBufferDumpData_instr_count_T_16 = io_toIbuffer_bits_enqEnable[6] + io_toIbuffer_bits_enqEnable[7]; // @[Bitwise.scala 48:55]
  wire [2:0] _fetchIBufferDumpData_instr_count_T_18 = _fetchIBufferDumpData_instr_count_T_14 +
    _fetchIBufferDumpData_instr_count_T_16; // @[Bitwise.scala 48:55]
  wire [3:0] _fetchIBufferDumpData_instr_count_T_20 = _fetchIBufferDumpData_instr_count_T_12 +
    _fetchIBufferDumpData_instr_count_T_18; // @[Bitwise.scala 48:55]
  reg [63:0] cnt; // @[ChiselDB.scala 133:22]
  reg [63:0] cnt_1; // @[ChiselDB.scala 133:22]
  PreDecode preDecoders_0 ( // @[IFU.scala 142:46]
    .io_in_data_0(preDecoders_0_io_in_data_0),
    .io_in_data_1(preDecoders_0_io_in_data_1),
    .io_in_data_2(preDecoders_0_io_in_data_2),
    .io_in_data_3(preDecoders_0_io_in_data_3),
    .io_in_data_4(preDecoders_0_io_in_data_4),
    .io_in_data_5(preDecoders_0_io_in_data_5),
    .io_in_data_6(preDecoders_0_io_in_data_6),
    .io_in_data_7(preDecoders_0_io_in_data_7),
    .io_in_data_8(preDecoders_0_io_in_data_8),
    .io_out_pd_0_isRVC(preDecoders_0_io_out_pd_0_isRVC),
    .io_out_pd_0_brType(preDecoders_0_io_out_pd_0_brType),
    .io_out_pd_0_isCall(preDecoders_0_io_out_pd_0_isCall),
    .io_out_pd_0_isRet(preDecoders_0_io_out_pd_0_isRet),
    .io_out_pd_1_valid(preDecoders_0_io_out_pd_1_valid),
    .io_out_pd_1_isRVC(preDecoders_0_io_out_pd_1_isRVC),
    .io_out_pd_1_brType(preDecoders_0_io_out_pd_1_brType),
    .io_out_pd_1_isCall(preDecoders_0_io_out_pd_1_isCall),
    .io_out_pd_1_isRet(preDecoders_0_io_out_pd_1_isRet),
    .io_out_pd_2_valid(preDecoders_0_io_out_pd_2_valid),
    .io_out_pd_2_isRVC(preDecoders_0_io_out_pd_2_isRVC),
    .io_out_pd_2_brType(preDecoders_0_io_out_pd_2_brType),
    .io_out_pd_2_isCall(preDecoders_0_io_out_pd_2_isCall),
    .io_out_pd_2_isRet(preDecoders_0_io_out_pd_2_isRet),
    .io_out_pd_3_valid(preDecoders_0_io_out_pd_3_valid),
    .io_out_pd_3_isRVC(preDecoders_0_io_out_pd_3_isRVC),
    .io_out_pd_3_brType(preDecoders_0_io_out_pd_3_brType),
    .io_out_pd_3_isCall(preDecoders_0_io_out_pd_3_isCall),
    .io_out_pd_3_isRet(preDecoders_0_io_out_pd_3_isRet),
    .io_out_pd_4_valid(preDecoders_0_io_out_pd_4_valid),
    .io_out_pd_4_isRVC(preDecoders_0_io_out_pd_4_isRVC),
    .io_out_pd_4_brType(preDecoders_0_io_out_pd_4_brType),
    .io_out_pd_4_isCall(preDecoders_0_io_out_pd_4_isCall),
    .io_out_pd_4_isRet(preDecoders_0_io_out_pd_4_isRet),
    .io_out_pd_5_valid(preDecoders_0_io_out_pd_5_valid),
    .io_out_pd_5_isRVC(preDecoders_0_io_out_pd_5_isRVC),
    .io_out_pd_5_brType(preDecoders_0_io_out_pd_5_brType),
    .io_out_pd_5_isCall(preDecoders_0_io_out_pd_5_isCall),
    .io_out_pd_5_isRet(preDecoders_0_io_out_pd_5_isRet),
    .io_out_pd_6_valid(preDecoders_0_io_out_pd_6_valid),
    .io_out_pd_6_isRVC(preDecoders_0_io_out_pd_6_isRVC),
    .io_out_pd_6_brType(preDecoders_0_io_out_pd_6_brType),
    .io_out_pd_6_isCall(preDecoders_0_io_out_pd_6_isCall),
    .io_out_pd_6_isRet(preDecoders_0_io_out_pd_6_isRet),
    .io_out_pd_7_valid(preDecoders_0_io_out_pd_7_valid),
    .io_out_pd_7_isRVC(preDecoders_0_io_out_pd_7_isRVC),
    .io_out_pd_7_brType(preDecoders_0_io_out_pd_7_brType),
    .io_out_pd_7_isCall(preDecoders_0_io_out_pd_7_isCall),
    .io_out_pd_7_isRet(preDecoders_0_io_out_pd_7_isRet),
    .io_out_hasHalfValid_2(preDecoders_0_io_out_hasHalfValid_2),
    .io_out_hasHalfValid_3(preDecoders_0_io_out_hasHalfValid_3),
    .io_out_hasHalfValid_4(preDecoders_0_io_out_hasHalfValid_4),
    .io_out_hasHalfValid_5(preDecoders_0_io_out_hasHalfValid_5),
    .io_out_hasHalfValid_6(preDecoders_0_io_out_hasHalfValid_6),
    .io_out_hasHalfValid_7(preDecoders_0_io_out_hasHalfValid_7),
    .io_out_instr_0(preDecoders_0_io_out_instr_0),
    .io_out_instr_1(preDecoders_0_io_out_instr_1),
    .io_out_instr_2(preDecoders_0_io_out_instr_2),
    .io_out_instr_3(preDecoders_0_io_out_instr_3),
    .io_out_instr_4(preDecoders_0_io_out_instr_4),
    .io_out_instr_5(preDecoders_0_io_out_instr_5),
    .io_out_instr_6(preDecoders_0_io_out_instr_6),
    .io_out_instr_7(preDecoders_0_io_out_instr_7),
    .io_out_jumpOffset_0(preDecoders_0_io_out_jumpOffset_0),
    .io_out_jumpOffset_1(preDecoders_0_io_out_jumpOffset_1),
    .io_out_jumpOffset_2(preDecoders_0_io_out_jumpOffset_2),
    .io_out_jumpOffset_3(preDecoders_0_io_out_jumpOffset_3),
    .io_out_jumpOffset_4(preDecoders_0_io_out_jumpOffset_4),
    .io_out_jumpOffset_5(preDecoders_0_io_out_jumpOffset_5),
    .io_out_jumpOffset_6(preDecoders_0_io_out_jumpOffset_6),
    .io_out_jumpOffset_7(preDecoders_0_io_out_jumpOffset_7)
  );
  PreDecode preDecoders_1 ( // @[IFU.scala 142:46]
    .io_in_data_0(preDecoders_1_io_in_data_0),
    .io_in_data_1(preDecoders_1_io_in_data_1),
    .io_in_data_2(preDecoders_1_io_in_data_2),
    .io_in_data_3(preDecoders_1_io_in_data_3),
    .io_in_data_4(preDecoders_1_io_in_data_4),
    .io_in_data_5(preDecoders_1_io_in_data_5),
    .io_in_data_6(preDecoders_1_io_in_data_6),
    .io_in_data_7(preDecoders_1_io_in_data_7),
    .io_in_data_8(preDecoders_1_io_in_data_8),
    .io_out_pd_0_isRVC(preDecoders_1_io_out_pd_0_isRVC),
    .io_out_pd_0_brType(preDecoders_1_io_out_pd_0_brType),
    .io_out_pd_0_isCall(preDecoders_1_io_out_pd_0_isCall),
    .io_out_pd_0_isRet(preDecoders_1_io_out_pd_0_isRet),
    .io_out_pd_1_valid(preDecoders_1_io_out_pd_1_valid),
    .io_out_pd_1_isRVC(preDecoders_1_io_out_pd_1_isRVC),
    .io_out_pd_1_brType(preDecoders_1_io_out_pd_1_brType),
    .io_out_pd_1_isCall(preDecoders_1_io_out_pd_1_isCall),
    .io_out_pd_1_isRet(preDecoders_1_io_out_pd_1_isRet),
    .io_out_pd_2_valid(preDecoders_1_io_out_pd_2_valid),
    .io_out_pd_2_isRVC(preDecoders_1_io_out_pd_2_isRVC),
    .io_out_pd_2_brType(preDecoders_1_io_out_pd_2_brType),
    .io_out_pd_2_isCall(preDecoders_1_io_out_pd_2_isCall),
    .io_out_pd_2_isRet(preDecoders_1_io_out_pd_2_isRet),
    .io_out_pd_3_valid(preDecoders_1_io_out_pd_3_valid),
    .io_out_pd_3_isRVC(preDecoders_1_io_out_pd_3_isRVC),
    .io_out_pd_3_brType(preDecoders_1_io_out_pd_3_brType),
    .io_out_pd_3_isCall(preDecoders_1_io_out_pd_3_isCall),
    .io_out_pd_3_isRet(preDecoders_1_io_out_pd_3_isRet),
    .io_out_pd_4_valid(preDecoders_1_io_out_pd_4_valid),
    .io_out_pd_4_isRVC(preDecoders_1_io_out_pd_4_isRVC),
    .io_out_pd_4_brType(preDecoders_1_io_out_pd_4_brType),
    .io_out_pd_4_isCall(preDecoders_1_io_out_pd_4_isCall),
    .io_out_pd_4_isRet(preDecoders_1_io_out_pd_4_isRet),
    .io_out_pd_5_valid(preDecoders_1_io_out_pd_5_valid),
    .io_out_pd_5_isRVC(preDecoders_1_io_out_pd_5_isRVC),
    .io_out_pd_5_brType(preDecoders_1_io_out_pd_5_brType),
    .io_out_pd_5_isCall(preDecoders_1_io_out_pd_5_isCall),
    .io_out_pd_5_isRet(preDecoders_1_io_out_pd_5_isRet),
    .io_out_pd_6_valid(preDecoders_1_io_out_pd_6_valid),
    .io_out_pd_6_isRVC(preDecoders_1_io_out_pd_6_isRVC),
    .io_out_pd_6_brType(preDecoders_1_io_out_pd_6_brType),
    .io_out_pd_6_isCall(preDecoders_1_io_out_pd_6_isCall),
    .io_out_pd_6_isRet(preDecoders_1_io_out_pd_6_isRet),
    .io_out_pd_7_valid(preDecoders_1_io_out_pd_7_valid),
    .io_out_pd_7_isRVC(preDecoders_1_io_out_pd_7_isRVC),
    .io_out_pd_7_brType(preDecoders_1_io_out_pd_7_brType),
    .io_out_pd_7_isCall(preDecoders_1_io_out_pd_7_isCall),
    .io_out_pd_7_isRet(preDecoders_1_io_out_pd_7_isRet),
    .io_out_hasHalfValid_2(preDecoders_1_io_out_hasHalfValid_2),
    .io_out_hasHalfValid_3(preDecoders_1_io_out_hasHalfValid_3),
    .io_out_hasHalfValid_4(preDecoders_1_io_out_hasHalfValid_4),
    .io_out_hasHalfValid_5(preDecoders_1_io_out_hasHalfValid_5),
    .io_out_hasHalfValid_6(preDecoders_1_io_out_hasHalfValid_6),
    .io_out_hasHalfValid_7(preDecoders_1_io_out_hasHalfValid_7),
    .io_out_instr_0(preDecoders_1_io_out_instr_0),
    .io_out_instr_1(preDecoders_1_io_out_instr_1),
    .io_out_instr_2(preDecoders_1_io_out_instr_2),
    .io_out_instr_3(preDecoders_1_io_out_instr_3),
    .io_out_instr_4(preDecoders_1_io_out_instr_4),
    .io_out_instr_5(preDecoders_1_io_out_instr_5),
    .io_out_instr_6(preDecoders_1_io_out_instr_6),
    .io_out_instr_7(preDecoders_1_io_out_instr_7),
    .io_out_jumpOffset_0(preDecoders_1_io_out_jumpOffset_0),
    .io_out_jumpOffset_1(preDecoders_1_io_out_jumpOffset_1),
    .io_out_jumpOffset_2(preDecoders_1_io_out_jumpOffset_2),
    .io_out_jumpOffset_3(preDecoders_1_io_out_jumpOffset_3),
    .io_out_jumpOffset_4(preDecoders_1_io_out_jumpOffset_4),
    .io_out_jumpOffset_5(preDecoders_1_io_out_jumpOffset_5),
    .io_out_jumpOffset_6(preDecoders_1_io_out_jumpOffset_6),
    .io_out_jumpOffset_7(preDecoders_1_io_out_jumpOffset_7)
  );
  PreDecode preDecoders_2 ( // @[IFU.scala 142:46]
    .io_in_data_0(preDecoders_2_io_in_data_0),
    .io_in_data_1(preDecoders_2_io_in_data_1),
    .io_in_data_2(preDecoders_2_io_in_data_2),
    .io_in_data_3(preDecoders_2_io_in_data_3),
    .io_in_data_4(preDecoders_2_io_in_data_4),
    .io_in_data_5(preDecoders_2_io_in_data_5),
    .io_in_data_6(preDecoders_2_io_in_data_6),
    .io_in_data_7(preDecoders_2_io_in_data_7),
    .io_in_data_8(preDecoders_2_io_in_data_8),
    .io_out_pd_0_isRVC(preDecoders_2_io_out_pd_0_isRVC),
    .io_out_pd_0_brType(preDecoders_2_io_out_pd_0_brType),
    .io_out_pd_0_isCall(preDecoders_2_io_out_pd_0_isCall),
    .io_out_pd_0_isRet(preDecoders_2_io_out_pd_0_isRet),
    .io_out_pd_1_valid(preDecoders_2_io_out_pd_1_valid),
    .io_out_pd_1_isRVC(preDecoders_2_io_out_pd_1_isRVC),
    .io_out_pd_1_brType(preDecoders_2_io_out_pd_1_brType),
    .io_out_pd_1_isCall(preDecoders_2_io_out_pd_1_isCall),
    .io_out_pd_1_isRet(preDecoders_2_io_out_pd_1_isRet),
    .io_out_pd_2_valid(preDecoders_2_io_out_pd_2_valid),
    .io_out_pd_2_isRVC(preDecoders_2_io_out_pd_2_isRVC),
    .io_out_pd_2_brType(preDecoders_2_io_out_pd_2_brType),
    .io_out_pd_2_isCall(preDecoders_2_io_out_pd_2_isCall),
    .io_out_pd_2_isRet(preDecoders_2_io_out_pd_2_isRet),
    .io_out_pd_3_valid(preDecoders_2_io_out_pd_3_valid),
    .io_out_pd_3_isRVC(preDecoders_2_io_out_pd_3_isRVC),
    .io_out_pd_3_brType(preDecoders_2_io_out_pd_3_brType),
    .io_out_pd_3_isCall(preDecoders_2_io_out_pd_3_isCall),
    .io_out_pd_3_isRet(preDecoders_2_io_out_pd_3_isRet),
    .io_out_pd_4_valid(preDecoders_2_io_out_pd_4_valid),
    .io_out_pd_4_isRVC(preDecoders_2_io_out_pd_4_isRVC),
    .io_out_pd_4_brType(preDecoders_2_io_out_pd_4_brType),
    .io_out_pd_4_isCall(preDecoders_2_io_out_pd_4_isCall),
    .io_out_pd_4_isRet(preDecoders_2_io_out_pd_4_isRet),
    .io_out_pd_5_valid(preDecoders_2_io_out_pd_5_valid),
    .io_out_pd_5_isRVC(preDecoders_2_io_out_pd_5_isRVC),
    .io_out_pd_5_brType(preDecoders_2_io_out_pd_5_brType),
    .io_out_pd_5_isCall(preDecoders_2_io_out_pd_5_isCall),
    .io_out_pd_5_isRet(preDecoders_2_io_out_pd_5_isRet),
    .io_out_pd_6_valid(preDecoders_2_io_out_pd_6_valid),
    .io_out_pd_6_isRVC(preDecoders_2_io_out_pd_6_isRVC),
    .io_out_pd_6_brType(preDecoders_2_io_out_pd_6_brType),
    .io_out_pd_6_isCall(preDecoders_2_io_out_pd_6_isCall),
    .io_out_pd_6_isRet(preDecoders_2_io_out_pd_6_isRet),
    .io_out_pd_7_valid(preDecoders_2_io_out_pd_7_valid),
    .io_out_pd_7_isRVC(preDecoders_2_io_out_pd_7_isRVC),
    .io_out_pd_7_brType(preDecoders_2_io_out_pd_7_brType),
    .io_out_pd_7_isCall(preDecoders_2_io_out_pd_7_isCall),
    .io_out_pd_7_isRet(preDecoders_2_io_out_pd_7_isRet),
    .io_out_hasHalfValid_2(preDecoders_2_io_out_hasHalfValid_2),
    .io_out_hasHalfValid_3(preDecoders_2_io_out_hasHalfValid_3),
    .io_out_hasHalfValid_4(preDecoders_2_io_out_hasHalfValid_4),
    .io_out_hasHalfValid_5(preDecoders_2_io_out_hasHalfValid_5),
    .io_out_hasHalfValid_6(preDecoders_2_io_out_hasHalfValid_6),
    .io_out_hasHalfValid_7(preDecoders_2_io_out_hasHalfValid_7),
    .io_out_instr_0(preDecoders_2_io_out_instr_0),
    .io_out_instr_1(preDecoders_2_io_out_instr_1),
    .io_out_instr_2(preDecoders_2_io_out_instr_2),
    .io_out_instr_3(preDecoders_2_io_out_instr_3),
    .io_out_instr_4(preDecoders_2_io_out_instr_4),
    .io_out_instr_5(preDecoders_2_io_out_instr_5),
    .io_out_instr_6(preDecoders_2_io_out_instr_6),
    .io_out_instr_7(preDecoders_2_io_out_instr_7),
    .io_out_jumpOffset_0(preDecoders_2_io_out_jumpOffset_0),
    .io_out_jumpOffset_1(preDecoders_2_io_out_jumpOffset_1),
    .io_out_jumpOffset_2(preDecoders_2_io_out_jumpOffset_2),
    .io_out_jumpOffset_3(preDecoders_2_io_out_jumpOffset_3),
    .io_out_jumpOffset_4(preDecoders_2_io_out_jumpOffset_4),
    .io_out_jumpOffset_5(preDecoders_2_io_out_jumpOffset_5),
    .io_out_jumpOffset_6(preDecoders_2_io_out_jumpOffset_6),
    .io_out_jumpOffset_7(preDecoders_2_io_out_jumpOffset_7)
  );
  PreDecode preDecoders_3 ( // @[IFU.scala 142:46]
    .io_in_data_0(preDecoders_3_io_in_data_0),
    .io_in_data_1(preDecoders_3_io_in_data_1),
    .io_in_data_2(preDecoders_3_io_in_data_2),
    .io_in_data_3(preDecoders_3_io_in_data_3),
    .io_in_data_4(preDecoders_3_io_in_data_4),
    .io_in_data_5(preDecoders_3_io_in_data_5),
    .io_in_data_6(preDecoders_3_io_in_data_6),
    .io_in_data_7(preDecoders_3_io_in_data_7),
    .io_in_data_8(preDecoders_3_io_in_data_8),
    .io_out_pd_0_isRVC(preDecoders_3_io_out_pd_0_isRVC),
    .io_out_pd_0_brType(preDecoders_3_io_out_pd_0_brType),
    .io_out_pd_0_isCall(preDecoders_3_io_out_pd_0_isCall),
    .io_out_pd_0_isRet(preDecoders_3_io_out_pd_0_isRet),
    .io_out_pd_1_valid(preDecoders_3_io_out_pd_1_valid),
    .io_out_pd_1_isRVC(preDecoders_3_io_out_pd_1_isRVC),
    .io_out_pd_1_brType(preDecoders_3_io_out_pd_1_brType),
    .io_out_pd_1_isCall(preDecoders_3_io_out_pd_1_isCall),
    .io_out_pd_1_isRet(preDecoders_3_io_out_pd_1_isRet),
    .io_out_pd_2_valid(preDecoders_3_io_out_pd_2_valid),
    .io_out_pd_2_isRVC(preDecoders_3_io_out_pd_2_isRVC),
    .io_out_pd_2_brType(preDecoders_3_io_out_pd_2_brType),
    .io_out_pd_2_isCall(preDecoders_3_io_out_pd_2_isCall),
    .io_out_pd_2_isRet(preDecoders_3_io_out_pd_2_isRet),
    .io_out_pd_3_valid(preDecoders_3_io_out_pd_3_valid),
    .io_out_pd_3_isRVC(preDecoders_3_io_out_pd_3_isRVC),
    .io_out_pd_3_brType(preDecoders_3_io_out_pd_3_brType),
    .io_out_pd_3_isCall(preDecoders_3_io_out_pd_3_isCall),
    .io_out_pd_3_isRet(preDecoders_3_io_out_pd_3_isRet),
    .io_out_pd_4_valid(preDecoders_3_io_out_pd_4_valid),
    .io_out_pd_4_isRVC(preDecoders_3_io_out_pd_4_isRVC),
    .io_out_pd_4_brType(preDecoders_3_io_out_pd_4_brType),
    .io_out_pd_4_isCall(preDecoders_3_io_out_pd_4_isCall),
    .io_out_pd_4_isRet(preDecoders_3_io_out_pd_4_isRet),
    .io_out_pd_5_valid(preDecoders_3_io_out_pd_5_valid),
    .io_out_pd_5_isRVC(preDecoders_3_io_out_pd_5_isRVC),
    .io_out_pd_5_brType(preDecoders_3_io_out_pd_5_brType),
    .io_out_pd_5_isCall(preDecoders_3_io_out_pd_5_isCall),
    .io_out_pd_5_isRet(preDecoders_3_io_out_pd_5_isRet),
    .io_out_pd_6_valid(preDecoders_3_io_out_pd_6_valid),
    .io_out_pd_6_isRVC(preDecoders_3_io_out_pd_6_isRVC),
    .io_out_pd_6_brType(preDecoders_3_io_out_pd_6_brType),
    .io_out_pd_6_isCall(preDecoders_3_io_out_pd_6_isCall),
    .io_out_pd_6_isRet(preDecoders_3_io_out_pd_6_isRet),
    .io_out_pd_7_valid(preDecoders_3_io_out_pd_7_valid),
    .io_out_pd_7_isRVC(preDecoders_3_io_out_pd_7_isRVC),
    .io_out_pd_7_brType(preDecoders_3_io_out_pd_7_brType),
    .io_out_pd_7_isCall(preDecoders_3_io_out_pd_7_isCall),
    .io_out_pd_7_isRet(preDecoders_3_io_out_pd_7_isRet),
    .io_out_hasHalfValid_2(preDecoders_3_io_out_hasHalfValid_2),
    .io_out_hasHalfValid_3(preDecoders_3_io_out_hasHalfValid_3),
    .io_out_hasHalfValid_4(preDecoders_3_io_out_hasHalfValid_4),
    .io_out_hasHalfValid_5(preDecoders_3_io_out_hasHalfValid_5),
    .io_out_hasHalfValid_6(preDecoders_3_io_out_hasHalfValid_6),
    .io_out_hasHalfValid_7(preDecoders_3_io_out_hasHalfValid_7),
    .io_out_instr_0(preDecoders_3_io_out_instr_0),
    .io_out_instr_1(preDecoders_3_io_out_instr_1),
    .io_out_instr_2(preDecoders_3_io_out_instr_2),
    .io_out_instr_3(preDecoders_3_io_out_instr_3),
    .io_out_instr_4(preDecoders_3_io_out_instr_4),
    .io_out_instr_5(preDecoders_3_io_out_instr_5),
    .io_out_instr_6(preDecoders_3_io_out_instr_6),
    .io_out_instr_7(preDecoders_3_io_out_instr_7),
    .io_out_jumpOffset_0(preDecoders_3_io_out_jumpOffset_0),
    .io_out_jumpOffset_1(preDecoders_3_io_out_jumpOffset_1),
    .io_out_jumpOffset_2(preDecoders_3_io_out_jumpOffset_2),
    .io_out_jumpOffset_3(preDecoders_3_io_out_jumpOffset_3),
    .io_out_jumpOffset_4(preDecoders_3_io_out_jumpOffset_4),
    .io_out_jumpOffset_5(preDecoders_3_io_out_jumpOffset_5),
    .io_out_jumpOffset_6(preDecoders_3_io_out_jumpOffset_6),
    .io_out_jumpOffset_7(preDecoders_3_io_out_jumpOffset_7)
  );
  PredChecker predChecker ( // @[IFU.scala 144:31]
    .clock(predChecker_clock),
    .io_in_ftqOffset_valid(predChecker_io_in_ftqOffset_valid),
    .io_in_ftqOffset_bits(predChecker_io_in_ftqOffset_bits),
    .io_in_jumpOffset_0(predChecker_io_in_jumpOffset_0),
    .io_in_jumpOffset_1(predChecker_io_in_jumpOffset_1),
    .io_in_jumpOffset_2(predChecker_io_in_jumpOffset_2),
    .io_in_jumpOffset_3(predChecker_io_in_jumpOffset_3),
    .io_in_jumpOffset_4(predChecker_io_in_jumpOffset_4),
    .io_in_jumpOffset_5(predChecker_io_in_jumpOffset_5),
    .io_in_jumpOffset_6(predChecker_io_in_jumpOffset_6),
    .io_in_jumpOffset_7(predChecker_io_in_jumpOffset_7),
    .io_in_target(predChecker_io_in_target),
    .io_in_instrRange_0(predChecker_io_in_instrRange_0),
    .io_in_instrRange_1(predChecker_io_in_instrRange_1),
    .io_in_instrRange_2(predChecker_io_in_instrRange_2),
    .io_in_instrRange_3(predChecker_io_in_instrRange_3),
    .io_in_instrRange_4(predChecker_io_in_instrRange_4),
    .io_in_instrRange_5(predChecker_io_in_instrRange_5),
    .io_in_instrRange_6(predChecker_io_in_instrRange_6),
    .io_in_instrRange_7(predChecker_io_in_instrRange_7),
    .io_in_instrValid_0(predChecker_io_in_instrValid_0),
    .io_in_instrValid_1(predChecker_io_in_instrValid_1),
    .io_in_instrValid_2(predChecker_io_in_instrValid_2),
    .io_in_instrValid_3(predChecker_io_in_instrValid_3),
    .io_in_instrValid_4(predChecker_io_in_instrValid_4),
    .io_in_instrValid_5(predChecker_io_in_instrValid_5),
    .io_in_instrValid_6(predChecker_io_in_instrValid_6),
    .io_in_instrValid_7(predChecker_io_in_instrValid_7),
    .io_in_pds_0_isRVC(predChecker_io_in_pds_0_isRVC),
    .io_in_pds_0_brType(predChecker_io_in_pds_0_brType),
    .io_in_pds_0_isRet(predChecker_io_in_pds_0_isRet),
    .io_in_pds_1_isRVC(predChecker_io_in_pds_1_isRVC),
    .io_in_pds_1_brType(predChecker_io_in_pds_1_brType),
    .io_in_pds_1_isRet(predChecker_io_in_pds_1_isRet),
    .io_in_pds_2_isRVC(predChecker_io_in_pds_2_isRVC),
    .io_in_pds_2_brType(predChecker_io_in_pds_2_brType),
    .io_in_pds_2_isRet(predChecker_io_in_pds_2_isRet),
    .io_in_pds_3_isRVC(predChecker_io_in_pds_3_isRVC),
    .io_in_pds_3_brType(predChecker_io_in_pds_3_brType),
    .io_in_pds_3_isRet(predChecker_io_in_pds_3_isRet),
    .io_in_pds_4_isRVC(predChecker_io_in_pds_4_isRVC),
    .io_in_pds_4_brType(predChecker_io_in_pds_4_brType),
    .io_in_pds_4_isRet(predChecker_io_in_pds_4_isRet),
    .io_in_pds_5_isRVC(predChecker_io_in_pds_5_isRVC),
    .io_in_pds_5_brType(predChecker_io_in_pds_5_brType),
    .io_in_pds_5_isRet(predChecker_io_in_pds_5_isRet),
    .io_in_pds_6_isRVC(predChecker_io_in_pds_6_isRVC),
    .io_in_pds_6_brType(predChecker_io_in_pds_6_brType),
    .io_in_pds_6_isRet(predChecker_io_in_pds_6_isRet),
    .io_in_pds_7_isRVC(predChecker_io_in_pds_7_isRVC),
    .io_in_pds_7_brType(predChecker_io_in_pds_7_brType),
    .io_in_pds_7_isRet(predChecker_io_in_pds_7_isRet),
    .io_in_pc_0(predChecker_io_in_pc_0),
    .io_in_pc_1(predChecker_io_in_pc_1),
    .io_in_pc_2(predChecker_io_in_pc_2),
    .io_in_pc_3(predChecker_io_in_pc_3),
    .io_in_pc_4(predChecker_io_in_pc_4),
    .io_in_pc_5(predChecker_io_in_pc_5),
    .io_in_pc_6(predChecker_io_in_pc_6),
    .io_in_pc_7(predChecker_io_in_pc_7),
    .io_out_stage1Out_fixedRange_0(predChecker_io_out_stage1Out_fixedRange_0),
    .io_out_stage1Out_fixedRange_1(predChecker_io_out_stage1Out_fixedRange_1),
    .io_out_stage1Out_fixedRange_2(predChecker_io_out_stage1Out_fixedRange_2),
    .io_out_stage1Out_fixedRange_3(predChecker_io_out_stage1Out_fixedRange_3),
    .io_out_stage1Out_fixedRange_4(predChecker_io_out_stage1Out_fixedRange_4),
    .io_out_stage1Out_fixedRange_5(predChecker_io_out_stage1Out_fixedRange_5),
    .io_out_stage1Out_fixedRange_6(predChecker_io_out_stage1Out_fixedRange_6),
    .io_out_stage1Out_fixedRange_7(predChecker_io_out_stage1Out_fixedRange_7),
    .io_out_stage1Out_fixedTaken_0(predChecker_io_out_stage1Out_fixedTaken_0),
    .io_out_stage1Out_fixedTaken_1(predChecker_io_out_stage1Out_fixedTaken_1),
    .io_out_stage1Out_fixedTaken_2(predChecker_io_out_stage1Out_fixedTaken_2),
    .io_out_stage1Out_fixedTaken_3(predChecker_io_out_stage1Out_fixedTaken_3),
    .io_out_stage1Out_fixedTaken_4(predChecker_io_out_stage1Out_fixedTaken_4),
    .io_out_stage1Out_fixedTaken_5(predChecker_io_out_stage1Out_fixedTaken_5),
    .io_out_stage1Out_fixedTaken_6(predChecker_io_out_stage1Out_fixedTaken_6),
    .io_out_stage1Out_fixedTaken_7(predChecker_io_out_stage1Out_fixedTaken_7),
    .io_out_stage2Out_fixedTarget_0(predChecker_io_out_stage2Out_fixedTarget_0),
    .io_out_stage2Out_fixedTarget_1(predChecker_io_out_stage2Out_fixedTarget_1),
    .io_out_stage2Out_fixedTarget_2(predChecker_io_out_stage2Out_fixedTarget_2),
    .io_out_stage2Out_fixedTarget_3(predChecker_io_out_stage2Out_fixedTarget_3),
    .io_out_stage2Out_fixedTarget_4(predChecker_io_out_stage2Out_fixedTarget_4),
    .io_out_stage2Out_fixedTarget_5(predChecker_io_out_stage2Out_fixedTarget_5),
    .io_out_stage2Out_fixedTarget_6(predChecker_io_out_stage2Out_fixedTarget_6),
    .io_out_stage2Out_fixedTarget_7(predChecker_io_out_stage2Out_fixedTarget_7),
    .io_out_stage2Out_fixedMissPred_0(predChecker_io_out_stage2Out_fixedMissPred_0),
    .io_out_stage2Out_fixedMissPred_1(predChecker_io_out_stage2Out_fixedMissPred_1),
    .io_out_stage2Out_fixedMissPred_2(predChecker_io_out_stage2Out_fixedMissPred_2),
    .io_out_stage2Out_fixedMissPred_3(predChecker_io_out_stage2Out_fixedMissPred_3),
    .io_out_stage2Out_fixedMissPred_4(predChecker_io_out_stage2Out_fixedMissPred_4),
    .io_out_stage2Out_fixedMissPred_5(predChecker_io_out_stage2Out_fixedMissPred_5),
    .io_out_stage2Out_fixedMissPred_6(predChecker_io_out_stage2Out_fixedMissPred_6),
    .io_out_stage2Out_fixedMissPred_7(predChecker_io_out_stage2Out_fixedMissPred_7),
    .io_out_stage2Out_faultType_0_value(predChecker_io_out_stage2Out_faultType_0_value),
    .io_out_stage2Out_faultType_1_value(predChecker_io_out_stage2Out_faultType_1_value),
    .io_out_stage2Out_faultType_2_value(predChecker_io_out_stage2Out_faultType_2_value),
    .io_out_stage2Out_faultType_3_value(predChecker_io_out_stage2Out_faultType_3_value),
    .io_out_stage2Out_faultType_4_value(predChecker_io_out_stage2Out_faultType_4_value),
    .io_out_stage2Out_faultType_5_value(predChecker_io_out_stage2Out_faultType_5_value),
    .io_out_stage2Out_faultType_6_value(predChecker_io_out_stage2Out_faultType_6_value),
    .io_out_stage2Out_faultType_7_value(predChecker_io_out_stage2Out_faultType_7_value)
  );
  FrontendTrigger frontendTrigger ( // @[IFU.scala 145:31]
    .clock(frontendTrigger_clock),
    .reset(frontendTrigger_reset),
    .io_frontendTrigger_t_valid(frontendTrigger_io_frontendTrigger_t_valid),
    .io_frontendTrigger_t_bits_addr(frontendTrigger_io_frontendTrigger_t_bits_addr),
    .io_frontendTrigger_t_bits_tdata_matchType(frontendTrigger_io_frontendTrigger_t_bits_tdata_matchType),
    .io_frontendTrigger_t_bits_tdata_select(frontendTrigger_io_frontendTrigger_t_bits_tdata_select),
    .io_frontendTrigger_t_bits_tdata_timing(frontendTrigger_io_frontendTrigger_t_bits_tdata_timing),
    .io_frontendTrigger_t_bits_tdata_chain(frontendTrigger_io_frontendTrigger_t_bits_tdata_chain),
    .io_frontendTrigger_t_bits_tdata_tdata2(frontendTrigger_io_frontendTrigger_t_bits_tdata_tdata2),
    .io_csrTriggerEnable_0(frontendTrigger_io_csrTriggerEnable_0),
    .io_csrTriggerEnable_1(frontendTrigger_io_csrTriggerEnable_1),
    .io_csrTriggerEnable_2(frontendTrigger_io_csrTriggerEnable_2),
    .io_csrTriggerEnable_3(frontendTrigger_io_csrTriggerEnable_3),
    .io_triggered_0_frontendHit_0(frontendTrigger_io_triggered_0_frontendHit_0),
    .io_triggered_0_frontendHit_1(frontendTrigger_io_triggered_0_frontendHit_1),
    .io_triggered_0_frontendHit_2(frontendTrigger_io_triggered_0_frontendHit_2),
    .io_triggered_0_frontendHit_3(frontendTrigger_io_triggered_0_frontendHit_3),
    .io_triggered_0_backendEn_0(frontendTrigger_io_triggered_0_backendEn_0),
    .io_triggered_0_backendEn_1(frontendTrigger_io_triggered_0_backendEn_1),
    .io_triggered_1_frontendHit_0(frontendTrigger_io_triggered_1_frontendHit_0),
    .io_triggered_1_frontendHit_1(frontendTrigger_io_triggered_1_frontendHit_1),
    .io_triggered_1_frontendHit_2(frontendTrigger_io_triggered_1_frontendHit_2),
    .io_triggered_1_frontendHit_3(frontendTrigger_io_triggered_1_frontendHit_3),
    .io_triggered_1_backendEn_0(frontendTrigger_io_triggered_1_backendEn_0),
    .io_triggered_1_backendEn_1(frontendTrigger_io_triggered_1_backendEn_1),
    .io_triggered_2_frontendHit_0(frontendTrigger_io_triggered_2_frontendHit_0),
    .io_triggered_2_frontendHit_1(frontendTrigger_io_triggered_2_frontendHit_1),
    .io_triggered_2_frontendHit_2(frontendTrigger_io_triggered_2_frontendHit_2),
    .io_triggered_2_frontendHit_3(frontendTrigger_io_triggered_2_frontendHit_3),
    .io_triggered_2_backendEn_0(frontendTrigger_io_triggered_2_backendEn_0),
    .io_triggered_2_backendEn_1(frontendTrigger_io_triggered_2_backendEn_1),
    .io_triggered_3_frontendHit_0(frontendTrigger_io_triggered_3_frontendHit_0),
    .io_triggered_3_frontendHit_1(frontendTrigger_io_triggered_3_frontendHit_1),
    .io_triggered_3_frontendHit_2(frontendTrigger_io_triggered_3_frontendHit_2),
    .io_triggered_3_frontendHit_3(frontendTrigger_io_triggered_3_frontendHit_3),
    .io_triggered_3_backendEn_0(frontendTrigger_io_triggered_3_backendEn_0),
    .io_triggered_3_backendEn_1(frontendTrigger_io_triggered_3_backendEn_1),
    .io_triggered_4_frontendHit_0(frontendTrigger_io_triggered_4_frontendHit_0),
    .io_triggered_4_frontendHit_1(frontendTrigger_io_triggered_4_frontendHit_1),
    .io_triggered_4_frontendHit_2(frontendTrigger_io_triggered_4_frontendHit_2),
    .io_triggered_4_frontendHit_3(frontendTrigger_io_triggered_4_frontendHit_3),
    .io_triggered_4_backendEn_0(frontendTrigger_io_triggered_4_backendEn_0),
    .io_triggered_4_backendEn_1(frontendTrigger_io_triggered_4_backendEn_1),
    .io_triggered_5_frontendHit_0(frontendTrigger_io_triggered_5_frontendHit_0),
    .io_triggered_5_frontendHit_1(frontendTrigger_io_triggered_5_frontendHit_1),
    .io_triggered_5_frontendHit_2(frontendTrigger_io_triggered_5_frontendHit_2),
    .io_triggered_5_frontendHit_3(frontendTrigger_io_triggered_5_frontendHit_3),
    .io_triggered_5_backendEn_0(frontendTrigger_io_triggered_5_backendEn_0),
    .io_triggered_5_backendEn_1(frontendTrigger_io_triggered_5_backendEn_1),
    .io_triggered_6_frontendHit_0(frontendTrigger_io_triggered_6_frontendHit_0),
    .io_triggered_6_frontendHit_1(frontendTrigger_io_triggered_6_frontendHit_1),
    .io_triggered_6_frontendHit_2(frontendTrigger_io_triggered_6_frontendHit_2),
    .io_triggered_6_frontendHit_3(frontendTrigger_io_triggered_6_frontendHit_3),
    .io_triggered_6_backendEn_0(frontendTrigger_io_triggered_6_backendEn_0),
    .io_triggered_6_backendEn_1(frontendTrigger_io_triggered_6_backendEn_1),
    .io_triggered_7_frontendHit_0(frontendTrigger_io_triggered_7_frontendHit_0),
    .io_triggered_7_frontendHit_1(frontendTrigger_io_triggered_7_frontendHit_1),
    .io_triggered_7_frontendHit_2(frontendTrigger_io_triggered_7_frontendHit_2),
    .io_triggered_7_frontendHit_3(frontendTrigger_io_triggered_7_frontendHit_3),
    .io_triggered_7_backendEn_0(frontendTrigger_io_triggered_7_backendEn_0),
    .io_triggered_7_backendEn_1(frontendTrigger_io_triggered_7_backendEn_1),
    .io_pds_0_isRVC(frontendTrigger_io_pds_0_isRVC),
    .io_pds_1_isRVC(frontendTrigger_io_pds_1_isRVC),
    .io_pds_2_isRVC(frontendTrigger_io_pds_2_isRVC),
    .io_pds_3_isRVC(frontendTrigger_io_pds_3_isRVC),
    .io_pds_4_isRVC(frontendTrigger_io_pds_4_isRVC),
    .io_pds_5_isRVC(frontendTrigger_io_pds_5_isRVC),
    .io_pds_6_isRVC(frontendTrigger_io_pds_6_isRVC),
    .io_pds_7_isRVC(frontendTrigger_io_pds_7_isRVC),
    .io_pc_0(frontendTrigger_io_pc_0),
    .io_pc_1(frontendTrigger_io_pc_1),
    .io_pc_2(frontendTrigger_io_pc_2),
    .io_pc_3(frontendTrigger_io_pc_3),
    .io_pc_4(frontendTrigger_io_pc_4),
    .io_pc_5(frontendTrigger_io_pc_5),
    .io_pc_6(frontendTrigger_io_pc_6),
    .io_pc_7(frontendTrigger_io_pc_7),
    .io_data_0(frontendTrigger_io_data_0),
    .io_data_1(frontendTrigger_io_data_1),
    .io_data_2(frontendTrigger_io_data_2),
    .io_data_3(frontendTrigger_io_data_3),
    .io_data_4(frontendTrigger_io_data_4),
    .io_data_5(frontendTrigger_io_data_5),
    .io_data_6(frontendTrigger_io_data_6),
    .io_data_7(frontendTrigger_io_data_7),
    .io_data_8(frontendTrigger_io_data_8)
  );
  RVCExpander f3_expd_instr_expander ( // @[IFU.scala 382:32]
    .io_in(f3_expd_instr_expander_io_in),
    .io_out_bits(f3_expd_instr_expander_io_out_bits)
  );
  RVCExpander f3_expd_instr_expander_1 ( // @[IFU.scala 382:32]
    .io_in(f3_expd_instr_expander_1_io_in),
    .io_out_bits(f3_expd_instr_expander_1_io_out_bits)
  );
  RVCExpander f3_expd_instr_expander_2 ( // @[IFU.scala 382:32]
    .io_in(f3_expd_instr_expander_2_io_in),
    .io_out_bits(f3_expd_instr_expander_2_io_out_bits)
  );
  RVCExpander f3_expd_instr_expander_3 ( // @[IFU.scala 382:32]
    .io_in(f3_expd_instr_expander_3_io_in),
    .io_out_bits(f3_expd_instr_expander_3_io_out_bits)
  );
  RVCExpander f3_expd_instr_expander_4 ( // @[IFU.scala 382:32]
    .io_in(f3_expd_instr_expander_4_io_in),
    .io_out_bits(f3_expd_instr_expander_4_io_out_bits)
  );
  RVCExpander f3_expd_instr_expander_5 ( // @[IFU.scala 382:32]
    .io_in(f3_expd_instr_expander_5_io_in),
    .io_out_bits(f3_expd_instr_expander_5_io_out_bits)
  );
  RVCExpander f3_expd_instr_expander_6 ( // @[IFU.scala 382:32]
    .io_in(f3_expd_instr_expander_6_io_in),
    .io_out_bits(f3_expd_instr_expander_6_io_out_bits)
  );
  RVCExpander f3_expd_instr_expander_7 ( // @[IFU.scala 382:32]
    .io_in(f3_expd_instr_expander_7_io_in),
    .io_out_bits(f3_expd_instr_expander_7_io_out_bits)
  );
  FetchToIBuffer0Writer #(.site("IFU0")) writer ( // @[ChiselDB.scala 132:24]
    .clock(writer_clock),
    .reset(writer_reset),
    .en(writer_en),
    .stamp(writer_stamp),
    .data_start_addr(writer_data_start_addr),
    .data_instr_count(writer_data_instr_count),
    .data_exception(writer_data_exception),
    .data_is_cache_hit(writer_data_is_cache_hit)
  );
  IfuWbToFtq0Writer #(.site("IFU0")) writer_1 ( // @[ChiselDB.scala 132:24]
    .clock(writer_1_clock),
    .reset(writer_1_reset),
    .en(writer_1_en),
    .stamp(writer_1_stamp),
    .data_start_addr(writer_1_data_start_addr),
    .data_is_miss_pred(writer_1_data_is_miss_pred),
    .data_miss_pred_offset(writer_1_data_miss_pred_offset),
    .data_checkJalFault(writer_1_data_checkJalFault),
    .data_checkRetFault(writer_1_data_checkRetFault),
    .data_checkTargetFault(writer_1_data_checkTargetFault),
    .data_checkNotCFIFault(writer_1_data_checkNotCFIFault),
    .data_checkInvalidTaken(writer_1_data_checkInvalidTaken)
  );
  assign io_ftqInter_fromFtq_req_ready = f1_ready & io_icacheInter_icacheReady; // @[IFU.scala 181:33]
  assign io_ftqInter_toFtq_pdWb_valid = wb_valid ? wb_valid : mmioFlushWb_valid; // @[IFU.scala 763:20]
  assign io_ftqInter_toFtq_pdWb_bits_pc_0 = wb_valid ? wb_pc_0 : f3_pc_0; // @[IFU.scala 763:20]
  assign io_ftqInter_toFtq_pdWb_bits_pc_1 = wb_valid ? wb_pc_1 : f3_pc_1; // @[IFU.scala 763:20]
  assign io_ftqInter_toFtq_pdWb_bits_pc_2 = wb_valid ? wb_pc_2 : f3_pc_2; // @[IFU.scala 763:20]
  assign io_ftqInter_toFtq_pdWb_bits_pc_3 = wb_valid ? wb_pc_3 : f3_pc_3; // @[IFU.scala 763:20]
  assign io_ftqInter_toFtq_pdWb_bits_pc_4 = wb_valid ? wb_pc_4 : f3_pc_4; // @[IFU.scala 763:20]
  assign io_ftqInter_toFtq_pdWb_bits_pc_5 = wb_valid ? wb_pc_5 : f3_pc_5; // @[IFU.scala 763:20]
  assign io_ftqInter_toFtq_pdWb_bits_pc_6 = wb_valid ? wb_pc_6 : f3_pc_6; // @[IFU.scala 763:20]
  assign io_ftqInter_toFtq_pdWb_bits_pc_7 = wb_valid ? wb_pc_7 : f3_pc_7; // @[IFU.scala 763:20]
  assign io_ftqInter_toFtq_pdWb_bits_pd_0_valid = wb_valid ? wb_instr_valid_0 : 1'h1; // @[IFU.scala 763:20]
  assign io_ftqInter_toFtq_pdWb_bits_pd_0_isRVC = wb_valid ? wb_pd_0_isRVC : mmioFlushWb_bits_pd_0_isRVC; // @[IFU.scala 763:20]
  assign io_ftqInter_toFtq_pdWb_bits_pd_0_brType = wb_valid ? wb_pd_0_brType : mmioFlushWb_bits_pd_0_brType; // @[IFU.scala 763:20]
  assign io_ftqInter_toFtq_pdWb_bits_pd_0_isCall = wb_valid ? wb_pd_0_isCall : mmioFlushWb_bits_pd_0_isCall; // @[IFU.scala 763:20]
  assign io_ftqInter_toFtq_pdWb_bits_pd_0_isRet = wb_valid ? wb_pd_0_isRet : mmioFlushWb_bits_pd_0_isRet; // @[IFU.scala 763:20]
  assign io_ftqInter_toFtq_pdWb_bits_pd_1_valid = wb_valid & wb_instr_valid_1; // @[IFU.scala 763:20]
  assign io_ftqInter_toFtq_pdWb_bits_pd_1_isRVC = wb_valid ? wb_pd_1_isRVC : f3_pd_1_isRVC; // @[IFU.scala 763:20]
  assign io_ftqInter_toFtq_pdWb_bits_pd_1_brType = wb_valid ? wb_pd_1_brType : f3_pd_1_brType; // @[IFU.scala 763:20]
  assign io_ftqInter_toFtq_pdWb_bits_pd_1_isCall = wb_valid ? wb_pd_1_isCall : f3_pd_1_isCall; // @[IFU.scala 763:20]
  assign io_ftqInter_toFtq_pdWb_bits_pd_1_isRet = wb_valid ? wb_pd_1_isRet : f3_pd_1_isRet; // @[IFU.scala 763:20]
  assign io_ftqInter_toFtq_pdWb_bits_pd_2_valid = wb_valid & wb_instr_valid_2; // @[IFU.scala 763:20]
  assign io_ftqInter_toFtq_pdWb_bits_pd_2_isRVC = wb_valid ? wb_pd_2_isRVC : f3_pd_2_isRVC; // @[IFU.scala 763:20]
  assign io_ftqInter_toFtq_pdWb_bits_pd_2_brType = wb_valid ? wb_pd_2_brType : f3_pd_2_brType; // @[IFU.scala 763:20]
  assign io_ftqInter_toFtq_pdWb_bits_pd_2_isCall = wb_valid ? wb_pd_2_isCall : f3_pd_2_isCall; // @[IFU.scala 763:20]
  assign io_ftqInter_toFtq_pdWb_bits_pd_2_isRet = wb_valid ? wb_pd_2_isRet : f3_pd_2_isRet; // @[IFU.scala 763:20]
  assign io_ftqInter_toFtq_pdWb_bits_pd_3_valid = wb_valid & wb_instr_valid_3; // @[IFU.scala 763:20]
  assign io_ftqInter_toFtq_pdWb_bits_pd_3_isRVC = wb_valid ? wb_pd_3_isRVC : f3_pd_3_isRVC; // @[IFU.scala 763:20]
  assign io_ftqInter_toFtq_pdWb_bits_pd_3_brType = wb_valid ? wb_pd_3_brType : f3_pd_3_brType; // @[IFU.scala 763:20]
  assign io_ftqInter_toFtq_pdWb_bits_pd_3_isCall = wb_valid ? wb_pd_3_isCall : f3_pd_3_isCall; // @[IFU.scala 763:20]
  assign io_ftqInter_toFtq_pdWb_bits_pd_3_isRet = wb_valid ? wb_pd_3_isRet : f3_pd_3_isRet; // @[IFU.scala 763:20]
  assign io_ftqInter_toFtq_pdWb_bits_pd_4_valid = wb_valid & wb_instr_valid_4; // @[IFU.scala 763:20]
  assign io_ftqInter_toFtq_pdWb_bits_pd_4_isRVC = wb_valid ? wb_pd_4_isRVC : f3_pd_4_isRVC; // @[IFU.scala 763:20]
  assign io_ftqInter_toFtq_pdWb_bits_pd_4_brType = wb_valid ? wb_pd_4_brType : f3_pd_4_brType; // @[IFU.scala 763:20]
  assign io_ftqInter_toFtq_pdWb_bits_pd_4_isCall = wb_valid ? wb_pd_4_isCall : f3_pd_4_isCall; // @[IFU.scala 763:20]
  assign io_ftqInter_toFtq_pdWb_bits_pd_4_isRet = wb_valid ? wb_pd_4_isRet : f3_pd_4_isRet; // @[IFU.scala 763:20]
  assign io_ftqInter_toFtq_pdWb_bits_pd_5_valid = wb_valid & wb_instr_valid_5; // @[IFU.scala 763:20]
  assign io_ftqInter_toFtq_pdWb_bits_pd_5_isRVC = wb_valid ? wb_pd_5_isRVC : f3_pd_5_isRVC; // @[IFU.scala 763:20]
  assign io_ftqInter_toFtq_pdWb_bits_pd_5_brType = wb_valid ? wb_pd_5_brType : f3_pd_5_brType; // @[IFU.scala 763:20]
  assign io_ftqInter_toFtq_pdWb_bits_pd_5_isCall = wb_valid ? wb_pd_5_isCall : f3_pd_5_isCall; // @[IFU.scala 763:20]
  assign io_ftqInter_toFtq_pdWb_bits_pd_5_isRet = wb_valid ? wb_pd_5_isRet : f3_pd_5_isRet; // @[IFU.scala 763:20]
  assign io_ftqInter_toFtq_pdWb_bits_pd_6_valid = wb_valid & wb_instr_valid_6; // @[IFU.scala 763:20]
  assign io_ftqInter_toFtq_pdWb_bits_pd_6_isRVC = wb_valid ? wb_pd_6_isRVC : f3_pd_6_isRVC; // @[IFU.scala 763:20]
  assign io_ftqInter_toFtq_pdWb_bits_pd_6_brType = wb_valid ? wb_pd_6_brType : f3_pd_6_brType; // @[IFU.scala 763:20]
  assign io_ftqInter_toFtq_pdWb_bits_pd_6_isCall = wb_valid ? wb_pd_6_isCall : f3_pd_6_isCall; // @[IFU.scala 763:20]
  assign io_ftqInter_toFtq_pdWb_bits_pd_6_isRet = wb_valid ? wb_pd_6_isRet : f3_pd_6_isRet; // @[IFU.scala 763:20]
  assign io_ftqInter_toFtq_pdWb_bits_pd_7_valid = wb_valid & wb_instr_valid_7; // @[IFU.scala 763:20]
  assign io_ftqInter_toFtq_pdWb_bits_pd_7_isRVC = wb_valid ? wb_pd_7_isRVC : f3_pd_7_isRVC; // @[IFU.scala 763:20]
  assign io_ftqInter_toFtq_pdWb_bits_pd_7_brType = wb_valid ? wb_pd_7_brType : f3_pd_7_brType; // @[IFU.scala 763:20]
  assign io_ftqInter_toFtq_pdWb_bits_pd_7_isCall = wb_valid ? wb_pd_7_isCall : f3_pd_7_isCall; // @[IFU.scala 763:20]
  assign io_ftqInter_toFtq_pdWb_bits_pd_7_isRet = wb_valid ? wb_pd_7_isRet : f3_pd_7_isRet; // @[IFU.scala 763:20]
  assign io_ftqInter_toFtq_pdWb_bits_ftqIdx_flag = wb_valid ? wb_ftq_req_ftqIdx_flag : f3_ftq_req_ftqIdx_flag; // @[IFU.scala 763:20]
  assign io_ftqInter_toFtq_pdWb_bits_ftqIdx_value = wb_valid ? wb_ftq_req_ftqIdx_value : f3_ftq_req_ftqIdx_value; // @[IFU.scala 763:20]
  assign io_ftqInter_toFtq_pdWb_bits_misOffset_valid = wb_valid ? checkFlushWb_bits_misOffset_valid : f3_req_is_mmio; // @[IFU.scala 763:20]
  assign io_ftqInter_toFtq_pdWb_bits_misOffset_bits = wb_valid ? checkFlushWb_bits_misOffset_bits : 3'h0; // @[IFU.scala 763:20]
  assign io_ftqInter_toFtq_pdWb_bits_cfiOffset_valid = wb_valid & checkFlushWb_bits_cfiOffset_valid; // @[IFU.scala 763:20]
  assign io_ftqInter_toFtq_pdWb_bits_target = wb_valid ? checkFlushWb_bits_target : mmioFlushWb_bits_target; // @[IFU.scala 763:20]
  assign io_ftqInter_toFtq_pdWb_bits_jalTarget = wb_valid ? checkFlushWb_bits_jalTarget : 39'h0; // @[IFU.scala 763:20]
  assign io_ftqInter_toFtq_pdWb_bits_instrRange_0 = wb_valid ? wb_instr_range[0] : 1'h1; // @[IFU.scala 763:20]
  assign io_ftqInter_toFtq_pdWb_bits_instrRange_1 = wb_valid & wb_instr_range[1]; // @[IFU.scala 763:20]
  assign io_ftqInter_toFtq_pdWb_bits_instrRange_2 = wb_valid & wb_instr_range[2]; // @[IFU.scala 763:20]
  assign io_ftqInter_toFtq_pdWb_bits_instrRange_3 = wb_valid & wb_instr_range[3]; // @[IFU.scala 763:20]
  assign io_ftqInter_toFtq_pdWb_bits_instrRange_4 = wb_valid & wb_instr_range[4]; // @[IFU.scala 763:20]
  assign io_ftqInter_toFtq_pdWb_bits_instrRange_5 = wb_valid & wb_instr_range[5]; // @[IFU.scala 763:20]
  assign io_ftqInter_toFtq_pdWb_bits_instrRange_6 = wb_valid & wb_instr_range[6]; // @[IFU.scala 763:20]
  assign io_ftqInter_toFtq_pdWb_bits_instrRange_7 = wb_valid & wb_instr_range[7]; // @[IFU.scala 763:20]
  assign io_icacheStop = ~f3_ready; // @[IFU.scala 250:20]
  assign io_toIbuffer_valid = f3_valid & (_T_21 | f3_mmio_can_go) & ~f3_flush; // @[IFU.scala 619:84]
  assign io_toIbuffer_bits_instrs_0 = f3_req_is_mmio ? _io_toIbuffer_bits_instrs_0_T_64_bits : f3_expd_instr_0; // @[IFU.scala 662:23 620:33 670:34]
  assign io_toIbuffer_bits_instrs_1 = f3_expd_instr_expander_1_io_out_bits; // @[IFU.scala 381:{34,34}]
  assign io_toIbuffer_bits_instrs_2 = f3_expd_instr_expander_2_io_out_bits; // @[IFU.scala 381:{34,34}]
  assign io_toIbuffer_bits_instrs_3 = f3_expd_instr_expander_3_io_out_bits; // @[IFU.scala 381:{34,34}]
  assign io_toIbuffer_bits_instrs_4 = f3_expd_instr_expander_4_io_out_bits; // @[IFU.scala 381:{34,34}]
  assign io_toIbuffer_bits_instrs_5 = f3_expd_instr_expander_5_io_out_bits; // @[IFU.scala 381:{34,34}]
  assign io_toIbuffer_bits_instrs_6 = f3_expd_instr_expander_6_io_out_bits; // @[IFU.scala 381:{34,34}]
  assign io_toIbuffer_bits_instrs_7 = f3_expd_instr_expander_7_io_out_bits; // @[IFU.scala 381:{34,34}]
  assign io_toIbuffer_bits_valid = f3_lastHalf_valid ? _io_toIbuffer_bits_valid_T_2 : _T_59; // @[IFU.scala 633:26 621:33 635:33]
  assign io_toIbuffer_bits_enqEnable = f3_req_is_mmio ? 8'h1 : _GEN_2077; // @[IFU.scala 662:23 683:35]
  assign io_toIbuffer_bits_pd_0_isRVC = f3_req_is_mmio ? currentIsRVC : f3_pd_0_isRVC; // @[IFU.scala 662:23 623:33 674:37]
  assign io_toIbuffer_bits_pd_0_brType = f3_req_is_mmio ? brType : f3_pd_0_brType; // @[IFU.scala 662:23 623:33 675:37]
  assign io_toIbuffer_bits_pd_0_isCall = f3_req_is_mmio ? isCall : f3_pd_0_isCall; // @[IFU.scala 662:23 623:33 676:37]
  assign io_toIbuffer_bits_pd_0_isRet = f3_req_is_mmio ? isRet : f3_pd_0_isRet; // @[IFU.scala 662:23 623:33 677:37]
  assign io_toIbuffer_bits_pd_1_isRVC = f3_pd_1_isRVC; // @[IFU.scala 623:33]
  assign io_toIbuffer_bits_pd_1_brType = f3_pd_1_brType; // @[IFU.scala 623:33]
  assign io_toIbuffer_bits_pd_1_isCall = f3_pd_1_isCall; // @[IFU.scala 623:33]
  assign io_toIbuffer_bits_pd_1_isRet = f3_pd_1_isRet; // @[IFU.scala 623:33]
  assign io_toIbuffer_bits_pd_2_isRVC = f3_pd_2_isRVC; // @[IFU.scala 623:33]
  assign io_toIbuffer_bits_pd_2_brType = f3_pd_2_brType; // @[IFU.scala 623:33]
  assign io_toIbuffer_bits_pd_2_isCall = f3_pd_2_isCall; // @[IFU.scala 623:33]
  assign io_toIbuffer_bits_pd_2_isRet = f3_pd_2_isRet; // @[IFU.scala 623:33]
  assign io_toIbuffer_bits_pd_3_isRVC = f3_pd_3_isRVC; // @[IFU.scala 623:33]
  assign io_toIbuffer_bits_pd_3_brType = f3_pd_3_brType; // @[IFU.scala 623:33]
  assign io_toIbuffer_bits_pd_3_isCall = f3_pd_3_isCall; // @[IFU.scala 623:33]
  assign io_toIbuffer_bits_pd_3_isRet = f3_pd_3_isRet; // @[IFU.scala 623:33]
  assign io_toIbuffer_bits_pd_4_isRVC = f3_pd_4_isRVC; // @[IFU.scala 623:33]
  assign io_toIbuffer_bits_pd_4_brType = f3_pd_4_brType; // @[IFU.scala 623:33]
  assign io_toIbuffer_bits_pd_4_isCall = f3_pd_4_isCall; // @[IFU.scala 623:33]
  assign io_toIbuffer_bits_pd_4_isRet = f3_pd_4_isRet; // @[IFU.scala 623:33]
  assign io_toIbuffer_bits_pd_5_isRVC = f3_pd_5_isRVC; // @[IFU.scala 623:33]
  assign io_toIbuffer_bits_pd_5_brType = f3_pd_5_brType; // @[IFU.scala 623:33]
  assign io_toIbuffer_bits_pd_5_isCall = f3_pd_5_isCall; // @[IFU.scala 623:33]
  assign io_toIbuffer_bits_pd_5_isRet = f3_pd_5_isRet; // @[IFU.scala 623:33]
  assign io_toIbuffer_bits_pd_6_isRVC = f3_pd_6_isRVC; // @[IFU.scala 623:33]
  assign io_toIbuffer_bits_pd_6_brType = f3_pd_6_brType; // @[IFU.scala 623:33]
  assign io_toIbuffer_bits_pd_6_isCall = f3_pd_6_isCall; // @[IFU.scala 623:33]
  assign io_toIbuffer_bits_pd_6_isRet = f3_pd_6_isRet; // @[IFU.scala 623:33]
  assign io_toIbuffer_bits_pd_7_isRVC = f3_pd_7_isRVC; // @[IFU.scala 623:33]
  assign io_toIbuffer_bits_pd_7_brType = f3_pd_7_brType; // @[IFU.scala 623:33]
  assign io_toIbuffer_bits_pd_7_isCall = f3_pd_7_isCall; // @[IFU.scala 623:33]
  assign io_toIbuffer_bits_pd_7_isRet = f3_pd_7_isRet; // @[IFU.scala 623:33]
  assign io_toIbuffer_bits_foldpc_0 = f3_foldpc_0; // @[IFU.scala 627:33]
  assign io_toIbuffer_bits_foldpc_1 = f3_foldpc_1; // @[IFU.scala 627:33]
  assign io_toIbuffer_bits_foldpc_2 = f3_foldpc_2; // @[IFU.scala 627:33]
  assign io_toIbuffer_bits_foldpc_3 = f3_foldpc_3; // @[IFU.scala 627:33]
  assign io_toIbuffer_bits_foldpc_4 = f3_foldpc_4; // @[IFU.scala 627:33]
  assign io_toIbuffer_bits_foldpc_5 = f3_foldpc_5; // @[IFU.scala 627:33]
  assign io_toIbuffer_bits_foldpc_6 = f3_foldpc_6; // @[IFU.scala 627:33]
  assign io_toIbuffer_bits_foldpc_7 = f3_foldpc_7; // @[IFU.scala 627:33]
  assign io_toIbuffer_bits_ftqPtr_flag = f3_ftq_req_ftqIdx_flag; // @[IFU.scala 624:33]
  assign io_toIbuffer_bits_ftqPtr_value = f3_ftq_req_ftqIdx_value; // @[IFU.scala 624:33]
  assign io_toIbuffer_bits_ftqOffset_0_valid = predChecker_io_out_stage1Out_fixedTaken_0 & _T_21; // @[IFU.scala 626:119]
  assign io_toIbuffer_bits_ftqOffset_1_valid = predChecker_io_out_stage1Out_fixedTaken_1 & _T_21; // @[IFU.scala 626:119]
  assign io_toIbuffer_bits_ftqOffset_2_valid = predChecker_io_out_stage1Out_fixedTaken_2 & _T_21; // @[IFU.scala 626:119]
  assign io_toIbuffer_bits_ftqOffset_3_valid = predChecker_io_out_stage1Out_fixedTaken_3 & _T_21; // @[IFU.scala 626:119]
  assign io_toIbuffer_bits_ftqOffset_4_valid = predChecker_io_out_stage1Out_fixedTaken_4 & _T_21; // @[IFU.scala 626:119]
  assign io_toIbuffer_bits_ftqOffset_5_valid = predChecker_io_out_stage1Out_fixedTaken_5 & _T_21; // @[IFU.scala 626:119]
  assign io_toIbuffer_bits_ftqOffset_6_valid = predChecker_io_out_stage1Out_fixedTaken_6 & _T_21; // @[IFU.scala 626:119]
  assign io_toIbuffer_bits_ftqOffset_7_valid = predChecker_io_out_stage1Out_fixedTaken_7 & _T_21; // @[IFU.scala 626:119]
  assign io_toIbuffer_bits_ipf_0 = f3_req_is_mmio ? mmio_resend_pf : f3_pf_vec_0 | f3_crossPageFault_0; // @[IFU.scala 662:23 680:30 628:33]
  assign io_toIbuffer_bits_ipf_1 = f3_pf_vec_1 | f3_crossPageFault_1; // @[IFU.scala 628:106]
  assign io_toIbuffer_bits_ipf_2 = f3_pf_vec_2 | f3_crossPageFault_2; // @[IFU.scala 628:106]
  assign io_toIbuffer_bits_ipf_3 = f3_pf_vec_3 | f3_crossPageFault_3; // @[IFU.scala 628:106]
  assign io_toIbuffer_bits_ipf_4 = f3_pf_vec_4 | f3_crossPageFault_4; // @[IFU.scala 628:106]
  assign io_toIbuffer_bits_ipf_5 = f3_pf_vec_5 | f3_crossPageFault_5; // @[IFU.scala 628:106]
  assign io_toIbuffer_bits_ipf_6 = f3_pf_vec_6 | f3_crossPageFault_6; // @[IFU.scala 628:106]
  assign io_toIbuffer_bits_ipf_7 = f3_pf_vec_7 | f3_crossPageFault_7; // @[IFU.scala 628:106]
  assign io_toIbuffer_bits_acf_0 = f3_req_is_mmio ? mmio_resend_af : f3_af_vec_0; // @[IFU.scala 662:23 679:30 629:33]
  assign io_toIbuffer_bits_acf_1 = f3_af_vec_1; // @[IFU.scala 629:33]
  assign io_toIbuffer_bits_acf_2 = f3_af_vec_2; // @[IFU.scala 629:33]
  assign io_toIbuffer_bits_acf_3 = f3_af_vec_3; // @[IFU.scala 629:33]
  assign io_toIbuffer_bits_acf_4 = f3_af_vec_4; // @[IFU.scala 629:33]
  assign io_toIbuffer_bits_acf_5 = f3_af_vec_5; // @[IFU.scala 629:33]
  assign io_toIbuffer_bits_acf_6 = f3_af_vec_6; // @[IFU.scala 629:33]
  assign io_toIbuffer_bits_acf_7 = f3_af_vec_7; // @[IFU.scala 629:33]
  assign io_toIbuffer_bits_crossPageIPFFix_0 = f3_req_is_mmio ? mmio_resend_pf : f3_crossPageFault_0; // @[IFU.scala 662:23 630:37 681:42]
  assign io_toIbuffer_bits_crossPageIPFFix_1 = f3_crossPageFault_1; // @[IFU.scala 630:37]
  assign io_toIbuffer_bits_crossPageIPFFix_2 = f3_crossPageFault_2; // @[IFU.scala 630:37]
  assign io_toIbuffer_bits_crossPageIPFFix_3 = f3_crossPageFault_3; // @[IFU.scala 630:37]
  assign io_toIbuffer_bits_crossPageIPFFix_4 = f3_crossPageFault_4; // @[IFU.scala 630:37]
  assign io_toIbuffer_bits_crossPageIPFFix_5 = f3_crossPageFault_5; // @[IFU.scala 630:37]
  assign io_toIbuffer_bits_crossPageIPFFix_6 = f3_crossPageFault_6; // @[IFU.scala 630:37]
  assign io_toIbuffer_bits_crossPageIPFFix_7 = f3_crossPageFault_7; // @[IFU.scala 630:37]
  assign io_toIbuffer_bits_triggered_0_frontendHit_0 = frontendTrigger_io_triggered_0_frontendHit_0; // @[IFU.scala 631:33]
  assign io_toIbuffer_bits_triggered_0_frontendHit_1 = frontendTrigger_io_triggered_0_frontendHit_1; // @[IFU.scala 631:33]
  assign io_toIbuffer_bits_triggered_0_frontendHit_2 = frontendTrigger_io_triggered_0_frontendHit_2; // @[IFU.scala 631:33]
  assign io_toIbuffer_bits_triggered_0_frontendHit_3 = frontendTrigger_io_triggered_0_frontendHit_3; // @[IFU.scala 631:33]
  assign io_toIbuffer_bits_triggered_0_backendEn_0 = frontendTrigger_io_triggered_0_backendEn_0; // @[IFU.scala 631:33]
  assign io_toIbuffer_bits_triggered_0_backendEn_1 = frontendTrigger_io_triggered_0_backendEn_1; // @[IFU.scala 631:33]
  assign io_toIbuffer_bits_triggered_1_frontendHit_0 = frontendTrigger_io_triggered_1_frontendHit_0; // @[IFU.scala 631:33]
  assign io_toIbuffer_bits_triggered_1_frontendHit_1 = frontendTrigger_io_triggered_1_frontendHit_1; // @[IFU.scala 631:33]
  assign io_toIbuffer_bits_triggered_1_frontendHit_2 = frontendTrigger_io_triggered_1_frontendHit_2; // @[IFU.scala 631:33]
  assign io_toIbuffer_bits_triggered_1_frontendHit_3 = frontendTrigger_io_triggered_1_frontendHit_3; // @[IFU.scala 631:33]
  assign io_toIbuffer_bits_triggered_1_backendEn_0 = frontendTrigger_io_triggered_1_backendEn_0; // @[IFU.scala 631:33]
  assign io_toIbuffer_bits_triggered_1_backendEn_1 = frontendTrigger_io_triggered_1_backendEn_1; // @[IFU.scala 631:33]
  assign io_toIbuffer_bits_triggered_2_frontendHit_0 = frontendTrigger_io_triggered_2_frontendHit_0; // @[IFU.scala 631:33]
  assign io_toIbuffer_bits_triggered_2_frontendHit_1 = frontendTrigger_io_triggered_2_frontendHit_1; // @[IFU.scala 631:33]
  assign io_toIbuffer_bits_triggered_2_frontendHit_2 = frontendTrigger_io_triggered_2_frontendHit_2; // @[IFU.scala 631:33]
  assign io_toIbuffer_bits_triggered_2_frontendHit_3 = frontendTrigger_io_triggered_2_frontendHit_3; // @[IFU.scala 631:33]
  assign io_toIbuffer_bits_triggered_2_backendEn_0 = frontendTrigger_io_triggered_2_backendEn_0; // @[IFU.scala 631:33]
  assign io_toIbuffer_bits_triggered_2_backendEn_1 = frontendTrigger_io_triggered_2_backendEn_1; // @[IFU.scala 631:33]
  assign io_toIbuffer_bits_triggered_3_frontendHit_0 = frontendTrigger_io_triggered_3_frontendHit_0; // @[IFU.scala 631:33]
  assign io_toIbuffer_bits_triggered_3_frontendHit_1 = frontendTrigger_io_triggered_3_frontendHit_1; // @[IFU.scala 631:33]
  assign io_toIbuffer_bits_triggered_3_frontendHit_2 = frontendTrigger_io_triggered_3_frontendHit_2; // @[IFU.scala 631:33]
  assign io_toIbuffer_bits_triggered_3_frontendHit_3 = frontendTrigger_io_triggered_3_frontendHit_3; // @[IFU.scala 631:33]
  assign io_toIbuffer_bits_triggered_3_backendEn_0 = frontendTrigger_io_triggered_3_backendEn_0; // @[IFU.scala 631:33]
  assign io_toIbuffer_bits_triggered_3_backendEn_1 = frontendTrigger_io_triggered_3_backendEn_1; // @[IFU.scala 631:33]
  assign io_toIbuffer_bits_triggered_4_frontendHit_0 = frontendTrigger_io_triggered_4_frontendHit_0; // @[IFU.scala 631:33]
  assign io_toIbuffer_bits_triggered_4_frontendHit_1 = frontendTrigger_io_triggered_4_frontendHit_1; // @[IFU.scala 631:33]
  assign io_toIbuffer_bits_triggered_4_frontendHit_2 = frontendTrigger_io_triggered_4_frontendHit_2; // @[IFU.scala 631:33]
  assign io_toIbuffer_bits_triggered_4_frontendHit_3 = frontendTrigger_io_triggered_4_frontendHit_3; // @[IFU.scala 631:33]
  assign io_toIbuffer_bits_triggered_4_backendEn_0 = frontendTrigger_io_triggered_4_backendEn_0; // @[IFU.scala 631:33]
  assign io_toIbuffer_bits_triggered_4_backendEn_1 = frontendTrigger_io_triggered_4_backendEn_1; // @[IFU.scala 631:33]
  assign io_toIbuffer_bits_triggered_5_frontendHit_0 = frontendTrigger_io_triggered_5_frontendHit_0; // @[IFU.scala 631:33]
  assign io_toIbuffer_bits_triggered_5_frontendHit_1 = frontendTrigger_io_triggered_5_frontendHit_1; // @[IFU.scala 631:33]
  assign io_toIbuffer_bits_triggered_5_frontendHit_2 = frontendTrigger_io_triggered_5_frontendHit_2; // @[IFU.scala 631:33]
  assign io_toIbuffer_bits_triggered_5_frontendHit_3 = frontendTrigger_io_triggered_5_frontendHit_3; // @[IFU.scala 631:33]
  assign io_toIbuffer_bits_triggered_5_backendEn_0 = frontendTrigger_io_triggered_5_backendEn_0; // @[IFU.scala 631:33]
  assign io_toIbuffer_bits_triggered_5_backendEn_1 = frontendTrigger_io_triggered_5_backendEn_1; // @[IFU.scala 631:33]
  assign io_toIbuffer_bits_triggered_6_frontendHit_0 = frontendTrigger_io_triggered_6_frontendHit_0; // @[IFU.scala 631:33]
  assign io_toIbuffer_bits_triggered_6_frontendHit_1 = frontendTrigger_io_triggered_6_frontendHit_1; // @[IFU.scala 631:33]
  assign io_toIbuffer_bits_triggered_6_frontendHit_2 = frontendTrigger_io_triggered_6_frontendHit_2; // @[IFU.scala 631:33]
  assign io_toIbuffer_bits_triggered_6_frontendHit_3 = frontendTrigger_io_triggered_6_frontendHit_3; // @[IFU.scala 631:33]
  assign io_toIbuffer_bits_triggered_6_backendEn_0 = frontendTrigger_io_triggered_6_backendEn_0; // @[IFU.scala 631:33]
  assign io_toIbuffer_bits_triggered_6_backendEn_1 = frontendTrigger_io_triggered_6_backendEn_1; // @[IFU.scala 631:33]
  assign io_toIbuffer_bits_triggered_7_frontendHit_0 = frontendTrigger_io_triggered_7_frontendHit_0; // @[IFU.scala 631:33]
  assign io_toIbuffer_bits_triggered_7_frontendHit_1 = frontendTrigger_io_triggered_7_frontendHit_1; // @[IFU.scala 631:33]
  assign io_toIbuffer_bits_triggered_7_frontendHit_2 = frontendTrigger_io_triggered_7_frontendHit_2; // @[IFU.scala 631:33]
  assign io_toIbuffer_bits_triggered_7_frontendHit_3 = frontendTrigger_io_triggered_7_frontendHit_3; // @[IFU.scala 631:33]
  assign io_toIbuffer_bits_triggered_7_backendEn_0 = frontendTrigger_io_triggered_7_backendEn_0; // @[IFU.scala 631:33]
  assign io_toIbuffer_bits_triggered_7_backendEn_1 = frontendTrigger_io_triggered_7_backendEn_1; // @[IFU.scala 631:33]
  assign io_uncacheInter_fromUncache_ready = 1'h1; // @[IFU.scala 544:23]
  assign io_uncacheInter_toUncache_valid = (mmio_state == 4'h2 | mmio_state == 4'h7) & f3_req_is_mmio; // @[IFU.scala 542:88]
  assign io_uncacheInter_toUncache_bits_addr = _io_uncacheInter_toUncache_valid_T_1 ? mmio_resend_addr : f3_pAddrs_0; // @[IFU.scala 543:29]
  assign io_iTLBInter_req_valid = mmio_state == 4'h4 & f3_req_is_mmio; // @[IFU.scala 546:64]
  assign io_iTLBInter_req_bits_vaddr = f3_resend_vaddr; // @[IFU.scala 548:34]
  assign io_pmp_req_bits_addr = mmio_resend_addr; // @[IFU.scala 559:25]
  assign io_mmioCommitRead_mmioFtqPtr_flag = io_mmioCommitRead_mmioFtqPtr_REG_flag; // @[IFU.scala 415:32]
  assign io_mmioCommitRead_mmioFtqPtr_value = io_mmioCommitRead_mmioFtqPtr_REG_value; // @[IFU.scala 415:32]
  assign io_perf_0_value = {{5'd0}, io_perf_0_value_REG_1}; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_1_value = {{5'd0}, io_perf_1_value_REG_1}; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_2_value = {{5'd0}, io_perf_2_value_REG_1}; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_3_value = {{5'd0}, io_perf_3_value_REG_1}; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_4_value = {{5'd0}, io_perf_4_value_REG_1}; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_5_value = {{5'd0}, io_perf_5_value_REG_1}; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_6_value = {{5'd0}, io_perf_6_value_REG_1}; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_7_value = {{5'd0}, io_perf_7_value_REG_1}; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_8_value = {{5'd0}, io_perf_8_value_REG_1}; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_9_value = {{5'd0}, io_perf_9_value_REG_1}; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_10_value = {{5'd0}, io_perf_10_value_REG_1}; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_11_value = {{5'd0}, io_perf_11_value_REG_1}; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_12_value = {{5'd0}, io_perf_12_value_REG_1}; // @[PerfCounterUtils.scala 188:17]
  assign preDecoders_0_io_in_data_0 = 6'h2f == f2_cut_ptr_0 ? f2_cut_data_dataVec__47 : _GEN_101; // @[IFU.scala 302:{19,19}]
  assign preDecoders_0_io_in_data_1 = 6'h2f == f2_cut_ptr_1 ? f2_cut_data_dataVec__47 : _GEN_149; // @[IFU.scala 302:{19,19}]
  assign preDecoders_0_io_in_data_2 = 6'h2f == f2_cut_ptr_2 ? f2_cut_data_dataVec__47 : _GEN_197; // @[IFU.scala 302:{19,19}]
  assign preDecoders_0_io_in_data_3 = 6'h2f == f2_cut_ptr_3 ? f2_cut_data_dataVec__47 : _GEN_245; // @[IFU.scala 302:{19,19}]
  assign preDecoders_0_io_in_data_4 = 6'h2f == f2_cut_ptr_4 ? f2_cut_data_dataVec__47 : _GEN_293; // @[IFU.scala 302:{19,19}]
  assign preDecoders_0_io_in_data_5 = 6'h2f == f2_cut_ptr_5 ? f2_cut_data_dataVec__47 : _GEN_341; // @[IFU.scala 302:{19,19}]
  assign preDecoders_0_io_in_data_6 = 6'h2f == f2_cut_ptr_6 ? f2_cut_data_dataVec__47 : _GEN_389; // @[IFU.scala 302:{19,19}]
  assign preDecoders_0_io_in_data_7 = 6'h2f == f2_cut_ptr_7 ? f2_cut_data_dataVec__47 : _GEN_437; // @[IFU.scala 302:{19,19}]
  assign preDecoders_0_io_in_data_8 = 6'h2f == f2_cut_ptr_8 ? f2_cut_data_dataVec__47 : _GEN_485; // @[IFU.scala 302:{19,19}]
  assign preDecoders_1_io_in_data_0 = 6'h2f == f2_cut_ptr_0 ? f2_cut_data_dataVec_1_47 : _GEN_533; // @[IFU.scala 302:{19,19}]
  assign preDecoders_1_io_in_data_1 = 6'h2f == f2_cut_ptr_1 ? f2_cut_data_dataVec_1_47 : _GEN_581; // @[IFU.scala 302:{19,19}]
  assign preDecoders_1_io_in_data_2 = 6'h2f == f2_cut_ptr_2 ? f2_cut_data_dataVec_1_47 : _GEN_629; // @[IFU.scala 302:{19,19}]
  assign preDecoders_1_io_in_data_3 = 6'h2f == f2_cut_ptr_3 ? f2_cut_data_dataVec_1_47 : _GEN_677; // @[IFU.scala 302:{19,19}]
  assign preDecoders_1_io_in_data_4 = 6'h2f == f2_cut_ptr_4 ? f2_cut_data_dataVec_1_47 : _GEN_725; // @[IFU.scala 302:{19,19}]
  assign preDecoders_1_io_in_data_5 = 6'h2f == f2_cut_ptr_5 ? f2_cut_data_dataVec_1_47 : _GEN_773; // @[IFU.scala 302:{19,19}]
  assign preDecoders_1_io_in_data_6 = 6'h2f == f2_cut_ptr_6 ? f2_cut_data_dataVec_1_47 : _GEN_821; // @[IFU.scala 302:{19,19}]
  assign preDecoders_1_io_in_data_7 = 6'h2f == f2_cut_ptr_7 ? f2_cut_data_dataVec_1_47 : _GEN_869; // @[IFU.scala 302:{19,19}]
  assign preDecoders_1_io_in_data_8 = 6'h2f == f2_cut_ptr_8 ? f2_cut_data_dataVec_1_47 : _GEN_917; // @[IFU.scala 302:{19,19}]
  assign preDecoders_2_io_in_data_0 = 6'h2f == f2_cut_ptr_0 ? f2_cut_data_dataVec_2_47 : _GEN_965; // @[IFU.scala 302:{19,19}]
  assign preDecoders_2_io_in_data_1 = 6'h2f == f2_cut_ptr_1 ? f2_cut_data_dataVec_2_47 : _GEN_1013; // @[IFU.scala 302:{19,19}]
  assign preDecoders_2_io_in_data_2 = 6'h2f == f2_cut_ptr_2 ? f2_cut_data_dataVec_2_47 : _GEN_1061; // @[IFU.scala 302:{19,19}]
  assign preDecoders_2_io_in_data_3 = 6'h2f == f2_cut_ptr_3 ? f2_cut_data_dataVec_2_47 : _GEN_1109; // @[IFU.scala 302:{19,19}]
  assign preDecoders_2_io_in_data_4 = 6'h2f == f2_cut_ptr_4 ? f2_cut_data_dataVec_2_47 : _GEN_1157; // @[IFU.scala 302:{19,19}]
  assign preDecoders_2_io_in_data_5 = 6'h2f == f2_cut_ptr_5 ? f2_cut_data_dataVec_2_47 : _GEN_1205; // @[IFU.scala 302:{19,19}]
  assign preDecoders_2_io_in_data_6 = 6'h2f == f2_cut_ptr_6 ? f2_cut_data_dataVec_2_47 : _GEN_1253; // @[IFU.scala 302:{19,19}]
  assign preDecoders_2_io_in_data_7 = 6'h2f == f2_cut_ptr_7 ? f2_cut_data_dataVec_2_47 : _GEN_1301; // @[IFU.scala 302:{19,19}]
  assign preDecoders_2_io_in_data_8 = 6'h2f == f2_cut_ptr_8 ? f2_cut_data_dataVec_2_47 : _GEN_1349; // @[IFU.scala 302:{19,19}]
  assign preDecoders_3_io_in_data_0 = 6'h2f == f2_cut_ptr_0 ? f2_cut_data_dataVec_3_47 : _GEN_1397; // @[IFU.scala 302:{19,19}]
  assign preDecoders_3_io_in_data_1 = 6'h2f == f2_cut_ptr_1 ? f2_cut_data_dataVec_3_47 : _GEN_1445; // @[IFU.scala 302:{19,19}]
  assign preDecoders_3_io_in_data_2 = 6'h2f == f2_cut_ptr_2 ? f2_cut_data_dataVec_3_47 : _GEN_1493; // @[IFU.scala 302:{19,19}]
  assign preDecoders_3_io_in_data_3 = 6'h2f == f2_cut_ptr_3 ? f2_cut_data_dataVec_3_47 : _GEN_1541; // @[IFU.scala 302:{19,19}]
  assign preDecoders_3_io_in_data_4 = 6'h2f == f2_cut_ptr_4 ? f2_cut_data_dataVec_3_47 : _GEN_1589; // @[IFU.scala 302:{19,19}]
  assign preDecoders_3_io_in_data_5 = 6'h2f == f2_cut_ptr_5 ? f2_cut_data_dataVec_3_47 : _GEN_1637; // @[IFU.scala 302:{19,19}]
  assign preDecoders_3_io_in_data_6 = 6'h2f == f2_cut_ptr_6 ? f2_cut_data_dataVec_3_47 : _GEN_1685; // @[IFU.scala 302:{19,19}]
  assign preDecoders_3_io_in_data_7 = 6'h2f == f2_cut_ptr_7 ? f2_cut_data_dataVec_3_47 : _GEN_1733; // @[IFU.scala 302:{19,19}]
  assign preDecoders_3_io_in_data_8 = 6'h2f == f2_cut_ptr_8 ? f2_cut_data_dataVec_3_47 : _GEN_1781; // @[IFU.scala 302:{19,19}]
  assign predChecker_clock = clock;
  assign predChecker_io_in_ftqOffset_valid = f3_ftq_req_ftqOffset_valid; // @[IFU.scala 570:25]
  assign predChecker_io_in_ftqOffset_bits = f3_ftq_req_ftqOffset_bits; // @[IFU.scala 570:25]
  assign predChecker_io_in_jumpOffset_0 = f3_jump_offset_0; // @[IFU.scala 571:25]
  assign predChecker_io_in_jumpOffset_1 = f3_jump_offset_1; // @[IFU.scala 571:25]
  assign predChecker_io_in_jumpOffset_2 = f3_jump_offset_2; // @[IFU.scala 571:25]
  assign predChecker_io_in_jumpOffset_3 = f3_jump_offset_3; // @[IFU.scala 571:25]
  assign predChecker_io_in_jumpOffset_4 = f3_jump_offset_4; // @[IFU.scala 571:25]
  assign predChecker_io_in_jumpOffset_5 = f3_jump_offset_5; // @[IFU.scala 571:25]
  assign predChecker_io_in_jumpOffset_6 = f3_jump_offset_6; // @[IFU.scala 571:25]
  assign predChecker_io_in_jumpOffset_7 = f3_jump_offset_7; // @[IFU.scala 571:25]
  assign predChecker_io_in_target = f3_ftq_req_nextStartAddr; // @[IFU.scala 572:25]
  assign predChecker_io_in_instrRange_0 = f3_instr_range[0]; // @[IFU.scala 573:51]
  assign predChecker_io_in_instrRange_1 = f3_instr_range[1]; // @[IFU.scala 573:51]
  assign predChecker_io_in_instrRange_2 = f3_instr_range[2]; // @[IFU.scala 573:51]
  assign predChecker_io_in_instrRange_3 = f3_instr_range[3]; // @[IFU.scala 573:51]
  assign predChecker_io_in_instrRange_4 = f3_instr_range[4]; // @[IFU.scala 573:51]
  assign predChecker_io_in_instrRange_5 = f3_instr_range[5]; // @[IFU.scala 573:51]
  assign predChecker_io_in_instrRange_6 = f3_instr_range[6]; // @[IFU.scala 573:51]
  assign predChecker_io_in_instrRange_7 = f3_instr_range[7]; // @[IFU.scala 573:51]
  assign predChecker_io_in_instrValid_0 = _T_59[0]; // @[IFU.scala 574:51]
  assign predChecker_io_in_instrValid_1 = _T_59[1]; // @[IFU.scala 574:51]
  assign predChecker_io_in_instrValid_2 = _T_59[2]; // @[IFU.scala 574:51]
  assign predChecker_io_in_instrValid_3 = _T_59[3]; // @[IFU.scala 574:51]
  assign predChecker_io_in_instrValid_4 = _T_59[4]; // @[IFU.scala 574:51]
  assign predChecker_io_in_instrValid_5 = _T_59[5]; // @[IFU.scala 574:51]
  assign predChecker_io_in_instrValid_6 = _T_59[6]; // @[IFU.scala 574:51]
  assign predChecker_io_in_instrValid_7 = _T_59[7]; // @[IFU.scala 574:51]
  assign predChecker_io_in_pds_0_isRVC = f3_pd_0_isRVC; // @[IFU.scala 575:25]
  assign predChecker_io_in_pds_0_brType = f3_pd_0_brType; // @[IFU.scala 575:25]
  assign predChecker_io_in_pds_0_isRet = f3_pd_0_isRet; // @[IFU.scala 575:25]
  assign predChecker_io_in_pds_1_isRVC = f3_pd_1_isRVC; // @[IFU.scala 575:25]
  assign predChecker_io_in_pds_1_brType = f3_pd_1_brType; // @[IFU.scala 575:25]
  assign predChecker_io_in_pds_1_isRet = f3_pd_1_isRet; // @[IFU.scala 575:25]
  assign predChecker_io_in_pds_2_isRVC = f3_pd_2_isRVC; // @[IFU.scala 575:25]
  assign predChecker_io_in_pds_2_brType = f3_pd_2_brType; // @[IFU.scala 575:25]
  assign predChecker_io_in_pds_2_isRet = f3_pd_2_isRet; // @[IFU.scala 575:25]
  assign predChecker_io_in_pds_3_isRVC = f3_pd_3_isRVC; // @[IFU.scala 575:25]
  assign predChecker_io_in_pds_3_brType = f3_pd_3_brType; // @[IFU.scala 575:25]
  assign predChecker_io_in_pds_3_isRet = f3_pd_3_isRet; // @[IFU.scala 575:25]
  assign predChecker_io_in_pds_4_isRVC = f3_pd_4_isRVC; // @[IFU.scala 575:25]
  assign predChecker_io_in_pds_4_brType = f3_pd_4_brType; // @[IFU.scala 575:25]
  assign predChecker_io_in_pds_4_isRet = f3_pd_4_isRet; // @[IFU.scala 575:25]
  assign predChecker_io_in_pds_5_isRVC = f3_pd_5_isRVC; // @[IFU.scala 575:25]
  assign predChecker_io_in_pds_5_brType = f3_pd_5_brType; // @[IFU.scala 575:25]
  assign predChecker_io_in_pds_5_isRet = f3_pd_5_isRet; // @[IFU.scala 575:25]
  assign predChecker_io_in_pds_6_isRVC = f3_pd_6_isRVC; // @[IFU.scala 575:25]
  assign predChecker_io_in_pds_6_brType = f3_pd_6_brType; // @[IFU.scala 575:25]
  assign predChecker_io_in_pds_6_isRet = f3_pd_6_isRet; // @[IFU.scala 575:25]
  assign predChecker_io_in_pds_7_isRVC = f3_pd_7_isRVC; // @[IFU.scala 575:25]
  assign predChecker_io_in_pds_7_brType = f3_pd_7_brType; // @[IFU.scala 575:25]
  assign predChecker_io_in_pds_7_isRet = f3_pd_7_isRet; // @[IFU.scala 575:25]
  assign predChecker_io_in_pc_0 = f3_pc_0; // @[IFU.scala 576:25]
  assign predChecker_io_in_pc_1 = f3_pc_1; // @[IFU.scala 576:25]
  assign predChecker_io_in_pc_2 = f3_pc_2; // @[IFU.scala 576:25]
  assign predChecker_io_in_pc_3 = f3_pc_3; // @[IFU.scala 576:25]
  assign predChecker_io_in_pc_4 = f3_pc_4; // @[IFU.scala 576:25]
  assign predChecker_io_in_pc_5 = f3_pc_5; // @[IFU.scala 576:25]
  assign predChecker_io_in_pc_6 = f3_pc_6; // @[IFU.scala 576:25]
  assign predChecker_io_in_pc_7 = f3_pc_7; // @[IFU.scala 576:25]
  assign frontendTrigger_clock = clock;
  assign frontendTrigger_reset = reset;
  assign frontendTrigger_io_frontendTrigger_t_valid = io_frontendTrigger_t_valid; // @[IFU.scala 612:39]
  assign frontendTrigger_io_frontendTrigger_t_bits_addr = io_frontendTrigger_t_bits_addr; // @[IFU.scala 612:39]
  assign frontendTrigger_io_frontendTrigger_t_bits_tdata_matchType = io_frontendTrigger_t_bits_tdata_matchType; // @[IFU.scala 612:39]
  assign frontendTrigger_io_frontendTrigger_t_bits_tdata_select = io_frontendTrigger_t_bits_tdata_select; // @[IFU.scala 612:39]
  assign frontendTrigger_io_frontendTrigger_t_bits_tdata_timing = io_frontendTrigger_t_bits_tdata_timing; // @[IFU.scala 612:39]
  assign frontendTrigger_io_frontendTrigger_t_bits_tdata_chain = io_frontendTrigger_t_bits_tdata_chain; // @[IFU.scala 612:39]
  assign frontendTrigger_io_frontendTrigger_t_bits_tdata_tdata2 = io_frontendTrigger_t_bits_tdata_tdata2; // @[IFU.scala 612:39]
  assign frontendTrigger_io_csrTriggerEnable_0 = io_csrTriggerEnable_0; // @[IFU.scala 613:39]
  assign frontendTrigger_io_csrTriggerEnable_1 = io_csrTriggerEnable_1; // @[IFU.scala 613:39]
  assign frontendTrigger_io_csrTriggerEnable_2 = io_csrTriggerEnable_2; // @[IFU.scala 613:39]
  assign frontendTrigger_io_csrTriggerEnable_3 = io_csrTriggerEnable_3; // @[IFU.scala 613:39]
  assign frontendTrigger_io_pds_0_isRVC = f3_pd_0_isRVC; // @[IFU.scala 608:27]
  assign frontendTrigger_io_pds_1_isRVC = f3_pd_1_isRVC; // @[IFU.scala 608:27]
  assign frontendTrigger_io_pds_2_isRVC = f3_pd_2_isRVC; // @[IFU.scala 608:27]
  assign frontendTrigger_io_pds_3_isRVC = f3_pd_3_isRVC; // @[IFU.scala 608:27]
  assign frontendTrigger_io_pds_4_isRVC = f3_pd_4_isRVC; // @[IFU.scala 608:27]
  assign frontendTrigger_io_pds_5_isRVC = f3_pd_5_isRVC; // @[IFU.scala 608:27]
  assign frontendTrigger_io_pds_6_isRVC = f3_pd_6_isRVC; // @[IFU.scala 608:27]
  assign frontendTrigger_io_pds_7_isRVC = f3_pd_7_isRVC; // @[IFU.scala 608:27]
  assign frontendTrigger_io_pc_0 = f3_pc_0; // @[IFU.scala 609:27]
  assign frontendTrigger_io_pc_1 = f3_pc_1; // @[IFU.scala 609:27]
  assign frontendTrigger_io_pc_2 = f3_pc_2; // @[IFU.scala 609:27]
  assign frontendTrigger_io_pc_3 = f3_pc_3; // @[IFU.scala 609:27]
  assign frontendTrigger_io_pc_4 = f3_pc_4; // @[IFU.scala 609:27]
  assign frontendTrigger_io_pc_5 = f3_pc_5; // @[IFU.scala 609:27]
  assign frontendTrigger_io_pc_6 = f3_pc_6; // @[IFU.scala 609:27]
  assign frontendTrigger_io_pc_7 = f3_pc_7; // @[IFU.scala 609:27]
  assign frontendTrigger_io_data_0 = f3_cut_data_0; // @[IFU.scala 610:29]
  assign frontendTrigger_io_data_1 = f3_cut_data_1; // @[IFU.scala 610:29]
  assign frontendTrigger_io_data_2 = f3_cut_data_2; // @[IFU.scala 610:29]
  assign frontendTrigger_io_data_3 = f3_cut_data_3; // @[IFU.scala 610:29]
  assign frontendTrigger_io_data_4 = f3_cut_data_4; // @[IFU.scala 610:29]
  assign frontendTrigger_io_data_5 = f3_cut_data_5; // @[IFU.scala 610:29]
  assign frontendTrigger_io_data_6 = f3_cut_data_6; // @[IFU.scala 610:29]
  assign frontendTrigger_io_data_7 = f3_cut_data_7; // @[IFU.scala 610:29]
  assign frontendTrigger_io_data_8 = f3_cut_data_8; // @[IFU.scala 610:29]
  assign f3_expd_instr_expander_io_in = f3_instr_0; // @[IFU.scala 383:20]
  assign f3_expd_instr_expander_1_io_in = f3_instr_1; // @[IFU.scala 383:20]
  assign f3_expd_instr_expander_2_io_in = f3_instr_2; // @[IFU.scala 383:20]
  assign f3_expd_instr_expander_3_io_in = f3_instr_3; // @[IFU.scala 383:20]
  assign f3_expd_instr_expander_4_io_in = f3_instr_4; // @[IFU.scala 383:20]
  assign f3_expd_instr_expander_5_io_in = f3_instr_5; // @[IFU.scala 383:20]
  assign f3_expd_instr_expander_6_io_in = f3_instr_6; // @[IFU.scala 383:20]
  assign f3_expd_instr_expander_7_io_in = f3_instr_7; // @[IFU.scala 383:20]
  assign writer_clock = clock; // @[ChiselDB.scala 135:21]
  assign writer_reset = reset; // @[ChiselDB.scala 136:21]
  assign writer_en = io_toIbuffer_ready & io_toIbuffer_valid; // @[Decoupled.scala 50:35]
  assign writer_stamp = cnt; // @[ChiselDB.scala 138:21]
  assign writer_data_start_addr = f3_ftq_req_startAddr; // @[IFU.scala 833:34 834:35]
  assign writer_data_instr_count = {{28'd0}, _fetchIBufferDumpData_instr_count_T_20}; // @[IFU.scala 833:34 835:36]
  assign writer_data_exception = _T_137 | _T_133 | _T_135; // @[IFU.scala 836:140]
  assign writer_data_is_cache_hit = f3_perf_info_hit; // @[IFU.scala 833:34 837:37]
  assign writer_1_clock = clock; // @[ChiselDB.scala 135:21]
  assign writer_1_reset = reset; // @[ChiselDB.scala 136:21]
  assign writer_1_en = wb_valid; // @[IFU.scala 748:26 749:39]
  assign writer_1_stamp = cnt_1; // @[ChiselDB.scala 138:21]
  assign writer_1_data_start_addr = wb_ftq_req_startAddr; // @[IFU.scala 839:32 840:33]
  assign writer_1_data_is_miss_pred = _checkFlushWb_bits_misOffset_valid_T_6 | wb_false_lastHalf; // @[IFU.scala 755:91]
  assign writer_1_data_miss_pred_offset = {{29'd0}, checkFlushWb_bits_misOffset_bits}; // @[IFU.scala 839:32 842:39]
  assign writer_1_data_checkJalFault = wb_valid & (_checkJalFault_T | _checkJalFault_T_1 | _checkJalFault_T_2 |
    _checkJalFault_T_3 | _checkJalFault_T_4 | _checkJalFault_T_5 | _checkJalFault_T_6 | _checkJalFault_T_7); // @[IFU.scala 769:33]
  assign writer_1_data_checkRetFault = wb_valid & (_checkRetFault_T | _checkRetFault_T_1 | _checkRetFault_T_2 |
    _checkRetFault_T_3 | _checkRetFault_T_4 | _checkRetFault_T_5 | _checkRetFault_T_6 | _checkRetFault_T_7); // @[IFU.scala 770:33]
  assign writer_1_data_checkTargetFault = wb_valid & (_checkTargetFault_T | _checkTargetFault_T_1 |
    _checkTargetFault_T_2 | _checkTargetFault_T_3 | _checkTargetFault_T_4 | _checkTargetFault_T_5 |
    _checkTargetFault_T_6 | _checkTargetFault_T_7); // @[IFU.scala 771:36]
  assign writer_1_data_checkNotCFIFault = wb_valid & (_checkNotCFIFault_T | _checkNotCFIFault_T_1 |
    _checkNotCFIFault_T_2 | _checkNotCFIFault_T_3 | _checkNotCFIFault_T_4 | _checkNotCFIFault_T_5 |
    _checkNotCFIFault_T_6 | _checkNotCFIFault_T_7); // @[IFU.scala 772:36]
  assign writer_1_data_checkInvalidTaken = wb_valid & (_checkInvalidTaken_T | _checkInvalidTaken_T_1 |
    _checkInvalidTaken_T_2 | _checkInvalidTaken_T_3 | _checkInvalidTaken_T_4 | _checkInvalidTaken_T_5 |
    _checkInvalidTaken_T_6 | _checkInvalidTaken_T_7); // @[IFU.scala 773:37]
  always @(posedge clock) begin
    wb_ftq_req_ftqIdx_flag <= f3_ftq_req_ftqIdx_flag; // @[IFU.scala 707:34]
    wb_ftq_req_ftqIdx_value <= f3_ftq_req_ftqIdx_value; // @[IFU.scala 707:34]
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_ftq_req_ftqIdx_flag <= f2_ftq_req_ftqIdx_flag; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_ftq_req_ftqIdx_value <= f2_ftq_req_ftqIdx_value; // @[Reg.scala 17:22]
    end
    wb_valid <= wb_valid_REG & _T_21 & _io_toIbuffer_valid_T_3; // @[IFU.scala 706:84]
    wb_false_lastHalf_REG <= ~_GEN_2047 & _GEN_2055 & _GEN_2063 & ~_GEN_2071 & _T_21; // @[IFU.scala 582:119]
    wb_lastIdx <= ~_f3_last_validIdx_T_13; // @[IFU.scala 585:38]
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_mmio <= f2_mmio; // @[Reg.scala 17:22]
    end
    mmio_redirect_REG <= io_uncacheInter_fromUncache_ready & io_uncacheInter_fromUncache_valid; // @[Decoupled.scala 50:35]
    if (f0_fire) begin // @[Reg.scala 17:18]
      f1_ftq_req_ftqIdx_flag <= io_ftqInter_fromFtq_req_bits_ftqIdx_flag; // @[Reg.scala 17:22]
    end
    if (f0_fire) begin // @[Reg.scala 17:18]
      f1_ftq_req_ftqIdx_value <= io_ftqInter_fromFtq_req_bits_ftqIdx_value; // @[Reg.scala 17:22]
    end
    if (f1_fire) begin // @[Reg.scala 17:18]
      f2_ftq_req_startAddr <= f1_ftq_req_startAddr; // @[Reg.scala 17:22]
    end
    if (f1_fire) begin // @[Reg.scala 17:18]
      f2_ftq_req_nextlineStart <= f1_ftq_req_nextlineStart; // @[Reg.scala 17:22]
    end
    if (f1_fire) begin // @[Reg.scala 17:18]
      f2_doubleLine <= f1_doubleLine; // @[Reg.scala 17:22]
    end
    if (f0_fire) begin // @[Reg.scala 17:18]
      f1_ftq_req_startAddr <= io_ftqInter_fromFtq_req_bits_startAddr; // @[Reg.scala 17:22]
    end
    if (f0_fire) begin // @[Reg.scala 17:18]
      f1_ftq_req_nextlineStart <= io_ftqInter_fromFtq_req_bits_nextlineStart; // @[Reg.scala 17:22]
    end
    if (f0_fire) begin // @[Reg.scala 17:18]
      f1_ftq_req_nextStartAddr <= io_ftqInter_fromFtq_req_bits_nextStartAddr; // @[Reg.scala 17:22]
    end
    if (f0_fire) begin // @[Reg.scala 17:18]
      f1_ftq_req_ftqOffset_valid <= io_ftqInter_fromFtq_req_bits_ftqOffset_valid; // @[Reg.scala 17:22]
    end
    if (f0_fire) begin // @[Reg.scala 17:18]
      f1_ftq_req_ftqOffset_bits <= io_ftqInter_fromFtq_req_bits_ftqOffset_bits; // @[Reg.scala 17:22]
    end
    if (f0_fire) begin // @[Reg.scala 17:18]
      f1_doubleLine <= f0_doubleLine; // @[Reg.scala 17:22]
    end
    if (f1_fire) begin // @[Reg.scala 17:18]
      f2_ftq_req_nextStartAddr <= f1_ftq_req_nextStartAddr; // @[Reg.scala 17:22]
    end
    if (f1_fire) begin // @[Reg.scala 17:18]
      f2_ftq_req_ftqIdx_flag <= f1_ftq_req_ftqIdx_flag; // @[Reg.scala 17:22]
    end
    if (f1_fire) begin // @[Reg.scala 17:18]
      f2_ftq_req_ftqIdx_value <= f1_ftq_req_ftqIdx_value; // @[Reg.scala 17:22]
    end
    if (f1_fire) begin // @[Reg.scala 17:18]
      f2_ftq_req_ftqOffset_valid <= f1_ftq_req_ftqOffset_valid; // @[Reg.scala 17:22]
    end
    if (f1_fire) begin // @[Reg.scala 17:18]
      f2_ftq_req_ftqOffset_bits <= f1_ftq_req_ftqOffset_bits; // @[Reg.scala 17:22]
    end
    if (f1_fire) begin // @[Reg.scala 17:18]
      f2_pc_0 <= f1_pc_0; // @[Reg.scala 17:22]
    end
    if (f1_fire) begin // @[Reg.scala 17:18]
      f2_pc_1 <= f1_pc_1; // @[Reg.scala 17:22]
    end
    if (f1_fire) begin // @[Reg.scala 17:18]
      f2_pc_2 <= f1_pc_2; // @[Reg.scala 17:22]
    end
    if (f1_fire) begin // @[Reg.scala 17:18]
      f2_pc_3 <= f1_pc_3; // @[Reg.scala 17:22]
    end
    if (f1_fire) begin // @[Reg.scala 17:18]
      f2_pc_4 <= f1_pc_4; // @[Reg.scala 17:22]
    end
    if (f1_fire) begin // @[Reg.scala 17:18]
      f2_pc_5 <= f1_pc_5; // @[Reg.scala 17:22]
    end
    if (f1_fire) begin // @[Reg.scala 17:18]
      f2_pc_6 <= f1_pc_6; // @[Reg.scala 17:22]
    end
    if (f1_fire) begin // @[Reg.scala 17:18]
      f2_pc_7 <= f1_pc_7; // @[Reg.scala 17:22]
    end
    if (f1_fire) begin // @[Reg.scala 17:18]
      f2_half_snpc_0 <= f1_pc_2; // @[Reg.scala 17:22]
    end
    if (f1_fire) begin // @[Reg.scala 17:18]
      f2_half_snpc_1 <= f1_pc_3; // @[Reg.scala 17:22]
    end
    if (f1_fire) begin // @[Reg.scala 17:18]
      f2_half_snpc_2 <= f1_pc_4; // @[Reg.scala 17:22]
    end
    if (f1_fire) begin // @[Reg.scala 17:18]
      f2_half_snpc_3 <= f1_pc_5; // @[Reg.scala 17:22]
    end
    if (f1_fire) begin // @[Reg.scala 17:18]
      f2_half_snpc_4 <= f1_pc_6; // @[Reg.scala 17:22]
    end
    if (f1_fire) begin // @[Reg.scala 17:18]
      f2_half_snpc_5 <= f1_pc_7; // @[Reg.scala 17:22]
    end
    if (f1_fire) begin // @[Reg.scala 17:18]
      f2_half_snpc_6 <= f1_half_snpc_6; // @[Reg.scala 17:22]
    end
    if (f1_fire) begin // @[Reg.scala 17:18]
      f2_half_snpc_7 <= f1_half_snpc_7; // @[Reg.scala 17:22]
    end
    if (f1_fire) begin // @[Reg.scala 17:18]
      f2_cut_ptr_0 <= f1_cut_ptr_0; // @[Reg.scala 17:22]
    end
    if (f1_fire) begin // @[Reg.scala 17:18]
      f2_cut_ptr_1 <= f1_cut_ptr_1; // @[Reg.scala 17:22]
    end
    if (f1_fire) begin // @[Reg.scala 17:18]
      f2_cut_ptr_2 <= f1_cut_ptr_2; // @[Reg.scala 17:22]
    end
    if (f1_fire) begin // @[Reg.scala 17:18]
      f2_cut_ptr_3 <= f1_cut_ptr_3; // @[Reg.scala 17:22]
    end
    if (f1_fire) begin // @[Reg.scala 17:18]
      f2_cut_ptr_4 <= f1_cut_ptr_4; // @[Reg.scala 17:22]
    end
    if (f1_fire) begin // @[Reg.scala 17:18]
      f2_cut_ptr_5 <= f1_cut_ptr_5; // @[Reg.scala 17:22]
    end
    if (f1_fire) begin // @[Reg.scala 17:18]
      f2_cut_ptr_6 <= f1_cut_ptr_6; // @[Reg.scala 17:22]
    end
    if (f1_fire) begin // @[Reg.scala 17:18]
      f2_cut_ptr_7 <= f1_cut_ptr_7; // @[Reg.scala 17:22]
    end
    if (f1_fire) begin // @[Reg.scala 17:18]
      f2_cut_ptr_8 <= f1_cut_ptr_8; // @[Reg.scala 17:22]
    end
    if (f1_fire) begin // @[Reg.scala 17:18]
      f2_resend_vaddr <= f1_pc_1; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_ftq_req_startAddr <= f2_ftq_req_startAddr; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_ftq_req_nextStartAddr <= f2_ftq_req_nextStartAddr; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_ftq_req_ftqOffset_valid <= f2_ftq_req_ftqOffset_valid; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_ftq_req_ftqOffset_bits <= f2_ftq_req_ftqOffset_bits; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_doubleLine <= f2_doubleLine; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      if (2'h3 == f2_predecod_ptr) begin // @[Reg.scala 17:22]
        if (6'h2f == f2_cut_ptr_0) begin // @[IFU.scala 302:19]
          f3_cut_data_0 <= f2_cut_data_dataVec_3_47; // @[IFU.scala 302:19]
        end else if (6'h2e == f2_cut_ptr_0) begin // @[IFU.scala 302:19]
          f3_cut_data_0 <= f2_cut_data_dataVec_3_46; // @[IFU.scala 302:19]
        end else begin
          f3_cut_data_0 <= _GEN_1396;
        end
      end else if (2'h2 == f2_predecod_ptr) begin // @[Reg.scala 17:22]
        if (6'h2f == f2_cut_ptr_0) begin // @[IFU.scala 302:19]
          f3_cut_data_0 <= f2_cut_data_dataVec_2_47; // @[IFU.scala 302:19]
        end else begin
          f3_cut_data_0 <= _GEN_965;
        end
      end else if (2'h1 == f2_predecod_ptr) begin // @[Reg.scala 17:22]
        f3_cut_data_0 <= f2_cut_data_result_1_0; // @[Reg.scala 17:22]
      end else begin
        f3_cut_data_0 <= f2_cut_data_result__0;
      end
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      if (2'h3 == f2_predecod_ptr) begin // @[Reg.scala 17:22]
        if (6'h2f == f2_cut_ptr_1) begin // @[IFU.scala 302:19]
          f3_cut_data_1 <= f2_cut_data_dataVec_3_47; // @[IFU.scala 302:19]
        end else if (6'h2e == f2_cut_ptr_1) begin // @[IFU.scala 302:19]
          f3_cut_data_1 <= f2_cut_data_dataVec_3_46; // @[IFU.scala 302:19]
        end else begin
          f3_cut_data_1 <= _GEN_1444;
        end
      end else if (2'h2 == f2_predecod_ptr) begin // @[Reg.scala 17:22]
        if (6'h2f == f2_cut_ptr_1) begin // @[IFU.scala 302:19]
          f3_cut_data_1 <= f2_cut_data_dataVec_2_47; // @[IFU.scala 302:19]
        end else begin
          f3_cut_data_1 <= _GEN_1013;
        end
      end else if (2'h1 == f2_predecod_ptr) begin // @[Reg.scala 17:22]
        f3_cut_data_1 <= f2_cut_data_result_1_1; // @[Reg.scala 17:22]
      end else begin
        f3_cut_data_1 <= f2_cut_data_result__1;
      end
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      if (2'h3 == f2_predecod_ptr) begin // @[Reg.scala 17:22]
        if (6'h2f == f2_cut_ptr_2) begin // @[IFU.scala 302:19]
          f3_cut_data_2 <= f2_cut_data_dataVec_3_47; // @[IFU.scala 302:19]
        end else if (6'h2e == f2_cut_ptr_2) begin // @[IFU.scala 302:19]
          f3_cut_data_2 <= f2_cut_data_dataVec_3_46; // @[IFU.scala 302:19]
        end else begin
          f3_cut_data_2 <= _GEN_1492;
        end
      end else if (2'h2 == f2_predecod_ptr) begin // @[Reg.scala 17:22]
        if (6'h2f == f2_cut_ptr_2) begin // @[IFU.scala 302:19]
          f3_cut_data_2 <= f2_cut_data_dataVec_2_47; // @[IFU.scala 302:19]
        end else begin
          f3_cut_data_2 <= _GEN_1061;
        end
      end else if (2'h1 == f2_predecod_ptr) begin // @[Reg.scala 17:22]
        f3_cut_data_2 <= f2_cut_data_result_1_2; // @[Reg.scala 17:22]
      end else begin
        f3_cut_data_2 <= f2_cut_data_result__2;
      end
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      if (2'h3 == f2_predecod_ptr) begin // @[Reg.scala 17:22]
        if (6'h2f == f2_cut_ptr_3) begin // @[IFU.scala 302:19]
          f3_cut_data_3 <= f2_cut_data_dataVec_3_47; // @[IFU.scala 302:19]
        end else if (6'h2e == f2_cut_ptr_3) begin // @[IFU.scala 302:19]
          f3_cut_data_3 <= f2_cut_data_dataVec_3_46; // @[IFU.scala 302:19]
        end else begin
          f3_cut_data_3 <= _GEN_1540;
        end
      end else if (2'h2 == f2_predecod_ptr) begin // @[Reg.scala 17:22]
        if (6'h2f == f2_cut_ptr_3) begin // @[IFU.scala 302:19]
          f3_cut_data_3 <= f2_cut_data_dataVec_2_47; // @[IFU.scala 302:19]
        end else begin
          f3_cut_data_3 <= _GEN_1109;
        end
      end else if (2'h1 == f2_predecod_ptr) begin // @[Reg.scala 17:22]
        f3_cut_data_3 <= f2_cut_data_result_1_3; // @[Reg.scala 17:22]
      end else begin
        f3_cut_data_3 <= f2_cut_data_result__3;
      end
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      if (2'h3 == f2_predecod_ptr) begin // @[Reg.scala 17:22]
        if (6'h2f == f2_cut_ptr_4) begin // @[IFU.scala 302:19]
          f3_cut_data_4 <= f2_cut_data_dataVec_3_47; // @[IFU.scala 302:19]
        end else if (6'h2e == f2_cut_ptr_4) begin // @[IFU.scala 302:19]
          f3_cut_data_4 <= f2_cut_data_dataVec_3_46; // @[IFU.scala 302:19]
        end else begin
          f3_cut_data_4 <= _GEN_1588;
        end
      end else if (2'h2 == f2_predecod_ptr) begin // @[Reg.scala 17:22]
        if (6'h2f == f2_cut_ptr_4) begin // @[IFU.scala 302:19]
          f3_cut_data_4 <= f2_cut_data_dataVec_2_47; // @[IFU.scala 302:19]
        end else begin
          f3_cut_data_4 <= _GEN_1157;
        end
      end else if (2'h1 == f2_predecod_ptr) begin // @[Reg.scala 17:22]
        f3_cut_data_4 <= f2_cut_data_result_1_4; // @[Reg.scala 17:22]
      end else begin
        f3_cut_data_4 <= f2_cut_data_result__4;
      end
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      if (2'h3 == f2_predecod_ptr) begin // @[Reg.scala 17:22]
        if (6'h2f == f2_cut_ptr_5) begin // @[IFU.scala 302:19]
          f3_cut_data_5 <= f2_cut_data_dataVec_3_47; // @[IFU.scala 302:19]
        end else if (6'h2e == f2_cut_ptr_5) begin // @[IFU.scala 302:19]
          f3_cut_data_5 <= f2_cut_data_dataVec_3_46; // @[IFU.scala 302:19]
        end else begin
          f3_cut_data_5 <= _GEN_1636;
        end
      end else if (2'h2 == f2_predecod_ptr) begin // @[Reg.scala 17:22]
        if (6'h2f == f2_cut_ptr_5) begin // @[IFU.scala 302:19]
          f3_cut_data_5 <= f2_cut_data_dataVec_2_47; // @[IFU.scala 302:19]
        end else begin
          f3_cut_data_5 <= _GEN_1205;
        end
      end else if (2'h1 == f2_predecod_ptr) begin // @[Reg.scala 17:22]
        f3_cut_data_5 <= f2_cut_data_result_1_5; // @[Reg.scala 17:22]
      end else begin
        f3_cut_data_5 <= f2_cut_data_result__5;
      end
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      if (2'h3 == f2_predecod_ptr) begin // @[Reg.scala 17:22]
        if (6'h2f == f2_cut_ptr_6) begin // @[IFU.scala 302:19]
          f3_cut_data_6 <= f2_cut_data_dataVec_3_47; // @[IFU.scala 302:19]
        end else if (6'h2e == f2_cut_ptr_6) begin // @[IFU.scala 302:19]
          f3_cut_data_6 <= f2_cut_data_dataVec_3_46; // @[IFU.scala 302:19]
        end else begin
          f3_cut_data_6 <= _GEN_1684;
        end
      end else if (2'h2 == f2_predecod_ptr) begin // @[Reg.scala 17:22]
        if (6'h2f == f2_cut_ptr_6) begin // @[IFU.scala 302:19]
          f3_cut_data_6 <= f2_cut_data_dataVec_2_47; // @[IFU.scala 302:19]
        end else begin
          f3_cut_data_6 <= _GEN_1253;
        end
      end else if (2'h1 == f2_predecod_ptr) begin // @[Reg.scala 17:22]
        f3_cut_data_6 <= f2_cut_data_result_1_6; // @[Reg.scala 17:22]
      end else begin
        f3_cut_data_6 <= f2_cut_data_result__6;
      end
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      if (2'h3 == f2_predecod_ptr) begin // @[Reg.scala 17:22]
        if (6'h2f == f2_cut_ptr_7) begin // @[IFU.scala 302:19]
          f3_cut_data_7 <= f2_cut_data_dataVec_3_47; // @[IFU.scala 302:19]
        end else if (6'h2e == f2_cut_ptr_7) begin // @[IFU.scala 302:19]
          f3_cut_data_7 <= f2_cut_data_dataVec_3_46; // @[IFU.scala 302:19]
        end else begin
          f3_cut_data_7 <= _GEN_1732;
        end
      end else if (2'h2 == f2_predecod_ptr) begin // @[Reg.scala 17:22]
        if (6'h2f == f2_cut_ptr_7) begin // @[IFU.scala 302:19]
          f3_cut_data_7 <= f2_cut_data_dataVec_2_47; // @[IFU.scala 302:19]
        end else begin
          f3_cut_data_7 <= _GEN_1301;
        end
      end else if (2'h1 == f2_predecod_ptr) begin // @[Reg.scala 17:22]
        f3_cut_data_7 <= f2_cut_data_result_1_7; // @[Reg.scala 17:22]
      end else begin
        f3_cut_data_7 <= f2_cut_data_result__7;
      end
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      if (2'h3 == f2_predecod_ptr) begin // @[Reg.scala 17:22]
        if (6'h2f == f2_cut_ptr_8) begin // @[IFU.scala 302:19]
          f3_cut_data_8 <= f2_cut_data_dataVec_3_47; // @[IFU.scala 302:19]
        end else if (6'h2e == f2_cut_ptr_8) begin // @[IFU.scala 302:19]
          f3_cut_data_8 <= f2_cut_data_dataVec_3_46; // @[IFU.scala 302:19]
        end else begin
          f3_cut_data_8 <= _GEN_1780;
        end
      end else if (2'h2 == f2_predecod_ptr) begin // @[Reg.scala 17:22]
        if (6'h2f == f2_cut_ptr_8) begin // @[IFU.scala 302:19]
          f3_cut_data_8 <= f2_cut_data_dataVec_2_47; // @[IFU.scala 302:19]
        end else begin
          f3_cut_data_8 <= _GEN_1349;
        end
      end else if (2'h1 == f2_predecod_ptr) begin // @[Reg.scala 17:22]
        f3_cut_data_8 <= f2_cut_data_result_1_8; // @[Reg.scala 17:22]
      end else begin
        f3_cut_data_8 <= f2_cut_data_result__8;
      end
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_instr_0 <= preDecoderOut_instr_0; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_instr_1 <= preDecoderOut_instr_1; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_instr_2 <= preDecoderOut_instr_2; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_instr_3 <= preDecoderOut_instr_3; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_instr_4 <= preDecoderOut_instr_4; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_instr_5 <= preDecoderOut_instr_5; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_instr_6 <= preDecoderOut_instr_6; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_instr_7 <= preDecoderOut_instr_7; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_pd_0_valid <= preDecoderOut_hasHalfValid_1; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_pd_0_isRVC <= preDecoderOut_pd_0_isRVC; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_pd_0_brType <= preDecoderOut_pd_0_brType; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_pd_0_isCall <= preDecoderOut_pd_0_isCall; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_pd_0_isRet <= preDecoderOut_pd_0_isRet; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_pd_1_valid <= preDecoderOut_pd_1_valid; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_pd_1_isRVC <= preDecoderOut_pd_1_isRVC; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_pd_1_brType <= preDecoderOut_pd_1_brType; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_pd_1_isCall <= preDecoderOut_pd_1_isCall; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_pd_1_isRet <= preDecoderOut_pd_1_isRet; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_pd_2_valid <= preDecoderOut_pd_2_valid; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_pd_2_isRVC <= preDecoderOut_pd_2_isRVC; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_pd_2_brType <= preDecoderOut_pd_2_brType; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_pd_2_isCall <= preDecoderOut_pd_2_isCall; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_pd_2_isRet <= preDecoderOut_pd_2_isRet; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_pd_3_valid <= preDecoderOut_pd_3_valid; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_pd_3_isRVC <= preDecoderOut_pd_3_isRVC; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_pd_3_brType <= preDecoderOut_pd_3_brType; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_pd_3_isCall <= preDecoderOut_pd_3_isCall; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_pd_3_isRet <= preDecoderOut_pd_3_isRet; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_pd_4_valid <= preDecoderOut_pd_4_valid; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_pd_4_isRVC <= preDecoderOut_pd_4_isRVC; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_pd_4_brType <= preDecoderOut_pd_4_brType; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_pd_4_isCall <= preDecoderOut_pd_4_isCall; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_pd_4_isRet <= preDecoderOut_pd_4_isRet; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_pd_5_valid <= preDecoderOut_pd_5_valid; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_pd_5_isRVC <= preDecoderOut_pd_5_isRVC; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_pd_5_brType <= preDecoderOut_pd_5_brType; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_pd_5_isCall <= preDecoderOut_pd_5_isCall; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_pd_5_isRet <= preDecoderOut_pd_5_isRet; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_pd_6_valid <= preDecoderOut_pd_6_valid; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_pd_6_isRVC <= preDecoderOut_pd_6_isRVC; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_pd_6_brType <= preDecoderOut_pd_6_brType; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_pd_6_isCall <= preDecoderOut_pd_6_isCall; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_pd_6_isRet <= preDecoderOut_pd_6_isRet; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_pd_7_valid <= preDecoderOut_pd_7_valid; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_pd_7_isRVC <= preDecoderOut_pd_7_isRVC; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_pd_7_brType <= preDecoderOut_pd_7_brType; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_pd_7_isCall <= preDecoderOut_pd_7_isCall; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_pd_7_isRet <= preDecoderOut_pd_7_isRet; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_jump_offset_0 <= preDecoderOut_jumpOffset_0; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_jump_offset_1 <= preDecoderOut_jumpOffset_1; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_jump_offset_2 <= preDecoderOut_jumpOffset_2; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_jump_offset_3 <= preDecoderOut_jumpOffset_3; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_jump_offset_4 <= preDecoderOut_jumpOffset_4; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_jump_offset_5 <= preDecoderOut_jumpOffset_5; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_jump_offset_6 <= preDecoderOut_jumpOffset_6; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_jump_offset_7 <= preDecoderOut_jumpOffset_7; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_af_vec_0 <= f2_af_vec_0; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_af_vec_1 <= f2_af_vec_1; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_af_vec_2 <= f2_af_vec_2; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_af_vec_3 <= f2_af_vec_3; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_af_vec_4 <= f2_af_vec_4; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_af_vec_5 <= f2_af_vec_5; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_af_vec_6 <= f2_af_vec_6; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_af_vec_7 <= f2_af_vec_7; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_pf_vec_0 <= f2_pf_vec_0; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_pf_vec_1 <= f2_pf_vec_1; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_pf_vec_2 <= f2_pf_vec_2; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_pf_vec_3 <= f2_pf_vec_3; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_pf_vec_4 <= f2_pf_vec_4; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_pf_vec_5 <= f2_pf_vec_5; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_pf_vec_6 <= f2_pf_vec_6; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_pf_vec_7 <= f2_pf_vec_7; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_pc_0 <= f2_pc_0; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_pc_1 <= f2_pc_1; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_pc_2 <= f2_pc_2; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_pc_3 <= f2_pc_3; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_pc_4 <= f2_pc_4; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_pc_5 <= f2_pc_5; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_pc_6 <= f2_pc_6; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_pc_7 <= f2_pc_7; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_half_snpc_0 <= f2_half_snpc_0; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_half_snpc_1 <= f2_half_snpc_1; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_half_snpc_2 <= f2_half_snpc_2; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_half_snpc_3 <= f2_half_snpc_3; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_half_snpc_4 <= f2_half_snpc_4; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_half_snpc_5 <= f2_half_snpc_5; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_half_snpc_6 <= f2_half_snpc_6; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_half_snpc_7 <= f2_half_snpc_7; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_instr_range <= f2_instr_range; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_foldpc_0 <= f2_foldpc_0; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_foldpc_1 <= f2_foldpc_1; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_foldpc_2 <= f2_foldpc_2; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_foldpc_3 <= f2_foldpc_3; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_foldpc_4 <= f2_foldpc_4; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_foldpc_5 <= f2_foldpc_5; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_foldpc_6 <= f2_foldpc_6; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_foldpc_7 <= f2_foldpc_7; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_crossPageFault_0 <= f2_crossPageFault_0; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_crossPageFault_1 <= f2_crossPageFault_1; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_crossPageFault_2 <= f2_crossPageFault_2; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_crossPageFault_3 <= f2_crossPageFault_3; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_crossPageFault_4 <= f2_crossPageFault_4; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_crossPageFault_5 <= f2_crossPageFault_5; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_crossPageFault_6 <= f2_crossPageFault_6; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_crossPageFault_7 <= f2_crossPageFault_7; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_hasHalfValid_1 <= preDecoderOut_hasHalfValid_1; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_hasHalfValid_2 <= preDecoderOut_hasHalfValid_2; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_hasHalfValid_3 <= preDecoderOut_hasHalfValid_3; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_hasHalfValid_4 <= preDecoderOut_hasHalfValid_4; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_hasHalfValid_5 <= preDecoderOut_hasHalfValid_5; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_hasHalfValid_6 <= preDecoderOut_hasHalfValid_6; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_hasHalfValid_7 <= preDecoderOut_hasHalfValid_7; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_pAddrs_0 <= io_icacheInter_resp_0_bits_paddr; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_resend_vaddr <= f2_resend_vaddr; // @[Reg.scala 17:22]
    end
    if (f3_ftq_flush_self | f3_ftq_flush_by_older) begin // @[IFU.scala 534:53]
      f3_mmio_data_0 <= 16'h0; // @[IFU.scala 539:24]
    end else if (!(4'h0 == mmio_state)) begin // @[IFU.scala 456:21]
      if (!(4'h1 == mmio_state)) begin // @[IFU.scala 456:21]
        if (!(4'h2 == mmio_state)) begin // @[IFU.scala 456:21]
          f3_mmio_data_0 <= _GEN_2008;
        end
      end
    end
    if (f3_ftq_flush_self | f3_ftq_flush_by_older) begin // @[IFU.scala 534:53]
      f3_mmio_data_1 <= 16'h0; // @[IFU.scala 539:24]
    end else if (!(4'h0 == mmio_state)) begin // @[IFU.scala 456:21]
      if (!(4'h1 == mmio_state)) begin // @[IFU.scala 456:21]
        if (!(4'h2 == mmio_state)) begin // @[IFU.scala 456:21]
          f3_mmio_data_1 <= _GEN_2009;
        end
      end
    end
    io_mmioCommitRead_mmioFtqPtr_REG_flag <= _io_mmioCommitRead_mmioFtqPtr_new_ptr_T_2[3]; // @[CircularQueuePtr.scala 39:59]
    io_mmioCommitRead_mmioFtqPtr_REG_value <= _io_mmioCommitRead_mmioFtqPtr_new_ptr_T_2[2:0]; // @[CircularQueuePtr.scala 39:59]
    f3_mmio_to_commit_next <= f3_req_is_mmio & _mmio_redirect_T; // @[IFU.scala 424:43]
    REG <= f2_fire & _T_26; // @[IFU.scala 450:24]
    mmioFlushWb_valid_REG <= io_uncacheInter_fromUncache_ready & io_uncacheInter_fromUncache_valid; // @[Decoupled.scala 50:35]
    wb_valid_REG <= f2_fire & _T_26; // @[IFU.scala 706:51]
    wb_ftq_req_startAddr <= f3_ftq_req_startAddr; // @[IFU.scala 707:34]
    wb_check_result_stage1_fixedTaken_0 <= predChecker_io_out_stage1Out_fixedTaken_0; // @[IFU.scala 709:41]
    wb_check_result_stage1_fixedTaken_1 <= predChecker_io_out_stage1Out_fixedTaken_1; // @[IFU.scala 709:41]
    wb_check_result_stage1_fixedTaken_2 <= predChecker_io_out_stage1Out_fixedTaken_2; // @[IFU.scala 709:41]
    wb_check_result_stage1_fixedTaken_3 <= predChecker_io_out_stage1Out_fixedTaken_3; // @[IFU.scala 709:41]
    wb_check_result_stage1_fixedTaken_4 <= predChecker_io_out_stage1Out_fixedTaken_4; // @[IFU.scala 709:41]
    wb_check_result_stage1_fixedTaken_5 <= predChecker_io_out_stage1Out_fixedTaken_5; // @[IFU.scala 709:41]
    wb_check_result_stage1_fixedTaken_6 <= predChecker_io_out_stage1Out_fixedTaken_6; // @[IFU.scala 709:41]
    wb_check_result_stage1_fixedTaken_7 <= predChecker_io_out_stage1Out_fixedTaken_7; // @[IFU.scala 709:41]
    wb_instr_range <= io_toIbuffer_bits_enqEnable; // @[IFU.scala 711:34]
    wb_pc_0 <= f3_pc_0; // @[IFU.scala 712:34]
    wb_pc_1 <= f3_pc_1; // @[IFU.scala 712:34]
    wb_pc_2 <= f3_pc_2; // @[IFU.scala 712:34]
    wb_pc_3 <= f3_pc_3; // @[IFU.scala 712:34]
    wb_pc_4 <= f3_pc_4; // @[IFU.scala 712:34]
    wb_pc_5 <= f3_pc_5; // @[IFU.scala 712:34]
    wb_pc_6 <= f3_pc_6; // @[IFU.scala 712:34]
    wb_pc_7 <= f3_pc_7; // @[IFU.scala 712:34]
    wb_pd_0_isRVC <= f3_pd_0_isRVC; // @[IFU.scala 713:34]
    wb_pd_0_brType <= f3_pd_0_brType; // @[IFU.scala 713:34]
    wb_pd_0_isCall <= f3_pd_0_isCall; // @[IFU.scala 713:34]
    wb_pd_0_isRet <= f3_pd_0_isRet; // @[IFU.scala 713:34]
    wb_pd_1_isRVC <= f3_pd_1_isRVC; // @[IFU.scala 713:34]
    wb_pd_1_brType <= f3_pd_1_brType; // @[IFU.scala 713:34]
    wb_pd_1_isCall <= f3_pd_1_isCall; // @[IFU.scala 713:34]
    wb_pd_1_isRet <= f3_pd_1_isRet; // @[IFU.scala 713:34]
    wb_pd_2_isRVC <= f3_pd_2_isRVC; // @[IFU.scala 713:34]
    wb_pd_2_brType <= f3_pd_2_brType; // @[IFU.scala 713:34]
    wb_pd_2_isCall <= f3_pd_2_isCall; // @[IFU.scala 713:34]
    wb_pd_2_isRet <= f3_pd_2_isRet; // @[IFU.scala 713:34]
    wb_pd_3_isRVC <= f3_pd_3_isRVC; // @[IFU.scala 713:34]
    wb_pd_3_brType <= f3_pd_3_brType; // @[IFU.scala 713:34]
    wb_pd_3_isCall <= f3_pd_3_isCall; // @[IFU.scala 713:34]
    wb_pd_3_isRet <= f3_pd_3_isRet; // @[IFU.scala 713:34]
    wb_pd_4_isRVC <= f3_pd_4_isRVC; // @[IFU.scala 713:34]
    wb_pd_4_brType <= f3_pd_4_brType; // @[IFU.scala 713:34]
    wb_pd_4_isCall <= f3_pd_4_isCall; // @[IFU.scala 713:34]
    wb_pd_4_isRet <= f3_pd_4_isRet; // @[IFU.scala 713:34]
    wb_pd_5_isRVC <= f3_pd_5_isRVC; // @[IFU.scala 713:34]
    wb_pd_5_brType <= f3_pd_5_brType; // @[IFU.scala 713:34]
    wb_pd_5_isCall <= f3_pd_5_isCall; // @[IFU.scala 713:34]
    wb_pd_5_isRet <= f3_pd_5_isRet; // @[IFU.scala 713:34]
    wb_pd_6_isRVC <= f3_pd_6_isRVC; // @[IFU.scala 713:34]
    wb_pd_6_brType <= f3_pd_6_brType; // @[IFU.scala 713:34]
    wb_pd_6_isCall <= f3_pd_6_isCall; // @[IFU.scala 713:34]
    wb_pd_6_isRet <= f3_pd_6_isRet; // @[IFU.scala 713:34]
    wb_pd_7_isRVC <= f3_pd_7_isRVC; // @[IFU.scala 713:34]
    wb_pd_7_brType <= f3_pd_7_brType; // @[IFU.scala 713:34]
    wb_pd_7_isCall <= f3_pd_7_isCall; // @[IFU.scala 713:34]
    wb_pd_7_isRet <= f3_pd_7_isRet; // @[IFU.scala 713:34]
    if (f3_lastHalf_valid) begin // @[IFU.scala 605:24]
      wb_instr_valid_0 <= 1'h0;
    end else begin
      wb_instr_valid_0 <= f3_pd_0_valid;
    end
    if (f3_lastHalf_valid) begin // @[IFU.scala 605:24]
      wb_instr_valid_1 <= f3_hasHalfValid_1;
    end else begin
      wb_instr_valid_1 <= f3_pd_1_valid;
    end
    if (f3_lastHalf_valid) begin // @[IFU.scala 605:24]
      wb_instr_valid_2 <= f3_hasHalfValid_2;
    end else begin
      wb_instr_valid_2 <= f3_pd_2_valid;
    end
    if (f3_lastHalf_valid) begin // @[IFU.scala 605:24]
      wb_instr_valid_3 <= f3_hasHalfValid_3;
    end else begin
      wb_instr_valid_3 <= f3_pd_3_valid;
    end
    if (f3_lastHalf_valid) begin // @[IFU.scala 605:24]
      wb_instr_valid_4 <= f3_hasHalfValid_4;
    end else begin
      wb_instr_valid_4 <= f3_pd_4_valid;
    end
    if (f3_lastHalf_valid) begin // @[IFU.scala 605:24]
      wb_instr_valid_5 <= f3_hasHalfValid_5;
    end else begin
      wb_instr_valid_5 <= f3_pd_5_valid;
    end
    if (f3_lastHalf_valid) begin // @[IFU.scala 605:24]
      wb_instr_valid_6 <= f3_hasHalfValid_6;
    end else begin
      wb_instr_valid_6 <= f3_pd_6_valid;
    end
    if (f3_lastHalf_valid) begin // @[IFU.scala 605:24]
      wb_instr_valid_7 <= f3_hasHalfValid_7;
    end else begin
      wb_instr_valid_7 <= f3_pd_7_valid;
    end
    if (3'h7 == f3_last_validIdx) begin // @[IFU.scala 719:34]
      wb_false_target <= f3_half_snpc_7; // @[IFU.scala 719:34]
    end else if (3'h6 == f3_last_validIdx) begin // @[IFU.scala 719:34]
      wb_false_target <= f3_half_snpc_6; // @[IFU.scala 719:34]
    end else if (3'h5 == f3_last_validIdx) begin // @[IFU.scala 719:34]
      wb_false_target <= f3_half_snpc_5; // @[IFU.scala 719:34]
    end else if (3'h4 == f3_last_validIdx) begin // @[IFU.scala 719:34]
      wb_false_target <= f3_half_snpc_4; // @[IFU.scala 719:34]
    end else begin
      wb_false_target <= _GEN_2093;
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_perf_info_only_0_hit <= io_icachePerfInfo_only_0_hit; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_perf_info_only_0_miss <= io_icachePerfInfo_only_0_miss; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_perf_info_hit_0_hit_1 <= io_icachePerfInfo_hit_0_hit_1; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_perf_info_hit_0_miss_1 <= io_icachePerfInfo_hit_0_miss_1; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_perf_info_miss_0_hit_1 <= io_icachePerfInfo_miss_0_hit_1; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_perf_info_miss_0_miss_1 <= io_icachePerfInfo_miss_0_miss_1; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_perf_info_hit_0_except_1 <= io_icachePerfInfo_hit_0_except_1; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_perf_info_miss_0_except_1 <= io_icachePerfInfo_miss_0_except_1; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_perf_info_except_0 <= io_icachePerfInfo_except_0; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_perf_info_bank_hit_1 <= io_icachePerfInfo_bank_hit_1; // @[Reg.scala 17:22]
    end
    if (f2_fire) begin // @[Reg.scala 17:18]
      f3_perf_info_hit <= io_icachePerfInfo_hit; // @[Reg.scala 17:22]
    end
    io_perf_0_value_REG <= checkFlushWb_bits_misOffset_valid & wb_valid; // @[IFU.scala 765:52]
    io_perf_0_value_REG_1 <= io_perf_0_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_1_value_REG <= io_toIbuffer_ready & io_toIbuffer_valid; // @[Decoupled.scala 50:35]
    io_perf_1_value_REG_1 <= io_perf_1_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_2_value_REG <= f3_fire & ~f3_perf_info_hit; // @[IFU.scala 798:59]
    io_perf_2_value_REG_1 <= io_perf_2_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_3_value_REG <= io_toIbuffer_ready & io_toIbuffer_valid; // @[Decoupled.scala 50:35]
    io_perf_3_value_REG_1 <= io_perf_3_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_4_value_REG <= f3_fire & f3_doubleLine; // @[IFU.scala 791:41]
    io_perf_4_value_REG_1 <= io_perf_4_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_5_value_REG <= f3_req_1 & f3_perf_info_bank_hit_1; // @[IFU.scala 793:58]
    io_perf_5_value_REG_1 <= io_perf_5_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_6_value_REG <= f3_req_1 & f3_perf_info_bank_hit_1; // @[IFU.scala 793:58]
    io_perf_6_value_REG_1 <= io_perf_6_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_7_value_REG <= f3_perf_info_only_0_hit & f3_fire; // @[IFU.scala 803:69]
    io_perf_7_value_REG_1 <= io_perf_7_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_8_value_REG <= f3_perf_info_only_0_miss & f3_fire; // @[IFU.scala 804:69]
    io_perf_8_value_REG_1 <= io_perf_8_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_9_value_REG <= f3_perf_info_hit_0_hit_1 & f3_fire; // @[IFU.scala 805:69]
    io_perf_9_value_REG_1 <= io_perf_9_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_10_value_REG <= f3_perf_info_hit_0_miss_1 & f3_fire; // @[IFU.scala 806:69]
    io_perf_10_value_REG_1 <= io_perf_10_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_11_value_REG <= f3_perf_info_miss_0_hit_1 & f3_fire; // @[IFU.scala 807:69]
    io_perf_11_value_REG_1 <= io_perf_11_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_12_value_REG <= f3_perf_info_miss_0_miss_1 & f3_fire; // @[IFU.scala 808:69]
    io_perf_12_value_REG_1 <= io_perf_12_value_REG; // @[PerfCounterUtils.scala 188:27]
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[IFU.scala 439:85]
      f3_valid <= 1'h0; // @[IFU.scala 439:95]
    end else if (f3_flush & ~f3_req_is_mmio) begin // @[IFU.scala 440:85]
      f3_valid <= 1'h0; // @[IFU.scala 440:95]
    end else if (mmioF3Flush & f3_req_is_mmio & ~f3_need_not_flush) begin
      f3_valid <= 1'h0;
    end else begin
      f3_valid <= _GEN_1960;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[IFU.scala 534:53]
      mmio_state <= 4'h0; // @[IFU.scala 535:16]
    end else if (f3_ftq_flush_self | f3_ftq_flush_by_older) begin // @[IFU.scala 456:21]
      mmio_state <= 4'h0; // @[IFU.scala 458:27 459:20 418:27]
    end else if (4'h0 == mmio_state) begin // @[IFU.scala 456:21]
      if (f3_req_is_mmio) begin // @[IFU.scala 464:27]
        mmio_state <= 4'h1; // @[IFU.scala 465:20]
      end
    end else if (4'h1 == mmio_state) begin // @[IFU.scala 456:21]
      if (is_first_instr) begin // @[IFU.scala 472:18]
        mmio_state <= 4'h2;
      end else begin
        mmio_state <= _mmio_state_T;
      end
    end else if (4'h2 == mmio_state) begin
      mmio_state <= _mmio_state_T_2;
    end else begin
      mmio_state <= _GEN_2006;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[IFU.scala 450:64]
      f3_mmio_use_seq_pc <= 1'h0; // @[IFU.scala 450:85]
    end else begin
      f3_mmio_use_seq_pc <= REG & f3_req_is_mmio | _GEN_1963;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[IFU.scala 214:35]
      f1_valid <= 1'h0; // @[IFU.scala 214:46]
    end else if (f1_flush) begin
      f1_valid <= 1'h0;
    end else begin
      f1_valid <= _GEN_11;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[IFU.scala 256:35]
      f2_valid <= 1'h0; // @[IFU.scala 256:45]
    end else if (f2_flush) begin
      f2_valid <= 1'h0;
    end else begin
      f2_valid <= _GEN_27;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[IFU.scala 252:63]
      f2_icache_all_resp_reg <= 1'h0; // @[IFU.scala 252:87]
    end else if (f2_flush) begin
      f2_icache_all_resp_reg <= 1'h0;
    end else begin
      f2_icache_all_resp_reg <= _GEN_24;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[IFU.scala 534:53]
      mmio_is_RVC <= 1'h0; // @[IFU.scala 536:17]
    end else if (f3_ftq_flush_self | f3_ftq_flush_by_older) begin // @[IFU.scala 456:21]
      mmio_is_RVC <= 1'h0; // @[IFU.scala 408:32]
    end else if (!(4'h0 == mmio_state)) begin // @[IFU.scala 456:21]
      if (!(4'h1 == mmio_state)) begin // @[IFU.scala 456:21]
        if (!(4'h2 == mmio_state)) begin
          mmio_is_RVC <= _GEN_2007;
        end
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[IFU.scala 534:53]
      mmio_resend_addr <= 36'h0; // @[IFU.scala 537:22]
    end else if (f3_ftq_flush_self | f3_ftq_flush_by_older) begin // @[IFU.scala 456:21]
      mmio_resend_addr <= 36'h0; // @[IFU.scala 409:32]
    end else if (!(4'h0 == mmio_state)) begin // @[IFU.scala 456:21]
      if (!(4'h1 == mmio_state)) begin // @[IFU.scala 456:21]
        if (!(4'h2 == mmio_state)) begin
          mmio_resend_addr <= _GEN_2010;
        end
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[IFU.scala 534:53]
      mmio_resend_af <= 1'h0; // @[IFU.scala 538:20]
    end else if (f3_ftq_flush_self | f3_ftq_flush_by_older) begin // @[IFU.scala 456:21]
      mmio_resend_af <= 1'h0; // @[IFU.scala 410:32]
    end else if (!(4'h0 == mmio_state)) begin // @[IFU.scala 456:21]
      if (!(4'h1 == mmio_state)) begin // @[IFU.scala 456:21]
        if (!(4'h2 == mmio_state)) begin
          mmio_resend_af <= _GEN_2011;
        end
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[IFU.scala 456:21]
      mmio_resend_pf <= 1'h0; // @[IFU.scala 411:32]
    end else if (!(4'h0 == mmio_state)) begin // @[IFU.scala 456:21]
      if (!(4'h1 == mmio_state)) begin // @[IFU.scala 456:21]
        if (!(4'h2 == mmio_state)) begin // @[IFU.scala 456:21]
          if (!(4'h3 == mmio_state)) begin
            mmio_resend_pf <= _GEN_2003;
          end
        end
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[IFU.scala 435:38]
      is_first_instr <= 1'h1; // @[IFU.scala 436:20]
    end else if (is_first_instr & mmio_commit) begin // @[IFU.scala 414:31]
      is_first_instr <= 1'h0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[IFU.scala 428:38]
      fromFtqRedirectReg_valid <= 1'h0; // @[IFU.scala 428:38]
    end else begin
      fromFtqRedirectReg_valid <= io_ftqInter_fromFtq_redirect_valid; // @[IFU.scala 428:38]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[IFU.scala 428:38]
      fromFtqRedirectReg_bits_ftqIdx_flag <= 1'h0; // @[IFU.scala 428:38]
    end else begin
      fromFtqRedirectReg_bits_ftqIdx_flag <= io_ftqInter_fromFtq_redirect_bits_ftqIdx_flag; // @[IFU.scala 428:38]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[IFU.scala 428:38]
      fromFtqRedirectReg_bits_ftqIdx_value <= 3'h0; // @[IFU.scala 428:38]
    end else begin
      fromFtqRedirectReg_bits_ftqIdx_value <= io_ftqInter_fromFtq_redirect_bits_ftqIdx_value; // @[IFU.scala 428:38]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[IFU.scala 428:38]
      fromFtqRedirectReg_bits_ftqOffset <= 3'h0; // @[IFU.scala 428:38]
    end else begin
      fromFtqRedirectReg_bits_ftqOffset <= io_ftqInter_fromFtq_redirect_bits_ftqOffset; // @[IFU.scala 428:38]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[IFU.scala 428:38]
      fromFtqRedirectReg_bits_level <= 1'h0; // @[IFU.scala 428:38]
    end else begin
      fromFtqRedirectReg_bits_level <= io_ftqInter_fromFtq_redirect_bits_level; // @[IFU.scala 428:38]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[IFU.scala 174:32]
      mmioF3Flush <= 1'h0;
    end else begin
      mmioF3Flush <= io_ftqInter_fromFtq_redirect_valid | wb_redirect & ~f3_wb_not_flush;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[IFU.scala 744:8]
      f3_lastHalf_valid <= 1'h0; // @[IFU.scala 745:23]
    end else if (_T_91) begin // @[IFU.scala 598:19]
      f3_lastHalf_valid <= 1'h0; // @[IFU.scala 599:23]
    end else if (f3_flush) begin // @[IFU.scala 600:24]
      f3_lastHalf_valid <= 1'h0; // @[IFU.scala 601:23]
    end else if (f3_fire) begin // @[IFU.scala 563:34]
      f3_lastHalf_valid <= f3_hasLastHalf & ~f3_lastHalf_disable;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[IFU.scala 737:8]
      f3_lastHalf_disable <= 1'h0; // @[IFU.scala 738:25]
    end else begin
      f3_lastHalf_disable <= _T_88 | _GEN_2072;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[IFU.scala 582:119]
      REG_1 <= 1'h0;
    end else begin
      REG_1 <= ~f3_pd_7_isRVC & predChecker_io_out_stage1Out_fixedRange_7 & f3_instr_valid_7 & ~
        predChecker_io_out_stage1Out_fixedTaken_7 & _T_21;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Decoupled.scala 50:35]
      REG_2 <= 1'h0;
    end else begin
      REG_2 <= io_toIbuffer_ready & io_toIbuffer_valid;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[IFU.scala 582:119]
      REG_3 <= 1'h0;
    end else begin
      REG_3 <= ~f3_pd_7_isRVC & predChecker_io_out_stage1Out_fixedRange_7 & f3_instr_valid_7 & ~
        predChecker_io_out_stage1Out_fixedTaken_7 & _T_21;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ChiselDB.scala 134:16]
      cnt <= 64'h0;
    end else begin
      cnt <= cnt + 64'h1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ChiselDB.scala 134:16]
      cnt_1 <= 64'h0;
    end else begin
      cnt_1 <= cnt_1 + 64'h1;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wb_ftq_req_ftqIdx_flag = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  wb_ftq_req_ftqIdx_value = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  f3_ftq_req_ftqIdx_flag = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  f3_ftq_req_ftqIdx_value = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  f3_valid = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  wb_valid = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  wb_false_lastHalf_REG = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  wb_lastIdx = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  f3_mmio = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  mmio_state = _RAND_9[3:0];
  _RAND_10 = {1{`RANDOM}};
  mmio_redirect_REG = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  f3_mmio_use_seq_pc = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  f1_ftq_req_ftqIdx_flag = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  f1_ftq_req_ftqIdx_value = _RAND_13[2:0];
  _RAND_14 = {1{`RANDOM}};
  f1_valid = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  f2_valid = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  f2_icache_all_resp_reg = _RAND_16[0:0];
  _RAND_17 = {2{`RANDOM}};
  f2_ftq_req_startAddr = _RAND_17[38:0];
  _RAND_18 = {2{`RANDOM}};
  f2_ftq_req_nextlineStart = _RAND_18[38:0];
  _RAND_19 = {1{`RANDOM}};
  f2_doubleLine = _RAND_19[0:0];
  _RAND_20 = {2{`RANDOM}};
  f1_ftq_req_startAddr = _RAND_20[38:0];
  _RAND_21 = {2{`RANDOM}};
  f1_ftq_req_nextlineStart = _RAND_21[38:0];
  _RAND_22 = {2{`RANDOM}};
  f1_ftq_req_nextStartAddr = _RAND_22[38:0];
  _RAND_23 = {1{`RANDOM}};
  f1_ftq_req_ftqOffset_valid = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  f1_ftq_req_ftqOffset_bits = _RAND_24[2:0];
  _RAND_25 = {1{`RANDOM}};
  f1_doubleLine = _RAND_25[0:0];
  _RAND_26 = {2{`RANDOM}};
  f2_ftq_req_nextStartAddr = _RAND_26[38:0];
  _RAND_27 = {1{`RANDOM}};
  f2_ftq_req_ftqIdx_flag = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  f2_ftq_req_ftqIdx_value = _RAND_28[2:0];
  _RAND_29 = {1{`RANDOM}};
  f2_ftq_req_ftqOffset_valid = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  f2_ftq_req_ftqOffset_bits = _RAND_30[2:0];
  _RAND_31 = {2{`RANDOM}};
  f2_pc_0 = _RAND_31[38:0];
  _RAND_32 = {2{`RANDOM}};
  f2_pc_1 = _RAND_32[38:0];
  _RAND_33 = {2{`RANDOM}};
  f2_pc_2 = _RAND_33[38:0];
  _RAND_34 = {2{`RANDOM}};
  f2_pc_3 = _RAND_34[38:0];
  _RAND_35 = {2{`RANDOM}};
  f2_pc_4 = _RAND_35[38:0];
  _RAND_36 = {2{`RANDOM}};
  f2_pc_5 = _RAND_36[38:0];
  _RAND_37 = {2{`RANDOM}};
  f2_pc_6 = _RAND_37[38:0];
  _RAND_38 = {2{`RANDOM}};
  f2_pc_7 = _RAND_38[38:0];
  _RAND_39 = {2{`RANDOM}};
  f2_half_snpc_0 = _RAND_39[38:0];
  _RAND_40 = {2{`RANDOM}};
  f2_half_snpc_1 = _RAND_40[38:0];
  _RAND_41 = {2{`RANDOM}};
  f2_half_snpc_2 = _RAND_41[38:0];
  _RAND_42 = {2{`RANDOM}};
  f2_half_snpc_3 = _RAND_42[38:0];
  _RAND_43 = {2{`RANDOM}};
  f2_half_snpc_4 = _RAND_43[38:0];
  _RAND_44 = {2{`RANDOM}};
  f2_half_snpc_5 = _RAND_44[38:0];
  _RAND_45 = {2{`RANDOM}};
  f2_half_snpc_6 = _RAND_45[38:0];
  _RAND_46 = {2{`RANDOM}};
  f2_half_snpc_7 = _RAND_46[38:0];
  _RAND_47 = {1{`RANDOM}};
  f2_cut_ptr_0 = _RAND_47[5:0];
  _RAND_48 = {1{`RANDOM}};
  f2_cut_ptr_1 = _RAND_48[5:0];
  _RAND_49 = {1{`RANDOM}};
  f2_cut_ptr_2 = _RAND_49[5:0];
  _RAND_50 = {1{`RANDOM}};
  f2_cut_ptr_3 = _RAND_50[5:0];
  _RAND_51 = {1{`RANDOM}};
  f2_cut_ptr_4 = _RAND_51[5:0];
  _RAND_52 = {1{`RANDOM}};
  f2_cut_ptr_5 = _RAND_52[5:0];
  _RAND_53 = {1{`RANDOM}};
  f2_cut_ptr_6 = _RAND_53[5:0];
  _RAND_54 = {1{`RANDOM}};
  f2_cut_ptr_7 = _RAND_54[5:0];
  _RAND_55 = {1{`RANDOM}};
  f2_cut_ptr_8 = _RAND_55[5:0];
  _RAND_56 = {2{`RANDOM}};
  f2_resend_vaddr = _RAND_56[38:0];
  _RAND_57 = {2{`RANDOM}};
  f3_ftq_req_startAddr = _RAND_57[38:0];
  _RAND_58 = {2{`RANDOM}};
  f3_ftq_req_nextStartAddr = _RAND_58[38:0];
  _RAND_59 = {1{`RANDOM}};
  f3_ftq_req_ftqOffset_valid = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  f3_ftq_req_ftqOffset_bits = _RAND_60[2:0];
  _RAND_61 = {1{`RANDOM}};
  f3_doubleLine = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  f3_cut_data_0 = _RAND_62[15:0];
  _RAND_63 = {1{`RANDOM}};
  f3_cut_data_1 = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  f3_cut_data_2 = _RAND_64[15:0];
  _RAND_65 = {1{`RANDOM}};
  f3_cut_data_3 = _RAND_65[15:0];
  _RAND_66 = {1{`RANDOM}};
  f3_cut_data_4 = _RAND_66[15:0];
  _RAND_67 = {1{`RANDOM}};
  f3_cut_data_5 = _RAND_67[15:0];
  _RAND_68 = {1{`RANDOM}};
  f3_cut_data_6 = _RAND_68[15:0];
  _RAND_69 = {1{`RANDOM}};
  f3_cut_data_7 = _RAND_69[15:0];
  _RAND_70 = {1{`RANDOM}};
  f3_cut_data_8 = _RAND_70[15:0];
  _RAND_71 = {1{`RANDOM}};
  f3_instr_0 = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  f3_instr_1 = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  f3_instr_2 = _RAND_73[31:0];
  _RAND_74 = {1{`RANDOM}};
  f3_instr_3 = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  f3_instr_4 = _RAND_75[31:0];
  _RAND_76 = {1{`RANDOM}};
  f3_instr_5 = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  f3_instr_6 = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  f3_instr_7 = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  f3_pd_0_valid = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  f3_pd_0_isRVC = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  f3_pd_0_brType = _RAND_81[1:0];
  _RAND_82 = {1{`RANDOM}};
  f3_pd_0_isCall = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  f3_pd_0_isRet = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  f3_pd_1_valid = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  f3_pd_1_isRVC = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  f3_pd_1_brType = _RAND_86[1:0];
  _RAND_87 = {1{`RANDOM}};
  f3_pd_1_isCall = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  f3_pd_1_isRet = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  f3_pd_2_valid = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  f3_pd_2_isRVC = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  f3_pd_2_brType = _RAND_91[1:0];
  _RAND_92 = {1{`RANDOM}};
  f3_pd_2_isCall = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  f3_pd_2_isRet = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  f3_pd_3_valid = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  f3_pd_3_isRVC = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  f3_pd_3_brType = _RAND_96[1:0];
  _RAND_97 = {1{`RANDOM}};
  f3_pd_3_isCall = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  f3_pd_3_isRet = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  f3_pd_4_valid = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  f3_pd_4_isRVC = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  f3_pd_4_brType = _RAND_101[1:0];
  _RAND_102 = {1{`RANDOM}};
  f3_pd_4_isCall = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  f3_pd_4_isRet = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  f3_pd_5_valid = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  f3_pd_5_isRVC = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  f3_pd_5_brType = _RAND_106[1:0];
  _RAND_107 = {1{`RANDOM}};
  f3_pd_5_isCall = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  f3_pd_5_isRet = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  f3_pd_6_valid = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  f3_pd_6_isRVC = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  f3_pd_6_brType = _RAND_111[1:0];
  _RAND_112 = {1{`RANDOM}};
  f3_pd_6_isCall = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  f3_pd_6_isRet = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  f3_pd_7_valid = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  f3_pd_7_isRVC = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  f3_pd_7_brType = _RAND_116[1:0];
  _RAND_117 = {1{`RANDOM}};
  f3_pd_7_isCall = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  f3_pd_7_isRet = _RAND_118[0:0];
  _RAND_119 = {2{`RANDOM}};
  f3_jump_offset_0 = _RAND_119[63:0];
  _RAND_120 = {2{`RANDOM}};
  f3_jump_offset_1 = _RAND_120[63:0];
  _RAND_121 = {2{`RANDOM}};
  f3_jump_offset_2 = _RAND_121[63:0];
  _RAND_122 = {2{`RANDOM}};
  f3_jump_offset_3 = _RAND_122[63:0];
  _RAND_123 = {2{`RANDOM}};
  f3_jump_offset_4 = _RAND_123[63:0];
  _RAND_124 = {2{`RANDOM}};
  f3_jump_offset_5 = _RAND_124[63:0];
  _RAND_125 = {2{`RANDOM}};
  f3_jump_offset_6 = _RAND_125[63:0];
  _RAND_126 = {2{`RANDOM}};
  f3_jump_offset_7 = _RAND_126[63:0];
  _RAND_127 = {1{`RANDOM}};
  f3_af_vec_0 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  f3_af_vec_1 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  f3_af_vec_2 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  f3_af_vec_3 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  f3_af_vec_4 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  f3_af_vec_5 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  f3_af_vec_6 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  f3_af_vec_7 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  f3_pf_vec_0 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  f3_pf_vec_1 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  f3_pf_vec_2 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  f3_pf_vec_3 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  f3_pf_vec_4 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  f3_pf_vec_5 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  f3_pf_vec_6 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  f3_pf_vec_7 = _RAND_142[0:0];
  _RAND_143 = {2{`RANDOM}};
  f3_pc_0 = _RAND_143[38:0];
  _RAND_144 = {2{`RANDOM}};
  f3_pc_1 = _RAND_144[38:0];
  _RAND_145 = {2{`RANDOM}};
  f3_pc_2 = _RAND_145[38:0];
  _RAND_146 = {2{`RANDOM}};
  f3_pc_3 = _RAND_146[38:0];
  _RAND_147 = {2{`RANDOM}};
  f3_pc_4 = _RAND_147[38:0];
  _RAND_148 = {2{`RANDOM}};
  f3_pc_5 = _RAND_148[38:0];
  _RAND_149 = {2{`RANDOM}};
  f3_pc_6 = _RAND_149[38:0];
  _RAND_150 = {2{`RANDOM}};
  f3_pc_7 = _RAND_150[38:0];
  _RAND_151 = {2{`RANDOM}};
  f3_half_snpc_0 = _RAND_151[38:0];
  _RAND_152 = {2{`RANDOM}};
  f3_half_snpc_1 = _RAND_152[38:0];
  _RAND_153 = {2{`RANDOM}};
  f3_half_snpc_2 = _RAND_153[38:0];
  _RAND_154 = {2{`RANDOM}};
  f3_half_snpc_3 = _RAND_154[38:0];
  _RAND_155 = {2{`RANDOM}};
  f3_half_snpc_4 = _RAND_155[38:0];
  _RAND_156 = {2{`RANDOM}};
  f3_half_snpc_5 = _RAND_156[38:0];
  _RAND_157 = {2{`RANDOM}};
  f3_half_snpc_6 = _RAND_157[38:0];
  _RAND_158 = {2{`RANDOM}};
  f3_half_snpc_7 = _RAND_158[38:0];
  _RAND_159 = {1{`RANDOM}};
  f3_instr_range = _RAND_159[7:0];
  _RAND_160 = {1{`RANDOM}};
  f3_foldpc_0 = _RAND_160[9:0];
  _RAND_161 = {1{`RANDOM}};
  f3_foldpc_1 = _RAND_161[9:0];
  _RAND_162 = {1{`RANDOM}};
  f3_foldpc_2 = _RAND_162[9:0];
  _RAND_163 = {1{`RANDOM}};
  f3_foldpc_3 = _RAND_163[9:0];
  _RAND_164 = {1{`RANDOM}};
  f3_foldpc_4 = _RAND_164[9:0];
  _RAND_165 = {1{`RANDOM}};
  f3_foldpc_5 = _RAND_165[9:0];
  _RAND_166 = {1{`RANDOM}};
  f3_foldpc_6 = _RAND_166[9:0];
  _RAND_167 = {1{`RANDOM}};
  f3_foldpc_7 = _RAND_167[9:0];
  _RAND_168 = {1{`RANDOM}};
  f3_crossPageFault_0 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  f3_crossPageFault_1 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  f3_crossPageFault_2 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  f3_crossPageFault_3 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  f3_crossPageFault_4 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  f3_crossPageFault_5 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  f3_crossPageFault_6 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  f3_crossPageFault_7 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  f3_hasHalfValid_1 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  f3_hasHalfValid_2 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  f3_hasHalfValid_3 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  f3_hasHalfValid_4 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  f3_hasHalfValid_5 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  f3_hasHalfValid_6 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  f3_hasHalfValid_7 = _RAND_182[0:0];
  _RAND_183 = {2{`RANDOM}};
  f3_pAddrs_0 = _RAND_183[35:0];
  _RAND_184 = {2{`RANDOM}};
  f3_resend_vaddr = _RAND_184[38:0];
  _RAND_185 = {1{`RANDOM}};
  f3_mmio_data_0 = _RAND_185[15:0];
  _RAND_186 = {1{`RANDOM}};
  f3_mmio_data_1 = _RAND_186[15:0];
  _RAND_187 = {1{`RANDOM}};
  mmio_is_RVC = _RAND_187[0:0];
  _RAND_188 = {2{`RANDOM}};
  mmio_resend_addr = _RAND_188[35:0];
  _RAND_189 = {1{`RANDOM}};
  mmio_resend_af = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  mmio_resend_pf = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  is_first_instr = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  io_mmioCommitRead_mmioFtqPtr_REG_flag = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  io_mmioCommitRead_mmioFtqPtr_REG_value = _RAND_193[2:0];
  _RAND_194 = {1{`RANDOM}};
  f3_mmio_to_commit_next = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  fromFtqRedirectReg_valid = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  fromFtqRedirectReg_bits_ftqIdx_flag = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  fromFtqRedirectReg_bits_ftqIdx_value = _RAND_197[2:0];
  _RAND_198 = {1{`RANDOM}};
  fromFtqRedirectReg_bits_ftqOffset = _RAND_198[2:0];
  _RAND_199 = {1{`RANDOM}};
  fromFtqRedirectReg_bits_level = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  mmioF3Flush = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  REG = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  f3_lastHalf_valid = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  f3_lastHalf_disable = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  mmioFlushWb_valid_REG = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  wb_valid_REG = _RAND_205[0:0];
  _RAND_206 = {2{`RANDOM}};
  wb_ftq_req_startAddr = _RAND_206[38:0];
  _RAND_207 = {1{`RANDOM}};
  wb_check_result_stage1_fixedTaken_0 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  wb_check_result_stage1_fixedTaken_1 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  wb_check_result_stage1_fixedTaken_2 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  wb_check_result_stage1_fixedTaken_3 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  wb_check_result_stage1_fixedTaken_4 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  wb_check_result_stage1_fixedTaken_5 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  wb_check_result_stage1_fixedTaken_6 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  wb_check_result_stage1_fixedTaken_7 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  wb_instr_range = _RAND_215[7:0];
  _RAND_216 = {2{`RANDOM}};
  wb_pc_0 = _RAND_216[38:0];
  _RAND_217 = {2{`RANDOM}};
  wb_pc_1 = _RAND_217[38:0];
  _RAND_218 = {2{`RANDOM}};
  wb_pc_2 = _RAND_218[38:0];
  _RAND_219 = {2{`RANDOM}};
  wb_pc_3 = _RAND_219[38:0];
  _RAND_220 = {2{`RANDOM}};
  wb_pc_4 = _RAND_220[38:0];
  _RAND_221 = {2{`RANDOM}};
  wb_pc_5 = _RAND_221[38:0];
  _RAND_222 = {2{`RANDOM}};
  wb_pc_6 = _RAND_222[38:0];
  _RAND_223 = {2{`RANDOM}};
  wb_pc_7 = _RAND_223[38:0];
  _RAND_224 = {1{`RANDOM}};
  wb_pd_0_isRVC = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  wb_pd_0_brType = _RAND_225[1:0];
  _RAND_226 = {1{`RANDOM}};
  wb_pd_0_isCall = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  wb_pd_0_isRet = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  wb_pd_1_isRVC = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  wb_pd_1_brType = _RAND_229[1:0];
  _RAND_230 = {1{`RANDOM}};
  wb_pd_1_isCall = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  wb_pd_1_isRet = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  wb_pd_2_isRVC = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  wb_pd_2_brType = _RAND_233[1:0];
  _RAND_234 = {1{`RANDOM}};
  wb_pd_2_isCall = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  wb_pd_2_isRet = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  wb_pd_3_isRVC = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  wb_pd_3_brType = _RAND_237[1:0];
  _RAND_238 = {1{`RANDOM}};
  wb_pd_3_isCall = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  wb_pd_3_isRet = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  wb_pd_4_isRVC = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  wb_pd_4_brType = _RAND_241[1:0];
  _RAND_242 = {1{`RANDOM}};
  wb_pd_4_isCall = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  wb_pd_4_isRet = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  wb_pd_5_isRVC = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  wb_pd_5_brType = _RAND_245[1:0];
  _RAND_246 = {1{`RANDOM}};
  wb_pd_5_isCall = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  wb_pd_5_isRet = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  wb_pd_6_isRVC = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  wb_pd_6_brType = _RAND_249[1:0];
  _RAND_250 = {1{`RANDOM}};
  wb_pd_6_isCall = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  wb_pd_6_isRet = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  wb_pd_7_isRVC = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  wb_pd_7_brType = _RAND_253[1:0];
  _RAND_254 = {1{`RANDOM}};
  wb_pd_7_isCall = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  wb_pd_7_isRet = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  wb_instr_valid_0 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  wb_instr_valid_1 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  wb_instr_valid_2 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  wb_instr_valid_3 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  wb_instr_valid_4 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  wb_instr_valid_5 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  wb_instr_valid_6 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  wb_instr_valid_7 = _RAND_263[0:0];
  _RAND_264 = {2{`RANDOM}};
  wb_false_target = _RAND_264[38:0];
  _RAND_265 = {1{`RANDOM}};
  REG_1 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  REG_2 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  REG_3 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  f3_perf_info_only_0_hit = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  f3_perf_info_only_0_miss = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  f3_perf_info_hit_0_hit_1 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  f3_perf_info_hit_0_miss_1 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  f3_perf_info_miss_0_hit_1 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  f3_perf_info_miss_0_miss_1 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  f3_perf_info_hit_0_except_1 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  f3_perf_info_miss_0_except_1 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  f3_perf_info_except_0 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  f3_perf_info_bank_hit_1 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  f3_perf_info_hit = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  io_perf_0_value_REG = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  io_perf_0_value_REG_1 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  io_perf_1_value_REG = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  io_perf_1_value_REG_1 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  io_perf_2_value_REG = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  io_perf_2_value_REG_1 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  io_perf_3_value_REG = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  io_perf_3_value_REG_1 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  io_perf_4_value_REG = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  io_perf_4_value_REG_1 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  io_perf_5_value_REG = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  io_perf_5_value_REG_1 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  io_perf_6_value_REG = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  io_perf_6_value_REG_1 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  io_perf_7_value_REG = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  io_perf_7_value_REG_1 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  io_perf_8_value_REG = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  io_perf_8_value_REG_1 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  io_perf_9_value_REG = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  io_perf_9_value_REG_1 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  io_perf_10_value_REG = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  io_perf_10_value_REG_1 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  io_perf_11_value_REG = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  io_perf_11_value_REG_1 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  io_perf_12_value_REG = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  io_perf_12_value_REG_1 = _RAND_304[0:0];
  _RAND_305 = {2{`RANDOM}};
  cnt = _RAND_305[63:0];
  _RAND_306 = {2{`RANDOM}};
  cnt_1 = _RAND_306[63:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    f3_valid = 1'h0;
  end
  if (reset) begin
    mmio_state = 4'h0;
  end
  if (reset) begin
    f3_mmio_use_seq_pc = 1'h0;
  end
  if (reset) begin
    f1_valid = 1'h0;
  end
  if (reset) begin
    f2_valid = 1'h0;
  end
  if (reset) begin
    f2_icache_all_resp_reg = 1'h0;
  end
  if (reset) begin
    mmio_is_RVC = 1'h0;
  end
  if (reset) begin
    mmio_resend_addr = 36'h0;
  end
  if (reset) begin
    mmio_resend_af = 1'h0;
  end
  if (reset) begin
    mmio_resend_pf = 1'h0;
  end
  if (reset) begin
    is_first_instr = 1'h1;
  end
  if (reset) begin
    fromFtqRedirectReg_valid = 1'h0;
  end
  if (reset) begin
    fromFtqRedirectReg_bits_ftqIdx_flag = 1'h0;
  end
  if (reset) begin
    fromFtqRedirectReg_bits_ftqIdx_value = 3'h0;
  end
  if (reset) begin
    fromFtqRedirectReg_bits_ftqOffset = 3'h0;
  end
  if (reset) begin
    fromFtqRedirectReg_bits_level = 1'h0;
  end
  if (reset) begin
    mmioF3Flush = 1'h0;
  end
  if (reset) begin
    f3_lastHalf_valid = 1'h0;
  end
  if (reset) begin
    f3_lastHalf_disable = 1'h0;
  end
  if (reset) begin
    REG_1 = 1'h0;
  end
  if (reset) begin
    REG_2 = 1'h0;
  end
  if (reset) begin
    REG_3 = 1'h0;
  end
  if (reset) begin
    cnt = 64'h0;
  end
  if (reset) begin
    cnt_1 = 64'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule

