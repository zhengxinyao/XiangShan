module FastArbiter_2(
  input        clock,
  input        reset,
  output       io_in_0_ready,
  input        io_in_0_valid,
  input  [9:0] io_in_0_bits_set,
  input  [2:0] io_in_0_bits_way,
  input        io_in_0_bits_data_dirty,
  input  [1:0] io_in_0_bits_data_state,
  input  [1:0] io_in_0_bits_data_clientStates_0,
  input  [1:0] io_in_0_bits_data_clientStates_1,
  output       io_in_1_ready,
  input        io_in_1_valid,
  input  [9:0] io_in_1_bits_set,
  input  [2:0] io_in_1_bits_way,
  input        io_in_1_bits_data_dirty,
  input  [1:0] io_in_1_bits_data_state,
  input  [1:0] io_in_1_bits_data_clientStates_0,
  input  [1:0] io_in_1_bits_data_clientStates_1,
  output       io_in_2_ready,
  input        io_in_2_valid,
  input  [9:0] io_in_2_bits_set,
  input  [2:0] io_in_2_bits_way,
  input        io_in_2_bits_data_dirty,
  input  [1:0] io_in_2_bits_data_state,
  input  [1:0] io_in_2_bits_data_clientStates_0,
  input  [1:0] io_in_2_bits_data_clientStates_1,
  output       io_in_3_ready,
  input        io_in_3_valid,
  input  [9:0] io_in_3_bits_set,
  input  [2:0] io_in_3_bits_way,
  input        io_in_3_bits_data_dirty,
  input  [1:0] io_in_3_bits_data_state,
  input  [1:0] io_in_3_bits_data_clientStates_0,
  input  [1:0] io_in_3_bits_data_clientStates_1,
  output       io_in_4_ready,
  input        io_in_4_valid,
  input  [9:0] io_in_4_bits_set,
  input  [2:0] io_in_4_bits_way,
  input        io_in_4_bits_data_dirty,
  input  [1:0] io_in_4_bits_data_state,
  input  [1:0] io_in_4_bits_data_clientStates_0,
  input  [1:0] io_in_4_bits_data_clientStates_1,
  output       io_in_5_ready,
  input        io_in_5_valid,
  input  [9:0] io_in_5_bits_set,
  input  [2:0] io_in_5_bits_way,
  input        io_in_5_bits_data_dirty,
  input  [1:0] io_in_5_bits_data_state,
  input  [1:0] io_in_5_bits_data_clientStates_0,
  input  [1:0] io_in_5_bits_data_clientStates_1,
  output       io_in_6_ready,
  input        io_in_6_valid,
  input  [9:0] io_in_6_bits_set,
  input  [2:0] io_in_6_bits_way,
  input        io_in_6_bits_data_dirty,
  input  [1:0] io_in_6_bits_data_state,
  input  [1:0] io_in_6_bits_data_clientStates_0,
  input  [1:0] io_in_6_bits_data_clientStates_1,
  output       io_in_7_ready,
  input        io_in_7_valid,
  input  [9:0] io_in_7_bits_set,
  input  [2:0] io_in_7_bits_way,
  input        io_in_7_bits_data_dirty,
  input  [1:0] io_in_7_bits_data_state,
  input  [1:0] io_in_7_bits_data_clientStates_0,
  input  [1:0] io_in_7_bits_data_clientStates_1,
  output       io_in_8_ready,
  input        io_in_8_valid,
  input  [9:0] io_in_8_bits_set,
  input  [2:0] io_in_8_bits_way,
  input        io_in_8_bits_data_dirty,
  input  [1:0] io_in_8_bits_data_state,
  input  [1:0] io_in_8_bits_data_clientStates_0,
  input  [1:0] io_in_8_bits_data_clientStates_1,
  output       io_in_9_ready,
  input        io_in_9_valid,
  input  [9:0] io_in_9_bits_set,
  input  [2:0] io_in_9_bits_way,
  input        io_in_9_bits_data_dirty,
  input  [1:0] io_in_9_bits_data_state,
  input  [1:0] io_in_9_bits_data_clientStates_0,
  input  [1:0] io_in_9_bits_data_clientStates_1,
  output       io_in_10_ready,
  input        io_in_10_valid,
  input  [9:0] io_in_10_bits_set,
  input  [2:0] io_in_10_bits_way,
  input        io_in_10_bits_data_dirty,
  input  [1:0] io_in_10_bits_data_state,
  input  [1:0] io_in_10_bits_data_clientStates_0,
  input  [1:0] io_in_10_bits_data_clientStates_1,
  output       io_in_11_ready,
  input        io_in_11_valid,
  input  [9:0] io_in_11_bits_set,
  input  [2:0] io_in_11_bits_way,
  input        io_in_11_bits_data_dirty,
  input  [1:0] io_in_11_bits_data_state,
  input  [1:0] io_in_11_bits_data_clientStates_0,
  input  [1:0] io_in_11_bits_data_clientStates_1,
  output       io_in_12_ready,
  input        io_in_12_valid,
  input  [9:0] io_in_12_bits_set,
  input  [2:0] io_in_12_bits_way,
  input        io_in_12_bits_data_dirty,
  input  [1:0] io_in_12_bits_data_state,
  input  [1:0] io_in_12_bits_data_clientStates_0,
  input  [1:0] io_in_12_bits_data_clientStates_1,
  output       io_in_13_ready,
  input        io_in_13_valid,
  input  [9:0] io_in_13_bits_set,
  input  [2:0] io_in_13_bits_way,
  input        io_in_13_bits_data_dirty,
  input  [1:0] io_in_13_bits_data_state,
  input  [1:0] io_in_13_bits_data_clientStates_0,
  input  [1:0] io_in_13_bits_data_clientStates_1,
  output       io_in_14_ready,
  input        io_in_14_valid,
  input  [9:0] io_in_14_bits_set,
  input  [2:0] io_in_14_bits_way,
  input        io_in_14_bits_data_dirty,
  input  [1:0] io_in_14_bits_data_state,
  input  [1:0] io_in_14_bits_data_clientStates_0,
  input  [1:0] io_in_14_bits_data_clientStates_1,
  output       io_in_15_ready,
  input        io_in_15_valid,
  input  [9:0] io_in_15_bits_set,
  input  [2:0] io_in_15_bits_way,
  input        io_in_15_bits_data_dirty,
  input  [1:0] io_in_15_bits_data_state,
  input  [1:0] io_in_15_bits_data_clientStates_0,
  input  [1:0] io_in_15_bits_data_clientStates_1,
  output       io_out_valid,
  output [9:0] io_out_bits_set,
  output [2:0] io_out_bits_way,
  output       io_out_bits_data_dirty,
  output [1:0] io_out_bits_data_state,
  output [1:0] io_out_bits_data_clientStates_0,
  output [1:0] io_out_bits_data_clientStates_1
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire [7:0] valids_lo = {io_in_7_valid,io_in_6_valid,io_in_5_valid,io_in_4_valid,io_in_3_valid,io_in_2_valid,
    io_in_1_valid,io_in_0_valid}; // @[FastArbiter.scala 36:50]
  wire [15:0] valids = {io_in_15_valid,io_in_14_valid,io_in_13_valid,io_in_12_valid,io_in_11_valid,io_in_10_valid,
    io_in_9_valid,io_in_8_valid,valids_lo}; // @[FastArbiter.scala 36:50]
  reg [15:0] rrGrantMask; // @[Reg.scala 28:20]
  reg [15:0] pendingMask; // @[Reg.scala 28:20]
  wire [15:0] _rrSelOH_T = rrGrantMask & pendingMask; // @[FastArbiter.scala 51:47]
  wire [1:0] rrSelOH_hi_hi_hi_6 = {_rrSelOH_T[0],_rrSelOH_T[1]}; // @[Cat.scala 31:58]
  wire [3:0] rrSelOH_hi_hi_10 = {_rrSelOH_T[0],_rrSelOH_T[1],_rrSelOH_T[2],_rrSelOH_T[3]}; // @[Cat.scala 31:58]
  wire [7:0] rrSelOH_hi_12 = {_rrSelOH_T[0],_rrSelOH_T[1],_rrSelOH_T[2],_rrSelOH_T[3],_rrSelOH_T[4],_rrSelOH_T[5],
    _rrSelOH_T[6],_rrSelOH_T[7]}; // @[Cat.scala 31:58]
  wire [6:0] rrSelOH_lo_11 = {_rrSelOH_T[8],_rrSelOH_T[9],_rrSelOH_T[10],_rrSelOH_T[11],_rrSelOH_T[12],_rrSelOH_T[13],
    _rrSelOH_T[14]}; // @[Cat.scala 31:58]
  wire [14:0] _rrSelOH_T_72 = {_rrSelOH_T[0],_rrSelOH_T[1],_rrSelOH_T[2],_rrSelOH_T[3],_rrSelOH_T[4],_rrSelOH_T[5],
    _rrSelOH_T[6],_rrSelOH_T[7],rrSelOH_lo_11}; // @[Cat.scala 31:58]
  wire  _rrSelOH_T_75 = _rrSelOH_T[15] & ~(|_rrSelOH_T_72); // @[FastArbiter.scala 28:24]
  wire [6:0] rrSelOH_hi_11 = {_rrSelOH_T[0],_rrSelOH_T[1],_rrSelOH_T[2],_rrSelOH_T[3],_rrSelOH_T[4],_rrSelOH_T[5],
    _rrSelOH_T[6]}; // @[Cat.scala 31:58]
  wire [6:0] rrSelOH_lo_10 = {_rrSelOH_T[7],_rrSelOH_T[8],_rrSelOH_T[9],_rrSelOH_T[10],_rrSelOH_T[11],_rrSelOH_T[12],
    _rrSelOH_T[13]}; // @[Cat.scala 31:58]
  wire [13:0] _rrSelOH_T_68 = {_rrSelOH_T[0],_rrSelOH_T[1],_rrSelOH_T[2],_rrSelOH_T[3],_rrSelOH_T[4],_rrSelOH_T[5],
    _rrSelOH_T[6],rrSelOH_lo_10}; // @[Cat.scala 31:58]
  wire  _rrSelOH_T_71 = _rrSelOH_T[14] & ~(|_rrSelOH_T_68); // @[FastArbiter.scala 28:24]
  wire [5:0] rrSelOH_lo_9 = {_rrSelOH_T[7],_rrSelOH_T[8],_rrSelOH_T[9],_rrSelOH_T[10],_rrSelOH_T[11],_rrSelOH_T[12]}; // @[Cat.scala 31:58]
  wire [12:0] _rrSelOH_T_64 = {_rrSelOH_T[0],_rrSelOH_T[1],_rrSelOH_T[2],_rrSelOH_T[3],_rrSelOH_T[4],_rrSelOH_T[5],
    _rrSelOH_T[6],rrSelOH_lo_9}; // @[Cat.scala 31:58]
  wire  _rrSelOH_T_67 = _rrSelOH_T[13] & ~(|_rrSelOH_T_64); // @[FastArbiter.scala 28:24]
  wire [2:0] rrSelOH_hi_hi_7 = {_rrSelOH_T[0],_rrSelOH_T[1],_rrSelOH_T[2]}; // @[Cat.scala 31:58]
  wire [5:0] rrSelOH_hi_9 = {_rrSelOH_T[0],_rrSelOH_T[1],_rrSelOH_T[2],_rrSelOH_T[3],_rrSelOH_T[4],_rrSelOH_T[5]}; // @[Cat.scala 31:58]
  wire [5:0] rrSelOH_lo_8 = {_rrSelOH_T[6],_rrSelOH_T[7],_rrSelOH_T[8],_rrSelOH_T[9],_rrSelOH_T[10],_rrSelOH_T[11]}; // @[Cat.scala 31:58]
  wire [11:0] _rrSelOH_T_60 = {_rrSelOH_T[0],_rrSelOH_T[1],_rrSelOH_T[2],_rrSelOH_T[3],_rrSelOH_T[4],_rrSelOH_T[5],
    rrSelOH_lo_8}; // @[Cat.scala 31:58]
  wire  _rrSelOH_T_63 = _rrSelOH_T[12] & ~(|_rrSelOH_T_60); // @[FastArbiter.scala 28:24]
  wire [4:0] rrSelOH_lo_7 = {_rrSelOH_T[6],_rrSelOH_T[7],_rrSelOH_T[8],_rrSelOH_T[9],_rrSelOH_T[10]}; // @[Cat.scala 31:58]
  wire [10:0] _rrSelOH_T_56 = {_rrSelOH_T[0],_rrSelOH_T[1],_rrSelOH_T[2],_rrSelOH_T[3],_rrSelOH_T[4],_rrSelOH_T[5],
    rrSelOH_lo_7}; // @[Cat.scala 31:58]
  wire  _rrSelOH_T_59 = _rrSelOH_T[11] & ~(|_rrSelOH_T_56); // @[FastArbiter.scala 28:24]
  wire [4:0] rrSelOH_hi_7 = {_rrSelOH_T[0],_rrSelOH_T[1],_rrSelOH_T[2],_rrSelOH_T[3],_rrSelOH_T[4]}; // @[Cat.scala 31:58]
  wire [9:0] _rrSelOH_T_52 = {_rrSelOH_T[0],_rrSelOH_T[1],_rrSelOH_T[2],_rrSelOH_T[3],_rrSelOH_T[4],_rrSelOH_T[5],
    _rrSelOH_T[6],_rrSelOH_T[7],_rrSelOH_T[8],_rrSelOH_T[9]}; // @[Cat.scala 31:58]
  wire  _rrSelOH_T_55 = _rrSelOH_T[10] & ~(|_rrSelOH_T_52); // @[FastArbiter.scala 28:24]
  wire [8:0] _rrSelOH_T_48 = {_rrSelOH_T[0],_rrSelOH_T[1],_rrSelOH_T[2],_rrSelOH_T[3],_rrSelOH_T[4],_rrSelOH_T[5],
    _rrSelOH_T[6],_rrSelOH_T[7],_rrSelOH_T[8]}; // @[Cat.scala 31:58]
  wire  _rrSelOH_T_51 = _rrSelOH_T[9] & ~(|_rrSelOH_T_48); // @[FastArbiter.scala 28:24]
  wire  _rrSelOH_T_47 = _rrSelOH_T[8] & ~(|rrSelOH_hi_12); // @[FastArbiter.scala 28:24]
  wire  _rrSelOH_T_43 = _rrSelOH_T[7] & ~(|rrSelOH_hi_11); // @[FastArbiter.scala 28:24]
  wire  _rrSelOH_T_39 = _rrSelOH_T[6] & ~(|rrSelOH_hi_9); // @[FastArbiter.scala 28:24]
  wire  _rrSelOH_T_35 = _rrSelOH_T[5] & ~(|rrSelOH_hi_7); // @[FastArbiter.scala 28:24]
  wire  _rrSelOH_T_31 = _rrSelOH_T[4] & ~(|rrSelOH_hi_hi_10); // @[FastArbiter.scala 28:24]
  wire  _rrSelOH_T_27 = _rrSelOH_T[3] & ~(|rrSelOH_hi_hi_7); // @[FastArbiter.scala 28:24]
  wire  _rrSelOH_T_23 = _rrSelOH_T[2] & ~(|rrSelOH_hi_hi_hi_6); // @[FastArbiter.scala 28:24]
  wire  _rrSelOH_T_19 = _rrSelOH_T[1] & ~(|_rrSelOH_T[0]); // @[FastArbiter.scala 28:24]
  wire [7:0] rrSelOH_lo_12 = {_rrSelOH_T_43,_rrSelOH_T_39,_rrSelOH_T_35,_rrSelOH_T_31,_rrSelOH_T_27,_rrSelOH_T_23,
    _rrSelOH_T_19,_rrSelOH_T[0]}; // @[FastArbiter.scala 51:80]
  wire [15:0] rrSelOH = {_rrSelOH_T_75,_rrSelOH_T_71,_rrSelOH_T_67,_rrSelOH_T_63,_rrSelOH_T_59,_rrSelOH_T_55,
    _rrSelOH_T_51,_rrSelOH_T_47,rrSelOH_lo_12}; // @[FastArbiter.scala 51:80]
  wire [15:0] _rrValid_T = rrSelOH & valids; // @[FastArbiter.scala 53:26]
  wire  rrValid = |_rrValid_T; // @[FastArbiter.scala 53:39]
  wire [1:0] firstOneOH_hi_hi_hi_6 = {valids[0],valids[1]}; // @[Cat.scala 31:58]
  wire [3:0] firstOneOH_hi_hi_10 = {valids[0],valids[1],valids[2],valids[3]}; // @[Cat.scala 31:58]
  wire [7:0] firstOneOH_hi_12 = {valids[0],valids[1],valids[2],valids[3],valids[4],valids[5],valids[6],valids[7]}; // @[Cat.scala 31:58]
  wire [6:0] firstOneOH_lo_11 = {valids[8],valids[9],valids[10],valids[11],valids[12],valids[13],valids[14]}; // @[Cat.scala 31:58]
  wire [14:0] _firstOneOH_T_71 = {valids[0],valids[1],valids[2],valids[3],valids[4],valids[5],valids[6],valids[7],
    firstOneOH_lo_11}; // @[Cat.scala 31:58]
  wire  _firstOneOH_T_74 = valids[15] & ~(|_firstOneOH_T_71); // @[FastArbiter.scala 28:24]
  wire [6:0] firstOneOH_hi_11 = {valids[0],valids[1],valids[2],valids[3],valids[4],valids[5],valids[6]}; // @[Cat.scala 31:58]
  wire [6:0] firstOneOH_lo_10 = {valids[7],valids[8],valids[9],valids[10],valids[11],valids[12],valids[13]}; // @[Cat.scala 31:58]
  wire [13:0] _firstOneOH_T_67 = {valids[0],valids[1],valids[2],valids[3],valids[4],valids[5],valids[6],firstOneOH_lo_10
    }; // @[Cat.scala 31:58]
  wire  _firstOneOH_T_70 = valids[14] & ~(|_firstOneOH_T_67); // @[FastArbiter.scala 28:24]
  wire [5:0] firstOneOH_lo_9 = {valids[7],valids[8],valids[9],valids[10],valids[11],valids[12]}; // @[Cat.scala 31:58]
  wire [12:0] _firstOneOH_T_63 = {valids[0],valids[1],valids[2],valids[3],valids[4],valids[5],valids[6],firstOneOH_lo_9}
    ; // @[Cat.scala 31:58]
  wire  _firstOneOH_T_66 = valids[13] & ~(|_firstOneOH_T_63); // @[FastArbiter.scala 28:24]
  wire [2:0] firstOneOH_hi_hi_7 = {valids[0],valids[1],valids[2]}; // @[Cat.scala 31:58]
  wire [5:0] firstOneOH_hi_9 = {valids[0],valids[1],valids[2],valids[3],valids[4],valids[5]}; // @[Cat.scala 31:58]
  wire [5:0] firstOneOH_lo_8 = {valids[6],valids[7],valids[8],valids[9],valids[10],valids[11]}; // @[Cat.scala 31:58]
  wire [11:0] _firstOneOH_T_59 = {valids[0],valids[1],valids[2],valids[3],valids[4],valids[5],firstOneOH_lo_8}; // @[Cat.scala 31:58]
  wire  _firstOneOH_T_62 = valids[12] & ~(|_firstOneOH_T_59); // @[FastArbiter.scala 28:24]
  wire [4:0] firstOneOH_lo_7 = {valids[6],valids[7],valids[8],valids[9],valids[10]}; // @[Cat.scala 31:58]
  wire [10:0] _firstOneOH_T_55 = {valids[0],valids[1],valids[2],valids[3],valids[4],valids[5],firstOneOH_lo_7}; // @[Cat.scala 31:58]
  wire  _firstOneOH_T_58 = valids[11] & ~(|_firstOneOH_T_55); // @[FastArbiter.scala 28:24]
  wire [4:0] firstOneOH_hi_7 = {valids[0],valids[1],valids[2],valids[3],valids[4]}; // @[Cat.scala 31:58]
  wire [9:0] _firstOneOH_T_51 = {valids[0],valids[1],valids[2],valids[3],valids[4],valids[5],valids[6],valids[7],valids[
    8],valids[9]}; // @[Cat.scala 31:58]
  wire  _firstOneOH_T_54 = valids[10] & ~(|_firstOneOH_T_51); // @[FastArbiter.scala 28:24]
  wire [8:0] _firstOneOH_T_47 = {valids[0],valids[1],valids[2],valids[3],valids[4],valids[5],valids[6],valids[7],valids[
    8]}; // @[Cat.scala 31:58]
  wire  _firstOneOH_T_50 = valids[9] & ~(|_firstOneOH_T_47); // @[FastArbiter.scala 28:24]
  wire  _firstOneOH_T_46 = valids[8] & ~(|firstOneOH_hi_12); // @[FastArbiter.scala 28:24]
  wire  _firstOneOH_T_42 = valids[7] & ~(|firstOneOH_hi_11); // @[FastArbiter.scala 28:24]
  wire  _firstOneOH_T_38 = valids[6] & ~(|firstOneOH_hi_9); // @[FastArbiter.scala 28:24]
  wire  _firstOneOH_T_34 = valids[5] & ~(|firstOneOH_hi_7); // @[FastArbiter.scala 28:24]
  wire  _firstOneOH_T_30 = valids[4] & ~(|firstOneOH_hi_hi_10); // @[FastArbiter.scala 28:24]
  wire  _firstOneOH_T_26 = valids[3] & ~(|firstOneOH_hi_hi_7); // @[FastArbiter.scala 28:24]
  wire  _firstOneOH_T_22 = valids[2] & ~(|firstOneOH_hi_hi_hi_6); // @[FastArbiter.scala 28:24]
  wire  _firstOneOH_T_18 = valids[1] & ~(|valids[0]); // @[FastArbiter.scala 28:24]
  wire [7:0] firstOneOH_lo_12 = {_firstOneOH_T_42,_firstOneOH_T_38,_firstOneOH_T_34,_firstOneOH_T_30,_firstOneOH_T_26,
    _firstOneOH_T_22,_firstOneOH_T_18,valids[0]}; // @[FastArbiter.scala 52:62]
  wire [15:0] firstOneOH = {_firstOneOH_T_74,_firstOneOH_T_70,_firstOneOH_T_66,_firstOneOH_T_62,_firstOneOH_T_58,
    _firstOneOH_T_54,_firstOneOH_T_50,_firstOneOH_T_46,firstOneOH_lo_12}; // @[FastArbiter.scala 52:62]
  wire [15:0] chosenOH = rrValid ? rrSelOH : firstOneOH; // @[FastArbiter.scala 54:18]
  wire [15:0] _pendingMask_T = ~chosenOH; // @[FastArbiter.scala 39:15]
  wire [15:0] _pendingMask_T_1 = valids & _pendingMask_T; // @[FastArbiter.scala 39:12]
  wire  _rrGrantMask_T_1 = |chosenOH[0]; // @[FastArbiter.scala 49:51]
  wire  _rrGrantMask_T_3 = |chosenOH[1:0]; // @[FastArbiter.scala 49:51]
  wire  _rrGrantMask_T_5 = |chosenOH[2:0]; // @[FastArbiter.scala 49:51]
  wire  _rrGrantMask_T_7 = |chosenOH[3:0]; // @[FastArbiter.scala 49:51]
  wire  _rrGrantMask_T_9 = |chosenOH[4:0]; // @[FastArbiter.scala 49:51]
  wire  _rrGrantMask_T_11 = |chosenOH[5:0]; // @[FastArbiter.scala 49:51]
  wire  _rrGrantMask_T_13 = |chosenOH[6:0]; // @[FastArbiter.scala 49:51]
  wire  _rrGrantMask_T_15 = |chosenOH[7:0]; // @[FastArbiter.scala 49:51]
  wire  _rrGrantMask_T_17 = |chosenOH[8:0]; // @[FastArbiter.scala 49:51]
  wire  _rrGrantMask_T_19 = |chosenOH[9:0]; // @[FastArbiter.scala 49:51]
  wire  _rrGrantMask_T_21 = |chosenOH[10:0]; // @[FastArbiter.scala 49:51]
  wire  _rrGrantMask_T_23 = |chosenOH[11:0]; // @[FastArbiter.scala 49:51]
  wire  _rrGrantMask_T_25 = |chosenOH[12:0]; // @[FastArbiter.scala 49:51]
  wire  _rrGrantMask_T_27 = |chosenOH[13:0]; // @[FastArbiter.scala 49:51]
  wire  _rrGrantMask_T_29 = |chosenOH[14:0]; // @[FastArbiter.scala 49:51]
  wire [7:0] rrGrantMask_lo = {_rrGrantMask_T_13,_rrGrantMask_T_11,_rrGrantMask_T_9,_rrGrantMask_T_7,_rrGrantMask_T_5,
    _rrGrantMask_T_3,_rrGrantMask_T_1,1'h0}; // @[FastArbiter.scala 50:12]
  wire [15:0] _rrGrantMask_T_30 = {_rrGrantMask_T_29,_rrGrantMask_T_27,_rrGrantMask_T_25,_rrGrantMask_T_23,
    _rrGrantMask_T_21,_rrGrantMask_T_19,_rrGrantMask_T_17,_rrGrantMask_T_15,rrGrantMask_lo}; // @[FastArbiter.scala 50:12]
  wire [1:0] _io_out_bits_T_16 = chosenOH[0] ? io_in_0_bits_data_clientStates_0 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_17 = chosenOH[1] ? io_in_1_bits_data_clientStates_0 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_18 = chosenOH[2] ? io_in_2_bits_data_clientStates_0 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_19 = chosenOH[3] ? io_in_3_bits_data_clientStates_0 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_20 = chosenOH[4] ? io_in_4_bits_data_clientStates_0 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_21 = chosenOH[5] ? io_in_5_bits_data_clientStates_0 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_22 = chosenOH[6] ? io_in_6_bits_data_clientStates_0 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_23 = chosenOH[7] ? io_in_7_bits_data_clientStates_0 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_24 = chosenOH[8] ? io_in_8_bits_data_clientStates_0 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_25 = chosenOH[9] ? io_in_9_bits_data_clientStates_0 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_26 = chosenOH[10] ? io_in_10_bits_data_clientStates_0 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_27 = chosenOH[11] ? io_in_11_bits_data_clientStates_0 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_28 = chosenOH[12] ? io_in_12_bits_data_clientStates_0 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_29 = chosenOH[13] ? io_in_13_bits_data_clientStates_0 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_30 = chosenOH[14] ? io_in_14_bits_data_clientStates_0 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_31 = chosenOH[15] ? io_in_15_bits_data_clientStates_0 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_32 = _io_out_bits_T_16 | _io_out_bits_T_17; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_33 = _io_out_bits_T_32 | _io_out_bits_T_18; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_34 = _io_out_bits_T_33 | _io_out_bits_T_19; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_35 = _io_out_bits_T_34 | _io_out_bits_T_20; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_36 = _io_out_bits_T_35 | _io_out_bits_T_21; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_37 = _io_out_bits_T_36 | _io_out_bits_T_22; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_38 = _io_out_bits_T_37 | _io_out_bits_T_23; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_39 = _io_out_bits_T_38 | _io_out_bits_T_24; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_40 = _io_out_bits_T_39 | _io_out_bits_T_25; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_41 = _io_out_bits_T_40 | _io_out_bits_T_26; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_42 = _io_out_bits_T_41 | _io_out_bits_T_27; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_43 = _io_out_bits_T_42 | _io_out_bits_T_28; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_44 = _io_out_bits_T_43 | _io_out_bits_T_29; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_45 = _io_out_bits_T_44 | _io_out_bits_T_30; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_47 = chosenOH[0] ? io_in_0_bits_data_clientStates_1 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_48 = chosenOH[1] ? io_in_1_bits_data_clientStates_1 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_49 = chosenOH[2] ? io_in_2_bits_data_clientStates_1 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_50 = chosenOH[3] ? io_in_3_bits_data_clientStates_1 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_51 = chosenOH[4] ? io_in_4_bits_data_clientStates_1 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_52 = chosenOH[5] ? io_in_5_bits_data_clientStates_1 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_53 = chosenOH[6] ? io_in_6_bits_data_clientStates_1 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_54 = chosenOH[7] ? io_in_7_bits_data_clientStates_1 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_55 = chosenOH[8] ? io_in_8_bits_data_clientStates_1 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_56 = chosenOH[9] ? io_in_9_bits_data_clientStates_1 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_57 = chosenOH[10] ? io_in_10_bits_data_clientStates_1 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_58 = chosenOH[11] ? io_in_11_bits_data_clientStates_1 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_59 = chosenOH[12] ? io_in_12_bits_data_clientStates_1 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_60 = chosenOH[13] ? io_in_13_bits_data_clientStates_1 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_61 = chosenOH[14] ? io_in_14_bits_data_clientStates_1 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_62 = chosenOH[15] ? io_in_15_bits_data_clientStates_1 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_63 = _io_out_bits_T_47 | _io_out_bits_T_48; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_64 = _io_out_bits_T_63 | _io_out_bits_T_49; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_65 = _io_out_bits_T_64 | _io_out_bits_T_50; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_66 = _io_out_bits_T_65 | _io_out_bits_T_51; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_67 = _io_out_bits_T_66 | _io_out_bits_T_52; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_68 = _io_out_bits_T_67 | _io_out_bits_T_53; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_69 = _io_out_bits_T_68 | _io_out_bits_T_54; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_70 = _io_out_bits_T_69 | _io_out_bits_T_55; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_71 = _io_out_bits_T_70 | _io_out_bits_T_56; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_72 = _io_out_bits_T_71 | _io_out_bits_T_57; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_73 = _io_out_bits_T_72 | _io_out_bits_T_58; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_74 = _io_out_bits_T_73 | _io_out_bits_T_59; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_75 = _io_out_bits_T_74 | _io_out_bits_T_60; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_76 = _io_out_bits_T_75 | _io_out_bits_T_61; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_78 = chosenOH[0] ? io_in_0_bits_data_state : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_79 = chosenOH[1] ? io_in_1_bits_data_state : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_80 = chosenOH[2] ? io_in_2_bits_data_state : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_81 = chosenOH[3] ? io_in_3_bits_data_state : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_82 = chosenOH[4] ? io_in_4_bits_data_state : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_83 = chosenOH[5] ? io_in_5_bits_data_state : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_84 = chosenOH[6] ? io_in_6_bits_data_state : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_85 = chosenOH[7] ? io_in_7_bits_data_state : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_86 = chosenOH[8] ? io_in_8_bits_data_state : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_87 = chosenOH[9] ? io_in_9_bits_data_state : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_88 = chosenOH[10] ? io_in_10_bits_data_state : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_89 = chosenOH[11] ? io_in_11_bits_data_state : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_90 = chosenOH[12] ? io_in_12_bits_data_state : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_91 = chosenOH[13] ? io_in_13_bits_data_state : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_92 = chosenOH[14] ? io_in_14_bits_data_state : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_93 = chosenOH[15] ? io_in_15_bits_data_state : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_94 = _io_out_bits_T_78 | _io_out_bits_T_79; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_95 = _io_out_bits_T_94 | _io_out_bits_T_80; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_96 = _io_out_bits_T_95 | _io_out_bits_T_81; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_97 = _io_out_bits_T_96 | _io_out_bits_T_82; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_98 = _io_out_bits_T_97 | _io_out_bits_T_83; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_99 = _io_out_bits_T_98 | _io_out_bits_T_84; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_100 = _io_out_bits_T_99 | _io_out_bits_T_85; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_101 = _io_out_bits_T_100 | _io_out_bits_T_86; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_102 = _io_out_bits_T_101 | _io_out_bits_T_87; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_103 = _io_out_bits_T_102 | _io_out_bits_T_88; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_104 = _io_out_bits_T_103 | _io_out_bits_T_89; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_105 = _io_out_bits_T_104 | _io_out_bits_T_90; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_106 = _io_out_bits_T_105 | _io_out_bits_T_91; // @[Mux.scala 27:73]
  wire [1:0] _io_out_bits_T_107 = _io_out_bits_T_106 | _io_out_bits_T_92; // @[Mux.scala 27:73]
  wire  _io_out_bits_T_124 = chosenOH[15] & io_in_15_bits_data_dirty; // @[Mux.scala 27:73]
  wire [2:0] _io_out_bits_T_140 = chosenOH[0] ? io_in_0_bits_way : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_out_bits_T_141 = chosenOH[1] ? io_in_1_bits_way : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_out_bits_T_142 = chosenOH[2] ? io_in_2_bits_way : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_out_bits_T_143 = chosenOH[3] ? io_in_3_bits_way : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_out_bits_T_144 = chosenOH[4] ? io_in_4_bits_way : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_out_bits_T_145 = chosenOH[5] ? io_in_5_bits_way : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_out_bits_T_146 = chosenOH[6] ? io_in_6_bits_way : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_out_bits_T_147 = chosenOH[7] ? io_in_7_bits_way : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_out_bits_T_148 = chosenOH[8] ? io_in_8_bits_way : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_out_bits_T_149 = chosenOH[9] ? io_in_9_bits_way : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_out_bits_T_150 = chosenOH[10] ? io_in_10_bits_way : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_out_bits_T_151 = chosenOH[11] ? io_in_11_bits_way : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_out_bits_T_152 = chosenOH[12] ? io_in_12_bits_way : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_out_bits_T_153 = chosenOH[13] ? io_in_13_bits_way : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_out_bits_T_154 = chosenOH[14] ? io_in_14_bits_way : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_out_bits_T_155 = chosenOH[15] ? io_in_15_bits_way : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_out_bits_T_156 = _io_out_bits_T_140 | _io_out_bits_T_141; // @[Mux.scala 27:73]
  wire [2:0] _io_out_bits_T_157 = _io_out_bits_T_156 | _io_out_bits_T_142; // @[Mux.scala 27:73]
  wire [2:0] _io_out_bits_T_158 = _io_out_bits_T_157 | _io_out_bits_T_143; // @[Mux.scala 27:73]
  wire [2:0] _io_out_bits_T_159 = _io_out_bits_T_158 | _io_out_bits_T_144; // @[Mux.scala 27:73]
  wire [2:0] _io_out_bits_T_160 = _io_out_bits_T_159 | _io_out_bits_T_145; // @[Mux.scala 27:73]
  wire [2:0] _io_out_bits_T_161 = _io_out_bits_T_160 | _io_out_bits_T_146; // @[Mux.scala 27:73]
  wire [2:0] _io_out_bits_T_162 = _io_out_bits_T_161 | _io_out_bits_T_147; // @[Mux.scala 27:73]
  wire [2:0] _io_out_bits_T_163 = _io_out_bits_T_162 | _io_out_bits_T_148; // @[Mux.scala 27:73]
  wire [2:0] _io_out_bits_T_164 = _io_out_bits_T_163 | _io_out_bits_T_149; // @[Mux.scala 27:73]
  wire [2:0] _io_out_bits_T_165 = _io_out_bits_T_164 | _io_out_bits_T_150; // @[Mux.scala 27:73]
  wire [2:0] _io_out_bits_T_166 = _io_out_bits_T_165 | _io_out_bits_T_151; // @[Mux.scala 27:73]
  wire [2:0] _io_out_bits_T_167 = _io_out_bits_T_166 | _io_out_bits_T_152; // @[Mux.scala 27:73]
  wire [2:0] _io_out_bits_T_168 = _io_out_bits_T_167 | _io_out_bits_T_153; // @[Mux.scala 27:73]
  wire [2:0] _io_out_bits_T_169 = _io_out_bits_T_168 | _io_out_bits_T_154; // @[Mux.scala 27:73]
  wire [9:0] _io_out_bits_T_171 = chosenOH[0] ? io_in_0_bits_set : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _io_out_bits_T_172 = chosenOH[1] ? io_in_1_bits_set : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _io_out_bits_T_173 = chosenOH[2] ? io_in_2_bits_set : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _io_out_bits_T_174 = chosenOH[3] ? io_in_3_bits_set : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _io_out_bits_T_175 = chosenOH[4] ? io_in_4_bits_set : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _io_out_bits_T_176 = chosenOH[5] ? io_in_5_bits_set : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _io_out_bits_T_177 = chosenOH[6] ? io_in_6_bits_set : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _io_out_bits_T_178 = chosenOH[7] ? io_in_7_bits_set : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _io_out_bits_T_179 = chosenOH[8] ? io_in_8_bits_set : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _io_out_bits_T_180 = chosenOH[9] ? io_in_9_bits_set : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _io_out_bits_T_181 = chosenOH[10] ? io_in_10_bits_set : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _io_out_bits_T_182 = chosenOH[11] ? io_in_11_bits_set : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _io_out_bits_T_183 = chosenOH[12] ? io_in_12_bits_set : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _io_out_bits_T_184 = chosenOH[13] ? io_in_13_bits_set : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _io_out_bits_T_185 = chosenOH[14] ? io_in_14_bits_set : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _io_out_bits_T_186 = chosenOH[15] ? io_in_15_bits_set : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _io_out_bits_T_187 = _io_out_bits_T_171 | _io_out_bits_T_172; // @[Mux.scala 27:73]
  wire [9:0] _io_out_bits_T_188 = _io_out_bits_T_187 | _io_out_bits_T_173; // @[Mux.scala 27:73]
  wire [9:0] _io_out_bits_T_189 = _io_out_bits_T_188 | _io_out_bits_T_174; // @[Mux.scala 27:73]
  wire [9:0] _io_out_bits_T_190 = _io_out_bits_T_189 | _io_out_bits_T_175; // @[Mux.scala 27:73]
  wire [9:0] _io_out_bits_T_191 = _io_out_bits_T_190 | _io_out_bits_T_176; // @[Mux.scala 27:73]
  wire [9:0] _io_out_bits_T_192 = _io_out_bits_T_191 | _io_out_bits_T_177; // @[Mux.scala 27:73]
  wire [9:0] _io_out_bits_T_193 = _io_out_bits_T_192 | _io_out_bits_T_178; // @[Mux.scala 27:73]
  wire [9:0] _io_out_bits_T_194 = _io_out_bits_T_193 | _io_out_bits_T_179; // @[Mux.scala 27:73]
  wire [9:0] _io_out_bits_T_195 = _io_out_bits_T_194 | _io_out_bits_T_180; // @[Mux.scala 27:73]
  wire [9:0] _io_out_bits_T_196 = _io_out_bits_T_195 | _io_out_bits_T_181; // @[Mux.scala 27:73]
  wire [9:0] _io_out_bits_T_197 = _io_out_bits_T_196 | _io_out_bits_T_182; // @[Mux.scala 27:73]
  wire [9:0] _io_out_bits_T_198 = _io_out_bits_T_197 | _io_out_bits_T_183; // @[Mux.scala 27:73]
  wire [9:0] _io_out_bits_T_199 = _io_out_bits_T_198 | _io_out_bits_T_184; // @[Mux.scala 27:73]
  wire [9:0] _io_out_bits_T_200 = _io_out_bits_T_199 | _io_out_bits_T_185; // @[Mux.scala 27:73]
  assign io_in_0_ready = chosenOH[0]; // @[FastArbiter.scala 59:42]
  assign io_in_1_ready = chosenOH[1]; // @[FastArbiter.scala 59:42]
  assign io_in_2_ready = chosenOH[2]; // @[FastArbiter.scala 59:42]
  assign io_in_3_ready = chosenOH[3]; // @[FastArbiter.scala 59:42]
  assign io_in_4_ready = chosenOH[4]; // @[FastArbiter.scala 59:42]
  assign io_in_5_ready = chosenOH[5]; // @[FastArbiter.scala 59:42]
  assign io_in_6_ready = chosenOH[6]; // @[FastArbiter.scala 59:42]
  assign io_in_7_ready = chosenOH[7]; // @[FastArbiter.scala 59:42]
  assign io_in_8_ready = chosenOH[8]; // @[FastArbiter.scala 59:42]
  assign io_in_9_ready = chosenOH[9]; // @[FastArbiter.scala 59:42]
  assign io_in_10_ready = chosenOH[10]; // @[FastArbiter.scala 59:42]
  assign io_in_11_ready = chosenOH[11]; // @[FastArbiter.scala 59:42]
  assign io_in_12_ready = chosenOH[12]; // @[FastArbiter.scala 59:42]
  assign io_in_13_ready = chosenOH[13]; // @[FastArbiter.scala 59:42]
  assign io_in_14_ready = chosenOH[14]; // @[FastArbiter.scala 59:42]
  assign io_in_15_ready = chosenOH[15]; // @[FastArbiter.scala 59:42]
  assign io_out_valid = |valids; // @[FastArbiter.scala 56:29]
  assign io_out_bits_set = _io_out_bits_T_200 | _io_out_bits_T_186; // @[Mux.scala 27:73]
  assign io_out_bits_way = _io_out_bits_T_169 | _io_out_bits_T_155; // @[Mux.scala 27:73]
  assign io_out_bits_data_dirty = chosenOH[0] & io_in_0_bits_data_dirty | chosenOH[1] & io_in_1_bits_data_dirty |
    chosenOH[2] & io_in_2_bits_data_dirty | chosenOH[3] & io_in_3_bits_data_dirty | chosenOH[4] &
    io_in_4_bits_data_dirty | chosenOH[5] & io_in_5_bits_data_dirty | chosenOH[6] & io_in_6_bits_data_dirty | chosenOH[7
    ] & io_in_7_bits_data_dirty | chosenOH[8] & io_in_8_bits_data_dirty | chosenOH[9] & io_in_9_bits_data_dirty |
    chosenOH[10] & io_in_10_bits_data_dirty | chosenOH[11] & io_in_11_bits_data_dirty | chosenOH[12] &
    io_in_12_bits_data_dirty | chosenOH[13] & io_in_13_bits_data_dirty | chosenOH[14] & io_in_14_bits_data_dirty |
    _io_out_bits_T_124; // @[Mux.scala 27:73]
  assign io_out_bits_data_state = _io_out_bits_T_107 | _io_out_bits_T_93; // @[Mux.scala 27:73]
  assign io_out_bits_data_clientStates_0 = _io_out_bits_T_45 | _io_out_bits_T_31; // @[Mux.scala 27:73]
  assign io_out_bits_data_clientStates_1 = _io_out_bits_T_76 | _io_out_bits_T_62; // @[Mux.scala 27:73]
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      rrGrantMask <= 16'h0; // @[Reg.scala 29:22]
    end else if (io_out_valid) begin // @[Reg.scala 28:20]
      rrGrantMask <= _rrGrantMask_T_30;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      pendingMask <= 16'h0; // @[Reg.scala 29:22]
    end else if (io_out_valid) begin // @[Reg.scala 28:20]
      pendingMask <= _pendingMask_T_1;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  rrGrantMask = _RAND_0[15:0];
  _RAND_1 = {1{`RANDOM}};
  pendingMask = _RAND_1[15:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    rrGrantMask = 16'h0;
  end
  if (reset) begin
    pendingMask = 16'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule

