module ICacheReplacePipe(
  input          clock,
  input          reset,
  output         io_pipe_req_ready,
  input          io_pipe_req_valid,
  input  [35:0]  io_pipe_req_bits_paddr,
  input  [38:0]  io_pipe_req_bits_vaddr,
  input  [2:0]   io_pipe_req_bits_param,
  input          io_pipe_req_bits_voluntary,
  input          io_pipe_req_bits_needData,
  input  [7:0]   io_pipe_req_bits_waymask,
  input  [4:0]   io_pipe_req_bits_id,
  input          io_meta_read_ready,
  output         io_meta_read_valid,
  output [5:0]   io_meta_read_bits_vSetIdx_0,
  input          io_data_read_ready,
  output         io_data_read_valid,
  output [5:0]   io_data_read_bits_0_vSetIdx_0,
  output [5:0]   io_data_read_bits_1_vSetIdx_0,
  output [5:0]   io_data_read_bits_2_vSetIdx_0,
  output [5:0]   io_data_read_bits_3_vSetIdx_0,
  output         io_error_source_tag,
  output         io_error_source_data,
  output         io_error_opType_probe,
  output         io_error_opType_release,
  output [35:0]  io_error_paddr,
  output         io_error_report_to_beu,
  output         io_error_valid,
  input  [1:0]   io_meta_response_metaData_0_0_coh_state,
  input  [23:0]  io_meta_response_metaData_0_0_tag,
  input  [1:0]   io_meta_response_metaData_0_1_coh_state,
  input  [23:0]  io_meta_response_metaData_0_1_tag,
  input  [1:0]   io_meta_response_metaData_0_2_coh_state,
  input  [23:0]  io_meta_response_metaData_0_2_tag,
  input  [1:0]   io_meta_response_metaData_0_3_coh_state,
  input  [23:0]  io_meta_response_metaData_0_3_tag,
  input  [1:0]   io_meta_response_metaData_0_4_coh_state,
  input  [23:0]  io_meta_response_metaData_0_4_tag,
  input  [1:0]   io_meta_response_metaData_0_5_coh_state,
  input  [23:0]  io_meta_response_metaData_0_5_tag,
  input  [1:0]   io_meta_response_metaData_0_6_coh_state,
  input  [23:0]  io_meta_response_metaData_0_6_tag,
  input  [1:0]   io_meta_response_metaData_0_7_coh_state,
  input  [23:0]  io_meta_response_metaData_0_7_tag,
  input          io_meta_response_errors_0_0,
  input          io_meta_response_errors_0_1,
  input          io_meta_response_errors_0_2,
  input          io_meta_response_errors_0_3,
  input          io_meta_response_errors_0_4,
  input          io_meta_response_errors_0_5,
  input          io_meta_response_errors_0_6,
  input          io_meta_response_errors_0_7,
  input  [511:0] io_data_response_datas_0_0,
  input  [511:0] io_data_response_datas_0_1,
  input  [511:0] io_data_response_datas_0_2,
  input  [511:0] io_data_response_datas_0_3,
  input  [511:0] io_data_response_datas_0_4,
  input  [511:0] io_data_response_datas_0_5,
  input  [511:0] io_data_response_datas_0_6,
  input  [511:0] io_data_response_datas_0_7,
  input  [31:0]  io_data_response_codes_0_0,
  input  [31:0]  io_data_response_codes_0_1,
  input  [31:0]  io_data_response_codes_0_2,
  input  [31:0]  io_data_response_codes_0_3,
  input  [31:0]  io_data_response_codes_0_4,
  input  [31:0]  io_data_response_codes_0_5,
  input  [31:0]  io_data_response_codes_0_6,
  input  [31:0]  io_data_response_codes_0_7,
  output         io_meta_write_valid,
  output [5:0]   io_meta_write_bits_virIdx,
  output [23:0]  io_meta_write_bits_phyTag,
  output [1:0]   io_meta_write_bits_coh_state,
  output [7:0]   io_meta_write_bits_waymask,
  output         io_meta_write_bits_bankIdx,
  input          io_release_req_ready,
  output         io_release_req_valid,
  output [35:0]  io_release_req_bits_addr,
  output [2:0]   io_release_req_bits_param,
  output         io_release_req_bits_voluntary,
  output         io_release_req_bits_hasData,
  output         io_release_req_bits_dirty,
  output [511:0] io_release_req_bits_data,
  input          io_release_finish,
  output         io_pipe_resp_valid,
  output [4:0]   io_pipe_resp_bits,
  output         io_status_r0_set_valid,
  output [5:0]   io_status_r0_set_bits,
  output         io_status_r1_set_valid,
  output [5:0]   io_status_r1_set_bits,
  output         io_status_r2_set_valid,
  output [5:0]   io_status_r2_set_bits,
  output         io_status_r3_set_valid,
  output [5:0]   io_status_r3_set_bits,
  input          io_csr_parity_enable
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [511:0] _RAND_45;
  reg [511:0] _RAND_46;
  reg [511:0] _RAND_47;
  reg [511:0] _RAND_48;
  reg [511:0] _RAND_49;
  reg [511:0] _RAND_50;
  reg [511:0] _RAND_51;
  reg [511:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [63:0] _RAND_62;
  reg [63:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [511:0] _RAND_69;
  reg [511:0] _RAND_70;
  reg [511:0] _RAND_71;
  reg [511:0] _RAND_72;
  reg [511:0] _RAND_73;
  reg [511:0] _RAND_74;
  reg [511:0] _RAND_75;
  reg [511:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [63:0] _RAND_382;
  reg [63:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [63:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [63:0] _RAND_396;
  reg [31:0] _RAND_397;
`endif // RANDOMIZE_REG_INIT
  wire  _r0_valid_T = io_pipe_req_ready & io_pipe_req_valid; // @[Decoupled.scala 50:35]
  reg  r0_valid; // @[ICache.scala 98:25]
  wire  _r0_ready_T = io_meta_read_ready & io_data_read_ready; // @[ReplacePipe.scala 91:34]
  reg  r2_valid; // @[ICache.scala 98:25]
  wire  _r2_ready_T = r2_valid & io_release_req_ready; // @[ReplacePipe.scala 157:29]
  wire  r2_ready = r2_valid & io_release_req_ready | ~r2_valid; // @[ReplacePipe.scala 157:54]
  reg  r1_valid; // @[ICache.scala 98:25]
  wire  r1_ready = r2_ready | ~r1_valid; // @[ReplacePipe.scala 118:25]
  wire  r0_ready = io_meta_read_ready & io_data_read_ready & r1_ready | ~r0_valid; // @[ReplacePipe.scala 91:69]
  wire  r0_fire = r0_valid & r0_ready; // @[ReplacePipe.scala 92:24]
  wire  _GEN_0 = r0_fire ? 1'h0 : r0_valid; // @[ICache.scala 101:{43,51} 98:25]
  reg [35:0] r0_req_paddr; // @[Reg.scala 16:16]
  reg [38:0] r0_req_vaddr; // @[Reg.scala 16:16]
  reg [2:0] r0_req_param; // @[Reg.scala 16:16]
  reg  r0_req_voluntary; // @[Reg.scala 16:16]
  reg  r0_req_needData; // @[Reg.scala 16:16]
  reg [7:0] r0_req_waymask; // @[Reg.scala 16:16]
  reg [4:0] r0_req_id; // @[Reg.scala 16:16]
  wire  r1_fire = r1_valid & r2_ready; // @[ReplacePipe.scala 119:24]
  wire  _GEN_10 = r1_fire ? 1'h0 : r1_valid; // @[ICache.scala 101:{43,51} 98:25]
  reg [35:0] r1_req_paddr; // @[Reg.scala 16:16]
  reg [38:0] r1_req_vaddr; // @[Reg.scala 16:16]
  reg [2:0] r1_req_param; // @[Reg.scala 16:16]
  reg  r1_req_voluntary; // @[Reg.scala 16:16]
  reg  r1_req_needData; // @[Reg.scala 16:16]
  reg [7:0] r1_req_waymask; // @[Reg.scala 16:16]
  reg [4:0] r1_req_id; // @[Reg.scala 16:16]
  reg  r1_meta_ptags_REG; // @[ReplacePipe.scala 124:113]
  reg [23:0] r1_meta_ptags_r0; // @[Reg.scala 16:16]
  reg [23:0] r1_meta_ptags_r1; // @[Reg.scala 16:16]
  reg [23:0] r1_meta_ptags_r2; // @[Reg.scala 16:16]
  reg [23:0] r1_meta_ptags_r3; // @[Reg.scala 16:16]
  reg [23:0] r1_meta_ptags_r4; // @[Reg.scala 16:16]
  reg [23:0] r1_meta_ptags_r5; // @[Reg.scala 16:16]
  reg [23:0] r1_meta_ptags_r6; // @[Reg.scala 16:16]
  reg [23:0] r1_meta_ptags_r7; // @[Reg.scala 16:16]
  wire [23:0] _GEN_20 = r1_meta_ptags_REG ? io_meta_response_metaData_0_0_tag : r1_meta_ptags_r0; // @[Reg.scala 16:16 17:{18,22}]
  wire [23:0] _GEN_21 = r1_meta_ptags_REG ? io_meta_response_metaData_0_1_tag : r1_meta_ptags_r1; // @[Reg.scala 16:16 17:{18,22}]
  wire [23:0] _GEN_22 = r1_meta_ptags_REG ? io_meta_response_metaData_0_2_tag : r1_meta_ptags_r2; // @[Reg.scala 16:16 17:{18,22}]
  wire [23:0] _GEN_23 = r1_meta_ptags_REG ? io_meta_response_metaData_0_3_tag : r1_meta_ptags_r3; // @[Reg.scala 16:16 17:{18,22}]
  wire [23:0] _GEN_24 = r1_meta_ptags_REG ? io_meta_response_metaData_0_4_tag : r1_meta_ptags_r4; // @[Reg.scala 16:16 17:{18,22}]
  wire [23:0] _GEN_25 = r1_meta_ptags_REG ? io_meta_response_metaData_0_5_tag : r1_meta_ptags_r5; // @[Reg.scala 16:16 17:{18,22}]
  wire [23:0] _GEN_26 = r1_meta_ptags_REG ? io_meta_response_metaData_0_6_tag : r1_meta_ptags_r6; // @[Reg.scala 16:16 17:{18,22}]
  wire [23:0] _GEN_27 = r1_meta_ptags_REG ? io_meta_response_metaData_0_7_tag : r1_meta_ptags_r7; // @[Reg.scala 16:16 17:{18,22}]
  reg  r1_meta_cohs_REG; // @[ReplacePipe.scala 125:113]
  reg [1:0] r1_meta_cohs_r0_state; // @[Reg.scala 16:16]
  reg [1:0] r1_meta_cohs_r1_state; // @[Reg.scala 16:16]
  reg [1:0] r1_meta_cohs_r2_state; // @[Reg.scala 16:16]
  reg [1:0] r1_meta_cohs_r3_state; // @[Reg.scala 16:16]
  reg [1:0] r1_meta_cohs_r4_state; // @[Reg.scala 16:16]
  reg [1:0] r1_meta_cohs_r5_state; // @[Reg.scala 16:16]
  reg [1:0] r1_meta_cohs_r6_state; // @[Reg.scala 16:16]
  reg [1:0] r1_meta_cohs_r7_state; // @[Reg.scala 16:16]
  wire [1:0] _GEN_28 = r1_meta_cohs_REG ? io_meta_response_metaData_0_0_coh_state : r1_meta_cohs_r0_state; // @[Reg.scala 16:16 17:{18,22}]
  wire [1:0] _GEN_29 = r1_meta_cohs_REG ? io_meta_response_metaData_0_1_coh_state : r1_meta_cohs_r1_state; // @[Reg.scala 16:16 17:{18,22}]
  wire [1:0] _GEN_30 = r1_meta_cohs_REG ? io_meta_response_metaData_0_2_coh_state : r1_meta_cohs_r2_state; // @[Reg.scala 16:16 17:{18,22}]
  wire [1:0] _GEN_31 = r1_meta_cohs_REG ? io_meta_response_metaData_0_3_coh_state : r1_meta_cohs_r3_state; // @[Reg.scala 16:16 17:{18,22}]
  wire [1:0] _GEN_32 = r1_meta_cohs_REG ? io_meta_response_metaData_0_4_coh_state : r1_meta_cohs_r4_state; // @[Reg.scala 16:16 17:{18,22}]
  wire [1:0] _GEN_33 = r1_meta_cohs_REG ? io_meta_response_metaData_0_5_coh_state : r1_meta_cohs_r5_state; // @[Reg.scala 16:16 17:{18,22}]
  wire [1:0] _GEN_34 = r1_meta_cohs_REG ? io_meta_response_metaData_0_6_coh_state : r1_meta_cohs_r6_state; // @[Reg.scala 16:16 17:{18,22}]
  wire [1:0] _GEN_35 = r1_meta_cohs_REG ? io_meta_response_metaData_0_7_coh_state : r1_meta_cohs_r7_state; // @[Reg.scala 16:16 17:{18,22}]
  reg  r1_meta_errors_REG; // @[ReplacePipe.scala 126:86]
  reg  r1_meta_errors_r0; // @[Reg.scala 16:16]
  reg  r1_meta_errors_r1; // @[Reg.scala 16:16]
  reg  r1_meta_errors_r2; // @[Reg.scala 16:16]
  reg  r1_meta_errors_r3; // @[Reg.scala 16:16]
  reg  r1_meta_errors_r4; // @[Reg.scala 16:16]
  reg  r1_meta_errors_r5; // @[Reg.scala 16:16]
  reg  r1_meta_errors_r6; // @[Reg.scala 16:16]
  reg  r1_meta_errors_r7; // @[Reg.scala 16:16]
  reg  r1_data_cacheline_REG; // @[ReplacePipe.scala 128:109]
  reg [511:0] r1_data_cacheline_r0; // @[Reg.scala 16:16]
  reg [511:0] r1_data_cacheline_r1; // @[Reg.scala 16:16]
  reg [511:0] r1_data_cacheline_r2; // @[Reg.scala 16:16]
  reg [511:0] r1_data_cacheline_r3; // @[Reg.scala 16:16]
  reg [511:0] r1_data_cacheline_r4; // @[Reg.scala 16:16]
  reg [511:0] r1_data_cacheline_r5; // @[Reg.scala 16:16]
  reg [511:0] r1_data_cacheline_r6; // @[Reg.scala 16:16]
  reg [511:0] r1_data_cacheline_r7; // @[Reg.scala 16:16]
  reg  r1_data_errorBits_REG; // @[ReplacePipe.scala 129:110]
  reg [31:0] r1_data_errorBits_r0; // @[Reg.scala 16:16]
  reg [31:0] r1_data_errorBits_r1; // @[Reg.scala 16:16]
  reg [31:0] r1_data_errorBits_r2; // @[Reg.scala 16:16]
  reg [31:0] r1_data_errorBits_r3; // @[Reg.scala 16:16]
  reg [31:0] r1_data_errorBits_r4; // @[Reg.scala 16:16]
  reg [31:0] r1_data_errorBits_r5; // @[Reg.scala 16:16]
  reg [31:0] r1_data_errorBits_r6; // @[Reg.scala 16:16]
  reg [31:0] r1_data_errorBits_r7; // @[Reg.scala 16:16]
  wire [23:0] probe_phy_tag = r1_req_paddr[35:12]; // @[L1Cache.scala 79:41]
  wire  _probe_hit_vec_T_1 = _GEN_28 > 2'h0; // @[Metadata.scala 49:45]
  wire  probe_hit_vec_0 = _GEN_20 == probe_phy_tag & _probe_hit_vec_T_1; // @[ReplacePipe.scala 134:120]
  wire  _probe_hit_vec_T_4 = _GEN_29 > 2'h0; // @[Metadata.scala 49:45]
  wire  probe_hit_vec_1 = _GEN_21 == probe_phy_tag & _probe_hit_vec_T_4; // @[ReplacePipe.scala 134:120]
  wire  _probe_hit_vec_T_7 = _GEN_30 > 2'h0; // @[Metadata.scala 49:45]
  wire  probe_hit_vec_2 = _GEN_22 == probe_phy_tag & _probe_hit_vec_T_7; // @[ReplacePipe.scala 134:120]
  wire  _probe_hit_vec_T_10 = _GEN_31 > 2'h0; // @[Metadata.scala 49:45]
  wire  probe_hit_vec_3 = _GEN_23 == probe_phy_tag & _probe_hit_vec_T_10; // @[ReplacePipe.scala 134:120]
  wire  _probe_hit_vec_T_13 = _GEN_32 > 2'h0; // @[Metadata.scala 49:45]
  wire  probe_hit_vec_4 = _GEN_24 == probe_phy_tag & _probe_hit_vec_T_13; // @[ReplacePipe.scala 134:120]
  wire  _probe_hit_vec_T_16 = _GEN_33 > 2'h0; // @[Metadata.scala 49:45]
  wire  probe_hit_vec_5 = _GEN_25 == probe_phy_tag & _probe_hit_vec_T_16; // @[ReplacePipe.scala 134:120]
  wire  _probe_hit_vec_T_19 = _GEN_34 > 2'h0; // @[Metadata.scala 49:45]
  wire  probe_hit_vec_6 = _GEN_26 == probe_phy_tag & _probe_hit_vec_T_19; // @[ReplacePipe.scala 134:120]
  wire  _probe_hit_vec_T_22 = _GEN_35 > 2'h0; // @[Metadata.scala 49:45]
  wire  probe_hit_vec_7 = _GEN_27 == probe_phy_tag & _probe_hit_vec_T_22; // @[ReplacePipe.scala 134:120]
  wire [1:0] _probe_hit_coh_T = probe_hit_vec_0 ? _GEN_28 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _probe_hit_coh_T_1 = probe_hit_vec_1 ? _GEN_29 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _probe_hit_coh_T_2 = probe_hit_vec_2 ? _GEN_30 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _probe_hit_coh_T_3 = probe_hit_vec_3 ? _GEN_31 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _probe_hit_coh_T_4 = probe_hit_vec_4 ? _GEN_32 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _probe_hit_coh_T_5 = probe_hit_vec_5 ? _GEN_33 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _probe_hit_coh_T_6 = probe_hit_vec_6 ? _GEN_34 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _probe_hit_coh_T_7 = probe_hit_vec_7 ? _GEN_35 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _probe_hit_coh_T_8 = _probe_hit_coh_T | _probe_hit_coh_T_1; // @[Mux.scala 27:73]
  wire [1:0] _probe_hit_coh_T_9 = _probe_hit_coh_T_8 | _probe_hit_coh_T_2; // @[Mux.scala 27:73]
  wire [1:0] _probe_hit_coh_T_10 = _probe_hit_coh_T_9 | _probe_hit_coh_T_3; // @[Mux.scala 27:73]
  wire [1:0] _probe_hit_coh_T_11 = _probe_hit_coh_T_10 | _probe_hit_coh_T_4; // @[Mux.scala 27:73]
  wire [1:0] _probe_hit_coh_T_12 = _probe_hit_coh_T_11 | _probe_hit_coh_T_5; // @[Mux.scala 27:73]
  wire [1:0] _probe_hit_coh_T_13 = _probe_hit_coh_T_12 | _probe_hit_coh_T_6; // @[Mux.scala 27:73]
  wire [1:0] probe_hit_coh_state = _probe_hit_coh_T_13 | _probe_hit_coh_T_7; // @[Mux.scala 27:73]
  wire [23:0] _T_8 = r1_req_waymask[0] ? _GEN_20 : 24'h0; // @[Mux.scala 27:73]
  wire [23:0] _T_9 = r1_req_waymask[1] ? _GEN_21 : 24'h0; // @[Mux.scala 27:73]
  wire [23:0] _T_10 = r1_req_waymask[2] ? _GEN_22 : 24'h0; // @[Mux.scala 27:73]
  wire [23:0] _T_11 = r1_req_waymask[3] ? _GEN_23 : 24'h0; // @[Mux.scala 27:73]
  wire [23:0] _T_12 = r1_req_waymask[4] ? _GEN_24 : 24'h0; // @[Mux.scala 27:73]
  wire [23:0] _T_13 = r1_req_waymask[5] ? _GEN_25 : 24'h0; // @[Mux.scala 27:73]
  wire [23:0] _T_14 = r1_req_waymask[6] ? _GEN_26 : 24'h0; // @[Mux.scala 27:73]
  wire [23:0] _T_15 = r1_req_waymask[7] ? _GEN_27 : 24'h0; // @[Mux.scala 27:73]
  wire [23:0] _T_16 = _T_8 | _T_9; // @[Mux.scala 27:73]
  wire [23:0] _T_17 = _T_16 | _T_10; // @[Mux.scala 27:73]
  wire [23:0] _T_18 = _T_17 | _T_11; // @[Mux.scala 27:73]
  wire [23:0] _T_19 = _T_18 | _T_12; // @[Mux.scala 27:73]
  wire [23:0] _T_20 = _T_19 | _T_13; // @[Mux.scala 27:73]
  wire [23:0] _T_21 = _T_20 | _T_14; // @[Mux.scala 27:73]
  wire [23:0] release_tag = _T_21 | _T_15; // @[Mux.scala 27:73]
  wire [1:0] _T_31 = r1_req_waymask[0] ? _GEN_28 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _T_32 = r1_req_waymask[1] ? _GEN_29 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _T_33 = r1_req_waymask[2] ? _GEN_30 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _T_34 = r1_req_waymask[3] ? _GEN_31 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _T_35 = r1_req_waymask[4] ? _GEN_32 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _T_36 = r1_req_waymask[5] ? _GEN_33 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _T_37 = r1_req_waymask[6] ? _GEN_34 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _T_38 = r1_req_waymask[7] ? _GEN_35 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _T_39 = _T_31 | _T_32; // @[Mux.scala 27:73]
  wire [1:0] _T_40 = _T_39 | _T_33; // @[Mux.scala 27:73]
  wire [1:0] _T_41 = _T_40 | _T_34; // @[Mux.scala 27:73]
  wire [1:0] _T_42 = _T_41 | _T_35; // @[Mux.scala 27:73]
  wire [1:0] _T_43 = _T_42 | _T_36; // @[Mux.scala 27:73]
  wire [1:0] _T_44 = _T_43 | _T_37; // @[Mux.scala 27:73]
  wire [1:0] release_coh_state = _T_44 | _T_38; // @[Mux.scala 27:73]
  wire [35:0] _release_addr_T_1 = {release_tag,r1_req_vaddr[11:0]}; // @[Cat.scala 31:58]
  wire [35:0] release_addr = {_release_addr_T_1[35:6], 6'h0}; // @[L1Cache.scala 84:59]
  wire  _GEN_60 = _r2_ready_T ? 1'h0 : r2_valid; // @[ICache.scala 101:{43,51} 98:25]
  reg [35:0] r2_req_paddr; // @[Reg.scala 16:16]
  reg [38:0] r2_req_vaddr; // @[Reg.scala 16:16]
  reg [2:0] r2_req_param; // @[Reg.scala 16:16]
  reg  r2_req_voluntary; // @[Reg.scala 16:16]
  reg  r2_req_needData; // @[Reg.scala 16:16]
  reg [7:0] r2_req_waymask; // @[Reg.scala 16:16]
  reg [4:0] r2_req_id; // @[Reg.scala 16:16]
  reg [511:0] r2_data_cacheline_0; // @[Reg.scala 16:16]
  reg [511:0] r2_data_cacheline_1; // @[Reg.scala 16:16]
  reg [511:0] r2_data_cacheline_2; // @[Reg.scala 16:16]
  reg [511:0] r2_data_cacheline_3; // @[Reg.scala 16:16]
  reg [511:0] r2_data_cacheline_4; // @[Reg.scala 16:16]
  reg [511:0] r2_data_cacheline_5; // @[Reg.scala 16:16]
  reg [511:0] r2_data_cacheline_6; // @[Reg.scala 16:16]
  reg [511:0] r2_data_cacheline_7; // @[Reg.scala 16:16]
  reg [23:0] r2_probe_hit_ptag; // @[Reg.scala 16:16]
  reg  r2_probe_hit_vec_0; // @[Reg.scala 16:16]
  reg  r2_probe_hit_vec_1; // @[Reg.scala 16:16]
  reg  r2_probe_hit_vec_2; // @[Reg.scala 16:16]
  reg  r2_probe_hit_vec_3; // @[Reg.scala 16:16]
  reg  r2_probe_hit_vec_4; // @[Reg.scala 16:16]
  reg  r2_probe_hit_vec_5; // @[Reg.scala 16:16]
  reg  r2_probe_hit_vec_6; // @[Reg.scala 16:16]
  reg  r2_probe_hit_vec_7; // @[Reg.scala 16:16]
  reg [1:0] r2_probe_hit_coh_state; // @[Reg.scala 16:16]
  wire [511:0] _r2_probe_hit_data_T = r2_probe_hit_vec_0 ? r2_data_cacheline_0 : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _r2_probe_hit_data_T_1 = r2_probe_hit_vec_1 ? r2_data_cacheline_1 : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _r2_probe_hit_data_T_2 = r2_probe_hit_vec_2 ? r2_data_cacheline_2 : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _r2_probe_hit_data_T_3 = r2_probe_hit_vec_3 ? r2_data_cacheline_3 : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _r2_probe_hit_data_T_4 = r2_probe_hit_vec_4 ? r2_data_cacheline_4 : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _r2_probe_hit_data_T_5 = r2_probe_hit_vec_5 ? r2_data_cacheline_5 : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _r2_probe_hit_data_T_6 = r2_probe_hit_vec_6 ? r2_data_cacheline_6 : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _r2_probe_hit_data_T_7 = r2_probe_hit_vec_7 ? r2_data_cacheline_7 : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _r2_probe_hit_data_T_8 = _r2_probe_hit_data_T | _r2_probe_hit_data_T_1; // @[Mux.scala 27:73]
  wire [511:0] _r2_probe_hit_data_T_9 = _r2_probe_hit_data_T_8 | _r2_probe_hit_data_T_2; // @[Mux.scala 27:73]
  wire [511:0] _r2_probe_hit_data_T_10 = _r2_probe_hit_data_T_9 | _r2_probe_hit_data_T_3; // @[Mux.scala 27:73]
  wire [511:0] _r2_probe_hit_data_T_11 = _r2_probe_hit_data_T_10 | _r2_probe_hit_data_T_4; // @[Mux.scala 27:73]
  wire [511:0] _r2_probe_hit_data_T_12 = _r2_probe_hit_data_T_11 | _r2_probe_hit_data_T_5; // @[Mux.scala 27:73]
  wire [511:0] _r2_probe_hit_data_T_13 = _r2_probe_hit_data_T_12 | _r2_probe_hit_data_T_6; // @[Mux.scala 27:73]
  wire [511:0] r2_probe_hit_data = _r2_probe_hit_data_T_13 | _r2_probe_hit_data_T_7; // @[Mux.scala 27:73]
  wire [4:0] _T_67 = {r2_req_param,r2_probe_hit_coh_state}; // @[Cat.scala 31:58]
  wire  _T_80 = 5'h8 == _T_67; // @[Misc.scala 55:20]
  wire [2:0] _T_82 = _T_80 ? 3'h5 : 3'h0; // @[Misc.scala 37:36]
  wire  _T_84 = 5'h9 == _T_67; // @[Misc.scala 55:20]
  wire [2:0] _T_86 = _T_84 ? 3'h2 : _T_82; // @[Misc.scala 37:36]
  wire  _T_88 = 5'ha == _T_67; // @[Misc.scala 55:20]
  wire [2:0] _T_90 = _T_88 ? 3'h1 : _T_86; // @[Misc.scala 37:36]
  wire  _T_92 = 5'hb == _T_67; // @[Misc.scala 55:20]
  wire [2:0] _T_94 = _T_92 ? 3'h1 : _T_90; // @[Misc.scala 37:36]
  wire  _T_96 = 5'h4 == _T_67; // @[Misc.scala 55:20]
  wire  _T_97 = _T_96 ? 1'h0 : _T_92; // @[Misc.scala 37:9]
  wire [2:0] _T_98 = _T_96 ? 3'h5 : _T_94; // @[Misc.scala 37:36]
  wire  _T_100 = 5'h5 == _T_67; // @[Misc.scala 55:20]
  wire  _T_101 = _T_100 ? 1'h0 : _T_97; // @[Misc.scala 37:9]
  wire [2:0] _T_102 = _T_100 ? 3'h4 : _T_98; // @[Misc.scala 37:36]
  wire [1:0] _T_103 = _T_100 ? 2'h1 : 2'h0; // @[Misc.scala 37:63]
  wire  _T_104 = 5'h6 == _T_67; // @[Misc.scala 55:20]
  wire  _T_105 = _T_104 ? 1'h0 : _T_101; // @[Misc.scala 37:9]
  wire [2:0] _T_106 = _T_104 ? 3'h0 : _T_102; // @[Misc.scala 37:36]
  wire [1:0] _T_107 = _T_104 ? 2'h1 : _T_103; // @[Misc.scala 37:63]
  wire  _T_108 = 5'h7 == _T_67; // @[Misc.scala 55:20]
  wire [2:0] _T_110 = _T_108 ? 3'h0 : _T_106; // @[Misc.scala 37:36]
  wire [1:0] _T_111 = _T_108 ? 2'h1 : _T_107; // @[Misc.scala 37:63]
  wire  _T_112 = 5'h0 == _T_67; // @[Misc.scala 55:20]
  wire  _T_113 = _T_112 ? 1'h0 : _T_108 | _T_105; // @[Misc.scala 37:9]
  wire [2:0] _T_114 = _T_112 ? 3'h5 : _T_110; // @[Misc.scala 37:36]
  wire [1:0] _T_115 = _T_112 ? 2'h0 : _T_111; // @[Misc.scala 37:63]
  wire  _T_116 = 5'h1 == _T_67; // @[Misc.scala 55:20]
  wire  _T_117 = _T_116 ? 1'h0 : _T_113; // @[Misc.scala 37:9]
  wire [2:0] _T_118 = _T_116 ? 3'h4 : _T_114; // @[Misc.scala 37:36]
  wire [1:0] _T_119 = _T_116 ? 2'h1 : _T_115; // @[Misc.scala 37:63]
  wire  _T_120 = 5'h2 == _T_67; // @[Misc.scala 55:20]
  wire  _T_121 = _T_120 ? 1'h0 : _T_117; // @[Misc.scala 37:9]
  wire [2:0] _T_122 = _T_120 ? 3'h3 : _T_118; // @[Misc.scala 37:36]
  wire [1:0] _T_123 = _T_120 ? 2'h2 : _T_119; // @[Misc.scala 37:63]
  wire  _T_124 = 5'h3 == _T_67; // @[Misc.scala 55:20]
  wire  probe_has_dirty_data = _T_124 | _T_121; // @[Misc.scala 37:9]
  wire [2:0] probe_shrink_param = _T_124 ? 3'h3 : _T_122; // @[Misc.scala 37:36]
  reg  r2_meta_errors_0; // @[Reg.scala 16:16]
  reg  r2_meta_errors_1; // @[Reg.scala 16:16]
  reg  r2_meta_errors_2; // @[Reg.scala 16:16]
  reg  r2_meta_errors_3; // @[Reg.scala 16:16]
  reg  r2_meta_errors_4; // @[Reg.scala 16:16]
  reg  r2_meta_errors_5; // @[Reg.scala 16:16]
  reg  r2_meta_errors_6; // @[Reg.scala 16:16]
  reg  r2_meta_errors_7; // @[Reg.scala 16:16]
  reg [31:0] r2_data_errorBits_0; // @[Reg.scala 16:16]
  reg [31:0] r2_data_errorBits_1; // @[Reg.scala 16:16]
  reg [31:0] r2_data_errorBits_2; // @[Reg.scala 16:16]
  reg [31:0] r2_data_errorBits_3; // @[Reg.scala 16:16]
  reg [31:0] r2_data_errorBits_4; // @[Reg.scala 16:16]
  reg [31:0] r2_data_errorBits_5; // @[Reg.scala 16:16]
  reg [31:0] r2_data_errorBits_6; // @[Reg.scala 16:16]
  reg [31:0] r2_data_errorBits_7; // @[Reg.scala 16:16]
  wire [4095:0] _read_datas_T = {r2_data_cacheline_7,r2_data_cacheline_6,r2_data_cacheline_5,r2_data_cacheline_4,
    r2_data_cacheline_3,r2_data_cacheline_2,r2_data_cacheline_1,r2_data_cacheline_0}; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_0_0 = _read_datas_T[15:0]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_0_1 = _read_datas_T[31:16]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_0_2 = _read_datas_T[47:32]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_0_3 = _read_datas_T[63:48]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_0_4 = _read_datas_T[79:64]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_0_5 = _read_datas_T[95:80]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_0_6 = _read_datas_T[111:96]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_0_7 = _read_datas_T[127:112]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_0_8 = _read_datas_T[143:128]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_0_9 = _read_datas_T[159:144]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_0_10 = _read_datas_T[175:160]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_0_11 = _read_datas_T[191:176]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_0_12 = _read_datas_T[207:192]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_0_13 = _read_datas_T[223:208]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_0_14 = _read_datas_T[239:224]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_0_15 = _read_datas_T[255:240]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_0_16 = _read_datas_T[271:256]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_0_17 = _read_datas_T[287:272]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_0_18 = _read_datas_T[303:288]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_0_19 = _read_datas_T[319:304]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_0_20 = _read_datas_T[335:320]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_0_21 = _read_datas_T[351:336]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_0_22 = _read_datas_T[367:352]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_0_23 = _read_datas_T[383:368]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_0_24 = _read_datas_T[399:384]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_0_25 = _read_datas_T[415:400]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_0_26 = _read_datas_T[431:416]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_0_27 = _read_datas_T[447:432]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_0_28 = _read_datas_T[463:448]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_0_29 = _read_datas_T[479:464]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_0_30 = _read_datas_T[495:480]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_0_31 = _read_datas_T[511:496]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_1_0 = _read_datas_T[527:512]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_1_1 = _read_datas_T[543:528]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_1_2 = _read_datas_T[559:544]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_1_3 = _read_datas_T[575:560]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_1_4 = _read_datas_T[591:576]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_1_5 = _read_datas_T[607:592]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_1_6 = _read_datas_T[623:608]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_1_7 = _read_datas_T[639:624]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_1_8 = _read_datas_T[655:640]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_1_9 = _read_datas_T[671:656]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_1_10 = _read_datas_T[687:672]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_1_11 = _read_datas_T[703:688]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_1_12 = _read_datas_T[719:704]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_1_13 = _read_datas_T[735:720]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_1_14 = _read_datas_T[751:736]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_1_15 = _read_datas_T[767:752]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_1_16 = _read_datas_T[783:768]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_1_17 = _read_datas_T[799:784]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_1_18 = _read_datas_T[815:800]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_1_19 = _read_datas_T[831:816]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_1_20 = _read_datas_T[847:832]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_1_21 = _read_datas_T[863:848]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_1_22 = _read_datas_T[879:864]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_1_23 = _read_datas_T[895:880]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_1_24 = _read_datas_T[911:896]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_1_25 = _read_datas_T[927:912]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_1_26 = _read_datas_T[943:928]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_1_27 = _read_datas_T[959:944]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_1_28 = _read_datas_T[975:960]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_1_29 = _read_datas_T[991:976]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_1_30 = _read_datas_T[1007:992]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_1_31 = _read_datas_T[1023:1008]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_2_0 = _read_datas_T[1039:1024]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_2_1 = _read_datas_T[1055:1040]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_2_2 = _read_datas_T[1071:1056]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_2_3 = _read_datas_T[1087:1072]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_2_4 = _read_datas_T[1103:1088]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_2_5 = _read_datas_T[1119:1104]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_2_6 = _read_datas_T[1135:1120]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_2_7 = _read_datas_T[1151:1136]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_2_8 = _read_datas_T[1167:1152]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_2_9 = _read_datas_T[1183:1168]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_2_10 = _read_datas_T[1199:1184]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_2_11 = _read_datas_T[1215:1200]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_2_12 = _read_datas_T[1231:1216]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_2_13 = _read_datas_T[1247:1232]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_2_14 = _read_datas_T[1263:1248]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_2_15 = _read_datas_T[1279:1264]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_2_16 = _read_datas_T[1295:1280]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_2_17 = _read_datas_T[1311:1296]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_2_18 = _read_datas_T[1327:1312]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_2_19 = _read_datas_T[1343:1328]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_2_20 = _read_datas_T[1359:1344]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_2_21 = _read_datas_T[1375:1360]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_2_22 = _read_datas_T[1391:1376]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_2_23 = _read_datas_T[1407:1392]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_2_24 = _read_datas_T[1423:1408]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_2_25 = _read_datas_T[1439:1424]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_2_26 = _read_datas_T[1455:1440]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_2_27 = _read_datas_T[1471:1456]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_2_28 = _read_datas_T[1487:1472]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_2_29 = _read_datas_T[1503:1488]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_2_30 = _read_datas_T[1519:1504]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_2_31 = _read_datas_T[1535:1520]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_3_0 = _read_datas_T[1551:1536]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_3_1 = _read_datas_T[1567:1552]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_3_2 = _read_datas_T[1583:1568]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_3_3 = _read_datas_T[1599:1584]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_3_4 = _read_datas_T[1615:1600]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_3_5 = _read_datas_T[1631:1616]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_3_6 = _read_datas_T[1647:1632]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_3_7 = _read_datas_T[1663:1648]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_3_8 = _read_datas_T[1679:1664]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_3_9 = _read_datas_T[1695:1680]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_3_10 = _read_datas_T[1711:1696]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_3_11 = _read_datas_T[1727:1712]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_3_12 = _read_datas_T[1743:1728]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_3_13 = _read_datas_T[1759:1744]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_3_14 = _read_datas_T[1775:1760]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_3_15 = _read_datas_T[1791:1776]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_3_16 = _read_datas_T[1807:1792]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_3_17 = _read_datas_T[1823:1808]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_3_18 = _read_datas_T[1839:1824]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_3_19 = _read_datas_T[1855:1840]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_3_20 = _read_datas_T[1871:1856]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_3_21 = _read_datas_T[1887:1872]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_3_22 = _read_datas_T[1903:1888]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_3_23 = _read_datas_T[1919:1904]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_3_24 = _read_datas_T[1935:1920]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_3_25 = _read_datas_T[1951:1936]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_3_26 = _read_datas_T[1967:1952]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_3_27 = _read_datas_T[1983:1968]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_3_28 = _read_datas_T[1999:1984]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_3_29 = _read_datas_T[2015:2000]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_3_30 = _read_datas_T[2031:2016]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_3_31 = _read_datas_T[2047:2032]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_4_0 = _read_datas_T[2063:2048]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_4_1 = _read_datas_T[2079:2064]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_4_2 = _read_datas_T[2095:2080]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_4_3 = _read_datas_T[2111:2096]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_4_4 = _read_datas_T[2127:2112]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_4_5 = _read_datas_T[2143:2128]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_4_6 = _read_datas_T[2159:2144]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_4_7 = _read_datas_T[2175:2160]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_4_8 = _read_datas_T[2191:2176]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_4_9 = _read_datas_T[2207:2192]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_4_10 = _read_datas_T[2223:2208]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_4_11 = _read_datas_T[2239:2224]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_4_12 = _read_datas_T[2255:2240]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_4_13 = _read_datas_T[2271:2256]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_4_14 = _read_datas_T[2287:2272]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_4_15 = _read_datas_T[2303:2288]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_4_16 = _read_datas_T[2319:2304]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_4_17 = _read_datas_T[2335:2320]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_4_18 = _read_datas_T[2351:2336]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_4_19 = _read_datas_T[2367:2352]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_4_20 = _read_datas_T[2383:2368]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_4_21 = _read_datas_T[2399:2384]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_4_22 = _read_datas_T[2415:2400]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_4_23 = _read_datas_T[2431:2416]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_4_24 = _read_datas_T[2447:2432]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_4_25 = _read_datas_T[2463:2448]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_4_26 = _read_datas_T[2479:2464]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_4_27 = _read_datas_T[2495:2480]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_4_28 = _read_datas_T[2511:2496]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_4_29 = _read_datas_T[2527:2512]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_4_30 = _read_datas_T[2543:2528]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_4_31 = _read_datas_T[2559:2544]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_5_0 = _read_datas_T[2575:2560]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_5_1 = _read_datas_T[2591:2576]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_5_2 = _read_datas_T[2607:2592]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_5_3 = _read_datas_T[2623:2608]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_5_4 = _read_datas_T[2639:2624]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_5_5 = _read_datas_T[2655:2640]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_5_6 = _read_datas_T[2671:2656]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_5_7 = _read_datas_T[2687:2672]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_5_8 = _read_datas_T[2703:2688]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_5_9 = _read_datas_T[2719:2704]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_5_10 = _read_datas_T[2735:2720]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_5_11 = _read_datas_T[2751:2736]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_5_12 = _read_datas_T[2767:2752]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_5_13 = _read_datas_T[2783:2768]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_5_14 = _read_datas_T[2799:2784]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_5_15 = _read_datas_T[2815:2800]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_5_16 = _read_datas_T[2831:2816]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_5_17 = _read_datas_T[2847:2832]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_5_18 = _read_datas_T[2863:2848]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_5_19 = _read_datas_T[2879:2864]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_5_20 = _read_datas_T[2895:2880]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_5_21 = _read_datas_T[2911:2896]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_5_22 = _read_datas_T[2927:2912]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_5_23 = _read_datas_T[2943:2928]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_5_24 = _read_datas_T[2959:2944]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_5_25 = _read_datas_T[2975:2960]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_5_26 = _read_datas_T[2991:2976]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_5_27 = _read_datas_T[3007:2992]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_5_28 = _read_datas_T[3023:3008]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_5_29 = _read_datas_T[3039:3024]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_5_30 = _read_datas_T[3055:3040]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_5_31 = _read_datas_T[3071:3056]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_6_0 = _read_datas_T[3087:3072]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_6_1 = _read_datas_T[3103:3088]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_6_2 = _read_datas_T[3119:3104]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_6_3 = _read_datas_T[3135:3120]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_6_4 = _read_datas_T[3151:3136]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_6_5 = _read_datas_T[3167:3152]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_6_6 = _read_datas_T[3183:3168]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_6_7 = _read_datas_T[3199:3184]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_6_8 = _read_datas_T[3215:3200]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_6_9 = _read_datas_T[3231:3216]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_6_10 = _read_datas_T[3247:3232]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_6_11 = _read_datas_T[3263:3248]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_6_12 = _read_datas_T[3279:3264]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_6_13 = _read_datas_T[3295:3280]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_6_14 = _read_datas_T[3311:3296]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_6_15 = _read_datas_T[3327:3312]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_6_16 = _read_datas_T[3343:3328]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_6_17 = _read_datas_T[3359:3344]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_6_18 = _read_datas_T[3375:3360]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_6_19 = _read_datas_T[3391:3376]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_6_20 = _read_datas_T[3407:3392]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_6_21 = _read_datas_T[3423:3408]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_6_22 = _read_datas_T[3439:3424]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_6_23 = _read_datas_T[3455:3440]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_6_24 = _read_datas_T[3471:3456]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_6_25 = _read_datas_T[3487:3472]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_6_26 = _read_datas_T[3503:3488]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_6_27 = _read_datas_T[3519:3504]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_6_28 = _read_datas_T[3535:3520]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_6_29 = _read_datas_T[3551:3536]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_6_30 = _read_datas_T[3567:3552]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_6_31 = _read_datas_T[3583:3568]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_7_0 = _read_datas_T[3599:3584]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_7_1 = _read_datas_T[3615:3600]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_7_2 = _read_datas_T[3631:3616]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_7_3 = _read_datas_T[3647:3632]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_7_4 = _read_datas_T[3663:3648]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_7_5 = _read_datas_T[3679:3664]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_7_6 = _read_datas_T[3695:3680]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_7_7 = _read_datas_T[3711:3696]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_7_8 = _read_datas_T[3727:3712]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_7_9 = _read_datas_T[3743:3728]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_7_10 = _read_datas_T[3759:3744]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_7_11 = _read_datas_T[3775:3760]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_7_12 = _read_datas_T[3791:3776]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_7_13 = _read_datas_T[3807:3792]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_7_14 = _read_datas_T[3823:3808]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_7_15 = _read_datas_T[3839:3824]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_7_16 = _read_datas_T[3855:3840]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_7_17 = _read_datas_T[3871:3856]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_7_18 = _read_datas_T[3887:3872]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_7_19 = _read_datas_T[3903:3888]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_7_20 = _read_datas_T[3919:3904]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_7_21 = _read_datas_T[3935:3920]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_7_22 = _read_datas_T[3951:3936]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_7_23 = _read_datas_T[3967:3952]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_7_24 = _read_datas_T[3983:3968]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_7_25 = _read_datas_T[3999:3984]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_7_26 = _read_datas_T[4015:4000]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_7_27 = _read_datas_T[4031:4016]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_7_28 = _read_datas_T[4047:4032]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_7_29 = _read_datas_T[4063:4048]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_7_30 = _read_datas_T[4079:4064]; // @[ReplacePipe.scala 178:46]
  wire [15:0] read_datas_7_31 = _read_datas_T[4095:4080]; // @[ReplacePipe.scala 178:46]
  wire [255:0] _read_codes_T = {r2_data_errorBits_7,r2_data_errorBits_6,r2_data_errorBits_5,r2_data_errorBits_4,
    r2_data_errorBits_3,r2_data_errorBits_2,r2_data_errorBits_1,r2_data_errorBits_0}; // @[ReplacePipe.scala 179:46]
  wire  read_codes_0_0 = _read_codes_T[0]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_0_1 = _read_codes_T[1]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_0_2 = _read_codes_T[2]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_0_3 = _read_codes_T[3]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_0_4 = _read_codes_T[4]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_0_5 = _read_codes_T[5]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_0_6 = _read_codes_T[6]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_0_7 = _read_codes_T[7]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_0_8 = _read_codes_T[8]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_0_9 = _read_codes_T[9]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_0_10 = _read_codes_T[10]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_0_11 = _read_codes_T[11]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_0_12 = _read_codes_T[12]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_0_13 = _read_codes_T[13]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_0_14 = _read_codes_T[14]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_0_15 = _read_codes_T[15]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_0_16 = _read_codes_T[16]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_0_17 = _read_codes_T[17]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_0_18 = _read_codes_T[18]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_0_19 = _read_codes_T[19]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_0_20 = _read_codes_T[20]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_0_21 = _read_codes_T[21]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_0_22 = _read_codes_T[22]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_0_23 = _read_codes_T[23]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_0_24 = _read_codes_T[24]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_0_25 = _read_codes_T[25]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_0_26 = _read_codes_T[26]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_0_27 = _read_codes_T[27]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_0_28 = _read_codes_T[28]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_0_29 = _read_codes_T[29]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_0_30 = _read_codes_T[30]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_0_31 = _read_codes_T[31]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_1_0 = _read_codes_T[32]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_1_1 = _read_codes_T[33]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_1_2 = _read_codes_T[34]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_1_3 = _read_codes_T[35]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_1_4 = _read_codes_T[36]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_1_5 = _read_codes_T[37]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_1_6 = _read_codes_T[38]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_1_7 = _read_codes_T[39]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_1_8 = _read_codes_T[40]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_1_9 = _read_codes_T[41]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_1_10 = _read_codes_T[42]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_1_11 = _read_codes_T[43]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_1_12 = _read_codes_T[44]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_1_13 = _read_codes_T[45]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_1_14 = _read_codes_T[46]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_1_15 = _read_codes_T[47]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_1_16 = _read_codes_T[48]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_1_17 = _read_codes_T[49]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_1_18 = _read_codes_T[50]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_1_19 = _read_codes_T[51]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_1_20 = _read_codes_T[52]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_1_21 = _read_codes_T[53]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_1_22 = _read_codes_T[54]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_1_23 = _read_codes_T[55]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_1_24 = _read_codes_T[56]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_1_25 = _read_codes_T[57]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_1_26 = _read_codes_T[58]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_1_27 = _read_codes_T[59]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_1_28 = _read_codes_T[60]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_1_29 = _read_codes_T[61]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_1_30 = _read_codes_T[62]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_1_31 = _read_codes_T[63]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_2_0 = _read_codes_T[64]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_2_1 = _read_codes_T[65]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_2_2 = _read_codes_T[66]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_2_3 = _read_codes_T[67]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_2_4 = _read_codes_T[68]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_2_5 = _read_codes_T[69]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_2_6 = _read_codes_T[70]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_2_7 = _read_codes_T[71]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_2_8 = _read_codes_T[72]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_2_9 = _read_codes_T[73]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_2_10 = _read_codes_T[74]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_2_11 = _read_codes_T[75]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_2_12 = _read_codes_T[76]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_2_13 = _read_codes_T[77]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_2_14 = _read_codes_T[78]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_2_15 = _read_codes_T[79]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_2_16 = _read_codes_T[80]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_2_17 = _read_codes_T[81]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_2_18 = _read_codes_T[82]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_2_19 = _read_codes_T[83]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_2_20 = _read_codes_T[84]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_2_21 = _read_codes_T[85]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_2_22 = _read_codes_T[86]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_2_23 = _read_codes_T[87]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_2_24 = _read_codes_T[88]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_2_25 = _read_codes_T[89]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_2_26 = _read_codes_T[90]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_2_27 = _read_codes_T[91]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_2_28 = _read_codes_T[92]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_2_29 = _read_codes_T[93]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_2_30 = _read_codes_T[94]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_2_31 = _read_codes_T[95]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_3_0 = _read_codes_T[96]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_3_1 = _read_codes_T[97]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_3_2 = _read_codes_T[98]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_3_3 = _read_codes_T[99]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_3_4 = _read_codes_T[100]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_3_5 = _read_codes_T[101]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_3_6 = _read_codes_T[102]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_3_7 = _read_codes_T[103]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_3_8 = _read_codes_T[104]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_3_9 = _read_codes_T[105]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_3_10 = _read_codes_T[106]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_3_11 = _read_codes_T[107]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_3_12 = _read_codes_T[108]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_3_13 = _read_codes_T[109]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_3_14 = _read_codes_T[110]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_3_15 = _read_codes_T[111]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_3_16 = _read_codes_T[112]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_3_17 = _read_codes_T[113]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_3_18 = _read_codes_T[114]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_3_19 = _read_codes_T[115]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_3_20 = _read_codes_T[116]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_3_21 = _read_codes_T[117]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_3_22 = _read_codes_T[118]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_3_23 = _read_codes_T[119]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_3_24 = _read_codes_T[120]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_3_25 = _read_codes_T[121]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_3_26 = _read_codes_T[122]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_3_27 = _read_codes_T[123]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_3_28 = _read_codes_T[124]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_3_29 = _read_codes_T[125]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_3_30 = _read_codes_T[126]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_3_31 = _read_codes_T[127]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_4_0 = _read_codes_T[128]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_4_1 = _read_codes_T[129]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_4_2 = _read_codes_T[130]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_4_3 = _read_codes_T[131]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_4_4 = _read_codes_T[132]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_4_5 = _read_codes_T[133]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_4_6 = _read_codes_T[134]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_4_7 = _read_codes_T[135]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_4_8 = _read_codes_T[136]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_4_9 = _read_codes_T[137]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_4_10 = _read_codes_T[138]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_4_11 = _read_codes_T[139]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_4_12 = _read_codes_T[140]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_4_13 = _read_codes_T[141]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_4_14 = _read_codes_T[142]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_4_15 = _read_codes_T[143]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_4_16 = _read_codes_T[144]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_4_17 = _read_codes_T[145]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_4_18 = _read_codes_T[146]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_4_19 = _read_codes_T[147]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_4_20 = _read_codes_T[148]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_4_21 = _read_codes_T[149]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_4_22 = _read_codes_T[150]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_4_23 = _read_codes_T[151]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_4_24 = _read_codes_T[152]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_4_25 = _read_codes_T[153]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_4_26 = _read_codes_T[154]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_4_27 = _read_codes_T[155]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_4_28 = _read_codes_T[156]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_4_29 = _read_codes_T[157]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_4_30 = _read_codes_T[158]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_4_31 = _read_codes_T[159]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_5_0 = _read_codes_T[160]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_5_1 = _read_codes_T[161]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_5_2 = _read_codes_T[162]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_5_3 = _read_codes_T[163]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_5_4 = _read_codes_T[164]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_5_5 = _read_codes_T[165]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_5_6 = _read_codes_T[166]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_5_7 = _read_codes_T[167]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_5_8 = _read_codes_T[168]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_5_9 = _read_codes_T[169]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_5_10 = _read_codes_T[170]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_5_11 = _read_codes_T[171]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_5_12 = _read_codes_T[172]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_5_13 = _read_codes_T[173]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_5_14 = _read_codes_T[174]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_5_15 = _read_codes_T[175]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_5_16 = _read_codes_T[176]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_5_17 = _read_codes_T[177]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_5_18 = _read_codes_T[178]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_5_19 = _read_codes_T[179]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_5_20 = _read_codes_T[180]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_5_21 = _read_codes_T[181]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_5_22 = _read_codes_T[182]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_5_23 = _read_codes_T[183]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_5_24 = _read_codes_T[184]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_5_25 = _read_codes_T[185]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_5_26 = _read_codes_T[186]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_5_27 = _read_codes_T[187]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_5_28 = _read_codes_T[188]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_5_29 = _read_codes_T[189]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_5_30 = _read_codes_T[190]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_5_31 = _read_codes_T[191]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_6_0 = _read_codes_T[192]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_6_1 = _read_codes_T[193]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_6_2 = _read_codes_T[194]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_6_3 = _read_codes_T[195]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_6_4 = _read_codes_T[196]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_6_5 = _read_codes_T[197]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_6_6 = _read_codes_T[198]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_6_7 = _read_codes_T[199]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_6_8 = _read_codes_T[200]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_6_9 = _read_codes_T[201]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_6_10 = _read_codes_T[202]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_6_11 = _read_codes_T[203]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_6_12 = _read_codes_T[204]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_6_13 = _read_codes_T[205]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_6_14 = _read_codes_T[206]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_6_15 = _read_codes_T[207]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_6_16 = _read_codes_T[208]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_6_17 = _read_codes_T[209]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_6_18 = _read_codes_T[210]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_6_19 = _read_codes_T[211]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_6_20 = _read_codes_T[212]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_6_21 = _read_codes_T[213]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_6_22 = _read_codes_T[214]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_6_23 = _read_codes_T[215]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_6_24 = _read_codes_T[216]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_6_25 = _read_codes_T[217]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_6_26 = _read_codes_T[218]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_6_27 = _read_codes_T[219]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_6_28 = _read_codes_T[220]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_6_29 = _read_codes_T[221]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_6_30 = _read_codes_T[222]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_6_31 = _read_codes_T[223]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_7_0 = _read_codes_T[224]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_7_1 = _read_codes_T[225]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_7_2 = _read_codes_T[226]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_7_3 = _read_codes_T[227]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_7_4 = _read_codes_T[228]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_7_5 = _read_codes_T[229]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_7_6 = _read_codes_T[230]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_7_7 = _read_codes_T[231]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_7_8 = _read_codes_T[232]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_7_9 = _read_codes_T[233]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_7_10 = _read_codes_T[234]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_7_11 = _read_codes_T[235]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_7_12 = _read_codes_T[236]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_7_13 = _read_codes_T[237]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_7_14 = _read_codes_T[238]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_7_15 = _read_codes_T[239]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_7_16 = _read_codes_T[240]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_7_17 = _read_codes_T[241]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_7_18 = _read_codes_T[242]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_7_19 = _read_codes_T[243]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_7_20 = _read_codes_T[244]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_7_21 = _read_codes_T[245]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_7_22 = _read_codes_T[246]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_7_23 = _read_codes_T[247]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_7_24 = _read_codes_T[248]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_7_25 = _read_codes_T[249]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_7_26 = _read_codes_T[250]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_7_27 = _read_codes_T[251]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_7_28 = _read_codes_T[252]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_7_29 = _read_codes_T[253]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_7_30 = _read_codes_T[254]; // @[ReplacePipe.scala 179:46]
  wire  read_codes_7_31 = _read_codes_T[255]; // @[ReplacePipe.scala 179:46]
  wire [16:0] data_full_wayBits_0_0 = {read_codes_0_0,read_datas_0_0}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_0_1 = {read_codes_0_1,read_datas_0_1}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_0_2 = {read_codes_0_2,read_datas_0_2}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_0_3 = {read_codes_0_3,read_datas_0_3}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_0_4 = {read_codes_0_4,read_datas_0_4}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_0_5 = {read_codes_0_5,read_datas_0_5}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_0_6 = {read_codes_0_6,read_datas_0_6}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_0_7 = {read_codes_0_7,read_datas_0_7}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_0_8 = {read_codes_0_8,read_datas_0_8}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_0_9 = {read_codes_0_9,read_datas_0_9}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_0_10 = {read_codes_0_10,read_datas_0_10}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_0_11 = {read_codes_0_11,read_datas_0_11}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_0_12 = {read_codes_0_12,read_datas_0_12}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_0_13 = {read_codes_0_13,read_datas_0_13}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_0_14 = {read_codes_0_14,read_datas_0_14}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_0_15 = {read_codes_0_15,read_datas_0_15}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_0_16 = {read_codes_0_16,read_datas_0_16}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_0_17 = {read_codes_0_17,read_datas_0_17}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_0_18 = {read_codes_0_18,read_datas_0_18}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_0_19 = {read_codes_0_19,read_datas_0_19}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_0_20 = {read_codes_0_20,read_datas_0_20}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_0_21 = {read_codes_0_21,read_datas_0_21}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_0_22 = {read_codes_0_22,read_datas_0_22}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_0_23 = {read_codes_0_23,read_datas_0_23}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_0_24 = {read_codes_0_24,read_datas_0_24}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_0_25 = {read_codes_0_25,read_datas_0_25}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_0_26 = {read_codes_0_26,read_datas_0_26}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_0_27 = {read_codes_0_27,read_datas_0_27}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_0_28 = {read_codes_0_28,read_datas_0_28}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_0_29 = {read_codes_0_29,read_datas_0_29}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_0_30 = {read_codes_0_30,read_datas_0_30}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_0_31 = {read_codes_0_31,read_datas_0_31}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_0 = {read_codes_1_0,read_datas_1_0}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_1 = {read_codes_1_1,read_datas_1_1}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_2 = {read_codes_1_2,read_datas_1_2}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_3 = {read_codes_1_3,read_datas_1_3}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_4 = {read_codes_1_4,read_datas_1_4}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_5 = {read_codes_1_5,read_datas_1_5}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_6 = {read_codes_1_6,read_datas_1_6}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_7 = {read_codes_1_7,read_datas_1_7}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_8 = {read_codes_1_8,read_datas_1_8}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_9 = {read_codes_1_9,read_datas_1_9}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_10 = {read_codes_1_10,read_datas_1_10}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_11 = {read_codes_1_11,read_datas_1_11}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_12 = {read_codes_1_12,read_datas_1_12}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_13 = {read_codes_1_13,read_datas_1_13}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_14 = {read_codes_1_14,read_datas_1_14}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_15 = {read_codes_1_15,read_datas_1_15}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_16 = {read_codes_1_16,read_datas_1_16}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_17 = {read_codes_1_17,read_datas_1_17}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_18 = {read_codes_1_18,read_datas_1_18}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_19 = {read_codes_1_19,read_datas_1_19}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_20 = {read_codes_1_20,read_datas_1_20}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_21 = {read_codes_1_21,read_datas_1_21}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_22 = {read_codes_1_22,read_datas_1_22}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_23 = {read_codes_1_23,read_datas_1_23}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_24 = {read_codes_1_24,read_datas_1_24}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_25 = {read_codes_1_25,read_datas_1_25}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_26 = {read_codes_1_26,read_datas_1_26}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_27 = {read_codes_1_27,read_datas_1_27}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_28 = {read_codes_1_28,read_datas_1_28}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_29 = {read_codes_1_29,read_datas_1_29}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_30 = {read_codes_1_30,read_datas_1_30}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_31 = {read_codes_1_31,read_datas_1_31}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_2_0 = {read_codes_2_0,read_datas_2_0}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_2_1 = {read_codes_2_1,read_datas_2_1}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_2_2 = {read_codes_2_2,read_datas_2_2}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_2_3 = {read_codes_2_3,read_datas_2_3}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_2_4 = {read_codes_2_4,read_datas_2_4}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_2_5 = {read_codes_2_5,read_datas_2_5}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_2_6 = {read_codes_2_6,read_datas_2_6}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_2_7 = {read_codes_2_7,read_datas_2_7}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_2_8 = {read_codes_2_8,read_datas_2_8}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_2_9 = {read_codes_2_9,read_datas_2_9}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_2_10 = {read_codes_2_10,read_datas_2_10}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_2_11 = {read_codes_2_11,read_datas_2_11}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_2_12 = {read_codes_2_12,read_datas_2_12}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_2_13 = {read_codes_2_13,read_datas_2_13}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_2_14 = {read_codes_2_14,read_datas_2_14}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_2_15 = {read_codes_2_15,read_datas_2_15}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_2_16 = {read_codes_2_16,read_datas_2_16}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_2_17 = {read_codes_2_17,read_datas_2_17}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_2_18 = {read_codes_2_18,read_datas_2_18}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_2_19 = {read_codes_2_19,read_datas_2_19}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_2_20 = {read_codes_2_20,read_datas_2_20}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_2_21 = {read_codes_2_21,read_datas_2_21}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_2_22 = {read_codes_2_22,read_datas_2_22}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_2_23 = {read_codes_2_23,read_datas_2_23}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_2_24 = {read_codes_2_24,read_datas_2_24}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_2_25 = {read_codes_2_25,read_datas_2_25}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_2_26 = {read_codes_2_26,read_datas_2_26}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_2_27 = {read_codes_2_27,read_datas_2_27}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_2_28 = {read_codes_2_28,read_datas_2_28}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_2_29 = {read_codes_2_29,read_datas_2_29}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_2_30 = {read_codes_2_30,read_datas_2_30}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_2_31 = {read_codes_2_31,read_datas_2_31}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_3_0 = {read_codes_3_0,read_datas_3_0}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_3_1 = {read_codes_3_1,read_datas_3_1}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_3_2 = {read_codes_3_2,read_datas_3_2}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_3_3 = {read_codes_3_3,read_datas_3_3}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_3_4 = {read_codes_3_4,read_datas_3_4}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_3_5 = {read_codes_3_5,read_datas_3_5}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_3_6 = {read_codes_3_6,read_datas_3_6}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_3_7 = {read_codes_3_7,read_datas_3_7}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_3_8 = {read_codes_3_8,read_datas_3_8}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_3_9 = {read_codes_3_9,read_datas_3_9}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_3_10 = {read_codes_3_10,read_datas_3_10}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_3_11 = {read_codes_3_11,read_datas_3_11}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_3_12 = {read_codes_3_12,read_datas_3_12}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_3_13 = {read_codes_3_13,read_datas_3_13}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_3_14 = {read_codes_3_14,read_datas_3_14}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_3_15 = {read_codes_3_15,read_datas_3_15}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_3_16 = {read_codes_3_16,read_datas_3_16}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_3_17 = {read_codes_3_17,read_datas_3_17}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_3_18 = {read_codes_3_18,read_datas_3_18}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_3_19 = {read_codes_3_19,read_datas_3_19}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_3_20 = {read_codes_3_20,read_datas_3_20}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_3_21 = {read_codes_3_21,read_datas_3_21}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_3_22 = {read_codes_3_22,read_datas_3_22}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_3_23 = {read_codes_3_23,read_datas_3_23}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_3_24 = {read_codes_3_24,read_datas_3_24}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_3_25 = {read_codes_3_25,read_datas_3_25}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_3_26 = {read_codes_3_26,read_datas_3_26}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_3_27 = {read_codes_3_27,read_datas_3_27}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_3_28 = {read_codes_3_28,read_datas_3_28}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_3_29 = {read_codes_3_29,read_datas_3_29}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_3_30 = {read_codes_3_30,read_datas_3_30}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_3_31 = {read_codes_3_31,read_datas_3_31}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_4_0 = {read_codes_4_0,read_datas_4_0}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_4_1 = {read_codes_4_1,read_datas_4_1}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_4_2 = {read_codes_4_2,read_datas_4_2}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_4_3 = {read_codes_4_3,read_datas_4_3}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_4_4 = {read_codes_4_4,read_datas_4_4}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_4_5 = {read_codes_4_5,read_datas_4_5}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_4_6 = {read_codes_4_6,read_datas_4_6}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_4_7 = {read_codes_4_7,read_datas_4_7}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_4_8 = {read_codes_4_8,read_datas_4_8}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_4_9 = {read_codes_4_9,read_datas_4_9}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_4_10 = {read_codes_4_10,read_datas_4_10}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_4_11 = {read_codes_4_11,read_datas_4_11}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_4_12 = {read_codes_4_12,read_datas_4_12}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_4_13 = {read_codes_4_13,read_datas_4_13}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_4_14 = {read_codes_4_14,read_datas_4_14}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_4_15 = {read_codes_4_15,read_datas_4_15}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_4_16 = {read_codes_4_16,read_datas_4_16}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_4_17 = {read_codes_4_17,read_datas_4_17}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_4_18 = {read_codes_4_18,read_datas_4_18}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_4_19 = {read_codes_4_19,read_datas_4_19}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_4_20 = {read_codes_4_20,read_datas_4_20}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_4_21 = {read_codes_4_21,read_datas_4_21}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_4_22 = {read_codes_4_22,read_datas_4_22}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_4_23 = {read_codes_4_23,read_datas_4_23}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_4_24 = {read_codes_4_24,read_datas_4_24}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_4_25 = {read_codes_4_25,read_datas_4_25}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_4_26 = {read_codes_4_26,read_datas_4_26}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_4_27 = {read_codes_4_27,read_datas_4_27}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_4_28 = {read_codes_4_28,read_datas_4_28}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_4_29 = {read_codes_4_29,read_datas_4_29}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_4_30 = {read_codes_4_30,read_datas_4_30}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_4_31 = {read_codes_4_31,read_datas_4_31}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_5_0 = {read_codes_5_0,read_datas_5_0}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_5_1 = {read_codes_5_1,read_datas_5_1}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_5_2 = {read_codes_5_2,read_datas_5_2}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_5_3 = {read_codes_5_3,read_datas_5_3}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_5_4 = {read_codes_5_4,read_datas_5_4}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_5_5 = {read_codes_5_5,read_datas_5_5}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_5_6 = {read_codes_5_6,read_datas_5_6}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_5_7 = {read_codes_5_7,read_datas_5_7}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_5_8 = {read_codes_5_8,read_datas_5_8}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_5_9 = {read_codes_5_9,read_datas_5_9}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_5_10 = {read_codes_5_10,read_datas_5_10}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_5_11 = {read_codes_5_11,read_datas_5_11}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_5_12 = {read_codes_5_12,read_datas_5_12}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_5_13 = {read_codes_5_13,read_datas_5_13}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_5_14 = {read_codes_5_14,read_datas_5_14}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_5_15 = {read_codes_5_15,read_datas_5_15}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_5_16 = {read_codes_5_16,read_datas_5_16}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_5_17 = {read_codes_5_17,read_datas_5_17}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_5_18 = {read_codes_5_18,read_datas_5_18}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_5_19 = {read_codes_5_19,read_datas_5_19}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_5_20 = {read_codes_5_20,read_datas_5_20}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_5_21 = {read_codes_5_21,read_datas_5_21}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_5_22 = {read_codes_5_22,read_datas_5_22}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_5_23 = {read_codes_5_23,read_datas_5_23}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_5_24 = {read_codes_5_24,read_datas_5_24}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_5_25 = {read_codes_5_25,read_datas_5_25}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_5_26 = {read_codes_5_26,read_datas_5_26}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_5_27 = {read_codes_5_27,read_datas_5_27}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_5_28 = {read_codes_5_28,read_datas_5_28}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_5_29 = {read_codes_5_29,read_datas_5_29}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_5_30 = {read_codes_5_30,read_datas_5_30}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_5_31 = {read_codes_5_31,read_datas_5_31}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_6_0 = {read_codes_6_0,read_datas_6_0}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_6_1 = {read_codes_6_1,read_datas_6_1}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_6_2 = {read_codes_6_2,read_datas_6_2}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_6_3 = {read_codes_6_3,read_datas_6_3}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_6_4 = {read_codes_6_4,read_datas_6_4}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_6_5 = {read_codes_6_5,read_datas_6_5}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_6_6 = {read_codes_6_6,read_datas_6_6}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_6_7 = {read_codes_6_7,read_datas_6_7}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_6_8 = {read_codes_6_8,read_datas_6_8}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_6_9 = {read_codes_6_9,read_datas_6_9}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_6_10 = {read_codes_6_10,read_datas_6_10}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_6_11 = {read_codes_6_11,read_datas_6_11}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_6_12 = {read_codes_6_12,read_datas_6_12}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_6_13 = {read_codes_6_13,read_datas_6_13}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_6_14 = {read_codes_6_14,read_datas_6_14}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_6_15 = {read_codes_6_15,read_datas_6_15}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_6_16 = {read_codes_6_16,read_datas_6_16}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_6_17 = {read_codes_6_17,read_datas_6_17}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_6_18 = {read_codes_6_18,read_datas_6_18}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_6_19 = {read_codes_6_19,read_datas_6_19}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_6_20 = {read_codes_6_20,read_datas_6_20}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_6_21 = {read_codes_6_21,read_datas_6_21}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_6_22 = {read_codes_6_22,read_datas_6_22}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_6_23 = {read_codes_6_23,read_datas_6_23}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_6_24 = {read_codes_6_24,read_datas_6_24}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_6_25 = {read_codes_6_25,read_datas_6_25}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_6_26 = {read_codes_6_26,read_datas_6_26}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_6_27 = {read_codes_6_27,read_datas_6_27}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_6_28 = {read_codes_6_28,read_datas_6_28}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_6_29 = {read_codes_6_29,read_datas_6_29}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_6_30 = {read_codes_6_30,read_datas_6_30}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_6_31 = {read_codes_6_31,read_datas_6_31}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_7_0 = {read_codes_7_0,read_datas_7_0}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_7_1 = {read_codes_7_1,read_datas_7_1}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_7_2 = {read_codes_7_2,read_datas_7_2}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_7_3 = {read_codes_7_3,read_datas_7_3}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_7_4 = {read_codes_7_4,read_datas_7_4}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_7_5 = {read_codes_7_5,read_datas_7_5}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_7_6 = {read_codes_7_6,read_datas_7_6}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_7_7 = {read_codes_7_7,read_datas_7_7}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_7_8 = {read_codes_7_8,read_datas_7_8}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_7_9 = {read_codes_7_9,read_datas_7_9}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_7_10 = {read_codes_7_10,read_datas_7_10}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_7_11 = {read_codes_7_11,read_datas_7_11}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_7_12 = {read_codes_7_12,read_datas_7_12}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_7_13 = {read_codes_7_13,read_datas_7_13}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_7_14 = {read_codes_7_14,read_datas_7_14}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_7_15 = {read_codes_7_15,read_datas_7_15}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_7_16 = {read_codes_7_16,read_datas_7_16}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_7_17 = {read_codes_7_17,read_datas_7_17}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_7_18 = {read_codes_7_18,read_datas_7_18}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_7_19 = {read_codes_7_19,read_datas_7_19}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_7_20 = {read_codes_7_20,read_datas_7_20}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_7_21 = {read_codes_7_21,read_datas_7_21}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_7_22 = {read_codes_7_22,read_datas_7_22}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_7_23 = {read_codes_7_23,read_datas_7_23}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_7_24 = {read_codes_7_24,read_datas_7_24}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_7_25 = {read_codes_7_25,read_datas_7_25}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_7_26 = {read_codes_7_26,read_datas_7_26}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_7_27 = {read_codes_7_27,read_datas_7_27}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_7_28 = {read_codes_7_28,read_datas_7_28}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_7_29 = {read_codes_7_29,read_datas_7_29}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_7_30 = {read_codes_7_30,read_datas_7_30}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_7_31 = {read_codes_7_31,read_datas_7_31}; // @[Cat.scala 31:58]
  reg  r2_data_errors_0_REG; // @[ReplacePipe.scala 186:65]
  reg  r2_data_errors_0_REG_1; // @[ReplacePipe.scala 186:57]
  reg  r2_data_errors_0_REG_2_0; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_0_REG_2_1; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_0_REG_2_2; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_0_REG_2_3; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_0_REG_2_4; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_0_REG_2_5; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_0_REG_2_6; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_0_REG_2_7; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_0_REG_2_8; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_0_REG_2_9; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_0_REG_2_10; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_0_REG_2_11; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_0_REG_2_12; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_0_REG_2_13; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_0_REG_2_14; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_0_REG_2_15; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_0_REG_2_16; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_0_REG_2_17; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_0_REG_2_18; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_0_REG_2_19; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_0_REG_2_20; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_0_REG_2_21; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_0_REG_2_22; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_0_REG_2_23; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_0_REG_2_24; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_0_REG_2_25; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_0_REG_2_26; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_0_REG_2_27; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_0_REG_2_28; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_0_REG_2_29; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_0_REG_2_30; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_0_REG_2_31; // @[ReplacePipe.scala 186:86]
  wire  _r2_data_errors_0_T_29 = r2_data_errors_0_REG_2_0 | r2_data_errors_0_REG_2_1 | r2_data_errors_0_REG_2_2 |
    r2_data_errors_0_REG_2_3 | r2_data_errors_0_REG_2_4 | r2_data_errors_0_REG_2_5 | r2_data_errors_0_REG_2_6 |
    r2_data_errors_0_REG_2_7 | r2_data_errors_0_REG_2_8 | r2_data_errors_0_REG_2_9 | r2_data_errors_0_REG_2_10 |
    r2_data_errors_0_REG_2_11 | r2_data_errors_0_REG_2_12 | r2_data_errors_0_REG_2_13 | r2_data_errors_0_REG_2_14 |
    r2_data_errors_0_REG_2_15 | r2_data_errors_0_REG_2_16 | r2_data_errors_0_REG_2_17 | r2_data_errors_0_REG_2_18 |
    r2_data_errors_0_REG_2_19 | r2_data_errors_0_REG_2_20 | r2_data_errors_0_REG_2_21 | r2_data_errors_0_REG_2_22 |
    r2_data_errors_0_REG_2_23 | r2_data_errors_0_REG_2_24 | r2_data_errors_0_REG_2_25 | r2_data_errors_0_REG_2_26 |
    r2_data_errors_0_REG_2_27 | r2_data_errors_0_REG_2_28 | r2_data_errors_0_REG_2_29 | r2_data_errors_0_REG_2_30; // @[ReplacePipe.scala 186:118]
  wire  r2_data_errors_0 = r2_data_errors_0_REG_1 & (_r2_data_errors_0_T_29 | r2_data_errors_0_REG_2_31); // @[ReplacePipe.scala 186:76]
  reg  r2_data_errors_1_REG; // @[ReplacePipe.scala 186:65]
  reg  r2_data_errors_1_REG_1; // @[ReplacePipe.scala 186:57]
  reg  r2_data_errors_1_REG_2_0; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_1_REG_2_1; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_1_REG_2_2; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_1_REG_2_3; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_1_REG_2_4; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_1_REG_2_5; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_1_REG_2_6; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_1_REG_2_7; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_1_REG_2_8; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_1_REG_2_9; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_1_REG_2_10; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_1_REG_2_11; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_1_REG_2_12; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_1_REG_2_13; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_1_REG_2_14; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_1_REG_2_15; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_1_REG_2_16; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_1_REG_2_17; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_1_REG_2_18; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_1_REG_2_19; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_1_REG_2_20; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_1_REG_2_21; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_1_REG_2_22; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_1_REG_2_23; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_1_REG_2_24; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_1_REG_2_25; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_1_REG_2_26; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_1_REG_2_27; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_1_REG_2_28; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_1_REG_2_29; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_1_REG_2_30; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_1_REG_2_31; // @[ReplacePipe.scala 186:86]
  wire  _r2_data_errors_1_T_29 = r2_data_errors_1_REG_2_0 | r2_data_errors_1_REG_2_1 | r2_data_errors_1_REG_2_2 |
    r2_data_errors_1_REG_2_3 | r2_data_errors_1_REG_2_4 | r2_data_errors_1_REG_2_5 | r2_data_errors_1_REG_2_6 |
    r2_data_errors_1_REG_2_7 | r2_data_errors_1_REG_2_8 | r2_data_errors_1_REG_2_9 | r2_data_errors_1_REG_2_10 |
    r2_data_errors_1_REG_2_11 | r2_data_errors_1_REG_2_12 | r2_data_errors_1_REG_2_13 | r2_data_errors_1_REG_2_14 |
    r2_data_errors_1_REG_2_15 | r2_data_errors_1_REG_2_16 | r2_data_errors_1_REG_2_17 | r2_data_errors_1_REG_2_18 |
    r2_data_errors_1_REG_2_19 | r2_data_errors_1_REG_2_20 | r2_data_errors_1_REG_2_21 | r2_data_errors_1_REG_2_22 |
    r2_data_errors_1_REG_2_23 | r2_data_errors_1_REG_2_24 | r2_data_errors_1_REG_2_25 | r2_data_errors_1_REG_2_26 |
    r2_data_errors_1_REG_2_27 | r2_data_errors_1_REG_2_28 | r2_data_errors_1_REG_2_29 | r2_data_errors_1_REG_2_30; // @[ReplacePipe.scala 186:118]
  wire  r2_data_errors_1 = r2_data_errors_1_REG_1 & (_r2_data_errors_1_T_29 | r2_data_errors_1_REG_2_31); // @[ReplacePipe.scala 186:76]
  reg  r2_data_errors_2_REG; // @[ReplacePipe.scala 186:65]
  reg  r2_data_errors_2_REG_1; // @[ReplacePipe.scala 186:57]
  reg  r2_data_errors_2_REG_2_0; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_2_REG_2_1; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_2_REG_2_2; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_2_REG_2_3; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_2_REG_2_4; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_2_REG_2_5; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_2_REG_2_6; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_2_REG_2_7; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_2_REG_2_8; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_2_REG_2_9; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_2_REG_2_10; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_2_REG_2_11; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_2_REG_2_12; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_2_REG_2_13; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_2_REG_2_14; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_2_REG_2_15; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_2_REG_2_16; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_2_REG_2_17; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_2_REG_2_18; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_2_REG_2_19; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_2_REG_2_20; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_2_REG_2_21; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_2_REG_2_22; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_2_REG_2_23; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_2_REG_2_24; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_2_REG_2_25; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_2_REG_2_26; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_2_REG_2_27; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_2_REG_2_28; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_2_REG_2_29; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_2_REG_2_30; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_2_REG_2_31; // @[ReplacePipe.scala 186:86]
  wire  _r2_data_errors_2_T_29 = r2_data_errors_2_REG_2_0 | r2_data_errors_2_REG_2_1 | r2_data_errors_2_REG_2_2 |
    r2_data_errors_2_REG_2_3 | r2_data_errors_2_REG_2_4 | r2_data_errors_2_REG_2_5 | r2_data_errors_2_REG_2_6 |
    r2_data_errors_2_REG_2_7 | r2_data_errors_2_REG_2_8 | r2_data_errors_2_REG_2_9 | r2_data_errors_2_REG_2_10 |
    r2_data_errors_2_REG_2_11 | r2_data_errors_2_REG_2_12 | r2_data_errors_2_REG_2_13 | r2_data_errors_2_REG_2_14 |
    r2_data_errors_2_REG_2_15 | r2_data_errors_2_REG_2_16 | r2_data_errors_2_REG_2_17 | r2_data_errors_2_REG_2_18 |
    r2_data_errors_2_REG_2_19 | r2_data_errors_2_REG_2_20 | r2_data_errors_2_REG_2_21 | r2_data_errors_2_REG_2_22 |
    r2_data_errors_2_REG_2_23 | r2_data_errors_2_REG_2_24 | r2_data_errors_2_REG_2_25 | r2_data_errors_2_REG_2_26 |
    r2_data_errors_2_REG_2_27 | r2_data_errors_2_REG_2_28 | r2_data_errors_2_REG_2_29 | r2_data_errors_2_REG_2_30; // @[ReplacePipe.scala 186:118]
  wire  r2_data_errors_2 = r2_data_errors_2_REG_1 & (_r2_data_errors_2_T_29 | r2_data_errors_2_REG_2_31); // @[ReplacePipe.scala 186:76]
  reg  r2_data_errors_3_REG; // @[ReplacePipe.scala 186:65]
  reg  r2_data_errors_3_REG_1; // @[ReplacePipe.scala 186:57]
  reg  r2_data_errors_3_REG_2_0; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_3_REG_2_1; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_3_REG_2_2; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_3_REG_2_3; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_3_REG_2_4; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_3_REG_2_5; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_3_REG_2_6; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_3_REG_2_7; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_3_REG_2_8; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_3_REG_2_9; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_3_REG_2_10; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_3_REG_2_11; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_3_REG_2_12; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_3_REG_2_13; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_3_REG_2_14; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_3_REG_2_15; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_3_REG_2_16; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_3_REG_2_17; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_3_REG_2_18; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_3_REG_2_19; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_3_REG_2_20; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_3_REG_2_21; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_3_REG_2_22; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_3_REG_2_23; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_3_REG_2_24; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_3_REG_2_25; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_3_REG_2_26; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_3_REG_2_27; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_3_REG_2_28; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_3_REG_2_29; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_3_REG_2_30; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_3_REG_2_31; // @[ReplacePipe.scala 186:86]
  wire  _r2_data_errors_3_T_29 = r2_data_errors_3_REG_2_0 | r2_data_errors_3_REG_2_1 | r2_data_errors_3_REG_2_2 |
    r2_data_errors_3_REG_2_3 | r2_data_errors_3_REG_2_4 | r2_data_errors_3_REG_2_5 | r2_data_errors_3_REG_2_6 |
    r2_data_errors_3_REG_2_7 | r2_data_errors_3_REG_2_8 | r2_data_errors_3_REG_2_9 | r2_data_errors_3_REG_2_10 |
    r2_data_errors_3_REG_2_11 | r2_data_errors_3_REG_2_12 | r2_data_errors_3_REG_2_13 | r2_data_errors_3_REG_2_14 |
    r2_data_errors_3_REG_2_15 | r2_data_errors_3_REG_2_16 | r2_data_errors_3_REG_2_17 | r2_data_errors_3_REG_2_18 |
    r2_data_errors_3_REG_2_19 | r2_data_errors_3_REG_2_20 | r2_data_errors_3_REG_2_21 | r2_data_errors_3_REG_2_22 |
    r2_data_errors_3_REG_2_23 | r2_data_errors_3_REG_2_24 | r2_data_errors_3_REG_2_25 | r2_data_errors_3_REG_2_26 |
    r2_data_errors_3_REG_2_27 | r2_data_errors_3_REG_2_28 | r2_data_errors_3_REG_2_29 | r2_data_errors_3_REG_2_30; // @[ReplacePipe.scala 186:118]
  wire  r2_data_errors_3 = r2_data_errors_3_REG_1 & (_r2_data_errors_3_T_29 | r2_data_errors_3_REG_2_31); // @[ReplacePipe.scala 186:76]
  reg  r2_data_errors_4_REG; // @[ReplacePipe.scala 186:65]
  reg  r2_data_errors_4_REG_1; // @[ReplacePipe.scala 186:57]
  reg  r2_data_errors_4_REG_2_0; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_4_REG_2_1; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_4_REG_2_2; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_4_REG_2_3; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_4_REG_2_4; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_4_REG_2_5; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_4_REG_2_6; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_4_REG_2_7; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_4_REG_2_8; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_4_REG_2_9; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_4_REG_2_10; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_4_REG_2_11; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_4_REG_2_12; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_4_REG_2_13; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_4_REG_2_14; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_4_REG_2_15; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_4_REG_2_16; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_4_REG_2_17; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_4_REG_2_18; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_4_REG_2_19; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_4_REG_2_20; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_4_REG_2_21; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_4_REG_2_22; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_4_REG_2_23; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_4_REG_2_24; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_4_REG_2_25; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_4_REG_2_26; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_4_REG_2_27; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_4_REG_2_28; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_4_REG_2_29; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_4_REG_2_30; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_4_REG_2_31; // @[ReplacePipe.scala 186:86]
  wire  _r2_data_errors_4_T_29 = r2_data_errors_4_REG_2_0 | r2_data_errors_4_REG_2_1 | r2_data_errors_4_REG_2_2 |
    r2_data_errors_4_REG_2_3 | r2_data_errors_4_REG_2_4 | r2_data_errors_4_REG_2_5 | r2_data_errors_4_REG_2_6 |
    r2_data_errors_4_REG_2_7 | r2_data_errors_4_REG_2_8 | r2_data_errors_4_REG_2_9 | r2_data_errors_4_REG_2_10 |
    r2_data_errors_4_REG_2_11 | r2_data_errors_4_REG_2_12 | r2_data_errors_4_REG_2_13 | r2_data_errors_4_REG_2_14 |
    r2_data_errors_4_REG_2_15 | r2_data_errors_4_REG_2_16 | r2_data_errors_4_REG_2_17 | r2_data_errors_4_REG_2_18 |
    r2_data_errors_4_REG_2_19 | r2_data_errors_4_REG_2_20 | r2_data_errors_4_REG_2_21 | r2_data_errors_4_REG_2_22 |
    r2_data_errors_4_REG_2_23 | r2_data_errors_4_REG_2_24 | r2_data_errors_4_REG_2_25 | r2_data_errors_4_REG_2_26 |
    r2_data_errors_4_REG_2_27 | r2_data_errors_4_REG_2_28 | r2_data_errors_4_REG_2_29 | r2_data_errors_4_REG_2_30; // @[ReplacePipe.scala 186:118]
  wire  r2_data_errors_4 = r2_data_errors_4_REG_1 & (_r2_data_errors_4_T_29 | r2_data_errors_4_REG_2_31); // @[ReplacePipe.scala 186:76]
  reg  r2_data_errors_5_REG; // @[ReplacePipe.scala 186:65]
  reg  r2_data_errors_5_REG_1; // @[ReplacePipe.scala 186:57]
  reg  r2_data_errors_5_REG_2_0; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_5_REG_2_1; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_5_REG_2_2; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_5_REG_2_3; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_5_REG_2_4; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_5_REG_2_5; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_5_REG_2_6; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_5_REG_2_7; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_5_REG_2_8; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_5_REG_2_9; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_5_REG_2_10; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_5_REG_2_11; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_5_REG_2_12; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_5_REG_2_13; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_5_REG_2_14; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_5_REG_2_15; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_5_REG_2_16; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_5_REG_2_17; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_5_REG_2_18; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_5_REG_2_19; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_5_REG_2_20; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_5_REG_2_21; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_5_REG_2_22; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_5_REG_2_23; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_5_REG_2_24; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_5_REG_2_25; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_5_REG_2_26; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_5_REG_2_27; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_5_REG_2_28; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_5_REG_2_29; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_5_REG_2_30; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_5_REG_2_31; // @[ReplacePipe.scala 186:86]
  wire  _r2_data_errors_5_T_29 = r2_data_errors_5_REG_2_0 | r2_data_errors_5_REG_2_1 | r2_data_errors_5_REG_2_2 |
    r2_data_errors_5_REG_2_3 | r2_data_errors_5_REG_2_4 | r2_data_errors_5_REG_2_5 | r2_data_errors_5_REG_2_6 |
    r2_data_errors_5_REG_2_7 | r2_data_errors_5_REG_2_8 | r2_data_errors_5_REG_2_9 | r2_data_errors_5_REG_2_10 |
    r2_data_errors_5_REG_2_11 | r2_data_errors_5_REG_2_12 | r2_data_errors_5_REG_2_13 | r2_data_errors_5_REG_2_14 |
    r2_data_errors_5_REG_2_15 | r2_data_errors_5_REG_2_16 | r2_data_errors_5_REG_2_17 | r2_data_errors_5_REG_2_18 |
    r2_data_errors_5_REG_2_19 | r2_data_errors_5_REG_2_20 | r2_data_errors_5_REG_2_21 | r2_data_errors_5_REG_2_22 |
    r2_data_errors_5_REG_2_23 | r2_data_errors_5_REG_2_24 | r2_data_errors_5_REG_2_25 | r2_data_errors_5_REG_2_26 |
    r2_data_errors_5_REG_2_27 | r2_data_errors_5_REG_2_28 | r2_data_errors_5_REG_2_29 | r2_data_errors_5_REG_2_30; // @[ReplacePipe.scala 186:118]
  wire  r2_data_errors_5 = r2_data_errors_5_REG_1 & (_r2_data_errors_5_T_29 | r2_data_errors_5_REG_2_31); // @[ReplacePipe.scala 186:76]
  reg  r2_data_errors_6_REG; // @[ReplacePipe.scala 186:65]
  reg  r2_data_errors_6_REG_1; // @[ReplacePipe.scala 186:57]
  reg  r2_data_errors_6_REG_2_0; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_6_REG_2_1; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_6_REG_2_2; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_6_REG_2_3; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_6_REG_2_4; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_6_REG_2_5; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_6_REG_2_6; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_6_REG_2_7; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_6_REG_2_8; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_6_REG_2_9; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_6_REG_2_10; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_6_REG_2_11; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_6_REG_2_12; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_6_REG_2_13; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_6_REG_2_14; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_6_REG_2_15; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_6_REG_2_16; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_6_REG_2_17; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_6_REG_2_18; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_6_REG_2_19; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_6_REG_2_20; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_6_REG_2_21; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_6_REG_2_22; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_6_REG_2_23; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_6_REG_2_24; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_6_REG_2_25; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_6_REG_2_26; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_6_REG_2_27; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_6_REG_2_28; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_6_REG_2_29; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_6_REG_2_30; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_6_REG_2_31; // @[ReplacePipe.scala 186:86]
  wire  _r2_data_errors_6_T_29 = r2_data_errors_6_REG_2_0 | r2_data_errors_6_REG_2_1 | r2_data_errors_6_REG_2_2 |
    r2_data_errors_6_REG_2_3 | r2_data_errors_6_REG_2_4 | r2_data_errors_6_REG_2_5 | r2_data_errors_6_REG_2_6 |
    r2_data_errors_6_REG_2_7 | r2_data_errors_6_REG_2_8 | r2_data_errors_6_REG_2_9 | r2_data_errors_6_REG_2_10 |
    r2_data_errors_6_REG_2_11 | r2_data_errors_6_REG_2_12 | r2_data_errors_6_REG_2_13 | r2_data_errors_6_REG_2_14 |
    r2_data_errors_6_REG_2_15 | r2_data_errors_6_REG_2_16 | r2_data_errors_6_REG_2_17 | r2_data_errors_6_REG_2_18 |
    r2_data_errors_6_REG_2_19 | r2_data_errors_6_REG_2_20 | r2_data_errors_6_REG_2_21 | r2_data_errors_6_REG_2_22 |
    r2_data_errors_6_REG_2_23 | r2_data_errors_6_REG_2_24 | r2_data_errors_6_REG_2_25 | r2_data_errors_6_REG_2_26 |
    r2_data_errors_6_REG_2_27 | r2_data_errors_6_REG_2_28 | r2_data_errors_6_REG_2_29 | r2_data_errors_6_REG_2_30; // @[ReplacePipe.scala 186:118]
  wire  r2_data_errors_6 = r2_data_errors_6_REG_1 & (_r2_data_errors_6_T_29 | r2_data_errors_6_REG_2_31); // @[ReplacePipe.scala 186:76]
  reg  r2_data_errors_7_REG; // @[ReplacePipe.scala 186:65]
  reg  r2_data_errors_7_REG_1; // @[ReplacePipe.scala 186:57]
  reg  r2_data_errors_7_REG_2_0; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_7_REG_2_1; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_7_REG_2_2; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_7_REG_2_3; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_7_REG_2_4; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_7_REG_2_5; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_7_REG_2_6; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_7_REG_2_7; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_7_REG_2_8; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_7_REG_2_9; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_7_REG_2_10; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_7_REG_2_11; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_7_REG_2_12; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_7_REG_2_13; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_7_REG_2_14; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_7_REG_2_15; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_7_REG_2_16; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_7_REG_2_17; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_7_REG_2_18; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_7_REG_2_19; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_7_REG_2_20; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_7_REG_2_21; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_7_REG_2_22; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_7_REG_2_23; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_7_REG_2_24; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_7_REG_2_25; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_7_REG_2_26; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_7_REG_2_27; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_7_REG_2_28; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_7_REG_2_29; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_7_REG_2_30; // @[ReplacePipe.scala 186:86]
  reg  r2_data_errors_7_REG_2_31; // @[ReplacePipe.scala 186:86]
  wire  _r2_data_errors_7_T_29 = r2_data_errors_7_REG_2_0 | r2_data_errors_7_REG_2_1 | r2_data_errors_7_REG_2_2 |
    r2_data_errors_7_REG_2_3 | r2_data_errors_7_REG_2_4 | r2_data_errors_7_REG_2_5 | r2_data_errors_7_REG_2_6 |
    r2_data_errors_7_REG_2_7 | r2_data_errors_7_REG_2_8 | r2_data_errors_7_REG_2_9 | r2_data_errors_7_REG_2_10 |
    r2_data_errors_7_REG_2_11 | r2_data_errors_7_REG_2_12 | r2_data_errors_7_REG_2_13 | r2_data_errors_7_REG_2_14 |
    r2_data_errors_7_REG_2_15 | r2_data_errors_7_REG_2_16 | r2_data_errors_7_REG_2_17 | r2_data_errors_7_REG_2_18 |
    r2_data_errors_7_REG_2_19 | r2_data_errors_7_REG_2_20 | r2_data_errors_7_REG_2_21 | r2_data_errors_7_REG_2_22 |
    r2_data_errors_7_REG_2_23 | r2_data_errors_7_REG_2_24 | r2_data_errors_7_REG_2_25 | r2_data_errors_7_REG_2_26 |
    r2_data_errors_7_REG_2_27 | r2_data_errors_7_REG_2_28 | r2_data_errors_7_REG_2_29 | r2_data_errors_7_REG_2_30; // @[ReplacePipe.scala 186:118]
  wire  r2_data_errors_7 = r2_data_errors_7_REG_1 & (_r2_data_errors_7_T_29 | r2_data_errors_7_REG_2_31); // @[ReplacePipe.scala 186:76]
  wire  r2_parity_data_error = (r2_data_errors_0 | r2_data_errors_1 | r2_data_errors_2 | r2_data_errors_3 |
    r2_data_errors_4 | r2_data_errors_5 | r2_data_errors_6 | r2_data_errors_7) & io_csr_parity_enable; // @[ReplacePipe.scala 189:58]
  reg  r2_parity_error_REG; // @[ReplacePipe.scala 190:37]
  wire  r2_parity_error = r2_parity_error_REG | r2_parity_data_error; // @[ReplacePipe.scala 190:60]
  reg  io_error_valid_REG; // @[ReplacePipe.scala 193:79]
  reg  io_error_valid_REG_1; // @[ReplacePipe.scala 193:71]
  reg  io_error_valid_REG_2; // @[ReplacePipe.scala 193:43]
  reg  io_error_report_to_beu_REG; // @[ReplacePipe.scala 194:79]
  reg  io_error_report_to_beu_REG_1; // @[ReplacePipe.scala 194:71]
  reg  io_error_report_to_beu_REG_2; // @[ReplacePipe.scala 194:43]
  reg [35:0] io_error_paddr_REG; // @[ReplacePipe.scala 195:51]
  reg [35:0] io_error_paddr_REG_1; // @[ReplacePipe.scala 195:43]
  reg  io_error_source_tag_REG; // @[ReplacePipe.scala 196:51]
  reg  io_error_source_tag_REG_1; // @[ReplacePipe.scala 196:43]
  reg  io_error_source_data_REG; // @[ReplacePipe.scala 197:43]
  reg  io_error_opType_release_REG; // @[ReplacePipe.scala 201:51]
  reg  io_error_opType_release_REG_1; // @[ReplacePipe.scala 201:43]
  wire  _io_error_opType_probe_T = ~r2_req_voluntary; // @[ReplacePipe.scala 39:17]
  reg  io_error_opType_probe_REG; // @[ReplacePipe.scala 202:51]
  reg  io_error_opType_probe_REG_1; // @[ReplacePipe.scala 202:43]
  reg [1:0] r2_release_coh_state; // @[Reg.scala 16:16]
  wire [511:0] _r2_release_data_T_8 = r2_req_waymask[0] ? r2_data_cacheline_0 : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _r2_release_data_T_9 = r2_req_waymask[1] ? r2_data_cacheline_1 : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _r2_release_data_T_10 = r2_req_waymask[2] ? r2_data_cacheline_2 : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _r2_release_data_T_11 = r2_req_waymask[3] ? r2_data_cacheline_3 : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _r2_release_data_T_12 = r2_req_waymask[4] ? r2_data_cacheline_4 : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _r2_release_data_T_13 = r2_req_waymask[5] ? r2_data_cacheline_5 : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _r2_release_data_T_14 = r2_req_waymask[6] ? r2_data_cacheline_6 : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _r2_release_data_T_15 = r2_req_waymask[7] ? r2_data_cacheline_7 : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _r2_release_data_T_16 = _r2_release_data_T_8 | _r2_release_data_T_9; // @[Mux.scala 27:73]
  wire [511:0] _r2_release_data_T_17 = _r2_release_data_T_16 | _r2_release_data_T_10; // @[Mux.scala 27:73]
  wire [511:0] _r2_release_data_T_18 = _r2_release_data_T_17 | _r2_release_data_T_11; // @[Mux.scala 27:73]
  wire [511:0] _r2_release_data_T_19 = _r2_release_data_T_18 | _r2_release_data_T_12; // @[Mux.scala 27:73]
  wire [511:0] _r2_release_data_T_20 = _r2_release_data_T_19 | _r2_release_data_T_13; // @[Mux.scala 27:73]
  wire [511:0] _r2_release_data_T_21 = _r2_release_data_T_20 | _r2_release_data_T_14; // @[Mux.scala 27:73]
  wire [511:0] r2_release_data = _r2_release_data_T_21 | _r2_release_data_T_15; // @[Mux.scala 27:73]
  reg [35:0] r2_release_addr; // @[Reg.scala 16:16]
  wire  _release_need_send_T_1 = r2_release_coh_state > 2'h0; // @[Metadata.scala 49:45]
  wire  release_need_send = r2_valid & r2_req_voluntary & _release_need_send_T_1; // @[ReplacePipe.scala 213:57]
  wire [3:0] _T_133 = {2'h2,r2_release_coh_state}; // @[Cat.scala 31:58]
  wire  _T_146 = 4'h8 == _T_133; // @[Misc.scala 55:20]
  wire [2:0] _T_148 = _T_146 ? 3'h5 : 3'h0; // @[Misc.scala 37:36]
  wire  _T_150 = 4'h9 == _T_133; // @[Misc.scala 55:20]
  wire [2:0] _T_152 = _T_150 ? 3'h2 : _T_148; // @[Misc.scala 37:36]
  wire  _T_154 = 4'ha == _T_133; // @[Misc.scala 55:20]
  wire [2:0] _T_156 = _T_154 ? 3'h1 : _T_152; // @[Misc.scala 37:36]
  wire  _T_158 = 4'hb == _T_133; // @[Misc.scala 55:20]
  wire [2:0] _T_160 = _T_158 ? 3'h1 : _T_156; // @[Misc.scala 37:36]
  wire  _T_162 = 4'h4 == _T_133; // @[Misc.scala 55:20]
  wire  _T_163 = _T_162 ? 1'h0 : _T_158; // @[Misc.scala 37:9]
  wire [2:0] _T_164 = _T_162 ? 3'h5 : _T_160; // @[Misc.scala 37:36]
  wire  _T_166 = 4'h5 == _T_133; // @[Misc.scala 55:20]
  wire  _T_167 = _T_166 ? 1'h0 : _T_163; // @[Misc.scala 37:9]
  wire [2:0] _T_168 = _T_166 ? 3'h4 : _T_164; // @[Misc.scala 37:36]
  wire  _T_170 = 4'h6 == _T_133; // @[Misc.scala 55:20]
  wire  _T_171 = _T_170 ? 1'h0 : _T_167; // @[Misc.scala 37:9]
  wire [2:0] _T_172 = _T_170 ? 3'h0 : _T_168; // @[Misc.scala 37:36]
  wire  _T_174 = 4'h7 == _T_133; // @[Misc.scala 55:20]
  wire [2:0] _T_176 = _T_174 ? 3'h0 : _T_172; // @[Misc.scala 37:36]
  wire  _T_178 = 4'h0 == _T_133; // @[Misc.scala 55:20]
  wire  _T_179 = _T_178 ? 1'h0 : _T_174 | _T_171; // @[Misc.scala 37:9]
  wire [2:0] _T_180 = _T_178 ? 3'h5 : _T_176; // @[Misc.scala 37:36]
  wire  _T_182 = 4'h1 == _T_133; // @[Misc.scala 55:20]
  wire  _T_183 = _T_182 ? 1'h0 : _T_179; // @[Misc.scala 37:9]
  wire [2:0] _T_184 = _T_182 ? 3'h4 : _T_180; // @[Misc.scala 37:36]
  wire  _T_186 = 4'h2 == _T_133; // @[Misc.scala 55:20]
  wire  _T_187 = _T_186 ? 1'h0 : _T_183; // @[Misc.scala 37:9]
  wire [2:0] _T_188 = _T_186 ? 3'h3 : _T_184; // @[Misc.scala 37:36]
  wire  _T_190 = 4'h3 == _T_133; // @[Misc.scala 55:20]
  wire  release_has_dirty_data = _T_190 | _T_187; // @[Misc.scala 37:9]
  wire [2:0] release_shrink_param = _T_190 ? 3'h3 : _T_188; // @[Misc.scala 37:36]
  wire  _r2_hasData_T_1 = r2_probe_hit_coh_state > 2'h0; // @[Metadata.scala 49:45]
  wire [3:0] r2_write_waymask_lo = {r2_probe_hit_vec_3,r2_probe_hit_vec_2,r2_probe_hit_vec_1,r2_probe_hit_vec_0}; // @[ReplacePipe.scala 225:63]
  wire [3:0] r2_write_waymask_hi = {r2_probe_hit_vec_7,r2_probe_hit_vec_6,r2_probe_hit_vec_5,r2_probe_hit_vec_4}; // @[ReplacePipe.scala 225:63]
  wire  _r3_valid_T = _r2_ready_T & r2_req_voluntary; // @[ReplacePipe.scala 255:66]
  reg  r3_valid; // @[ICache.scala 98:25]
  reg  r3_fire_REG; // @[ReplacePipe.scala 258:40]
  reg  r3_release_need_send; // @[Reg.scala 16:16]
  wire  r3_fire = r3_valid & r3_fire_REG & r3_release_need_send | r3_valid & ~r3_release_need_send; // @[ReplacePipe.scala 258:85]
  wire  _GEN_107 = r3_fire ? 1'h0 : r3_valid; // @[ICache.scala 101:{43,51} 98:25]
  reg [38:0] r3_req_vaddr; // @[Reg.scala 16:16]
  reg [4:0] r3_req_id; // @[Reg.scala 16:16]
  assign io_pipe_req_ready = _r0_ready_T & r1_ready; // @[ReplacePipe.scala 106:65]
  assign io_meta_read_valid = r0_valid; // @[ReplacePipe.scala 101:30]
  assign io_meta_read_bits_vSetIdx_0 = r0_req_vaddr[11:6]; // @[L1Cache.scala 81:33]
  assign io_data_read_valid = r0_valid; // @[ReplacePipe.scala 95:37]
  assign io_data_read_bits_0_vSetIdx_0 = r0_req_vaddr[11:6]; // @[L1Cache.scala 81:33]
  assign io_data_read_bits_1_vSetIdx_0 = r0_req_vaddr[11:6]; // @[L1Cache.scala 81:33]
  assign io_data_read_bits_2_vSetIdx_0 = r0_req_vaddr[11:6]; // @[L1Cache.scala 81:33]
  assign io_data_read_bits_3_vSetIdx_0 = r0_req_vaddr[11:6]; // @[L1Cache.scala 81:33]
  assign io_error_source_tag = io_error_source_tag_REG_1; // @[ReplacePipe.scala 196:33]
  assign io_error_source_data = io_error_source_data_REG; // @[ReplacePipe.scala 197:33]
  assign io_error_opType_probe = io_error_opType_probe_REG_1; // @[ReplacePipe.scala 202:33]
  assign io_error_opType_release = io_error_opType_release_REG_1; // @[ReplacePipe.scala 201:33]
  assign io_error_paddr = io_error_paddr_REG_1; // @[ReplacePipe.scala 195:33]
  assign io_error_report_to_beu = io_error_report_to_beu_REG_2; // @[ReplacePipe.scala 194:33]
  assign io_error_valid = io_error_valid_REG_2; // @[ReplacePipe.scala 193:33]
  assign io_meta_write_valid = _r2_ready_T & _io_error_opType_probe_T; // @[ReplacePipe.scala 228:34]
  assign io_meta_write_bits_virIdx = r2_req_vaddr[11:6]; // @[L1Cache.scala 81:33]
  assign io_meta_write_bits_phyTag = r2_probe_hit_ptag; // @[ICacheBundle.scala 61:18]
  assign io_meta_write_bits_coh_state = _T_124 ? 2'h2 : _T_123; // @[Misc.scala 37:63]
  assign io_meta_write_bits_waymask = {r2_write_waymask_hi,r2_write_waymask_lo}; // @[ReplacePipe.scala 229:123]
  assign io_meta_write_bits_bankIdx = r2_req_vaddr[6]; // @[ReplacePipe.scala 229:152]
  assign io_release_req_valid = r2_valid & (_io_error_opType_probe_T | release_need_send); // @[ReplacePipe.scala 232:45]
  assign io_release_req_bits_addr = _io_error_opType_probe_T ? r2_req_paddr : r2_release_addr; // @[ReplacePipe.scala 218:21]
  assign io_release_req_bits_param = _io_error_opType_probe_T ? probe_shrink_param : release_shrink_param; // @[ReplacePipe.scala 219:21]
  assign io_release_req_bits_voluntary = r2_req_voluntary; // @[ReplacePipe.scala 235:33]
  assign io_release_req_bits_hasData = _io_error_opType_probe_T & _r2_hasData_T_1 & (r2_req_needData |
    probe_has_dirty_data) | r2_req_voluntary; // @[ReplacePipe.scala 220:110]
  assign io_release_req_bits_dirty = release_has_dirty_data | probe_has_dirty_data; // @[ReplacePipe.scala 238:59]
  assign io_release_req_bits_data = _io_error_opType_probe_T ? r2_probe_hit_data : r2_release_data; // @[ReplacePipe.scala 221:21]
  assign io_pipe_resp_valid = r3_valid & r3_fire_REG & r3_release_need_send | r3_valid & ~r3_release_need_send; // @[ReplacePipe.scala 258:85]
  assign io_pipe_resp_bits = r3_req_id; // @[ReplacePipe.scala 263:22]
  assign io_status_r0_set_valid = r0_valid; // @[ReplacePipe.scala 108:26]
  assign io_status_r0_set_bits = r0_req_vaddr[11:6]; // @[L1Cache.scala 81:33]
  assign io_status_r1_set_valid = r1_valid; // @[ReplacePipe.scala 146:26]
  assign io_status_r1_set_bits = r1_req_vaddr[11:6]; // @[L1Cache.scala 81:33]
  assign io_status_r2_set_valid = r2_valid; // @[ReplacePipe.scala 246:26]
  assign io_status_r2_set_bits = r2_req_vaddr[11:6]; // @[L1Cache.scala 81:33]
  assign io_status_r3_set_valid = r3_valid; // @[ReplacePipe.scala 265:26]
  assign io_status_r3_set_bits = r3_req_vaddr[11:6]; // @[L1Cache.scala 81:33]
  always @(posedge clock) begin
    if (_r0_valid_T) begin // @[Reg.scala 17:18]
      r0_req_paddr <= io_pipe_req_bits_paddr; // @[Reg.scala 17:22]
    end
    if (_r0_valid_T) begin // @[Reg.scala 17:18]
      r0_req_vaddr <= io_pipe_req_bits_vaddr; // @[Reg.scala 17:22]
    end
    if (_r0_valid_T) begin // @[Reg.scala 17:18]
      r0_req_param <= io_pipe_req_bits_param; // @[Reg.scala 17:22]
    end
    if (_r0_valid_T) begin // @[Reg.scala 17:18]
      r0_req_voluntary <= io_pipe_req_bits_voluntary; // @[Reg.scala 17:22]
    end
    if (_r0_valid_T) begin // @[Reg.scala 17:18]
      r0_req_needData <= io_pipe_req_bits_needData; // @[Reg.scala 17:22]
    end
    if (_r0_valid_T) begin // @[Reg.scala 17:18]
      r0_req_waymask <= io_pipe_req_bits_waymask; // @[Reg.scala 17:22]
    end
    if (_r0_valid_T) begin // @[Reg.scala 17:18]
      r0_req_id <= io_pipe_req_bits_id; // @[Reg.scala 17:22]
    end
    if (r0_fire) begin // @[Reg.scala 17:18]
      r1_req_paddr <= r0_req_paddr; // @[Reg.scala 17:22]
    end
    if (r0_fire) begin // @[Reg.scala 17:18]
      r1_req_vaddr <= r0_req_vaddr; // @[Reg.scala 17:22]
    end
    if (r0_fire) begin // @[Reg.scala 17:18]
      r1_req_param <= r0_req_param; // @[Reg.scala 17:22]
    end
    if (r0_fire) begin // @[Reg.scala 17:18]
      r1_req_voluntary <= r0_req_voluntary; // @[Reg.scala 17:22]
    end
    if (r0_fire) begin // @[Reg.scala 17:18]
      r1_req_needData <= r0_req_needData; // @[Reg.scala 17:22]
    end
    if (r0_fire) begin // @[Reg.scala 17:18]
      r1_req_waymask <= r0_req_waymask; // @[Reg.scala 17:22]
    end
    if (r0_fire) begin // @[Reg.scala 17:18]
      r1_req_id <= r0_req_id; // @[Reg.scala 17:22]
    end
    r1_meta_ptags_REG <= r0_valid & r0_ready; // @[ReplacePipe.scala 92:24]
    if (r1_meta_ptags_REG) begin // @[Reg.scala 17:18]
      r1_meta_ptags_r0 <= io_meta_response_metaData_0_0_tag; // @[Reg.scala 17:22]
    end
    if (r1_meta_ptags_REG) begin // @[Reg.scala 17:18]
      r1_meta_ptags_r1 <= io_meta_response_metaData_0_1_tag; // @[Reg.scala 17:22]
    end
    if (r1_meta_ptags_REG) begin // @[Reg.scala 17:18]
      r1_meta_ptags_r2 <= io_meta_response_metaData_0_2_tag; // @[Reg.scala 17:22]
    end
    if (r1_meta_ptags_REG) begin // @[Reg.scala 17:18]
      r1_meta_ptags_r3 <= io_meta_response_metaData_0_3_tag; // @[Reg.scala 17:22]
    end
    if (r1_meta_ptags_REG) begin // @[Reg.scala 17:18]
      r1_meta_ptags_r4 <= io_meta_response_metaData_0_4_tag; // @[Reg.scala 17:22]
    end
    if (r1_meta_ptags_REG) begin // @[Reg.scala 17:18]
      r1_meta_ptags_r5 <= io_meta_response_metaData_0_5_tag; // @[Reg.scala 17:22]
    end
    if (r1_meta_ptags_REG) begin // @[Reg.scala 17:18]
      r1_meta_ptags_r6 <= io_meta_response_metaData_0_6_tag; // @[Reg.scala 17:22]
    end
    if (r1_meta_ptags_REG) begin // @[Reg.scala 17:18]
      r1_meta_ptags_r7 <= io_meta_response_metaData_0_7_tag; // @[Reg.scala 17:22]
    end
    r1_meta_cohs_REG <= r0_valid & r0_ready; // @[ReplacePipe.scala 92:24]
    if (r1_meta_cohs_REG) begin // @[Reg.scala 17:18]
      r1_meta_cohs_r0_state <= io_meta_response_metaData_0_0_coh_state; // @[Reg.scala 17:22]
    end
    if (r1_meta_cohs_REG) begin // @[Reg.scala 17:18]
      r1_meta_cohs_r1_state <= io_meta_response_metaData_0_1_coh_state; // @[Reg.scala 17:22]
    end
    if (r1_meta_cohs_REG) begin // @[Reg.scala 17:18]
      r1_meta_cohs_r2_state <= io_meta_response_metaData_0_2_coh_state; // @[Reg.scala 17:22]
    end
    if (r1_meta_cohs_REG) begin // @[Reg.scala 17:18]
      r1_meta_cohs_r3_state <= io_meta_response_metaData_0_3_coh_state; // @[Reg.scala 17:22]
    end
    if (r1_meta_cohs_REG) begin // @[Reg.scala 17:18]
      r1_meta_cohs_r4_state <= io_meta_response_metaData_0_4_coh_state; // @[Reg.scala 17:22]
    end
    if (r1_meta_cohs_REG) begin // @[Reg.scala 17:18]
      r1_meta_cohs_r5_state <= io_meta_response_metaData_0_5_coh_state; // @[Reg.scala 17:22]
    end
    if (r1_meta_cohs_REG) begin // @[Reg.scala 17:18]
      r1_meta_cohs_r6_state <= io_meta_response_metaData_0_6_coh_state; // @[Reg.scala 17:22]
    end
    if (r1_meta_cohs_REG) begin // @[Reg.scala 17:18]
      r1_meta_cohs_r7_state <= io_meta_response_metaData_0_7_coh_state; // @[Reg.scala 17:22]
    end
    r1_meta_errors_REG <= r0_valid & r0_ready; // @[ReplacePipe.scala 92:24]
    if (r1_meta_errors_REG) begin // @[Reg.scala 17:18]
      r1_meta_errors_r0 <= io_meta_response_errors_0_0; // @[Reg.scala 17:22]
    end
    if (r1_meta_errors_REG) begin // @[Reg.scala 17:18]
      r1_meta_errors_r1 <= io_meta_response_errors_0_1; // @[Reg.scala 17:22]
    end
    if (r1_meta_errors_REG) begin // @[Reg.scala 17:18]
      r1_meta_errors_r2 <= io_meta_response_errors_0_2; // @[Reg.scala 17:22]
    end
    if (r1_meta_errors_REG) begin // @[Reg.scala 17:18]
      r1_meta_errors_r3 <= io_meta_response_errors_0_3; // @[Reg.scala 17:22]
    end
    if (r1_meta_errors_REG) begin // @[Reg.scala 17:18]
      r1_meta_errors_r4 <= io_meta_response_errors_0_4; // @[Reg.scala 17:22]
    end
    if (r1_meta_errors_REG) begin // @[Reg.scala 17:18]
      r1_meta_errors_r5 <= io_meta_response_errors_0_5; // @[Reg.scala 17:22]
    end
    if (r1_meta_errors_REG) begin // @[Reg.scala 17:18]
      r1_meta_errors_r6 <= io_meta_response_errors_0_6; // @[Reg.scala 17:22]
    end
    if (r1_meta_errors_REG) begin // @[Reg.scala 17:18]
      r1_meta_errors_r7 <= io_meta_response_errors_0_7; // @[Reg.scala 17:22]
    end
    r1_data_cacheline_REG <= r0_valid & r0_ready; // @[ReplacePipe.scala 92:24]
    if (r1_data_cacheline_REG) begin // @[Reg.scala 17:18]
      r1_data_cacheline_r0 <= io_data_response_datas_0_0; // @[Reg.scala 17:22]
    end
    if (r1_data_cacheline_REG) begin // @[Reg.scala 17:18]
      r1_data_cacheline_r1 <= io_data_response_datas_0_1; // @[Reg.scala 17:22]
    end
    if (r1_data_cacheline_REG) begin // @[Reg.scala 17:18]
      r1_data_cacheline_r2 <= io_data_response_datas_0_2; // @[Reg.scala 17:22]
    end
    if (r1_data_cacheline_REG) begin // @[Reg.scala 17:18]
      r1_data_cacheline_r3 <= io_data_response_datas_0_3; // @[Reg.scala 17:22]
    end
    if (r1_data_cacheline_REG) begin // @[Reg.scala 17:18]
      r1_data_cacheline_r4 <= io_data_response_datas_0_4; // @[Reg.scala 17:22]
    end
    if (r1_data_cacheline_REG) begin // @[Reg.scala 17:18]
      r1_data_cacheline_r5 <= io_data_response_datas_0_5; // @[Reg.scala 17:22]
    end
    if (r1_data_cacheline_REG) begin // @[Reg.scala 17:18]
      r1_data_cacheline_r6 <= io_data_response_datas_0_6; // @[Reg.scala 17:22]
    end
    if (r1_data_cacheline_REG) begin // @[Reg.scala 17:18]
      r1_data_cacheline_r7 <= io_data_response_datas_0_7; // @[Reg.scala 17:22]
    end
    r1_data_errorBits_REG <= r0_valid & r0_ready; // @[ReplacePipe.scala 92:24]
    if (r1_data_errorBits_REG) begin // @[Reg.scala 17:18]
      r1_data_errorBits_r0 <= io_data_response_codes_0_0; // @[Reg.scala 17:22]
    end
    if (r1_data_errorBits_REG) begin // @[Reg.scala 17:18]
      r1_data_errorBits_r1 <= io_data_response_codes_0_1; // @[Reg.scala 17:22]
    end
    if (r1_data_errorBits_REG) begin // @[Reg.scala 17:18]
      r1_data_errorBits_r2 <= io_data_response_codes_0_2; // @[Reg.scala 17:22]
    end
    if (r1_data_errorBits_REG) begin // @[Reg.scala 17:18]
      r1_data_errorBits_r3 <= io_data_response_codes_0_3; // @[Reg.scala 17:22]
    end
    if (r1_data_errorBits_REG) begin // @[Reg.scala 17:18]
      r1_data_errorBits_r4 <= io_data_response_codes_0_4; // @[Reg.scala 17:22]
    end
    if (r1_data_errorBits_REG) begin // @[Reg.scala 17:18]
      r1_data_errorBits_r5 <= io_data_response_codes_0_5; // @[Reg.scala 17:22]
    end
    if (r1_data_errorBits_REG) begin // @[Reg.scala 17:18]
      r1_data_errorBits_r6 <= io_data_response_codes_0_6; // @[Reg.scala 17:22]
    end
    if (r1_data_errorBits_REG) begin // @[Reg.scala 17:18]
      r1_data_errorBits_r7 <= io_data_response_codes_0_7; // @[Reg.scala 17:22]
    end
    if (r1_fire) begin // @[Reg.scala 17:18]
      r2_req_paddr <= r1_req_paddr; // @[Reg.scala 17:22]
    end
    if (r1_fire) begin // @[Reg.scala 17:18]
      r2_req_vaddr <= r1_req_vaddr; // @[Reg.scala 17:22]
    end
    if (r1_fire) begin // @[Reg.scala 17:18]
      r2_req_param <= r1_req_param; // @[Reg.scala 17:22]
    end
    if (r1_fire) begin // @[Reg.scala 17:18]
      r2_req_voluntary <= r1_req_voluntary; // @[Reg.scala 17:22]
    end
    if (r1_fire) begin // @[Reg.scala 17:18]
      r2_req_needData <= r1_req_needData; // @[Reg.scala 17:22]
    end
    if (r1_fire) begin // @[Reg.scala 17:18]
      r2_req_waymask <= r1_req_waymask; // @[Reg.scala 17:22]
    end
    if (r1_fire) begin // @[Reg.scala 17:18]
      r2_req_id <= r1_req_id; // @[Reg.scala 17:22]
    end
    if (r1_fire) begin // @[Reg.scala 17:18]
      if (r1_data_cacheline_REG) begin // @[Reg.scala 17:18]
        r2_data_cacheline_0 <= io_data_response_datas_0_0; // @[Reg.scala 17:22]
      end else begin
        r2_data_cacheline_0 <= r1_data_cacheline_r0; // @[Reg.scala 16:16]
      end
    end
    if (r1_fire) begin // @[Reg.scala 17:18]
      if (r1_data_cacheline_REG) begin // @[Reg.scala 17:18]
        r2_data_cacheline_1 <= io_data_response_datas_0_1; // @[Reg.scala 17:22]
      end else begin
        r2_data_cacheline_1 <= r1_data_cacheline_r1; // @[Reg.scala 16:16]
      end
    end
    if (r1_fire) begin // @[Reg.scala 17:18]
      if (r1_data_cacheline_REG) begin // @[Reg.scala 17:18]
        r2_data_cacheline_2 <= io_data_response_datas_0_2; // @[Reg.scala 17:22]
      end else begin
        r2_data_cacheline_2 <= r1_data_cacheline_r2; // @[Reg.scala 16:16]
      end
    end
    if (r1_fire) begin // @[Reg.scala 17:18]
      if (r1_data_cacheline_REG) begin // @[Reg.scala 17:18]
        r2_data_cacheline_3 <= io_data_response_datas_0_3; // @[Reg.scala 17:22]
      end else begin
        r2_data_cacheline_3 <= r1_data_cacheline_r3; // @[Reg.scala 16:16]
      end
    end
    if (r1_fire) begin // @[Reg.scala 17:18]
      if (r1_data_cacheline_REG) begin // @[Reg.scala 17:18]
        r2_data_cacheline_4 <= io_data_response_datas_0_4; // @[Reg.scala 17:22]
      end else begin
        r2_data_cacheline_4 <= r1_data_cacheline_r4; // @[Reg.scala 16:16]
      end
    end
    if (r1_fire) begin // @[Reg.scala 17:18]
      if (r1_data_cacheline_REG) begin // @[Reg.scala 17:18]
        r2_data_cacheline_5 <= io_data_response_datas_0_5; // @[Reg.scala 17:22]
      end else begin
        r2_data_cacheline_5 <= r1_data_cacheline_r5; // @[Reg.scala 16:16]
      end
    end
    if (r1_fire) begin // @[Reg.scala 17:18]
      if (r1_data_cacheline_REG) begin // @[Reg.scala 17:18]
        r2_data_cacheline_6 <= io_data_response_datas_0_6; // @[Reg.scala 17:22]
      end else begin
        r2_data_cacheline_6 <= r1_data_cacheline_r6; // @[Reg.scala 16:16]
      end
    end
    if (r1_fire) begin // @[Reg.scala 17:18]
      if (r1_data_cacheline_REG) begin // @[Reg.scala 17:18]
        r2_data_cacheline_7 <= io_data_response_datas_0_7; // @[Reg.scala 17:22]
      end else begin
        r2_data_cacheline_7 <= r1_data_cacheline_r7; // @[Reg.scala 16:16]
      end
    end
    if (r1_fire) begin // @[Reg.scala 17:18]
      r2_probe_hit_ptag <= probe_phy_tag; // @[Reg.scala 17:22]
    end
    if (r1_fire) begin // @[Reg.scala 17:18]
      r2_probe_hit_vec_0 <= probe_hit_vec_0; // @[Reg.scala 17:22]
    end
    if (r1_fire) begin // @[Reg.scala 17:18]
      r2_probe_hit_vec_1 <= probe_hit_vec_1; // @[Reg.scala 17:22]
    end
    if (r1_fire) begin // @[Reg.scala 17:18]
      r2_probe_hit_vec_2 <= probe_hit_vec_2; // @[Reg.scala 17:22]
    end
    if (r1_fire) begin // @[Reg.scala 17:18]
      r2_probe_hit_vec_3 <= probe_hit_vec_3; // @[Reg.scala 17:22]
    end
    if (r1_fire) begin // @[Reg.scala 17:18]
      r2_probe_hit_vec_4 <= probe_hit_vec_4; // @[Reg.scala 17:22]
    end
    if (r1_fire) begin // @[Reg.scala 17:18]
      r2_probe_hit_vec_5 <= probe_hit_vec_5; // @[Reg.scala 17:22]
    end
    if (r1_fire) begin // @[Reg.scala 17:18]
      r2_probe_hit_vec_6 <= probe_hit_vec_6; // @[Reg.scala 17:22]
    end
    if (r1_fire) begin // @[Reg.scala 17:18]
      r2_probe_hit_vec_7 <= probe_hit_vec_7; // @[Reg.scala 17:22]
    end
    if (r1_fire) begin // @[Reg.scala 17:18]
      r2_probe_hit_coh_state <= probe_hit_coh_state; // @[Reg.scala 17:22]
    end
    if (r1_fire) begin // @[Reg.scala 17:18]
      if (r1_meta_errors_REG) begin // @[Reg.scala 17:18]
        r2_meta_errors_0 <= io_meta_response_errors_0_0; // @[Reg.scala 17:22]
      end else begin
        r2_meta_errors_0 <= r1_meta_errors_r0; // @[Reg.scala 16:16]
      end
    end
    if (r1_fire) begin // @[Reg.scala 17:18]
      if (r1_meta_errors_REG) begin // @[Reg.scala 17:18]
        r2_meta_errors_1 <= io_meta_response_errors_0_1; // @[Reg.scala 17:22]
      end else begin
        r2_meta_errors_1 <= r1_meta_errors_r1; // @[Reg.scala 16:16]
      end
    end
    if (r1_fire) begin // @[Reg.scala 17:18]
      if (r1_meta_errors_REG) begin // @[Reg.scala 17:18]
        r2_meta_errors_2 <= io_meta_response_errors_0_2; // @[Reg.scala 17:22]
      end else begin
        r2_meta_errors_2 <= r1_meta_errors_r2; // @[Reg.scala 16:16]
      end
    end
    if (r1_fire) begin // @[Reg.scala 17:18]
      if (r1_meta_errors_REG) begin // @[Reg.scala 17:18]
        r2_meta_errors_3 <= io_meta_response_errors_0_3; // @[Reg.scala 17:22]
      end else begin
        r2_meta_errors_3 <= r1_meta_errors_r3; // @[Reg.scala 16:16]
      end
    end
    if (r1_fire) begin // @[Reg.scala 17:18]
      if (r1_meta_errors_REG) begin // @[Reg.scala 17:18]
        r2_meta_errors_4 <= io_meta_response_errors_0_4; // @[Reg.scala 17:22]
      end else begin
        r2_meta_errors_4 <= r1_meta_errors_r4; // @[Reg.scala 16:16]
      end
    end
    if (r1_fire) begin // @[Reg.scala 17:18]
      if (r1_meta_errors_REG) begin // @[Reg.scala 17:18]
        r2_meta_errors_5 <= io_meta_response_errors_0_5; // @[Reg.scala 17:22]
      end else begin
        r2_meta_errors_5 <= r1_meta_errors_r5; // @[Reg.scala 16:16]
      end
    end
    if (r1_fire) begin // @[Reg.scala 17:18]
      if (r1_meta_errors_REG) begin // @[Reg.scala 17:18]
        r2_meta_errors_6 <= io_meta_response_errors_0_6; // @[Reg.scala 17:22]
      end else begin
        r2_meta_errors_6 <= r1_meta_errors_r6; // @[Reg.scala 16:16]
      end
    end
    if (r1_fire) begin // @[Reg.scala 17:18]
      if (r1_meta_errors_REG) begin // @[Reg.scala 17:18]
        r2_meta_errors_7 <= io_meta_response_errors_0_7; // @[Reg.scala 17:22]
      end else begin
        r2_meta_errors_7 <= r1_meta_errors_r7; // @[Reg.scala 16:16]
      end
    end
    if (r1_fire) begin // @[Reg.scala 17:18]
      if (r1_data_errorBits_REG) begin // @[Reg.scala 17:18]
        r2_data_errorBits_0 <= io_data_response_codes_0_0; // @[Reg.scala 17:22]
      end else begin
        r2_data_errorBits_0 <= r1_data_errorBits_r0; // @[Reg.scala 16:16]
      end
    end
    if (r1_fire) begin // @[Reg.scala 17:18]
      if (r1_data_errorBits_REG) begin // @[Reg.scala 17:18]
        r2_data_errorBits_1 <= io_data_response_codes_0_1; // @[Reg.scala 17:22]
      end else begin
        r2_data_errorBits_1 <= r1_data_errorBits_r1; // @[Reg.scala 16:16]
      end
    end
    if (r1_fire) begin // @[Reg.scala 17:18]
      if (r1_data_errorBits_REG) begin // @[Reg.scala 17:18]
        r2_data_errorBits_2 <= io_data_response_codes_0_2; // @[Reg.scala 17:22]
      end else begin
        r2_data_errorBits_2 <= r1_data_errorBits_r2; // @[Reg.scala 16:16]
      end
    end
    if (r1_fire) begin // @[Reg.scala 17:18]
      if (r1_data_errorBits_REG) begin // @[Reg.scala 17:18]
        r2_data_errorBits_3 <= io_data_response_codes_0_3; // @[Reg.scala 17:22]
      end else begin
        r2_data_errorBits_3 <= r1_data_errorBits_r3; // @[Reg.scala 16:16]
      end
    end
    if (r1_fire) begin // @[Reg.scala 17:18]
      if (r1_data_errorBits_REG) begin // @[Reg.scala 17:18]
        r2_data_errorBits_4 <= io_data_response_codes_0_4; // @[Reg.scala 17:22]
      end else begin
        r2_data_errorBits_4 <= r1_data_errorBits_r4; // @[Reg.scala 16:16]
      end
    end
    if (r1_fire) begin // @[Reg.scala 17:18]
      if (r1_data_errorBits_REG) begin // @[Reg.scala 17:18]
        r2_data_errorBits_5 <= io_data_response_codes_0_5; // @[Reg.scala 17:22]
      end else begin
        r2_data_errorBits_5 <= r1_data_errorBits_r5; // @[Reg.scala 16:16]
      end
    end
    if (r1_fire) begin // @[Reg.scala 17:18]
      if (r1_data_errorBits_REG) begin // @[Reg.scala 17:18]
        r2_data_errorBits_6 <= io_data_response_codes_0_6; // @[Reg.scala 17:22]
      end else begin
        r2_data_errorBits_6 <= r1_data_errorBits_r6; // @[Reg.scala 16:16]
      end
    end
    if (r1_fire) begin // @[Reg.scala 17:18]
      if (r1_data_errorBits_REG) begin // @[Reg.scala 17:18]
        r2_data_errorBits_7 <= io_data_response_codes_0_7; // @[Reg.scala 17:22]
      end else begin
        r2_data_errorBits_7 <= r1_data_errorBits_r7; // @[Reg.scala 16:16]
      end
    end
    r2_data_errors_0_REG <= r1_valid & r2_ready; // @[ReplacePipe.scala 119:24]
    r2_data_errors_0_REG_1 <= r2_data_errors_0_REG; // @[ReplacePipe.scala 186:57]
    r2_data_errors_0_REG_2_0 <= ^data_full_wayBits_0_0; // @[ECC.scala 87:27]
    r2_data_errors_0_REG_2_1 <= ^data_full_wayBits_0_1; // @[ECC.scala 87:27]
    r2_data_errors_0_REG_2_2 <= ^data_full_wayBits_0_2; // @[ECC.scala 87:27]
    r2_data_errors_0_REG_2_3 <= ^data_full_wayBits_0_3; // @[ECC.scala 87:27]
    r2_data_errors_0_REG_2_4 <= ^data_full_wayBits_0_4; // @[ECC.scala 87:27]
    r2_data_errors_0_REG_2_5 <= ^data_full_wayBits_0_5; // @[ECC.scala 87:27]
    r2_data_errors_0_REG_2_6 <= ^data_full_wayBits_0_6; // @[ECC.scala 87:27]
    r2_data_errors_0_REG_2_7 <= ^data_full_wayBits_0_7; // @[ECC.scala 87:27]
    r2_data_errors_0_REG_2_8 <= ^data_full_wayBits_0_8; // @[ECC.scala 87:27]
    r2_data_errors_0_REG_2_9 <= ^data_full_wayBits_0_9; // @[ECC.scala 87:27]
    r2_data_errors_0_REG_2_10 <= ^data_full_wayBits_0_10; // @[ECC.scala 87:27]
    r2_data_errors_0_REG_2_11 <= ^data_full_wayBits_0_11; // @[ECC.scala 87:27]
    r2_data_errors_0_REG_2_12 <= ^data_full_wayBits_0_12; // @[ECC.scala 87:27]
    r2_data_errors_0_REG_2_13 <= ^data_full_wayBits_0_13; // @[ECC.scala 87:27]
    r2_data_errors_0_REG_2_14 <= ^data_full_wayBits_0_14; // @[ECC.scala 87:27]
    r2_data_errors_0_REG_2_15 <= ^data_full_wayBits_0_15; // @[ECC.scala 87:27]
    r2_data_errors_0_REG_2_16 <= ^data_full_wayBits_0_16; // @[ECC.scala 87:27]
    r2_data_errors_0_REG_2_17 <= ^data_full_wayBits_0_17; // @[ECC.scala 87:27]
    r2_data_errors_0_REG_2_18 <= ^data_full_wayBits_0_18; // @[ECC.scala 87:27]
    r2_data_errors_0_REG_2_19 <= ^data_full_wayBits_0_19; // @[ECC.scala 87:27]
    r2_data_errors_0_REG_2_20 <= ^data_full_wayBits_0_20; // @[ECC.scala 87:27]
    r2_data_errors_0_REG_2_21 <= ^data_full_wayBits_0_21; // @[ECC.scala 87:27]
    r2_data_errors_0_REG_2_22 <= ^data_full_wayBits_0_22; // @[ECC.scala 87:27]
    r2_data_errors_0_REG_2_23 <= ^data_full_wayBits_0_23; // @[ECC.scala 87:27]
    r2_data_errors_0_REG_2_24 <= ^data_full_wayBits_0_24; // @[ECC.scala 87:27]
    r2_data_errors_0_REG_2_25 <= ^data_full_wayBits_0_25; // @[ECC.scala 87:27]
    r2_data_errors_0_REG_2_26 <= ^data_full_wayBits_0_26; // @[ECC.scala 87:27]
    r2_data_errors_0_REG_2_27 <= ^data_full_wayBits_0_27; // @[ECC.scala 87:27]
    r2_data_errors_0_REG_2_28 <= ^data_full_wayBits_0_28; // @[ECC.scala 87:27]
    r2_data_errors_0_REG_2_29 <= ^data_full_wayBits_0_29; // @[ECC.scala 87:27]
    r2_data_errors_0_REG_2_30 <= ^data_full_wayBits_0_30; // @[ECC.scala 87:27]
    r2_data_errors_0_REG_2_31 <= ^data_full_wayBits_0_31; // @[ECC.scala 87:27]
    r2_data_errors_1_REG <= r1_valid & r2_ready; // @[ReplacePipe.scala 119:24]
    r2_data_errors_1_REG_1 <= r2_data_errors_1_REG; // @[ReplacePipe.scala 186:57]
    r2_data_errors_1_REG_2_0 <= ^data_full_wayBits_1_0; // @[ECC.scala 87:27]
    r2_data_errors_1_REG_2_1 <= ^data_full_wayBits_1_1; // @[ECC.scala 87:27]
    r2_data_errors_1_REG_2_2 <= ^data_full_wayBits_1_2; // @[ECC.scala 87:27]
    r2_data_errors_1_REG_2_3 <= ^data_full_wayBits_1_3; // @[ECC.scala 87:27]
    r2_data_errors_1_REG_2_4 <= ^data_full_wayBits_1_4; // @[ECC.scala 87:27]
    r2_data_errors_1_REG_2_5 <= ^data_full_wayBits_1_5; // @[ECC.scala 87:27]
    r2_data_errors_1_REG_2_6 <= ^data_full_wayBits_1_6; // @[ECC.scala 87:27]
    r2_data_errors_1_REG_2_7 <= ^data_full_wayBits_1_7; // @[ECC.scala 87:27]
    r2_data_errors_1_REG_2_8 <= ^data_full_wayBits_1_8; // @[ECC.scala 87:27]
    r2_data_errors_1_REG_2_9 <= ^data_full_wayBits_1_9; // @[ECC.scala 87:27]
    r2_data_errors_1_REG_2_10 <= ^data_full_wayBits_1_10; // @[ECC.scala 87:27]
    r2_data_errors_1_REG_2_11 <= ^data_full_wayBits_1_11; // @[ECC.scala 87:27]
    r2_data_errors_1_REG_2_12 <= ^data_full_wayBits_1_12; // @[ECC.scala 87:27]
    r2_data_errors_1_REG_2_13 <= ^data_full_wayBits_1_13; // @[ECC.scala 87:27]
    r2_data_errors_1_REG_2_14 <= ^data_full_wayBits_1_14; // @[ECC.scala 87:27]
    r2_data_errors_1_REG_2_15 <= ^data_full_wayBits_1_15; // @[ECC.scala 87:27]
    r2_data_errors_1_REG_2_16 <= ^data_full_wayBits_1_16; // @[ECC.scala 87:27]
    r2_data_errors_1_REG_2_17 <= ^data_full_wayBits_1_17; // @[ECC.scala 87:27]
    r2_data_errors_1_REG_2_18 <= ^data_full_wayBits_1_18; // @[ECC.scala 87:27]
    r2_data_errors_1_REG_2_19 <= ^data_full_wayBits_1_19; // @[ECC.scala 87:27]
    r2_data_errors_1_REG_2_20 <= ^data_full_wayBits_1_20; // @[ECC.scala 87:27]
    r2_data_errors_1_REG_2_21 <= ^data_full_wayBits_1_21; // @[ECC.scala 87:27]
    r2_data_errors_1_REG_2_22 <= ^data_full_wayBits_1_22; // @[ECC.scala 87:27]
    r2_data_errors_1_REG_2_23 <= ^data_full_wayBits_1_23; // @[ECC.scala 87:27]
    r2_data_errors_1_REG_2_24 <= ^data_full_wayBits_1_24; // @[ECC.scala 87:27]
    r2_data_errors_1_REG_2_25 <= ^data_full_wayBits_1_25; // @[ECC.scala 87:27]
    r2_data_errors_1_REG_2_26 <= ^data_full_wayBits_1_26; // @[ECC.scala 87:27]
    r2_data_errors_1_REG_2_27 <= ^data_full_wayBits_1_27; // @[ECC.scala 87:27]
    r2_data_errors_1_REG_2_28 <= ^data_full_wayBits_1_28; // @[ECC.scala 87:27]
    r2_data_errors_1_REG_2_29 <= ^data_full_wayBits_1_29; // @[ECC.scala 87:27]
    r2_data_errors_1_REG_2_30 <= ^data_full_wayBits_1_30; // @[ECC.scala 87:27]
    r2_data_errors_1_REG_2_31 <= ^data_full_wayBits_1_31; // @[ECC.scala 87:27]
    r2_data_errors_2_REG <= r1_valid & r2_ready; // @[ReplacePipe.scala 119:24]
    r2_data_errors_2_REG_1 <= r2_data_errors_2_REG; // @[ReplacePipe.scala 186:57]
    r2_data_errors_2_REG_2_0 <= ^data_full_wayBits_2_0; // @[ECC.scala 87:27]
    r2_data_errors_2_REG_2_1 <= ^data_full_wayBits_2_1; // @[ECC.scala 87:27]
    r2_data_errors_2_REG_2_2 <= ^data_full_wayBits_2_2; // @[ECC.scala 87:27]
    r2_data_errors_2_REG_2_3 <= ^data_full_wayBits_2_3; // @[ECC.scala 87:27]
    r2_data_errors_2_REG_2_4 <= ^data_full_wayBits_2_4; // @[ECC.scala 87:27]
    r2_data_errors_2_REG_2_5 <= ^data_full_wayBits_2_5; // @[ECC.scala 87:27]
    r2_data_errors_2_REG_2_6 <= ^data_full_wayBits_2_6; // @[ECC.scala 87:27]
    r2_data_errors_2_REG_2_7 <= ^data_full_wayBits_2_7; // @[ECC.scala 87:27]
    r2_data_errors_2_REG_2_8 <= ^data_full_wayBits_2_8; // @[ECC.scala 87:27]
    r2_data_errors_2_REG_2_9 <= ^data_full_wayBits_2_9; // @[ECC.scala 87:27]
    r2_data_errors_2_REG_2_10 <= ^data_full_wayBits_2_10; // @[ECC.scala 87:27]
    r2_data_errors_2_REG_2_11 <= ^data_full_wayBits_2_11; // @[ECC.scala 87:27]
    r2_data_errors_2_REG_2_12 <= ^data_full_wayBits_2_12; // @[ECC.scala 87:27]
    r2_data_errors_2_REG_2_13 <= ^data_full_wayBits_2_13; // @[ECC.scala 87:27]
    r2_data_errors_2_REG_2_14 <= ^data_full_wayBits_2_14; // @[ECC.scala 87:27]
    r2_data_errors_2_REG_2_15 <= ^data_full_wayBits_2_15; // @[ECC.scala 87:27]
    r2_data_errors_2_REG_2_16 <= ^data_full_wayBits_2_16; // @[ECC.scala 87:27]
    r2_data_errors_2_REG_2_17 <= ^data_full_wayBits_2_17; // @[ECC.scala 87:27]
    r2_data_errors_2_REG_2_18 <= ^data_full_wayBits_2_18; // @[ECC.scala 87:27]
    r2_data_errors_2_REG_2_19 <= ^data_full_wayBits_2_19; // @[ECC.scala 87:27]
    r2_data_errors_2_REG_2_20 <= ^data_full_wayBits_2_20; // @[ECC.scala 87:27]
    r2_data_errors_2_REG_2_21 <= ^data_full_wayBits_2_21; // @[ECC.scala 87:27]
    r2_data_errors_2_REG_2_22 <= ^data_full_wayBits_2_22; // @[ECC.scala 87:27]
    r2_data_errors_2_REG_2_23 <= ^data_full_wayBits_2_23; // @[ECC.scala 87:27]
    r2_data_errors_2_REG_2_24 <= ^data_full_wayBits_2_24; // @[ECC.scala 87:27]
    r2_data_errors_2_REG_2_25 <= ^data_full_wayBits_2_25; // @[ECC.scala 87:27]
    r2_data_errors_2_REG_2_26 <= ^data_full_wayBits_2_26; // @[ECC.scala 87:27]
    r2_data_errors_2_REG_2_27 <= ^data_full_wayBits_2_27; // @[ECC.scala 87:27]
    r2_data_errors_2_REG_2_28 <= ^data_full_wayBits_2_28; // @[ECC.scala 87:27]
    r2_data_errors_2_REG_2_29 <= ^data_full_wayBits_2_29; // @[ECC.scala 87:27]
    r2_data_errors_2_REG_2_30 <= ^data_full_wayBits_2_30; // @[ECC.scala 87:27]
    r2_data_errors_2_REG_2_31 <= ^data_full_wayBits_2_31; // @[ECC.scala 87:27]
    r2_data_errors_3_REG <= r1_valid & r2_ready; // @[ReplacePipe.scala 119:24]
    r2_data_errors_3_REG_1 <= r2_data_errors_3_REG; // @[ReplacePipe.scala 186:57]
    r2_data_errors_3_REG_2_0 <= ^data_full_wayBits_3_0; // @[ECC.scala 87:27]
    r2_data_errors_3_REG_2_1 <= ^data_full_wayBits_3_1; // @[ECC.scala 87:27]
    r2_data_errors_3_REG_2_2 <= ^data_full_wayBits_3_2; // @[ECC.scala 87:27]
    r2_data_errors_3_REG_2_3 <= ^data_full_wayBits_3_3; // @[ECC.scala 87:27]
    r2_data_errors_3_REG_2_4 <= ^data_full_wayBits_3_4; // @[ECC.scala 87:27]
    r2_data_errors_3_REG_2_5 <= ^data_full_wayBits_3_5; // @[ECC.scala 87:27]
    r2_data_errors_3_REG_2_6 <= ^data_full_wayBits_3_6; // @[ECC.scala 87:27]
    r2_data_errors_3_REG_2_7 <= ^data_full_wayBits_3_7; // @[ECC.scala 87:27]
    r2_data_errors_3_REG_2_8 <= ^data_full_wayBits_3_8; // @[ECC.scala 87:27]
    r2_data_errors_3_REG_2_9 <= ^data_full_wayBits_3_9; // @[ECC.scala 87:27]
    r2_data_errors_3_REG_2_10 <= ^data_full_wayBits_3_10; // @[ECC.scala 87:27]
    r2_data_errors_3_REG_2_11 <= ^data_full_wayBits_3_11; // @[ECC.scala 87:27]
    r2_data_errors_3_REG_2_12 <= ^data_full_wayBits_3_12; // @[ECC.scala 87:27]
    r2_data_errors_3_REG_2_13 <= ^data_full_wayBits_3_13; // @[ECC.scala 87:27]
    r2_data_errors_3_REG_2_14 <= ^data_full_wayBits_3_14; // @[ECC.scala 87:27]
    r2_data_errors_3_REG_2_15 <= ^data_full_wayBits_3_15; // @[ECC.scala 87:27]
    r2_data_errors_3_REG_2_16 <= ^data_full_wayBits_3_16; // @[ECC.scala 87:27]
    r2_data_errors_3_REG_2_17 <= ^data_full_wayBits_3_17; // @[ECC.scala 87:27]
    r2_data_errors_3_REG_2_18 <= ^data_full_wayBits_3_18; // @[ECC.scala 87:27]
    r2_data_errors_3_REG_2_19 <= ^data_full_wayBits_3_19; // @[ECC.scala 87:27]
    r2_data_errors_3_REG_2_20 <= ^data_full_wayBits_3_20; // @[ECC.scala 87:27]
    r2_data_errors_3_REG_2_21 <= ^data_full_wayBits_3_21; // @[ECC.scala 87:27]
    r2_data_errors_3_REG_2_22 <= ^data_full_wayBits_3_22; // @[ECC.scala 87:27]
    r2_data_errors_3_REG_2_23 <= ^data_full_wayBits_3_23; // @[ECC.scala 87:27]
    r2_data_errors_3_REG_2_24 <= ^data_full_wayBits_3_24; // @[ECC.scala 87:27]
    r2_data_errors_3_REG_2_25 <= ^data_full_wayBits_3_25; // @[ECC.scala 87:27]
    r2_data_errors_3_REG_2_26 <= ^data_full_wayBits_3_26; // @[ECC.scala 87:27]
    r2_data_errors_3_REG_2_27 <= ^data_full_wayBits_3_27; // @[ECC.scala 87:27]
    r2_data_errors_3_REG_2_28 <= ^data_full_wayBits_3_28; // @[ECC.scala 87:27]
    r2_data_errors_3_REG_2_29 <= ^data_full_wayBits_3_29; // @[ECC.scala 87:27]
    r2_data_errors_3_REG_2_30 <= ^data_full_wayBits_3_30; // @[ECC.scala 87:27]
    r2_data_errors_3_REG_2_31 <= ^data_full_wayBits_3_31; // @[ECC.scala 87:27]
    r2_data_errors_4_REG <= r1_valid & r2_ready; // @[ReplacePipe.scala 119:24]
    r2_data_errors_4_REG_1 <= r2_data_errors_4_REG; // @[ReplacePipe.scala 186:57]
    r2_data_errors_4_REG_2_0 <= ^data_full_wayBits_4_0; // @[ECC.scala 87:27]
    r2_data_errors_4_REG_2_1 <= ^data_full_wayBits_4_1; // @[ECC.scala 87:27]
    r2_data_errors_4_REG_2_2 <= ^data_full_wayBits_4_2; // @[ECC.scala 87:27]
    r2_data_errors_4_REG_2_3 <= ^data_full_wayBits_4_3; // @[ECC.scala 87:27]
    r2_data_errors_4_REG_2_4 <= ^data_full_wayBits_4_4; // @[ECC.scala 87:27]
    r2_data_errors_4_REG_2_5 <= ^data_full_wayBits_4_5; // @[ECC.scala 87:27]
    r2_data_errors_4_REG_2_6 <= ^data_full_wayBits_4_6; // @[ECC.scala 87:27]
    r2_data_errors_4_REG_2_7 <= ^data_full_wayBits_4_7; // @[ECC.scala 87:27]
    r2_data_errors_4_REG_2_8 <= ^data_full_wayBits_4_8; // @[ECC.scala 87:27]
    r2_data_errors_4_REG_2_9 <= ^data_full_wayBits_4_9; // @[ECC.scala 87:27]
    r2_data_errors_4_REG_2_10 <= ^data_full_wayBits_4_10; // @[ECC.scala 87:27]
    r2_data_errors_4_REG_2_11 <= ^data_full_wayBits_4_11; // @[ECC.scala 87:27]
    r2_data_errors_4_REG_2_12 <= ^data_full_wayBits_4_12; // @[ECC.scala 87:27]
    r2_data_errors_4_REG_2_13 <= ^data_full_wayBits_4_13; // @[ECC.scala 87:27]
    r2_data_errors_4_REG_2_14 <= ^data_full_wayBits_4_14; // @[ECC.scala 87:27]
    r2_data_errors_4_REG_2_15 <= ^data_full_wayBits_4_15; // @[ECC.scala 87:27]
    r2_data_errors_4_REG_2_16 <= ^data_full_wayBits_4_16; // @[ECC.scala 87:27]
    r2_data_errors_4_REG_2_17 <= ^data_full_wayBits_4_17; // @[ECC.scala 87:27]
    r2_data_errors_4_REG_2_18 <= ^data_full_wayBits_4_18; // @[ECC.scala 87:27]
    r2_data_errors_4_REG_2_19 <= ^data_full_wayBits_4_19; // @[ECC.scala 87:27]
    r2_data_errors_4_REG_2_20 <= ^data_full_wayBits_4_20; // @[ECC.scala 87:27]
    r2_data_errors_4_REG_2_21 <= ^data_full_wayBits_4_21; // @[ECC.scala 87:27]
    r2_data_errors_4_REG_2_22 <= ^data_full_wayBits_4_22; // @[ECC.scala 87:27]
    r2_data_errors_4_REG_2_23 <= ^data_full_wayBits_4_23; // @[ECC.scala 87:27]
    r2_data_errors_4_REG_2_24 <= ^data_full_wayBits_4_24; // @[ECC.scala 87:27]
    r2_data_errors_4_REG_2_25 <= ^data_full_wayBits_4_25; // @[ECC.scala 87:27]
    r2_data_errors_4_REG_2_26 <= ^data_full_wayBits_4_26; // @[ECC.scala 87:27]
    r2_data_errors_4_REG_2_27 <= ^data_full_wayBits_4_27; // @[ECC.scala 87:27]
    r2_data_errors_4_REG_2_28 <= ^data_full_wayBits_4_28; // @[ECC.scala 87:27]
    r2_data_errors_4_REG_2_29 <= ^data_full_wayBits_4_29; // @[ECC.scala 87:27]
    r2_data_errors_4_REG_2_30 <= ^data_full_wayBits_4_30; // @[ECC.scala 87:27]
    r2_data_errors_4_REG_2_31 <= ^data_full_wayBits_4_31; // @[ECC.scala 87:27]
    r2_data_errors_5_REG <= r1_valid & r2_ready; // @[ReplacePipe.scala 119:24]
    r2_data_errors_5_REG_1 <= r2_data_errors_5_REG; // @[ReplacePipe.scala 186:57]
    r2_data_errors_5_REG_2_0 <= ^data_full_wayBits_5_0; // @[ECC.scala 87:27]
    r2_data_errors_5_REG_2_1 <= ^data_full_wayBits_5_1; // @[ECC.scala 87:27]
    r2_data_errors_5_REG_2_2 <= ^data_full_wayBits_5_2; // @[ECC.scala 87:27]
    r2_data_errors_5_REG_2_3 <= ^data_full_wayBits_5_3; // @[ECC.scala 87:27]
    r2_data_errors_5_REG_2_4 <= ^data_full_wayBits_5_4; // @[ECC.scala 87:27]
    r2_data_errors_5_REG_2_5 <= ^data_full_wayBits_5_5; // @[ECC.scala 87:27]
    r2_data_errors_5_REG_2_6 <= ^data_full_wayBits_5_6; // @[ECC.scala 87:27]
    r2_data_errors_5_REG_2_7 <= ^data_full_wayBits_5_7; // @[ECC.scala 87:27]
    r2_data_errors_5_REG_2_8 <= ^data_full_wayBits_5_8; // @[ECC.scala 87:27]
    r2_data_errors_5_REG_2_9 <= ^data_full_wayBits_5_9; // @[ECC.scala 87:27]
    r2_data_errors_5_REG_2_10 <= ^data_full_wayBits_5_10; // @[ECC.scala 87:27]
    r2_data_errors_5_REG_2_11 <= ^data_full_wayBits_5_11; // @[ECC.scala 87:27]
    r2_data_errors_5_REG_2_12 <= ^data_full_wayBits_5_12; // @[ECC.scala 87:27]
    r2_data_errors_5_REG_2_13 <= ^data_full_wayBits_5_13; // @[ECC.scala 87:27]
    r2_data_errors_5_REG_2_14 <= ^data_full_wayBits_5_14; // @[ECC.scala 87:27]
    r2_data_errors_5_REG_2_15 <= ^data_full_wayBits_5_15; // @[ECC.scala 87:27]
    r2_data_errors_5_REG_2_16 <= ^data_full_wayBits_5_16; // @[ECC.scala 87:27]
    r2_data_errors_5_REG_2_17 <= ^data_full_wayBits_5_17; // @[ECC.scala 87:27]
    r2_data_errors_5_REG_2_18 <= ^data_full_wayBits_5_18; // @[ECC.scala 87:27]
    r2_data_errors_5_REG_2_19 <= ^data_full_wayBits_5_19; // @[ECC.scala 87:27]
    r2_data_errors_5_REG_2_20 <= ^data_full_wayBits_5_20; // @[ECC.scala 87:27]
    r2_data_errors_5_REG_2_21 <= ^data_full_wayBits_5_21; // @[ECC.scala 87:27]
    r2_data_errors_5_REG_2_22 <= ^data_full_wayBits_5_22; // @[ECC.scala 87:27]
    r2_data_errors_5_REG_2_23 <= ^data_full_wayBits_5_23; // @[ECC.scala 87:27]
    r2_data_errors_5_REG_2_24 <= ^data_full_wayBits_5_24; // @[ECC.scala 87:27]
    r2_data_errors_5_REG_2_25 <= ^data_full_wayBits_5_25; // @[ECC.scala 87:27]
    r2_data_errors_5_REG_2_26 <= ^data_full_wayBits_5_26; // @[ECC.scala 87:27]
    r2_data_errors_5_REG_2_27 <= ^data_full_wayBits_5_27; // @[ECC.scala 87:27]
    r2_data_errors_5_REG_2_28 <= ^data_full_wayBits_5_28; // @[ECC.scala 87:27]
    r2_data_errors_5_REG_2_29 <= ^data_full_wayBits_5_29; // @[ECC.scala 87:27]
    r2_data_errors_5_REG_2_30 <= ^data_full_wayBits_5_30; // @[ECC.scala 87:27]
    r2_data_errors_5_REG_2_31 <= ^data_full_wayBits_5_31; // @[ECC.scala 87:27]
    r2_data_errors_6_REG <= r1_valid & r2_ready; // @[ReplacePipe.scala 119:24]
    r2_data_errors_6_REG_1 <= r2_data_errors_6_REG; // @[ReplacePipe.scala 186:57]
    r2_data_errors_6_REG_2_0 <= ^data_full_wayBits_6_0; // @[ECC.scala 87:27]
    r2_data_errors_6_REG_2_1 <= ^data_full_wayBits_6_1; // @[ECC.scala 87:27]
    r2_data_errors_6_REG_2_2 <= ^data_full_wayBits_6_2; // @[ECC.scala 87:27]
    r2_data_errors_6_REG_2_3 <= ^data_full_wayBits_6_3; // @[ECC.scala 87:27]
    r2_data_errors_6_REG_2_4 <= ^data_full_wayBits_6_4; // @[ECC.scala 87:27]
    r2_data_errors_6_REG_2_5 <= ^data_full_wayBits_6_5; // @[ECC.scala 87:27]
    r2_data_errors_6_REG_2_6 <= ^data_full_wayBits_6_6; // @[ECC.scala 87:27]
    r2_data_errors_6_REG_2_7 <= ^data_full_wayBits_6_7; // @[ECC.scala 87:27]
    r2_data_errors_6_REG_2_8 <= ^data_full_wayBits_6_8; // @[ECC.scala 87:27]
    r2_data_errors_6_REG_2_9 <= ^data_full_wayBits_6_9; // @[ECC.scala 87:27]
    r2_data_errors_6_REG_2_10 <= ^data_full_wayBits_6_10; // @[ECC.scala 87:27]
    r2_data_errors_6_REG_2_11 <= ^data_full_wayBits_6_11; // @[ECC.scala 87:27]
    r2_data_errors_6_REG_2_12 <= ^data_full_wayBits_6_12; // @[ECC.scala 87:27]
    r2_data_errors_6_REG_2_13 <= ^data_full_wayBits_6_13; // @[ECC.scala 87:27]
    r2_data_errors_6_REG_2_14 <= ^data_full_wayBits_6_14; // @[ECC.scala 87:27]
    r2_data_errors_6_REG_2_15 <= ^data_full_wayBits_6_15; // @[ECC.scala 87:27]
    r2_data_errors_6_REG_2_16 <= ^data_full_wayBits_6_16; // @[ECC.scala 87:27]
    r2_data_errors_6_REG_2_17 <= ^data_full_wayBits_6_17; // @[ECC.scala 87:27]
    r2_data_errors_6_REG_2_18 <= ^data_full_wayBits_6_18; // @[ECC.scala 87:27]
    r2_data_errors_6_REG_2_19 <= ^data_full_wayBits_6_19; // @[ECC.scala 87:27]
    r2_data_errors_6_REG_2_20 <= ^data_full_wayBits_6_20; // @[ECC.scala 87:27]
    r2_data_errors_6_REG_2_21 <= ^data_full_wayBits_6_21; // @[ECC.scala 87:27]
    r2_data_errors_6_REG_2_22 <= ^data_full_wayBits_6_22; // @[ECC.scala 87:27]
    r2_data_errors_6_REG_2_23 <= ^data_full_wayBits_6_23; // @[ECC.scala 87:27]
    r2_data_errors_6_REG_2_24 <= ^data_full_wayBits_6_24; // @[ECC.scala 87:27]
    r2_data_errors_6_REG_2_25 <= ^data_full_wayBits_6_25; // @[ECC.scala 87:27]
    r2_data_errors_6_REG_2_26 <= ^data_full_wayBits_6_26; // @[ECC.scala 87:27]
    r2_data_errors_6_REG_2_27 <= ^data_full_wayBits_6_27; // @[ECC.scala 87:27]
    r2_data_errors_6_REG_2_28 <= ^data_full_wayBits_6_28; // @[ECC.scala 87:27]
    r2_data_errors_6_REG_2_29 <= ^data_full_wayBits_6_29; // @[ECC.scala 87:27]
    r2_data_errors_6_REG_2_30 <= ^data_full_wayBits_6_30; // @[ECC.scala 87:27]
    r2_data_errors_6_REG_2_31 <= ^data_full_wayBits_6_31; // @[ECC.scala 87:27]
    r2_data_errors_7_REG <= r1_valid & r2_ready; // @[ReplacePipe.scala 119:24]
    r2_data_errors_7_REG_1 <= r2_data_errors_7_REG; // @[ReplacePipe.scala 186:57]
    r2_data_errors_7_REG_2_0 <= ^data_full_wayBits_7_0; // @[ECC.scala 87:27]
    r2_data_errors_7_REG_2_1 <= ^data_full_wayBits_7_1; // @[ECC.scala 87:27]
    r2_data_errors_7_REG_2_2 <= ^data_full_wayBits_7_2; // @[ECC.scala 87:27]
    r2_data_errors_7_REG_2_3 <= ^data_full_wayBits_7_3; // @[ECC.scala 87:27]
    r2_data_errors_7_REG_2_4 <= ^data_full_wayBits_7_4; // @[ECC.scala 87:27]
    r2_data_errors_7_REG_2_5 <= ^data_full_wayBits_7_5; // @[ECC.scala 87:27]
    r2_data_errors_7_REG_2_6 <= ^data_full_wayBits_7_6; // @[ECC.scala 87:27]
    r2_data_errors_7_REG_2_7 <= ^data_full_wayBits_7_7; // @[ECC.scala 87:27]
    r2_data_errors_7_REG_2_8 <= ^data_full_wayBits_7_8; // @[ECC.scala 87:27]
    r2_data_errors_7_REG_2_9 <= ^data_full_wayBits_7_9; // @[ECC.scala 87:27]
    r2_data_errors_7_REG_2_10 <= ^data_full_wayBits_7_10; // @[ECC.scala 87:27]
    r2_data_errors_7_REG_2_11 <= ^data_full_wayBits_7_11; // @[ECC.scala 87:27]
    r2_data_errors_7_REG_2_12 <= ^data_full_wayBits_7_12; // @[ECC.scala 87:27]
    r2_data_errors_7_REG_2_13 <= ^data_full_wayBits_7_13; // @[ECC.scala 87:27]
    r2_data_errors_7_REG_2_14 <= ^data_full_wayBits_7_14; // @[ECC.scala 87:27]
    r2_data_errors_7_REG_2_15 <= ^data_full_wayBits_7_15; // @[ECC.scala 87:27]
    r2_data_errors_7_REG_2_16 <= ^data_full_wayBits_7_16; // @[ECC.scala 87:27]
    r2_data_errors_7_REG_2_17 <= ^data_full_wayBits_7_17; // @[ECC.scala 87:27]
    r2_data_errors_7_REG_2_18 <= ^data_full_wayBits_7_18; // @[ECC.scala 87:27]
    r2_data_errors_7_REG_2_19 <= ^data_full_wayBits_7_19; // @[ECC.scala 87:27]
    r2_data_errors_7_REG_2_20 <= ^data_full_wayBits_7_20; // @[ECC.scala 87:27]
    r2_data_errors_7_REG_2_21 <= ^data_full_wayBits_7_21; // @[ECC.scala 87:27]
    r2_data_errors_7_REG_2_22 <= ^data_full_wayBits_7_22; // @[ECC.scala 87:27]
    r2_data_errors_7_REG_2_23 <= ^data_full_wayBits_7_23; // @[ECC.scala 87:27]
    r2_data_errors_7_REG_2_24 <= ^data_full_wayBits_7_24; // @[ECC.scala 87:27]
    r2_data_errors_7_REG_2_25 <= ^data_full_wayBits_7_25; // @[ECC.scala 87:27]
    r2_data_errors_7_REG_2_26 <= ^data_full_wayBits_7_26; // @[ECC.scala 87:27]
    r2_data_errors_7_REG_2_27 <= ^data_full_wayBits_7_27; // @[ECC.scala 87:27]
    r2_data_errors_7_REG_2_28 <= ^data_full_wayBits_7_28; // @[ECC.scala 87:27]
    r2_data_errors_7_REG_2_29 <= ^data_full_wayBits_7_29; // @[ECC.scala 87:27]
    r2_data_errors_7_REG_2_30 <= ^data_full_wayBits_7_30; // @[ECC.scala 87:27]
    r2_data_errors_7_REG_2_31 <= ^data_full_wayBits_7_31; // @[ECC.scala 87:27]
    r2_parity_error_REG <= (r2_meta_errors_0 | r2_meta_errors_1 | r2_meta_errors_2 | r2_meta_errors_3 | r2_meta_errors_4
       | r2_meta_errors_5 | r2_meta_errors_6 | r2_meta_errors_7) & io_csr_parity_enable; // @[ReplacePipe.scala 188:58]
    io_error_valid_REG <= r1_valid & r2_ready; // @[ReplacePipe.scala 119:24]
    io_error_valid_REG_1 <= io_error_valid_REG; // @[ReplacePipe.scala 193:71]
    io_error_valid_REG_2 <= r2_parity_error & io_error_valid_REG_1; // @[ReplacePipe.scala 193:60]
    io_error_report_to_beu_REG <= r1_valid & r2_ready; // @[ReplacePipe.scala 119:24]
    io_error_report_to_beu_REG_1 <= io_error_report_to_beu_REG; // @[ReplacePipe.scala 194:71]
    io_error_report_to_beu_REG_2 <= r2_parity_error & io_error_report_to_beu_REG_1; // @[ReplacePipe.scala 194:60]
    io_error_paddr_REG <= r2_req_paddr; // @[ReplacePipe.scala 195:51]
    io_error_paddr_REG_1 <= io_error_paddr_REG; // @[ReplacePipe.scala 195:43]
    io_error_source_tag_REG <= (r2_meta_errors_0 | r2_meta_errors_1 | r2_meta_errors_2 | r2_meta_errors_3 |
      r2_meta_errors_4 | r2_meta_errors_5 | r2_meta_errors_6 | r2_meta_errors_7) & io_csr_parity_enable; // @[ReplacePipe.scala 188:58]
    io_error_source_tag_REG_1 <= io_error_source_tag_REG; // @[ReplacePipe.scala 196:43]
    io_error_source_data_REG <= (r2_data_errors_0 | r2_data_errors_1 | r2_data_errors_2 | r2_data_errors_3 |
      r2_data_errors_4 | r2_data_errors_5 | r2_data_errors_6 | r2_data_errors_7) & io_csr_parity_enable; // @[ReplacePipe.scala 189:58]
    io_error_opType_release_REG <= r2_req_voluntary; // @[ReplacePipe.scala 201:51]
    io_error_opType_release_REG_1 <= io_error_opType_release_REG; // @[ReplacePipe.scala 201:43]
    io_error_opType_probe_REG <= ~r2_req_voluntary; // @[ReplacePipe.scala 39:17]
    io_error_opType_probe_REG_1 <= io_error_opType_probe_REG; // @[ReplacePipe.scala 202:43]
    if (r1_fire) begin // @[Reg.scala 17:18]
      r2_release_coh_state <= release_coh_state; // @[Reg.scala 17:22]
    end
    if (r1_fire) begin // @[Reg.scala 17:18]
      r2_release_addr <= release_addr; // @[Reg.scala 17:22]
    end
    r3_fire_REG <= io_release_finish; // @[ReplacePipe.scala 258:40]
    if (_r3_valid_T) begin // @[Reg.scala 17:18]
      r3_release_need_send <= release_need_send; // @[Reg.scala 17:22]
    end
    if (_r3_valid_T) begin // @[Reg.scala 17:18]
      r3_req_vaddr <= r2_req_vaddr; // @[Reg.scala 17:22]
    end
    if (_r3_valid_T) begin // @[Reg.scala 17:18]
      r3_req_id <= r2_req_id; // @[Reg.scala 17:22]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ICache.scala 100:42]
      r0_valid <= 1'h0; // @[ICache.scala 100:50]
    end else begin
      r0_valid <= _r0_valid_T | _GEN_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ICache.scala 100:42]
      r2_valid <= 1'h0; // @[ICache.scala 100:50]
    end else begin
      r2_valid <= r1_fire | _GEN_60;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ICache.scala 100:42]
      r1_valid <= 1'h0; // @[ICache.scala 100:50]
    end else begin
      r1_valid <= r0_fire | _GEN_10;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ICache.scala 100:42]
      r3_valid <= 1'h0; // @[ICache.scala 100:50]
    end else begin
      r3_valid <= _r3_valid_T | _GEN_107;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r0_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  r2_valid = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  r1_valid = _RAND_2[0:0];
  _RAND_3 = {2{`RANDOM}};
  r0_req_paddr = _RAND_3[35:0];
  _RAND_4 = {2{`RANDOM}};
  r0_req_vaddr = _RAND_4[38:0];
  _RAND_5 = {1{`RANDOM}};
  r0_req_param = _RAND_5[2:0];
  _RAND_6 = {1{`RANDOM}};
  r0_req_voluntary = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  r0_req_needData = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  r0_req_waymask = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  r0_req_id = _RAND_9[4:0];
  _RAND_10 = {2{`RANDOM}};
  r1_req_paddr = _RAND_10[35:0];
  _RAND_11 = {2{`RANDOM}};
  r1_req_vaddr = _RAND_11[38:0];
  _RAND_12 = {1{`RANDOM}};
  r1_req_param = _RAND_12[2:0];
  _RAND_13 = {1{`RANDOM}};
  r1_req_voluntary = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  r1_req_needData = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  r1_req_waymask = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  r1_req_id = _RAND_16[4:0];
  _RAND_17 = {1{`RANDOM}};
  r1_meta_ptags_REG = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  r1_meta_ptags_r0 = _RAND_18[23:0];
  _RAND_19 = {1{`RANDOM}};
  r1_meta_ptags_r1 = _RAND_19[23:0];
  _RAND_20 = {1{`RANDOM}};
  r1_meta_ptags_r2 = _RAND_20[23:0];
  _RAND_21 = {1{`RANDOM}};
  r1_meta_ptags_r3 = _RAND_21[23:0];
  _RAND_22 = {1{`RANDOM}};
  r1_meta_ptags_r4 = _RAND_22[23:0];
  _RAND_23 = {1{`RANDOM}};
  r1_meta_ptags_r5 = _RAND_23[23:0];
  _RAND_24 = {1{`RANDOM}};
  r1_meta_ptags_r6 = _RAND_24[23:0];
  _RAND_25 = {1{`RANDOM}};
  r1_meta_ptags_r7 = _RAND_25[23:0];
  _RAND_26 = {1{`RANDOM}};
  r1_meta_cohs_REG = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  r1_meta_cohs_r0_state = _RAND_27[1:0];
  _RAND_28 = {1{`RANDOM}};
  r1_meta_cohs_r1_state = _RAND_28[1:0];
  _RAND_29 = {1{`RANDOM}};
  r1_meta_cohs_r2_state = _RAND_29[1:0];
  _RAND_30 = {1{`RANDOM}};
  r1_meta_cohs_r3_state = _RAND_30[1:0];
  _RAND_31 = {1{`RANDOM}};
  r1_meta_cohs_r4_state = _RAND_31[1:0];
  _RAND_32 = {1{`RANDOM}};
  r1_meta_cohs_r5_state = _RAND_32[1:0];
  _RAND_33 = {1{`RANDOM}};
  r1_meta_cohs_r6_state = _RAND_33[1:0];
  _RAND_34 = {1{`RANDOM}};
  r1_meta_cohs_r7_state = _RAND_34[1:0];
  _RAND_35 = {1{`RANDOM}};
  r1_meta_errors_REG = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  r1_meta_errors_r0 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  r1_meta_errors_r1 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  r1_meta_errors_r2 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  r1_meta_errors_r3 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  r1_meta_errors_r4 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  r1_meta_errors_r5 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  r1_meta_errors_r6 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  r1_meta_errors_r7 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  r1_data_cacheline_REG = _RAND_44[0:0];
  _RAND_45 = {16{`RANDOM}};
  r1_data_cacheline_r0 = _RAND_45[511:0];
  _RAND_46 = {16{`RANDOM}};
  r1_data_cacheline_r1 = _RAND_46[511:0];
  _RAND_47 = {16{`RANDOM}};
  r1_data_cacheline_r2 = _RAND_47[511:0];
  _RAND_48 = {16{`RANDOM}};
  r1_data_cacheline_r3 = _RAND_48[511:0];
  _RAND_49 = {16{`RANDOM}};
  r1_data_cacheline_r4 = _RAND_49[511:0];
  _RAND_50 = {16{`RANDOM}};
  r1_data_cacheline_r5 = _RAND_50[511:0];
  _RAND_51 = {16{`RANDOM}};
  r1_data_cacheline_r6 = _RAND_51[511:0];
  _RAND_52 = {16{`RANDOM}};
  r1_data_cacheline_r7 = _RAND_52[511:0];
  _RAND_53 = {1{`RANDOM}};
  r1_data_errorBits_REG = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  r1_data_errorBits_r0 = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  r1_data_errorBits_r1 = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  r1_data_errorBits_r2 = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  r1_data_errorBits_r3 = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  r1_data_errorBits_r4 = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  r1_data_errorBits_r5 = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  r1_data_errorBits_r6 = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  r1_data_errorBits_r7 = _RAND_61[31:0];
  _RAND_62 = {2{`RANDOM}};
  r2_req_paddr = _RAND_62[35:0];
  _RAND_63 = {2{`RANDOM}};
  r2_req_vaddr = _RAND_63[38:0];
  _RAND_64 = {1{`RANDOM}};
  r2_req_param = _RAND_64[2:0];
  _RAND_65 = {1{`RANDOM}};
  r2_req_voluntary = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  r2_req_needData = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  r2_req_waymask = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  r2_req_id = _RAND_68[4:0];
  _RAND_69 = {16{`RANDOM}};
  r2_data_cacheline_0 = _RAND_69[511:0];
  _RAND_70 = {16{`RANDOM}};
  r2_data_cacheline_1 = _RAND_70[511:0];
  _RAND_71 = {16{`RANDOM}};
  r2_data_cacheline_2 = _RAND_71[511:0];
  _RAND_72 = {16{`RANDOM}};
  r2_data_cacheline_3 = _RAND_72[511:0];
  _RAND_73 = {16{`RANDOM}};
  r2_data_cacheline_4 = _RAND_73[511:0];
  _RAND_74 = {16{`RANDOM}};
  r2_data_cacheline_5 = _RAND_74[511:0];
  _RAND_75 = {16{`RANDOM}};
  r2_data_cacheline_6 = _RAND_75[511:0];
  _RAND_76 = {16{`RANDOM}};
  r2_data_cacheline_7 = _RAND_76[511:0];
  _RAND_77 = {1{`RANDOM}};
  r2_probe_hit_ptag = _RAND_77[23:0];
  _RAND_78 = {1{`RANDOM}};
  r2_probe_hit_vec_0 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  r2_probe_hit_vec_1 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  r2_probe_hit_vec_2 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  r2_probe_hit_vec_3 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  r2_probe_hit_vec_4 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  r2_probe_hit_vec_5 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  r2_probe_hit_vec_6 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  r2_probe_hit_vec_7 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  r2_probe_hit_coh_state = _RAND_86[1:0];
  _RAND_87 = {1{`RANDOM}};
  r2_meta_errors_0 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  r2_meta_errors_1 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  r2_meta_errors_2 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  r2_meta_errors_3 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  r2_meta_errors_4 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  r2_meta_errors_5 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  r2_meta_errors_6 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  r2_meta_errors_7 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  r2_data_errorBits_0 = _RAND_95[31:0];
  _RAND_96 = {1{`RANDOM}};
  r2_data_errorBits_1 = _RAND_96[31:0];
  _RAND_97 = {1{`RANDOM}};
  r2_data_errorBits_2 = _RAND_97[31:0];
  _RAND_98 = {1{`RANDOM}};
  r2_data_errorBits_3 = _RAND_98[31:0];
  _RAND_99 = {1{`RANDOM}};
  r2_data_errorBits_4 = _RAND_99[31:0];
  _RAND_100 = {1{`RANDOM}};
  r2_data_errorBits_5 = _RAND_100[31:0];
  _RAND_101 = {1{`RANDOM}};
  r2_data_errorBits_6 = _RAND_101[31:0];
  _RAND_102 = {1{`RANDOM}};
  r2_data_errorBits_7 = _RAND_102[31:0];
  _RAND_103 = {1{`RANDOM}};
  r2_data_errors_0_REG = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  r2_data_errors_0_REG_1 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  r2_data_errors_0_REG_2_0 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  r2_data_errors_0_REG_2_1 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  r2_data_errors_0_REG_2_2 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  r2_data_errors_0_REG_2_3 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  r2_data_errors_0_REG_2_4 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  r2_data_errors_0_REG_2_5 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  r2_data_errors_0_REG_2_6 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  r2_data_errors_0_REG_2_7 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  r2_data_errors_0_REG_2_8 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  r2_data_errors_0_REG_2_9 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  r2_data_errors_0_REG_2_10 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  r2_data_errors_0_REG_2_11 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  r2_data_errors_0_REG_2_12 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  r2_data_errors_0_REG_2_13 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  r2_data_errors_0_REG_2_14 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  r2_data_errors_0_REG_2_15 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  r2_data_errors_0_REG_2_16 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  r2_data_errors_0_REG_2_17 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  r2_data_errors_0_REG_2_18 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  r2_data_errors_0_REG_2_19 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  r2_data_errors_0_REG_2_20 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  r2_data_errors_0_REG_2_21 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  r2_data_errors_0_REG_2_22 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  r2_data_errors_0_REG_2_23 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  r2_data_errors_0_REG_2_24 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  r2_data_errors_0_REG_2_25 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  r2_data_errors_0_REG_2_26 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  r2_data_errors_0_REG_2_27 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  r2_data_errors_0_REG_2_28 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  r2_data_errors_0_REG_2_29 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  r2_data_errors_0_REG_2_30 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  r2_data_errors_0_REG_2_31 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  r2_data_errors_1_REG = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  r2_data_errors_1_REG_1 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  r2_data_errors_1_REG_2_0 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  r2_data_errors_1_REG_2_1 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  r2_data_errors_1_REG_2_2 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  r2_data_errors_1_REG_2_3 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  r2_data_errors_1_REG_2_4 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  r2_data_errors_1_REG_2_5 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  r2_data_errors_1_REG_2_6 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  r2_data_errors_1_REG_2_7 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  r2_data_errors_1_REG_2_8 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  r2_data_errors_1_REG_2_9 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  r2_data_errors_1_REG_2_10 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  r2_data_errors_1_REG_2_11 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  r2_data_errors_1_REG_2_12 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  r2_data_errors_1_REG_2_13 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  r2_data_errors_1_REG_2_14 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  r2_data_errors_1_REG_2_15 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  r2_data_errors_1_REG_2_16 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  r2_data_errors_1_REG_2_17 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  r2_data_errors_1_REG_2_18 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  r2_data_errors_1_REG_2_19 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  r2_data_errors_1_REG_2_20 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  r2_data_errors_1_REG_2_21 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  r2_data_errors_1_REG_2_22 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  r2_data_errors_1_REG_2_23 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  r2_data_errors_1_REG_2_24 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  r2_data_errors_1_REG_2_25 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  r2_data_errors_1_REG_2_26 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  r2_data_errors_1_REG_2_27 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  r2_data_errors_1_REG_2_28 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  r2_data_errors_1_REG_2_29 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  r2_data_errors_1_REG_2_30 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  r2_data_errors_1_REG_2_31 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  r2_data_errors_2_REG = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  r2_data_errors_2_REG_1 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  r2_data_errors_2_REG_2_0 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  r2_data_errors_2_REG_2_1 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  r2_data_errors_2_REG_2_2 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  r2_data_errors_2_REG_2_3 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  r2_data_errors_2_REG_2_4 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  r2_data_errors_2_REG_2_5 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  r2_data_errors_2_REG_2_6 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  r2_data_errors_2_REG_2_7 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  r2_data_errors_2_REG_2_8 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  r2_data_errors_2_REG_2_9 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  r2_data_errors_2_REG_2_10 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  r2_data_errors_2_REG_2_11 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  r2_data_errors_2_REG_2_12 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  r2_data_errors_2_REG_2_13 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  r2_data_errors_2_REG_2_14 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  r2_data_errors_2_REG_2_15 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  r2_data_errors_2_REG_2_16 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  r2_data_errors_2_REG_2_17 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  r2_data_errors_2_REG_2_18 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  r2_data_errors_2_REG_2_19 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  r2_data_errors_2_REG_2_20 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  r2_data_errors_2_REG_2_21 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  r2_data_errors_2_REG_2_22 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  r2_data_errors_2_REG_2_23 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  r2_data_errors_2_REG_2_24 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  r2_data_errors_2_REG_2_25 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  r2_data_errors_2_REG_2_26 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  r2_data_errors_2_REG_2_27 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  r2_data_errors_2_REG_2_28 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  r2_data_errors_2_REG_2_29 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  r2_data_errors_2_REG_2_30 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  r2_data_errors_2_REG_2_31 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  r2_data_errors_3_REG = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  r2_data_errors_3_REG_1 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  r2_data_errors_3_REG_2_0 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  r2_data_errors_3_REG_2_1 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  r2_data_errors_3_REG_2_2 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  r2_data_errors_3_REG_2_3 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  r2_data_errors_3_REG_2_4 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  r2_data_errors_3_REG_2_5 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  r2_data_errors_3_REG_2_6 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  r2_data_errors_3_REG_2_7 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  r2_data_errors_3_REG_2_8 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  r2_data_errors_3_REG_2_9 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  r2_data_errors_3_REG_2_10 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  r2_data_errors_3_REG_2_11 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  r2_data_errors_3_REG_2_12 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  r2_data_errors_3_REG_2_13 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  r2_data_errors_3_REG_2_14 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  r2_data_errors_3_REG_2_15 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  r2_data_errors_3_REG_2_16 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  r2_data_errors_3_REG_2_17 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  r2_data_errors_3_REG_2_18 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  r2_data_errors_3_REG_2_19 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  r2_data_errors_3_REG_2_20 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  r2_data_errors_3_REG_2_21 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  r2_data_errors_3_REG_2_22 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  r2_data_errors_3_REG_2_23 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  r2_data_errors_3_REG_2_24 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  r2_data_errors_3_REG_2_25 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  r2_data_errors_3_REG_2_26 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  r2_data_errors_3_REG_2_27 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  r2_data_errors_3_REG_2_28 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  r2_data_errors_3_REG_2_29 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  r2_data_errors_3_REG_2_30 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  r2_data_errors_3_REG_2_31 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  r2_data_errors_4_REG = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  r2_data_errors_4_REG_1 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  r2_data_errors_4_REG_2_0 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  r2_data_errors_4_REG_2_1 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  r2_data_errors_4_REG_2_2 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  r2_data_errors_4_REG_2_3 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  r2_data_errors_4_REG_2_4 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  r2_data_errors_4_REG_2_5 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  r2_data_errors_4_REG_2_6 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  r2_data_errors_4_REG_2_7 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  r2_data_errors_4_REG_2_8 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  r2_data_errors_4_REG_2_9 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  r2_data_errors_4_REG_2_10 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  r2_data_errors_4_REG_2_11 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  r2_data_errors_4_REG_2_12 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  r2_data_errors_4_REG_2_13 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  r2_data_errors_4_REG_2_14 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  r2_data_errors_4_REG_2_15 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  r2_data_errors_4_REG_2_16 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  r2_data_errors_4_REG_2_17 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  r2_data_errors_4_REG_2_18 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  r2_data_errors_4_REG_2_19 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  r2_data_errors_4_REG_2_20 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  r2_data_errors_4_REG_2_21 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  r2_data_errors_4_REG_2_22 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  r2_data_errors_4_REG_2_23 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  r2_data_errors_4_REG_2_24 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  r2_data_errors_4_REG_2_25 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  r2_data_errors_4_REG_2_26 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  r2_data_errors_4_REG_2_27 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  r2_data_errors_4_REG_2_28 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  r2_data_errors_4_REG_2_29 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  r2_data_errors_4_REG_2_30 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  r2_data_errors_4_REG_2_31 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  r2_data_errors_5_REG = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  r2_data_errors_5_REG_1 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  r2_data_errors_5_REG_2_0 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  r2_data_errors_5_REG_2_1 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  r2_data_errors_5_REG_2_2 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  r2_data_errors_5_REG_2_3 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  r2_data_errors_5_REG_2_4 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  r2_data_errors_5_REG_2_5 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  r2_data_errors_5_REG_2_6 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  r2_data_errors_5_REG_2_7 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  r2_data_errors_5_REG_2_8 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  r2_data_errors_5_REG_2_9 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  r2_data_errors_5_REG_2_10 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  r2_data_errors_5_REG_2_11 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  r2_data_errors_5_REG_2_12 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  r2_data_errors_5_REG_2_13 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  r2_data_errors_5_REG_2_14 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  r2_data_errors_5_REG_2_15 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  r2_data_errors_5_REG_2_16 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  r2_data_errors_5_REG_2_17 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  r2_data_errors_5_REG_2_18 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  r2_data_errors_5_REG_2_19 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  r2_data_errors_5_REG_2_20 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  r2_data_errors_5_REG_2_21 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  r2_data_errors_5_REG_2_22 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  r2_data_errors_5_REG_2_23 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  r2_data_errors_5_REG_2_24 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  r2_data_errors_5_REG_2_25 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  r2_data_errors_5_REG_2_26 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  r2_data_errors_5_REG_2_27 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  r2_data_errors_5_REG_2_28 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  r2_data_errors_5_REG_2_29 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  r2_data_errors_5_REG_2_30 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  r2_data_errors_5_REG_2_31 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  r2_data_errors_6_REG = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  r2_data_errors_6_REG_1 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  r2_data_errors_6_REG_2_0 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  r2_data_errors_6_REG_2_1 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  r2_data_errors_6_REG_2_2 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  r2_data_errors_6_REG_2_3 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  r2_data_errors_6_REG_2_4 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  r2_data_errors_6_REG_2_5 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  r2_data_errors_6_REG_2_6 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  r2_data_errors_6_REG_2_7 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  r2_data_errors_6_REG_2_8 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  r2_data_errors_6_REG_2_9 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  r2_data_errors_6_REG_2_10 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  r2_data_errors_6_REG_2_11 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  r2_data_errors_6_REG_2_12 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  r2_data_errors_6_REG_2_13 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  r2_data_errors_6_REG_2_14 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  r2_data_errors_6_REG_2_15 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  r2_data_errors_6_REG_2_16 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  r2_data_errors_6_REG_2_17 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  r2_data_errors_6_REG_2_18 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  r2_data_errors_6_REG_2_19 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  r2_data_errors_6_REG_2_20 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  r2_data_errors_6_REG_2_21 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  r2_data_errors_6_REG_2_22 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  r2_data_errors_6_REG_2_23 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  r2_data_errors_6_REG_2_24 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  r2_data_errors_6_REG_2_25 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  r2_data_errors_6_REG_2_26 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  r2_data_errors_6_REG_2_27 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  r2_data_errors_6_REG_2_28 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  r2_data_errors_6_REG_2_29 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  r2_data_errors_6_REG_2_30 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  r2_data_errors_6_REG_2_31 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  r2_data_errors_7_REG = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  r2_data_errors_7_REG_1 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  r2_data_errors_7_REG_2_0 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  r2_data_errors_7_REG_2_1 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  r2_data_errors_7_REG_2_2 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  r2_data_errors_7_REG_2_3 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  r2_data_errors_7_REG_2_4 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  r2_data_errors_7_REG_2_5 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  r2_data_errors_7_REG_2_6 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  r2_data_errors_7_REG_2_7 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  r2_data_errors_7_REG_2_8 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  r2_data_errors_7_REG_2_9 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  r2_data_errors_7_REG_2_10 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  r2_data_errors_7_REG_2_11 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  r2_data_errors_7_REG_2_12 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  r2_data_errors_7_REG_2_13 = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  r2_data_errors_7_REG_2_14 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  r2_data_errors_7_REG_2_15 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  r2_data_errors_7_REG_2_16 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  r2_data_errors_7_REG_2_17 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  r2_data_errors_7_REG_2_18 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  r2_data_errors_7_REG_2_19 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  r2_data_errors_7_REG_2_20 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  r2_data_errors_7_REG_2_21 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  r2_data_errors_7_REG_2_22 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  r2_data_errors_7_REG_2_23 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  r2_data_errors_7_REG_2_24 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  r2_data_errors_7_REG_2_25 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  r2_data_errors_7_REG_2_26 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  r2_data_errors_7_REG_2_27 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  r2_data_errors_7_REG_2_28 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  r2_data_errors_7_REG_2_29 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  r2_data_errors_7_REG_2_30 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  r2_data_errors_7_REG_2_31 = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  r2_parity_error_REG = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  io_error_valid_REG = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  io_error_valid_REG_1 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  io_error_valid_REG_2 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  io_error_report_to_beu_REG = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  io_error_report_to_beu_REG_1 = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  io_error_report_to_beu_REG_2 = _RAND_381[0:0];
  _RAND_382 = {2{`RANDOM}};
  io_error_paddr_REG = _RAND_382[35:0];
  _RAND_383 = {2{`RANDOM}};
  io_error_paddr_REG_1 = _RAND_383[35:0];
  _RAND_384 = {1{`RANDOM}};
  io_error_source_tag_REG = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  io_error_source_tag_REG_1 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  io_error_source_data_REG = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  io_error_opType_release_REG = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  io_error_opType_release_REG_1 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  io_error_opType_probe_REG = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  io_error_opType_probe_REG_1 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  r2_release_coh_state = _RAND_391[1:0];
  _RAND_392 = {2{`RANDOM}};
  r2_release_addr = _RAND_392[35:0];
  _RAND_393 = {1{`RANDOM}};
  r3_valid = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  r3_fire_REG = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  r3_release_need_send = _RAND_395[0:0];
  _RAND_396 = {2{`RANDOM}};
  r3_req_vaddr = _RAND_396[38:0];
  _RAND_397 = {1{`RANDOM}};
  r3_req_id = _RAND_397[4:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    r0_valid = 1'h0;
  end
  if (reset) begin
    r2_valid = 1'h0;
  end
  if (reset) begin
    r1_valid = 1'h0;
  end
  if (reset) begin
    r3_valid = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule

