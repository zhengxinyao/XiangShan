module Rob(
  input        clock,
  input        reset,
  input  [7:0] io_hartId,
  input        io_redirect_valid,
  input        io_redirect_bits_robIdx_flag,
  input  [4:0] io_redirect_bits_robIdx_value,
  input        io_redirect_bits_level,
  output       io_enq_canAccept,
  output       io_enq_isEmpty,
  input        io_enq_needAlloc_0,
  input        io_enq_req_0_valid,
  input        io_enq_req_0_bits_cf_exceptionVec_1,
  input        io_enq_req_0_bits_cf_exceptionVec_2,
  input        io_enq_req_0_bits_cf_exceptionVec_12,
  input        io_enq_req_0_bits_cf_trigger_frontendHit_0,
  input        io_enq_req_0_bits_cf_trigger_frontendHit_1,
  input        io_enq_req_0_bits_cf_trigger_frontendHit_2,
  input        io_enq_req_0_bits_cf_trigger_frontendHit_3,
  input        io_enq_req_0_bits_cf_pd_isRVC,
  input        io_enq_req_0_bits_cf_crossPageIPFFix,
  input        io_enq_req_0_bits_cf_loadWaitBit,
  input        io_enq_req_0_bits_cf_ftqPtr_flag,
  input  [2:0] io_enq_req_0_bits_cf_ftqPtr_value,
  input  [2:0] io_enq_req_0_bits_cf_ftqOffset,
  input  [4:0] io_enq_req_0_bits_ctrl_ldest,
  input  [3:0] io_enq_req_0_bits_ctrl_fuType,
  input  [6:0] io_enq_req_0_bits_ctrl_fuOpType,
  input        io_enq_req_0_bits_ctrl_rfWen,
  input        io_enq_req_0_bits_ctrl_fpWen,
  input        io_enq_req_0_bits_ctrl_isXSTrap,
  input        io_enq_req_0_bits_ctrl_noSpecExec,
  input        io_enq_req_0_bits_ctrl_blockBackward,
  input        io_enq_req_0_bits_ctrl_flushPipe,
  input  [2:0] io_enq_req_0_bits_ctrl_commitType,
  input        io_enq_req_0_bits_ctrl_fpu_wflags,
  input        io_enq_req_0_bits_ctrl_isMove,
  input        io_enq_req_0_bits_ctrl_singleStep,
  input  [5:0] io_enq_req_0_bits_pdest,
  input  [5:0] io_enq_req_0_bits_old_pdest,
  input        io_enq_req_0_bits_robIdx_flag,
  input  [4:0] io_enq_req_0_bits_robIdx_value,
  input        io_enq_req_0_bits_eliminatedMove,
  input        io_enq_req_1_valid,
  input        io_enq_req_1_bits_cf_exceptionVec_1,
  input        io_enq_req_1_bits_cf_exceptionVec_2,
  input        io_enq_req_1_bits_cf_exceptionVec_12,
  input        io_enq_req_1_bits_cf_trigger_frontendHit_0,
  input        io_enq_req_1_bits_cf_trigger_frontendHit_1,
  input        io_enq_req_1_bits_cf_trigger_frontendHit_2,
  input        io_enq_req_1_bits_cf_trigger_frontendHit_3,
  input        io_enq_req_1_bits_cf_pd_isRVC,
  input        io_enq_req_1_bits_cf_crossPageIPFFix,
  input        io_enq_req_1_bits_cf_loadWaitBit,
  input        io_enq_req_1_bits_cf_ftqPtr_flag,
  input  [2:0] io_enq_req_1_bits_cf_ftqPtr_value,
  input  [2:0] io_enq_req_1_bits_cf_ftqOffset,
  input  [4:0] io_enq_req_1_bits_ctrl_ldest,
  input  [3:0] io_enq_req_1_bits_ctrl_fuType,
  input  [6:0] io_enq_req_1_bits_ctrl_fuOpType,
  input        io_enq_req_1_bits_ctrl_rfWen,
  input        io_enq_req_1_bits_ctrl_fpWen,
  input        io_enq_req_1_bits_ctrl_isXSTrap,
  input        io_enq_req_1_bits_ctrl_noSpecExec,
  input        io_enq_req_1_bits_ctrl_blockBackward,
  input        io_enq_req_1_bits_ctrl_flushPipe,
  input  [2:0] io_enq_req_1_bits_ctrl_commitType,
  input        io_enq_req_1_bits_ctrl_fpu_wflags,
  input        io_enq_req_1_bits_ctrl_isMove,
  input        io_enq_req_1_bits_ctrl_singleStep,
  input  [5:0] io_enq_req_1_bits_pdest,
  input  [5:0] io_enq_req_1_bits_old_pdest,
  input        io_enq_req_1_bits_robIdx_flag,
  input  [4:0] io_enq_req_1_bits_robIdx_value,
  input        io_enq_req_1_bits_eliminatedMove,
  output       io_flushOut_valid,
  output       io_flushOut_bits_robIdx_flag,
  output [4:0] io_flushOut_bits_robIdx_value,
  output       io_flushOut_bits_ftqIdx_flag,
  output [2:0] io_flushOut_bits_ftqIdx_value,
  output [2:0] io_flushOut_bits_ftqOffset,
  output       io_flushOut_bits_level,
  output       io_exception_valid,
  output       io_exception_bits_uop_cf_exceptionVec_0,
  output       io_exception_bits_uop_cf_exceptionVec_1,
  output       io_exception_bits_uop_cf_exceptionVec_2,
  output       io_exception_bits_uop_cf_exceptionVec_3,
  output       io_exception_bits_uop_cf_exceptionVec_4,
  output       io_exception_bits_uop_cf_exceptionVec_5,
  output       io_exception_bits_uop_cf_exceptionVec_6,
  output       io_exception_bits_uop_cf_exceptionVec_7,
  output       io_exception_bits_uop_cf_exceptionVec_8,
  output       io_exception_bits_uop_cf_exceptionVec_9,
  output       io_exception_bits_uop_cf_exceptionVec_11,
  output       io_exception_bits_uop_cf_exceptionVec_12,
  output       io_exception_bits_uop_cf_exceptionVec_13,
  output       io_exception_bits_uop_cf_exceptionVec_15,
  output       io_exception_bits_uop_cf_trigger_frontendHit_0,
  output       io_exception_bits_uop_cf_trigger_frontendHit_1,
  output       io_exception_bits_uop_cf_trigger_frontendHit_2,
  output       io_exception_bits_uop_cf_trigger_frontendHit_3,
  output       io_exception_bits_uop_cf_trigger_backendHit_0,
  output       io_exception_bits_uop_cf_trigger_backendHit_1,
  output       io_exception_bits_uop_cf_trigger_backendHit_2,
  output       io_exception_bits_uop_cf_trigger_backendHit_3,
  output       io_exception_bits_uop_cf_trigger_backendHit_4,
  output       io_exception_bits_uop_cf_trigger_backendHit_5,
  output       io_exception_bits_uop_cf_crossPageIPFFix,
  output [2:0] io_exception_bits_uop_ctrl_commitType,
  output       io_exception_bits_uop_ctrl_singleStep,
  output       io_exception_bits_isInterrupt,
  input        io_writeback_1_0_valid,
  input  [4:0] io_writeback_1_0_bits_uop_robIdx_value,
  input        io_writeback_1_0_bits_redirectValid,
  input        io_writeback_1_0_bits_redirect_cfiUpdate_isMisPred,
  input        io_writeback_1_1_valid,
  input  [4:0] io_writeback_1_1_bits_uop_robIdx_value,
  input        io_writeback_1_1_bits_redirectValid,
  input        io_writeback_1_1_bits_redirect_cfiUpdate_isMisPred,
  input        io_writeback_1_2_valid,
  input        io_writeback_1_2_bits_uop_cf_exceptionVec_4,
  input        io_writeback_1_2_bits_uop_cf_exceptionVec_5,
  input        io_writeback_1_2_bits_uop_cf_exceptionVec_13,
  input        io_writeback_1_2_bits_uop_cf_trigger_backendHit_0,
  input        io_writeback_1_2_bits_uop_cf_trigger_backendHit_1,
  input        io_writeback_1_2_bits_uop_cf_trigger_backendHit_2,
  input        io_writeback_1_2_bits_uop_cf_trigger_backendHit_3,
  input        io_writeback_1_2_bits_uop_cf_trigger_backendHit_4,
  input        io_writeback_1_2_bits_uop_cf_trigger_backendHit_5,
  input        io_writeback_1_2_bits_uop_ctrl_flushPipe,
  input        io_writeback_1_2_bits_uop_ctrl_replayInst,
  input  [4:0] io_writeback_1_2_bits_uop_robIdx_value,
  input        io_writeback_1_2_bits_debug_isMMIO,
  input        io_writeback_1_3_valid,
  input        io_writeback_1_3_bits_uop_cf_exceptionVec_4,
  input        io_writeback_1_3_bits_uop_cf_exceptionVec_5,
  input        io_writeback_1_3_bits_uop_cf_exceptionVec_13,
  input        io_writeback_1_3_bits_uop_cf_trigger_backendHit_0,
  input        io_writeback_1_3_bits_uop_cf_trigger_backendHit_1,
  input        io_writeback_1_3_bits_uop_cf_trigger_backendHit_2,
  input        io_writeback_1_3_bits_uop_cf_trigger_backendHit_3,
  input        io_writeback_1_3_bits_uop_cf_trigger_backendHit_4,
  input        io_writeback_1_3_bits_uop_cf_trigger_backendHit_5,
  input        io_writeback_1_3_bits_uop_ctrl_flushPipe,
  input        io_writeback_1_3_bits_uop_ctrl_replayInst,
  input  [4:0] io_writeback_1_3_bits_uop_robIdx_value,
  input        io_writeback_1_3_bits_debug_isMMIO,
  input        io_writeback_1_4_valid,
  input        io_writeback_1_4_bits_uop_cf_exceptionVec_2,
  input        io_writeback_1_4_bits_uop_cf_exceptionVec_3,
  input        io_writeback_1_4_bits_uop_cf_exceptionVec_8,
  input        io_writeback_1_4_bits_uop_cf_exceptionVec_9,
  input        io_writeback_1_4_bits_uop_cf_exceptionVec_11,
  input        io_writeback_1_4_bits_uop_ctrl_flushPipe,
  input  [4:0] io_writeback_1_4_bits_uop_robIdx_value,
  input        io_writeback_1_4_bits_redirectValid,
  input        io_writeback_1_4_bits_redirect_cfiUpdate_isMisPred,
  input        io_writeback_1_4_bits_debug_isPerfCnt,
  input        io_writeback_1_5_valid,
  input        io_writeback_1_5_bits_uop_cf_trigger_backendHit_0,
  input        io_writeback_1_5_bits_uop_cf_trigger_backendHit_1,
  input        io_writeback_1_5_bits_uop_cf_trigger_backendHit_2,
  input        io_writeback_1_5_bits_uop_cf_trigger_backendHit_3,
  input        io_writeback_1_5_bits_uop_cf_trigger_backendHit_4,
  input        io_writeback_1_5_bits_uop_cf_trigger_backendHit_5,
  input  [4:0] io_writeback_1_5_bits_uop_robIdx_value,
  input        io_writeback_1_6_valid,
  input        io_writeback_1_6_bits_uop_cf_exceptionVec_2,
  input        io_writeback_1_6_bits_uop_cf_exceptionVec_3,
  input        io_writeback_1_6_bits_uop_cf_exceptionVec_8,
  input        io_writeback_1_6_bits_uop_cf_exceptionVec_9,
  input        io_writeback_1_6_bits_uop_cf_exceptionVec_11,
  input        io_writeback_1_6_bits_uop_ctrl_flushPipe,
  input  [4:0] io_writeback_1_6_bits_uop_robIdx_value,
  input        io_writeback_1_6_bits_redirectValid,
  input        io_writeback_1_6_bits_redirect_cfiUpdate_isMisPred,
  input        io_writeback_1_6_bits_debug_isPerfCnt,
  input        io_writeback_1_7_valid,
  input        io_writeback_1_7_bits_uop_cf_exceptionVec_4,
  input        io_writeback_1_7_bits_uop_cf_exceptionVec_5,
  input        io_writeback_1_7_bits_uop_cf_exceptionVec_6,
  input        io_writeback_1_7_bits_uop_cf_exceptionVec_7,
  input        io_writeback_1_7_bits_uop_cf_exceptionVec_13,
  input        io_writeback_1_7_bits_uop_cf_exceptionVec_15,
  input        io_writeback_1_7_bits_uop_cf_trigger_backendHit_0,
  input        io_writeback_1_7_bits_uop_cf_trigger_backendHit_1,
  input        io_writeback_1_7_bits_uop_cf_trigger_backendHit_2,
  input        io_writeback_1_7_bits_uop_cf_trigger_backendHit_3,
  input        io_writeback_1_7_bits_uop_cf_trigger_backendHit_4,
  input        io_writeback_1_7_bits_uop_cf_trigger_backendHit_5,
  input  [4:0] io_writeback_1_7_bits_uop_robIdx_value,
  input        io_writeback_1_7_bits_redirectValid,
  input        io_writeback_1_7_bits_redirect_cfiUpdate_isMisPred,
  input        io_writeback_1_7_bits_debug_isMMIO,
  input        io_writeback_1_7_bits_debug_isPerfCnt,
  input        io_writeback_1_8_valid,
  input        io_writeback_1_8_bits_uop_cf_exceptionVec_4,
  input        io_writeback_1_8_bits_uop_cf_exceptionVec_5,
  input        io_writeback_1_8_bits_uop_cf_exceptionVec_6,
  input        io_writeback_1_8_bits_uop_cf_exceptionVec_7,
  input        io_writeback_1_8_bits_uop_cf_exceptionVec_13,
  input        io_writeback_1_8_bits_uop_cf_exceptionVec_15,
  input        io_writeback_1_8_bits_uop_cf_trigger_backendHit_0,
  input        io_writeback_1_8_bits_uop_cf_trigger_backendHit_1,
  input        io_writeback_1_8_bits_uop_cf_trigger_backendHit_2,
  input        io_writeback_1_8_bits_uop_cf_trigger_backendHit_3,
  input        io_writeback_1_8_bits_uop_cf_trigger_backendHit_4,
  input        io_writeback_1_8_bits_uop_cf_trigger_backendHit_5,
  input  [4:0] io_writeback_1_8_bits_uop_robIdx_value,
  input        io_writeback_1_8_bits_redirectValid,
  input        io_writeback_1_8_bits_redirect_cfiUpdate_isMisPred,
  input        io_writeback_1_8_bits_debug_isMMIO,
  input        io_writeback_1_8_bits_debug_isPerfCnt,
  input        io_writeback_1_9_valid,
  input  [4:0] io_writeback_1_9_bits_uop_robIdx_value,
  input        io_writeback_1_10_valid,
  input  [4:0] io_writeback_1_10_bits_uop_robIdx_value,
  input        io_writeback_0_3_valid,
  input        io_writeback_0_3_bits_uop_cf_exceptionVec_2,
  input        io_writeback_0_3_bits_uop_cf_exceptionVec_3,
  input        io_writeback_0_3_bits_uop_cf_exceptionVec_8,
  input        io_writeback_0_3_bits_uop_cf_exceptionVec_9,
  input        io_writeback_0_3_bits_uop_cf_exceptionVec_11,
  input        io_writeback_0_3_bits_uop_ctrl_flushPipe,
  input        io_writeback_0_3_bits_uop_robIdx_flag,
  input  [4:0] io_writeback_0_3_bits_uop_robIdx_value,
  input  [4:0] io_writeback_0_3_bits_fflags,
  input        io_writeback_0_4_valid,
  input  [4:0] io_writeback_0_4_bits_uop_robIdx_value,
  input  [4:0] io_writeback_0_4_bits_fflags,
  input        io_writeback_0_5_valid,
  input  [4:0] io_writeback_0_5_bits_uop_robIdx_value,
  input  [4:0] io_writeback_0_5_bits_fflags,
  input        io_writeback_0_6_valid,
  input        io_writeback_0_6_bits_uop_cf_exceptionVec_4,
  input        io_writeback_0_6_bits_uop_cf_exceptionVec_5,
  input        io_writeback_0_6_bits_uop_cf_exceptionVec_13,
  input        io_writeback_0_6_bits_uop_cf_trigger_backendHit_0,
  input        io_writeback_0_6_bits_uop_cf_trigger_backendHit_1,
  input        io_writeback_0_6_bits_uop_cf_trigger_backendHit_2,
  input        io_writeback_0_6_bits_uop_cf_trigger_backendHit_3,
  input        io_writeback_0_6_bits_uop_cf_trigger_backendHit_4,
  input        io_writeback_0_6_bits_uop_cf_trigger_backendHit_5,
  input        io_writeback_0_6_bits_uop_ctrl_flushPipe,
  input        io_writeback_0_6_bits_uop_ctrl_replayInst,
  input        io_writeback_0_6_bits_uop_robIdx_flag,
  input  [4:0] io_writeback_0_6_bits_uop_robIdx_value,
  input        io_writeback_0_7_valid,
  input        io_writeback_0_7_bits_uop_cf_exceptionVec_4,
  input        io_writeback_0_7_bits_uop_cf_exceptionVec_5,
  input        io_writeback_0_7_bits_uop_cf_exceptionVec_13,
  input        io_writeback_0_7_bits_uop_cf_trigger_backendHit_0,
  input        io_writeback_0_7_bits_uop_cf_trigger_backendHit_1,
  input        io_writeback_0_7_bits_uop_cf_trigger_backendHit_2,
  input        io_writeback_0_7_bits_uop_cf_trigger_backendHit_3,
  input        io_writeback_0_7_bits_uop_cf_trigger_backendHit_4,
  input        io_writeback_0_7_bits_uop_cf_trigger_backendHit_5,
  input        io_writeback_0_7_bits_uop_ctrl_flushPipe,
  input        io_writeback_0_7_bits_uop_ctrl_replayInst,
  input        io_writeback_0_7_bits_uop_robIdx_flag,
  input  [4:0] io_writeback_0_7_bits_uop_robIdx_value,
  input        io_writeback_0_8_valid,
  input        io_writeback_0_8_bits_uop_cf_exceptionVec_4,
  input        io_writeback_0_8_bits_uop_cf_exceptionVec_5,
  input        io_writeback_0_8_bits_uop_cf_exceptionVec_6,
  input        io_writeback_0_8_bits_uop_cf_exceptionVec_7,
  input        io_writeback_0_8_bits_uop_cf_exceptionVec_13,
  input        io_writeback_0_8_bits_uop_cf_exceptionVec_15,
  input        io_writeback_0_8_bits_uop_cf_trigger_backendHit_0,
  input        io_writeback_0_8_bits_uop_cf_trigger_backendHit_1,
  input        io_writeback_0_8_bits_uop_cf_trigger_backendHit_2,
  input        io_writeback_0_8_bits_uop_cf_trigger_backendHit_3,
  input        io_writeback_0_8_bits_uop_cf_trigger_backendHit_4,
  input        io_writeback_0_8_bits_uop_cf_trigger_backendHit_5,
  input        io_writeback_0_8_bits_uop_robIdx_flag,
  input  [4:0] io_writeback_0_8_bits_uop_robIdx_value,
  input        io_writeback_0_9_valid,
  input        io_writeback_0_9_bits_uop_cf_exceptionVec_6,
  input        io_writeback_0_9_bits_uop_cf_exceptionVec_7,
  input        io_writeback_0_9_bits_uop_cf_exceptionVec_15,
  input        io_writeback_0_9_bits_uop_cf_trigger_backendHit_0,
  input        io_writeback_0_9_bits_uop_cf_trigger_backendHit_1,
  input        io_writeback_0_9_bits_uop_cf_trigger_backendHit_4,
  input        io_writeback_0_9_bits_uop_robIdx_flag,
  input  [4:0] io_writeback_0_9_bits_uop_robIdx_value,
  output       io_commits_isCommit,
  output       io_commits_commitValid_0,
  output       io_commits_commitValid_1,
  output       io_commits_isWalk,
  output       io_commits_walkValid_0,
  output       io_commits_walkValid_1,
  output [4:0] io_commits_info_0_ldest,
  output       io_commits_info_0_rfWen,
  output       io_commits_info_0_fpWen,
  output       io_commits_info_0_wflags,
  output [2:0] io_commits_info_0_commitType,
  output [5:0] io_commits_info_0_pdest,
  output [5:0] io_commits_info_0_old_pdest,
  output       io_commits_info_0_ftqIdx_flag,
  output [2:0] io_commits_info_0_ftqIdx_value,
  output [2:0] io_commits_info_0_ftqOffset,
  output       io_commits_info_0_isMove,
  output [4:0] io_commits_info_1_ldest,
  output       io_commits_info_1_rfWen,
  output       io_commits_info_1_fpWen,
  output       io_commits_info_1_wflags,
  output [2:0] io_commits_info_1_commitType,
  output [5:0] io_commits_info_1_pdest,
  output [5:0] io_commits_info_1_old_pdest,
  output       io_commits_info_1_ftqIdx_flag,
  output [2:0] io_commits_info_1_ftqIdx_value,
  output [2:0] io_commits_info_1_ftqOffset,
  output       io_commits_info_1_isMove,
  output [1:0] io_lsq_scommit,
  output       io_lsq_pendingld,
  output       io_lsq_pendingst,
  output       io_lsq_commit,
  input        io_lsq_isMMIO_0,
  input        io_lsq_isMMIO_1,
  input  [4:0] io_lsq_uop_0_robIdx_value,
  input  [4:0] io_lsq_uop_1_robIdx_value,
  input        io_csr_intrBitSet,
  input        io_csr_wfiEvent,
  output       io_csr_fflags_valid,
  output [4:0] io_csr_fflags_bits,
  output       io_csr_dirty_fs,
  output [2:0] io_csr_perfinfo_retiredInstr,
  output       io_cpu_halt,
  input        io_wfi_enable,
  output [5:0] io_perf_0_value,
  output [5:0] io_perf_1_value,
  output [5:0] io_perf_2_value,
  output [5:0] io_perf_3_value,
  output [5:0] io_perf_4_value,
  output [5:0] io_perf_5_value,
  output [5:0] io_perf_6_value,
  output [5:0] io_perf_7_value,
  output [5:0] io_perf_8_value,
  output [5:0] io_perf_9_value,
  output [5:0] io_perf_10_value,
  output [5:0] io_perf_11_value,
  output [5:0] io_perf_12_value,
  output [5:0] io_perf_13_value,
  output [5:0] io_perf_14_value,
  output [5:0] io_perf_15_value,
  output [5:0] io_perf_16_value,
  output [5:0] io_perf_17_value
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [63:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [63:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
`endif // RANDOMIZE_REG_INIT
  reg  writebacked [0:31]; // @[Rob.scala 428:24]
  wire  writebacked_exceptionEnable_MPORT_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_exceptionEnable_MPORT_addr; // @[Rob.scala 428:24]
  wire  writebacked_exceptionEnable_MPORT_data; // @[Rob.scala 428:24]
  wire  writebacked_isFlushPipe_MPORT_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_isFlushPipe_MPORT_addr; // @[Rob.scala 428:24]
  wire  writebacked_isFlushPipe_MPORT_data; // @[Rob.scala 428:24]
  wire  writebacked_commit_wMPORT_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_commit_wMPORT_addr; // @[Rob.scala 428:24]
  wire  writebacked_commit_wMPORT_data; // @[Rob.scala 428:24]
  wire  writebacked_commit_wMPORT_2_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_commit_wMPORT_2_addr; // @[Rob.scala 428:24]
  wire  writebacked_commit_wMPORT_2_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_113_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_113_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_113_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_114_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_114_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_114_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_115_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_115_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_115_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_116_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_116_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_116_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_117_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_117_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_117_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_118_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_118_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_118_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_119_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_119_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_119_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_120_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_120_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_120_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_121_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_121_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_121_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_122_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_122_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_122_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_123_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_123_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_123_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_124_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_124_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_124_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_125_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_125_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_125_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_126_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_126_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_126_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_127_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_127_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_127_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_128_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_128_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_128_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_129_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_129_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_129_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_130_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_130_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_130_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_131_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_131_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_131_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_132_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_132_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_132_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_133_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_133_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_133_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_134_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_134_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_134_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_135_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_135_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_135_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_136_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_136_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_136_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_137_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_137_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_137_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_138_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_138_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_138_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_139_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_139_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_139_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_140_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_140_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_140_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_141_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_141_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_141_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_142_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_142_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_142_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_143_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_143_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_143_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_144_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_144_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_144_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_145_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_145_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_145_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_146_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_146_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_146_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_147_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_147_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_147_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_148_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_148_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_148_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_149_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_149_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_149_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_150_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_150_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_150_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_151_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_151_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_151_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_152_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_152_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_152_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_153_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_153_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_153_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_154_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_154_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_154_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_155_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_155_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_155_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_156_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_156_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_156_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_157_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_157_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_157_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_158_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_158_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_158_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_159_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_159_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_159_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_160_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_160_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_160_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_161_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_161_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_161_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_162_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_162_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_162_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_163_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_163_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_163_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_164_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_164_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_164_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_165_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_165_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_165_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_166_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_166_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_166_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_167_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_167_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_167_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_168_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_168_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_168_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_169_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_169_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_169_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_170_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_170_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_170_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_171_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_171_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_171_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_172_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_172_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_172_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_173_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_173_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_173_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_174_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_174_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_174_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_175_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_175_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_175_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_176_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_176_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_176_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_178_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_178_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_178_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_179_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_179_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_179_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_181_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_181_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_181_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_182_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_182_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_182_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_184_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_184_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_184_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_185_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_185_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_185_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_187_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_187_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_187_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_188_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_188_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_188_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_190_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_190_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_190_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_191_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_191_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_191_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_193_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_193_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_193_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_194_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_194_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_194_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_196_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_196_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_196_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_197_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_197_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_197_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_199_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_199_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_199_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_200_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_200_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_200_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_202_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_202_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_202_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_203_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_203_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_203_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_205_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_205_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_205_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_206_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_206_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_206_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_208_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_208_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_208_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_209_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_209_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_209_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_211_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_211_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_211_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_212_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_212_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_212_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_214_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_214_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_214_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_215_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_215_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_215_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_217_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_217_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_217_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_218_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_218_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_218_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_220_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_220_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_220_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_221_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_221_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_221_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_223_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_223_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_223_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_224_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_224_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_224_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_226_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_226_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_226_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_227_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_227_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_227_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_229_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_229_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_229_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_230_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_230_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_230_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_232_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_232_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_232_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_233_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_233_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_233_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_235_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_235_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_235_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_236_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_236_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_236_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_238_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_238_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_238_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_239_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_239_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_239_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_241_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_241_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_241_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_242_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_242_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_242_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_244_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_244_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_244_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_245_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_245_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_245_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_247_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_247_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_247_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_248_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_248_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_248_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_250_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_250_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_250_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_251_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_251_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_251_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_253_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_253_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_253_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_254_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_254_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_254_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_256_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_256_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_256_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_257_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_257_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_257_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_259_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_259_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_259_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_260_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_260_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_260_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_262_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_262_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_262_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_263_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_263_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_263_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_265_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_265_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_265_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_266_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_266_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_266_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_268_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_268_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_268_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_269_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_269_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_269_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_271_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_271_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_271_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_272_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_272_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_272_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_273_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_273_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_273_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_274_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_274_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_274_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_275_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_275_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_275_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_276_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_276_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_276_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_277_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_277_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_277_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_278_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_278_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_278_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_279_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_279_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_279_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_280_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_280_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_280_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_281_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_281_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_281_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_282_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_282_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_282_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_283_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_283_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_283_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_284_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_284_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_284_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_285_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_285_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_285_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_286_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_286_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_286_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_287_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_287_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_287_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_288_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_288_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_288_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_289_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_289_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_289_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_290_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_290_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_290_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_291_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_291_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_291_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_292_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_292_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_292_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_293_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_293_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_293_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_294_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_294_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_294_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_295_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_295_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_295_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_296_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_296_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_296_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_297_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_297_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_297_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_298_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_298_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_298_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_299_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_299_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_299_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_300_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_300_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_300_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_301_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_301_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_301_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_302_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_302_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_302_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_303_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_303_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_303_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_304_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_304_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_304_data; // @[Rob.scala 428:24]
  wire  writebacked_deqNotWritebacked_MPORT_en; // @[Rob.scala 428:24]
  wire [4:0] writebacked_deqNotWritebacked_MPORT_addr; // @[Rob.scala 428:24]
  wire  writebacked_deqNotWritebacked_MPORT_data; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_92_data; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_92_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_92_mask; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_92_en; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_94_data; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_94_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_94_mask; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_94_en; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_96_data; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_96_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_96_mask; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_96_en; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_98_data; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_98_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_98_mask; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_98_en; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_99_data; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_99_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_99_mask; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_99_en; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_100_data; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_100_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_100_mask; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_100_en; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_101_data; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_101_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_101_mask; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_101_en; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_102_data; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_102_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_102_mask; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_102_en; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_103_data; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_103_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_103_mask; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_103_en; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_104_data; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_104_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_104_mask; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_104_en; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_105_data; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_105_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_105_mask; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_105_en; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_106_data; // @[Rob.scala 428:24]
  wire [4:0] writebacked_MPORT_106_addr; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_106_mask; // @[Rob.scala 428:24]
  wire  writebacked_MPORT_106_en; // @[Rob.scala 428:24]
  reg  store_data_writebacked [0:31]; // @[Rob.scala 429:35]
  wire  store_data_writebacked_commit_wMPORT_1_en; // @[Rob.scala 429:35]
  wire [4:0] store_data_writebacked_commit_wMPORT_1_addr; // @[Rob.scala 429:35]
  wire  store_data_writebacked_commit_wMPORT_1_data; // @[Rob.scala 429:35]
  wire  store_data_writebacked_commit_wMPORT_3_en; // @[Rob.scala 429:35]
  wire [4:0] store_data_writebacked_commit_wMPORT_3_addr; // @[Rob.scala 429:35]
  wire  store_data_writebacked_commit_wMPORT_3_data; // @[Rob.scala 429:35]
  wire  store_data_writebacked_MPORT_93_data; // @[Rob.scala 429:35]
  wire [4:0] store_data_writebacked_MPORT_93_addr; // @[Rob.scala 429:35]
  wire  store_data_writebacked_MPORT_93_mask; // @[Rob.scala 429:35]
  wire  store_data_writebacked_MPORT_93_en; // @[Rob.scala 429:35]
  wire  store_data_writebacked_MPORT_95_data; // @[Rob.scala 429:35]
  wire [4:0] store_data_writebacked_MPORT_95_addr; // @[Rob.scala 429:35]
  wire  store_data_writebacked_MPORT_95_mask; // @[Rob.scala 429:35]
  wire  store_data_writebacked_MPORT_95_en; // @[Rob.scala 429:35]
  wire  store_data_writebacked_MPORT_97_data; // @[Rob.scala 429:35]
  wire [4:0] store_data_writebacked_MPORT_97_addr; // @[Rob.scala 429:35]
  wire  store_data_writebacked_MPORT_97_mask; // @[Rob.scala 429:35]
  wire  store_data_writebacked_MPORT_97_en; // @[Rob.scala 429:35]
  wire  store_data_writebacked_MPORT_107_data; // @[Rob.scala 429:35]
  wire [4:0] store_data_writebacked_MPORT_107_addr; // @[Rob.scala 429:35]
  wire  store_data_writebacked_MPORT_107_mask; // @[Rob.scala 429:35]
  wire  store_data_writebacked_MPORT_107_en; // @[Rob.scala 429:35]
  wire  store_data_writebacked_MPORT_108_data; // @[Rob.scala 429:35]
  wire [4:0] store_data_writebacked_MPORT_108_addr; // @[Rob.scala 429:35]
  wire  store_data_writebacked_MPORT_108_mask; // @[Rob.scala 429:35]
  wire  store_data_writebacked_MPORT_108_en; // @[Rob.scala 429:35]
  reg  interrupt_safe [0:31]; // @[Rob.scala 436:27]
  wire  interrupt_safe_intrEnable_MPORT_en; // @[Rob.scala 436:27]
  wire [4:0] interrupt_safe_intrEnable_MPORT_addr; // @[Rob.scala 436:27]
  wire  interrupt_safe_intrEnable_MPORT_data; // @[Rob.scala 436:27]
  wire  interrupt_safe_deqPtrGenModule_io_interrupt_safe_MPORT_en; // @[Rob.scala 436:27]
  wire [4:0] interrupt_safe_deqPtrGenModule_io_interrupt_safe_MPORT_addr; // @[Rob.scala 436:27]
  wire  interrupt_safe_deqPtrGenModule_io_interrupt_safe_MPORT_data; // @[Rob.scala 436:27]
  wire  interrupt_safe_MPORT_111_data; // @[Rob.scala 436:27]
  wire [4:0] interrupt_safe_MPORT_111_addr; // @[Rob.scala 436:27]
  wire  interrupt_safe_MPORT_111_mask; // @[Rob.scala 436:27]
  wire  interrupt_safe_MPORT_111_en; // @[Rob.scala 436:27]
  wire  interrupt_safe_MPORT_112_data; // @[Rob.scala 436:27]
  wire [4:0] interrupt_safe_MPORT_112_addr; // @[Rob.scala 436:27]
  wire  interrupt_safe_MPORT_112_mask; // @[Rob.scala 436:27]
  wire  interrupt_safe_MPORT_112_en; // @[Rob.scala 436:27]
  reg  debug_microOp_cf_loadWaitBit [0:31]; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_debug_deqUop_en; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_debug_deqUop_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_debug_deqUop_data; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_commitDebugUop_0_en; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_commitDebugUop_0_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_commitDebugUop_0_data; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_commitDebugUop_1_en; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_commitDebugUop_1_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_commitDebugUop_1_data; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_1_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_1_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_1_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_1_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_2_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_2_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_2_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_2_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_3_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_3_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_3_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_3_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_4_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_4_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_4_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_4_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_5_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_5_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_5_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_5_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_6_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_6_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_6_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_6_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_7_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_7_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_7_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_7_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_8_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_8_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_8_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_8_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_9_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_9_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_9_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_9_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_10_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_10_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_10_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_10_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_11_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_11_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_11_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_11_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_12_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_12_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_12_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_12_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_13_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_13_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_13_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_13_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_14_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_14_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_14_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_14_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_15_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_15_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_15_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_15_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_16_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_16_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_16_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_16_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_17_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_17_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_17_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_17_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_18_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_18_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_18_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_18_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_19_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_19_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_19_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_19_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_20_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_20_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_20_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_20_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_21_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_21_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_21_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_21_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_22_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_22_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_22_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_22_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_23_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_23_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_23_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_23_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_24_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_24_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_24_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_24_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_25_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_25_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_25_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_25_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_26_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_26_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_26_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_26_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_27_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_27_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_27_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_27_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_28_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_28_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_28_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_28_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_29_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_29_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_29_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_29_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_30_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_30_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_30_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_30_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_31_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_31_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_31_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_31_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_32_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_32_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_32_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_32_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_33_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_33_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_33_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_33_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_34_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_34_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_34_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_34_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_35_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_35_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_35_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_35_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_36_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_36_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_36_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_36_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_37_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_37_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_37_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_37_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_38_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_38_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_38_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_38_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_39_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_39_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_39_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_39_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_40_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_40_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_40_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_40_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_41_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_41_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_41_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_41_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_42_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_42_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_42_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_42_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_43_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_43_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_43_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_43_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_44_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_44_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_44_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_44_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_45_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_45_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_45_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_45_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_46_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_46_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_46_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_46_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_47_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_47_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_47_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_47_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_48_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_48_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_48_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_48_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_49_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_49_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_49_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_49_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_50_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_50_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_50_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_50_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_51_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_51_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_51_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_51_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_52_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_52_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_52_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_52_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_53_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_53_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_53_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_53_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_54_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_54_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_54_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_54_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_55_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_55_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_55_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_55_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_56_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_56_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_56_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_56_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_57_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_57_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_57_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_57_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_58_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_58_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_58_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_58_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_59_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_59_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_59_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_59_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_60_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_60_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_60_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_60_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_61_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_61_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_61_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_61_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_62_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_62_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_62_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_62_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_63_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_63_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_63_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_63_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_64_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_64_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_64_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_64_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_65_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_65_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_65_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_65_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_66_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_66_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_66_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_66_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_67_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_67_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_67_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_67_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_68_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_68_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_68_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_68_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_69_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_69_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_69_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_69_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_70_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_70_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_70_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_70_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_71_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_71_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_71_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_71_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_72_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_72_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_72_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_72_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_73_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_73_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_73_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_73_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_74_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_74_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_74_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_74_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_75_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_75_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_75_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_75_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_76_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_76_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_76_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_76_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_77_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_77_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_77_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_77_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_78_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_78_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_78_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_78_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_79_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_79_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_79_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_79_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_80_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_80_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_80_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_80_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_81_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_81_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_81_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_81_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_82_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_82_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_82_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_82_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_83_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_83_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_83_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_83_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_84_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_84_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_84_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_84_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_85_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_85_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_85_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_85_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_86_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_86_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_86_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_86_en; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_87_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_cf_loadWaitBit_MPORT_87_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_87_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_cf_loadWaitBit_MPORT_87_en; // @[Rob.scala 440:26]
  reg  debug_microOp_ctrl_isMove [0:31]; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_debug_deqUop_en; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_debug_deqUop_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_debug_deqUop_data; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_commitDebugUop_0_en; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_commitDebugUop_0_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_commitDebugUop_0_data; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_commitDebugUop_1_en; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_commitDebugUop_1_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_commitDebugUop_1_data; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_1_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_1_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_1_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_1_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_2_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_2_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_2_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_2_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_3_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_3_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_3_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_3_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_4_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_4_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_4_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_4_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_5_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_5_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_5_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_5_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_6_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_6_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_6_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_6_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_7_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_7_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_7_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_7_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_8_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_8_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_8_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_8_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_9_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_9_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_9_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_9_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_10_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_10_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_10_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_10_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_11_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_11_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_11_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_11_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_12_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_12_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_12_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_12_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_13_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_13_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_13_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_13_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_14_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_14_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_14_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_14_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_15_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_15_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_15_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_15_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_16_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_16_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_16_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_16_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_17_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_17_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_17_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_17_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_18_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_18_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_18_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_18_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_19_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_19_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_19_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_19_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_20_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_20_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_20_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_20_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_21_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_21_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_21_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_21_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_22_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_22_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_22_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_22_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_23_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_23_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_23_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_23_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_24_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_24_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_24_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_24_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_25_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_25_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_25_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_25_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_26_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_26_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_26_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_26_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_27_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_27_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_27_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_27_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_28_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_28_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_28_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_28_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_29_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_29_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_29_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_29_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_30_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_30_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_30_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_30_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_31_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_31_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_31_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_31_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_32_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_32_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_32_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_32_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_33_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_33_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_33_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_33_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_34_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_34_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_34_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_34_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_35_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_35_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_35_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_35_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_36_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_36_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_36_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_36_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_37_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_37_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_37_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_37_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_38_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_38_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_38_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_38_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_39_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_39_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_39_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_39_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_40_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_40_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_40_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_40_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_41_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_41_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_41_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_41_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_42_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_42_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_42_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_42_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_43_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_43_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_43_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_43_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_44_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_44_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_44_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_44_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_45_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_45_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_45_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_45_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_46_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_46_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_46_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_46_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_47_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_47_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_47_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_47_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_48_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_48_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_48_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_48_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_49_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_49_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_49_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_49_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_50_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_50_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_50_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_50_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_51_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_51_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_51_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_51_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_52_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_52_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_52_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_52_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_53_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_53_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_53_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_53_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_54_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_54_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_54_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_54_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_55_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_55_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_55_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_55_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_56_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_56_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_56_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_56_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_57_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_57_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_57_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_57_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_58_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_58_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_58_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_58_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_59_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_59_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_59_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_59_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_60_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_60_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_60_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_60_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_61_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_61_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_61_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_61_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_62_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_62_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_62_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_62_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_63_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_63_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_63_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_63_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_64_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_64_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_64_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_64_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_65_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_65_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_65_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_65_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_66_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_66_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_66_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_66_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_67_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_67_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_67_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_67_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_68_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_68_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_68_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_68_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_69_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_69_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_69_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_69_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_70_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_70_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_70_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_70_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_71_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_71_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_71_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_71_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_72_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_72_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_72_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_72_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_73_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_73_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_73_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_73_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_74_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_74_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_74_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_74_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_75_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_75_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_75_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_75_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_76_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_76_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_76_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_76_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_77_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_77_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_77_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_77_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_78_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_78_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_78_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_78_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_79_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_79_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_79_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_79_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_80_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_80_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_80_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_80_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_81_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_81_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_81_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_81_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_82_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_82_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_82_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_82_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_83_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_83_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_83_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_83_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_84_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_84_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_84_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_84_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_85_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_85_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_85_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_85_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_86_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_86_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_86_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_86_en; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_87_data; // @[Rob.scala 440:26]
  wire [4:0] debug_microOp_ctrl_isMove_MPORT_87_addr; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_87_mask; // @[Rob.scala 440:26]
  wire  debug_microOp_ctrl_isMove_MPORT_87_en; // @[Rob.scala 440:26]
  wire  dispatchData_clock; // @[Rob.scala 477:28]
  wire [4:0] dispatchData_io_raddr_0; // @[Rob.scala 477:28]
  wire [4:0] dispatchData_io_raddr_1; // @[Rob.scala 477:28]
  wire [4:0] dispatchData_io_rdata_0_ldest; // @[Rob.scala 477:28]
  wire  dispatchData_io_rdata_0_rfWen; // @[Rob.scala 477:28]
  wire  dispatchData_io_rdata_0_fpWen; // @[Rob.scala 477:28]
  wire  dispatchData_io_rdata_0_wflags; // @[Rob.scala 477:28]
  wire [2:0] dispatchData_io_rdata_0_commitType; // @[Rob.scala 477:28]
  wire [5:0] dispatchData_io_rdata_0_pdest; // @[Rob.scala 477:28]
  wire [5:0] dispatchData_io_rdata_0_old_pdest; // @[Rob.scala 477:28]
  wire  dispatchData_io_rdata_0_ftqIdx_flag; // @[Rob.scala 477:28]
  wire [2:0] dispatchData_io_rdata_0_ftqIdx_value; // @[Rob.scala 477:28]
  wire [2:0] dispatchData_io_rdata_0_ftqOffset; // @[Rob.scala 477:28]
  wire  dispatchData_io_rdata_0_isMove; // @[Rob.scala 477:28]
  wire [4:0] dispatchData_io_rdata_1_ldest; // @[Rob.scala 477:28]
  wire  dispatchData_io_rdata_1_rfWen; // @[Rob.scala 477:28]
  wire  dispatchData_io_rdata_1_fpWen; // @[Rob.scala 477:28]
  wire  dispatchData_io_rdata_1_wflags; // @[Rob.scala 477:28]
  wire [2:0] dispatchData_io_rdata_1_commitType; // @[Rob.scala 477:28]
  wire [5:0] dispatchData_io_rdata_1_pdest; // @[Rob.scala 477:28]
  wire [5:0] dispatchData_io_rdata_1_old_pdest; // @[Rob.scala 477:28]
  wire  dispatchData_io_rdata_1_ftqIdx_flag; // @[Rob.scala 477:28]
  wire [2:0] dispatchData_io_rdata_1_ftqIdx_value; // @[Rob.scala 477:28]
  wire [2:0] dispatchData_io_rdata_1_ftqOffset; // @[Rob.scala 477:28]
  wire  dispatchData_io_rdata_1_isMove; // @[Rob.scala 477:28]
  wire  dispatchData_io_wen_0; // @[Rob.scala 477:28]
  wire  dispatchData_io_wen_1; // @[Rob.scala 477:28]
  wire [4:0] dispatchData_io_waddr_0; // @[Rob.scala 477:28]
  wire [4:0] dispatchData_io_waddr_1; // @[Rob.scala 477:28]
  wire [4:0] dispatchData_io_wdata_0_ldest; // @[Rob.scala 477:28]
  wire  dispatchData_io_wdata_0_rfWen; // @[Rob.scala 477:28]
  wire  dispatchData_io_wdata_0_fpWen; // @[Rob.scala 477:28]
  wire  dispatchData_io_wdata_0_wflags; // @[Rob.scala 477:28]
  wire [2:0] dispatchData_io_wdata_0_commitType; // @[Rob.scala 477:28]
  wire [5:0] dispatchData_io_wdata_0_pdest; // @[Rob.scala 477:28]
  wire [5:0] dispatchData_io_wdata_0_old_pdest; // @[Rob.scala 477:28]
  wire  dispatchData_io_wdata_0_ftqIdx_flag; // @[Rob.scala 477:28]
  wire [2:0] dispatchData_io_wdata_0_ftqIdx_value; // @[Rob.scala 477:28]
  wire [2:0] dispatchData_io_wdata_0_ftqOffset; // @[Rob.scala 477:28]
  wire  dispatchData_io_wdata_0_isMove; // @[Rob.scala 477:28]
  wire [4:0] dispatchData_io_wdata_1_ldest; // @[Rob.scala 477:28]
  wire  dispatchData_io_wdata_1_rfWen; // @[Rob.scala 477:28]
  wire  dispatchData_io_wdata_1_fpWen; // @[Rob.scala 477:28]
  wire  dispatchData_io_wdata_1_wflags; // @[Rob.scala 477:28]
  wire [2:0] dispatchData_io_wdata_1_commitType; // @[Rob.scala 477:28]
  wire [5:0] dispatchData_io_wdata_1_pdest; // @[Rob.scala 477:28]
  wire [5:0] dispatchData_io_wdata_1_old_pdest; // @[Rob.scala 477:28]
  wire  dispatchData_io_wdata_1_ftqIdx_flag; // @[Rob.scala 477:28]
  wire [2:0] dispatchData_io_wdata_1_ftqIdx_value; // @[Rob.scala 477:28]
  wire [2:0] dispatchData_io_wdata_1_ftqOffset; // @[Rob.scala 477:28]
  wire  dispatchData_io_wdata_1_isMove; // @[Rob.scala 477:28]
  wire  exceptionGen_clock; // @[Rob.scala 480:28]
  wire  exceptionGen_reset; // @[Rob.scala 480:28]
  wire  exceptionGen_io_redirect_valid; // @[Rob.scala 480:28]
  wire  exceptionGen_io_redirect_bits_robIdx_flag; // @[Rob.scala 480:28]
  wire [4:0] exceptionGen_io_redirect_bits_robIdx_value; // @[Rob.scala 480:28]
  wire  exceptionGen_io_redirect_bits_level; // @[Rob.scala 480:28]
  wire  exceptionGen_io_flush; // @[Rob.scala 480:28]
  wire  exceptionGen_io_enq_0_valid; // @[Rob.scala 480:28]
  wire  exceptionGen_io_enq_0_bits_robIdx_flag; // @[Rob.scala 480:28]
  wire [4:0] exceptionGen_io_enq_0_bits_robIdx_value; // @[Rob.scala 480:28]
  wire  exceptionGen_io_enq_0_bits_exceptionVec_1; // @[Rob.scala 480:28]
  wire  exceptionGen_io_enq_0_bits_exceptionVec_2; // @[Rob.scala 480:28]
  wire  exceptionGen_io_enq_0_bits_exceptionVec_12; // @[Rob.scala 480:28]
  wire  exceptionGen_io_enq_0_bits_flushPipe; // @[Rob.scala 480:28]
  wire  exceptionGen_io_enq_0_bits_singleStep; // @[Rob.scala 480:28]
  wire  exceptionGen_io_enq_0_bits_crossPageIPFFix; // @[Rob.scala 480:28]
  wire  exceptionGen_io_enq_0_bits_trigger_frontendHit_0; // @[Rob.scala 480:28]
  wire  exceptionGen_io_enq_0_bits_trigger_frontendHit_1; // @[Rob.scala 480:28]
  wire  exceptionGen_io_enq_0_bits_trigger_frontendHit_2; // @[Rob.scala 480:28]
  wire  exceptionGen_io_enq_0_bits_trigger_frontendHit_3; // @[Rob.scala 480:28]
  wire  exceptionGen_io_enq_1_valid; // @[Rob.scala 480:28]
  wire  exceptionGen_io_enq_1_bits_robIdx_flag; // @[Rob.scala 480:28]
  wire [4:0] exceptionGen_io_enq_1_bits_robIdx_value; // @[Rob.scala 480:28]
  wire  exceptionGen_io_enq_1_bits_exceptionVec_1; // @[Rob.scala 480:28]
  wire  exceptionGen_io_enq_1_bits_exceptionVec_2; // @[Rob.scala 480:28]
  wire  exceptionGen_io_enq_1_bits_exceptionVec_12; // @[Rob.scala 480:28]
  wire  exceptionGen_io_enq_1_bits_flushPipe; // @[Rob.scala 480:28]
  wire  exceptionGen_io_enq_1_bits_singleStep; // @[Rob.scala 480:28]
  wire  exceptionGen_io_enq_1_bits_crossPageIPFFix; // @[Rob.scala 480:28]
  wire  exceptionGen_io_enq_1_bits_trigger_frontendHit_0; // @[Rob.scala 480:28]
  wire  exceptionGen_io_enq_1_bits_trigger_frontendHit_1; // @[Rob.scala 480:28]
  wire  exceptionGen_io_enq_1_bits_trigger_frontendHit_2; // @[Rob.scala 480:28]
  wire  exceptionGen_io_enq_1_bits_trigger_frontendHit_3; // @[Rob.scala 480:28]
  wire  exceptionGen_io_wb_0_valid; // @[Rob.scala 480:28]
  wire  exceptionGen_io_wb_0_bits_robIdx_flag; // @[Rob.scala 480:28]
  wire [4:0] exceptionGen_io_wb_0_bits_robIdx_value; // @[Rob.scala 480:28]
  wire  exceptionGen_io_wb_0_bits_exceptionVec_2; // @[Rob.scala 480:28]
  wire  exceptionGen_io_wb_0_bits_exceptionVec_3; // @[Rob.scala 480:28]
  wire  exceptionGen_io_wb_0_bits_exceptionVec_8; // @[Rob.scala 480:28]
  wire  exceptionGen_io_wb_0_bits_exceptionVec_9; // @[Rob.scala 480:28]
  wire  exceptionGen_io_wb_0_bits_exceptionVec_11; // @[Rob.scala 480:28]
  wire  exceptionGen_io_wb_0_bits_flushPipe; // @[Rob.scala 480:28]
  wire  exceptionGen_io_wb_1_valid; // @[Rob.scala 480:28]
  wire  exceptionGen_io_wb_1_bits_robIdx_flag; // @[Rob.scala 480:28]
  wire [4:0] exceptionGen_io_wb_1_bits_robIdx_value; // @[Rob.scala 480:28]
  wire  exceptionGen_io_wb_1_bits_exceptionVec_4; // @[Rob.scala 480:28]
  wire  exceptionGen_io_wb_1_bits_exceptionVec_5; // @[Rob.scala 480:28]
  wire  exceptionGen_io_wb_1_bits_exceptionVec_13; // @[Rob.scala 480:28]
  wire  exceptionGen_io_wb_1_bits_flushPipe; // @[Rob.scala 480:28]
  wire  exceptionGen_io_wb_1_bits_replayInst; // @[Rob.scala 480:28]
  wire  exceptionGen_io_wb_1_bits_trigger_backendHit_0; // @[Rob.scala 480:28]
  wire  exceptionGen_io_wb_1_bits_trigger_backendHit_1; // @[Rob.scala 480:28]
  wire  exceptionGen_io_wb_1_bits_trigger_backendHit_2; // @[Rob.scala 480:28]
  wire  exceptionGen_io_wb_1_bits_trigger_backendHit_3; // @[Rob.scala 480:28]
  wire  exceptionGen_io_wb_1_bits_trigger_backendHit_4; // @[Rob.scala 480:28]
  wire  exceptionGen_io_wb_1_bits_trigger_backendHit_5; // @[Rob.scala 480:28]
  wire  exceptionGen_io_wb_2_valid; // @[Rob.scala 480:28]
  wire  exceptionGen_io_wb_2_bits_robIdx_flag; // @[Rob.scala 480:28]
  wire [4:0] exceptionGen_io_wb_2_bits_robIdx_value; // @[Rob.scala 480:28]
  wire  exceptionGen_io_wb_2_bits_exceptionVec_4; // @[Rob.scala 480:28]
  wire  exceptionGen_io_wb_2_bits_exceptionVec_5; // @[Rob.scala 480:28]
  wire  exceptionGen_io_wb_2_bits_exceptionVec_13; // @[Rob.scala 480:28]
  wire  exceptionGen_io_wb_2_bits_flushPipe; // @[Rob.scala 480:28]
  wire  exceptionGen_io_wb_2_bits_replayInst; // @[Rob.scala 480:28]
  wire  exceptionGen_io_wb_2_bits_trigger_backendHit_0; // @[Rob.scala 480:28]
  wire  exceptionGen_io_wb_2_bits_trigger_backendHit_1; // @[Rob.scala 480:28]
  wire  exceptionGen_io_wb_2_bits_trigger_backendHit_2; // @[Rob.scala 480:28]
  wire  exceptionGen_io_wb_2_bits_trigger_backendHit_3; // @[Rob.scala 480:28]
  wire  exceptionGen_io_wb_2_bits_trigger_backendHit_4; // @[Rob.scala 480:28]
  wire  exceptionGen_io_wb_2_bits_trigger_backendHit_5; // @[Rob.scala 480:28]
  wire  exceptionGen_io_wb_3_valid; // @[Rob.scala 480:28]
  wire  exceptionGen_io_wb_3_bits_robIdx_flag; // @[Rob.scala 480:28]
  wire [4:0] exceptionGen_io_wb_3_bits_robIdx_value; // @[Rob.scala 480:28]
  wire  exceptionGen_io_wb_3_bits_exceptionVec_4; // @[Rob.scala 480:28]
  wire  exceptionGen_io_wb_3_bits_exceptionVec_5; // @[Rob.scala 480:28]
  wire  exceptionGen_io_wb_3_bits_exceptionVec_6; // @[Rob.scala 480:28]
  wire  exceptionGen_io_wb_3_bits_exceptionVec_7; // @[Rob.scala 480:28]
  wire  exceptionGen_io_wb_3_bits_exceptionVec_13; // @[Rob.scala 480:28]
  wire  exceptionGen_io_wb_3_bits_exceptionVec_15; // @[Rob.scala 480:28]
  wire  exceptionGen_io_wb_3_bits_trigger_backendHit_0; // @[Rob.scala 480:28]
  wire  exceptionGen_io_wb_3_bits_trigger_backendHit_1; // @[Rob.scala 480:28]
  wire  exceptionGen_io_wb_3_bits_trigger_backendHit_2; // @[Rob.scala 480:28]
  wire  exceptionGen_io_wb_3_bits_trigger_backendHit_3; // @[Rob.scala 480:28]
  wire  exceptionGen_io_wb_3_bits_trigger_backendHit_4; // @[Rob.scala 480:28]
  wire  exceptionGen_io_wb_3_bits_trigger_backendHit_5; // @[Rob.scala 480:28]
  wire  exceptionGen_io_wb_4_valid; // @[Rob.scala 480:28]
  wire  exceptionGen_io_wb_4_bits_robIdx_flag; // @[Rob.scala 480:28]
  wire [4:0] exceptionGen_io_wb_4_bits_robIdx_value; // @[Rob.scala 480:28]
  wire  exceptionGen_io_wb_4_bits_exceptionVec_6; // @[Rob.scala 480:28]
  wire  exceptionGen_io_wb_4_bits_exceptionVec_7; // @[Rob.scala 480:28]
  wire  exceptionGen_io_wb_4_bits_exceptionVec_15; // @[Rob.scala 480:28]
  wire  exceptionGen_io_wb_4_bits_trigger_backendHit_0; // @[Rob.scala 480:28]
  wire  exceptionGen_io_wb_4_bits_trigger_backendHit_1; // @[Rob.scala 480:28]
  wire  exceptionGen_io_wb_4_bits_trigger_backendHit_4; // @[Rob.scala 480:28]
  wire  exceptionGen_io_out_valid; // @[Rob.scala 480:28]
  wire [4:0] exceptionGen_io_out_bits_robIdx_value; // @[Rob.scala 480:28]
  wire  exceptionGen_io_state_valid; // @[Rob.scala 480:28]
  wire  exceptionGen_io_state_bits_robIdx_flag; // @[Rob.scala 480:28]
  wire [4:0] exceptionGen_io_state_bits_robIdx_value; // @[Rob.scala 480:28]
  wire  exceptionGen_io_state_bits_exceptionVec_0; // @[Rob.scala 480:28]
  wire  exceptionGen_io_state_bits_exceptionVec_1; // @[Rob.scala 480:28]
  wire  exceptionGen_io_state_bits_exceptionVec_2; // @[Rob.scala 480:28]
  wire  exceptionGen_io_state_bits_exceptionVec_3; // @[Rob.scala 480:28]
  wire  exceptionGen_io_state_bits_exceptionVec_4; // @[Rob.scala 480:28]
  wire  exceptionGen_io_state_bits_exceptionVec_5; // @[Rob.scala 480:28]
  wire  exceptionGen_io_state_bits_exceptionVec_6; // @[Rob.scala 480:28]
  wire  exceptionGen_io_state_bits_exceptionVec_7; // @[Rob.scala 480:28]
  wire  exceptionGen_io_state_bits_exceptionVec_8; // @[Rob.scala 480:28]
  wire  exceptionGen_io_state_bits_exceptionVec_9; // @[Rob.scala 480:28]
  wire  exceptionGen_io_state_bits_exceptionVec_10; // @[Rob.scala 480:28]
  wire  exceptionGen_io_state_bits_exceptionVec_11; // @[Rob.scala 480:28]
  wire  exceptionGen_io_state_bits_exceptionVec_12; // @[Rob.scala 480:28]
  wire  exceptionGen_io_state_bits_exceptionVec_13; // @[Rob.scala 480:28]
  wire  exceptionGen_io_state_bits_exceptionVec_14; // @[Rob.scala 480:28]
  wire  exceptionGen_io_state_bits_exceptionVec_15; // @[Rob.scala 480:28]
  wire  exceptionGen_io_state_bits_flushPipe; // @[Rob.scala 480:28]
  wire  exceptionGen_io_state_bits_replayInst; // @[Rob.scala 480:28]
  wire  exceptionGen_io_state_bits_singleStep; // @[Rob.scala 480:28]
  wire  exceptionGen_io_state_bits_crossPageIPFFix; // @[Rob.scala 480:28]
  wire  exceptionGen_io_state_bits_trigger_frontendHit_0; // @[Rob.scala 480:28]
  wire  exceptionGen_io_state_bits_trigger_frontendHit_1; // @[Rob.scala 480:28]
  wire  exceptionGen_io_state_bits_trigger_frontendHit_2; // @[Rob.scala 480:28]
  wire  exceptionGen_io_state_bits_trigger_frontendHit_3; // @[Rob.scala 480:28]
  wire  exceptionGen_io_state_bits_trigger_backendHit_0; // @[Rob.scala 480:28]
  wire  exceptionGen_io_state_bits_trigger_backendHit_1; // @[Rob.scala 480:28]
  wire  exceptionGen_io_state_bits_trigger_backendHit_2; // @[Rob.scala 480:28]
  wire  exceptionGen_io_state_bits_trigger_backendHit_3; // @[Rob.scala 480:28]
  wire  exceptionGen_io_state_bits_trigger_backendHit_4; // @[Rob.scala 480:28]
  wire  exceptionGen_io_state_bits_trigger_backendHit_5; // @[Rob.scala 480:28]
  wire  deqPtrGenModule_clock; // @[Rob.scala 774:31]
  wire  deqPtrGenModule_reset; // @[Rob.scala 774:31]
  wire [1:0] deqPtrGenModule_io_state; // @[Rob.scala 774:31]
  wire  deqPtrGenModule_io_deq_v_0; // @[Rob.scala 774:31]
  wire  deqPtrGenModule_io_deq_v_1; // @[Rob.scala 774:31]
  wire  deqPtrGenModule_io_deq_w0; // @[Rob.scala 774:31]
  wire  deqPtrGenModule_io_deq_w1; // @[Rob.scala 774:31]
  wire  deqPtrGenModule_io_exception_state_valid; // @[Rob.scala 774:31]
  wire  deqPtrGenModule_io_exception_state_bits_robIdx_flag; // @[Rob.scala 774:31]
  wire [4:0] deqPtrGenModule_io_exception_state_bits_robIdx_value; // @[Rob.scala 774:31]
  wire  deqPtrGenModule_io_exception_state_bits_exceptionVec_0; // @[Rob.scala 774:31]
  wire  deqPtrGenModule_io_exception_state_bits_exceptionVec_1; // @[Rob.scala 774:31]
  wire  deqPtrGenModule_io_exception_state_bits_exceptionVec_2; // @[Rob.scala 774:31]
  wire  deqPtrGenModule_io_exception_state_bits_exceptionVec_3; // @[Rob.scala 774:31]
  wire  deqPtrGenModule_io_exception_state_bits_exceptionVec_4; // @[Rob.scala 774:31]
  wire  deqPtrGenModule_io_exception_state_bits_exceptionVec_5; // @[Rob.scala 774:31]
  wire  deqPtrGenModule_io_exception_state_bits_exceptionVec_6; // @[Rob.scala 774:31]
  wire  deqPtrGenModule_io_exception_state_bits_exceptionVec_7; // @[Rob.scala 774:31]
  wire  deqPtrGenModule_io_exception_state_bits_exceptionVec_8; // @[Rob.scala 774:31]
  wire  deqPtrGenModule_io_exception_state_bits_exceptionVec_9; // @[Rob.scala 774:31]
  wire  deqPtrGenModule_io_exception_state_bits_exceptionVec_10; // @[Rob.scala 774:31]
  wire  deqPtrGenModule_io_exception_state_bits_exceptionVec_11; // @[Rob.scala 774:31]
  wire  deqPtrGenModule_io_exception_state_bits_exceptionVec_12; // @[Rob.scala 774:31]
  wire  deqPtrGenModule_io_exception_state_bits_exceptionVec_13; // @[Rob.scala 774:31]
  wire  deqPtrGenModule_io_exception_state_bits_exceptionVec_14; // @[Rob.scala 774:31]
  wire  deqPtrGenModule_io_exception_state_bits_exceptionVec_15; // @[Rob.scala 774:31]
  wire  deqPtrGenModule_io_exception_state_bits_replayInst; // @[Rob.scala 774:31]
  wire  deqPtrGenModule_io_exception_state_bits_singleStep; // @[Rob.scala 774:31]
  wire  deqPtrGenModule_io_exception_state_bits_trigger_frontendHit_0; // @[Rob.scala 774:31]
  wire  deqPtrGenModule_io_exception_state_bits_trigger_frontendHit_1; // @[Rob.scala 774:31]
  wire  deqPtrGenModule_io_exception_state_bits_trigger_frontendHit_2; // @[Rob.scala 774:31]
  wire  deqPtrGenModule_io_exception_state_bits_trigger_frontendHit_3; // @[Rob.scala 774:31]
  wire  deqPtrGenModule_io_exception_state_bits_trigger_backendHit_0; // @[Rob.scala 774:31]
  wire  deqPtrGenModule_io_exception_state_bits_trigger_backendHit_1; // @[Rob.scala 774:31]
  wire  deqPtrGenModule_io_exception_state_bits_trigger_backendHit_2; // @[Rob.scala 774:31]
  wire  deqPtrGenModule_io_exception_state_bits_trigger_backendHit_3; // @[Rob.scala 774:31]
  wire  deqPtrGenModule_io_exception_state_bits_trigger_backendHit_4; // @[Rob.scala 774:31]
  wire  deqPtrGenModule_io_exception_state_bits_trigger_backendHit_5; // @[Rob.scala 774:31]
  wire  deqPtrGenModule_io_intrBitSetReg; // @[Rob.scala 774:31]
  wire  deqPtrGenModule_io_hasNoSpecExec; // @[Rob.scala 774:31]
  wire  deqPtrGenModule_io_interrupt_safe; // @[Rob.scala 774:31]
  wire  deqPtrGenModule_io_blockCommit; // @[Rob.scala 774:31]
  wire  deqPtrGenModule_io_out_0_flag; // @[Rob.scala 774:31]
  wire [4:0] deqPtrGenModule_io_out_0_value; // @[Rob.scala 774:31]
  wire  deqPtrGenModule_io_out_1_flag; // @[Rob.scala 774:31]
  wire [4:0] deqPtrGenModule_io_out_1_value; // @[Rob.scala 774:31]
  wire  deqPtrGenModule_io_next_out_0_flag; // @[Rob.scala 774:31]
  wire [4:0] deqPtrGenModule_io_next_out_0_value; // @[Rob.scala 774:31]
  wire  deqPtrGenModule_io_next_out_1_flag; // @[Rob.scala 774:31]
  wire [4:0] deqPtrGenModule_io_next_out_1_value; // @[Rob.scala 774:31]
  wire  enqPtrGenModule_clock; // @[Rob.scala 786:31]
  wire  enqPtrGenModule_reset; // @[Rob.scala 786:31]
  wire  enqPtrGenModule_io_redirect_valid; // @[Rob.scala 786:31]
  wire  enqPtrGenModule_io_redirect_bits_robIdx_flag; // @[Rob.scala 786:31]
  wire [4:0] enqPtrGenModule_io_redirect_bits_robIdx_value; // @[Rob.scala 786:31]
  wire  enqPtrGenModule_io_redirect_bits_level; // @[Rob.scala 786:31]
  wire  enqPtrGenModule_io_allowEnqueue; // @[Rob.scala 786:31]
  wire  enqPtrGenModule_io_hasBlockBackward; // @[Rob.scala 786:31]
  wire  enqPtrGenModule_io_enq_0; // @[Rob.scala 786:31]
  wire  enqPtrGenModule_io_enq_1; // @[Rob.scala 786:31]
  wire  enqPtrGenModule_io_out_0_flag; // @[Rob.scala 786:31]
  wire [4:0] enqPtrGenModule_io_out_0_value; // @[Rob.scala 786:31]
  wire [4:0] enqPtrGenModule_io_out_1_value; // @[Rob.scala 786:31]
  wire  fflagsDataModule_clock; // @[Rob.scala 1007:32]
  wire [4:0] fflagsDataModule_io_raddr_0; // @[Rob.scala 1007:32]
  wire [4:0] fflagsDataModule_io_raddr_1; // @[Rob.scala 1007:32]
  wire [4:0] fflagsDataModule_io_rdata_0; // @[Rob.scala 1007:32]
  wire [4:0] fflagsDataModule_io_rdata_1; // @[Rob.scala 1007:32]
  wire  fflagsDataModule_io_wen_0; // @[Rob.scala 1007:32]
  wire  fflagsDataModule_io_wen_1; // @[Rob.scala 1007:32]
  wire  fflagsDataModule_io_wen_2; // @[Rob.scala 1007:32]
  wire [4:0] fflagsDataModule_io_waddr_0; // @[Rob.scala 1007:32]
  wire [4:0] fflagsDataModule_io_waddr_1; // @[Rob.scala 1007:32]
  wire [4:0] fflagsDataModule_io_waddr_2; // @[Rob.scala 1007:32]
  wire [4:0] fflagsDataModule_io_wdata_0; // @[Rob.scala 1007:32]
  wire [4:0] fflagsDataModule_io_wdata_1; // @[Rob.scala 1007:32]
  wire [4:0] fflagsDataModule_io_wdata_2; // @[Rob.scala 1007:32]
  reg  dt_eliminatedMove [0:31]; // @[Rob.scala 1212:32]
  wire  dt_eliminatedMove_eliminatedMove_en; // @[Rob.scala 1212:32]
  wire [4:0] dt_eliminatedMove_eliminatedMove_addr; // @[Rob.scala 1212:32]
  wire  dt_eliminatedMove_eliminatedMove_data; // @[Rob.scala 1212:32]
  wire  dt_eliminatedMove_eliminatedMove_1_en; // @[Rob.scala 1212:32]
  wire [4:0] dt_eliminatedMove_eliminatedMove_1_addr; // @[Rob.scala 1212:32]
  wire  dt_eliminatedMove_eliminatedMove_1_data; // @[Rob.scala 1212:32]
  wire  dt_eliminatedMove_MPORT_305_data; // @[Rob.scala 1212:32]
  wire [4:0] dt_eliminatedMove_MPORT_305_addr; // @[Rob.scala 1212:32]
  wire  dt_eliminatedMove_MPORT_305_mask; // @[Rob.scala 1212:32]
  wire  dt_eliminatedMove_MPORT_305_en; // @[Rob.scala 1212:32]
  wire  dt_eliminatedMove_MPORT_307_data; // @[Rob.scala 1212:32]
  wire [4:0] dt_eliminatedMove_MPORT_307_addr; // @[Rob.scala 1212:32]
  wire  dt_eliminatedMove_MPORT_307_mask; // @[Rob.scala 1212:32]
  wire  dt_eliminatedMove_MPORT_307_en; // @[Rob.scala 1212:32]
  reg  dt_isRVC [0:31]; // @[Rob.scala 1213:23]
  wire  dt_isRVC_isRVC_en; // @[Rob.scala 1213:23]
  wire [4:0] dt_isRVC_isRVC_addr; // @[Rob.scala 1213:23]
  wire  dt_isRVC_isRVC_data; // @[Rob.scala 1213:23]
  wire  dt_isRVC_isRVC_1_en; // @[Rob.scala 1213:23]
  wire [4:0] dt_isRVC_isRVC_1_addr; // @[Rob.scala 1213:23]
  wire  dt_isRVC_isRVC_1_data; // @[Rob.scala 1213:23]
  wire  dt_isRVC_MPORT_306_data; // @[Rob.scala 1213:23]
  wire [4:0] dt_isRVC_MPORT_306_addr; // @[Rob.scala 1213:23]
  wire  dt_isRVC_MPORT_306_mask; // @[Rob.scala 1213:23]
  wire  dt_isRVC_MPORT_306_en; // @[Rob.scala 1213:23]
  wire  dt_isRVC_MPORT_308_data; // @[Rob.scala 1213:23]
  wire [4:0] dt_isRVC_MPORT_308_addr; // @[Rob.scala 1213:23]
  wire  dt_isRVC_MPORT_308_mask; // @[Rob.scala 1213:23]
  wire  dt_isRVC_MPORT_308_en; // @[Rob.scala 1213:23]
  wire  difftest_io_clock; // @[Rob.scala 1235:28]
  wire [7:0] difftest_io_coreid; // @[Rob.scala 1235:28]
  wire [7:0] difftest_io_index; // @[Rob.scala 1235:28]
  wire  difftest_io_valid; // @[Rob.scala 1235:28]
  wire [7:0] difftest_io_special; // @[Rob.scala 1235:28]
  wire  difftest_io_skip; // @[Rob.scala 1235:28]
  wire  difftest_io_isRVC; // @[Rob.scala 1235:28]
  wire  difftest_io_rfwen; // @[Rob.scala 1235:28]
  wire  difftest_io_fpwen; // @[Rob.scala 1235:28]
  wire [31:0] difftest_io_wpdest; // @[Rob.scala 1235:28]
  wire [7:0] difftest_io_wdest; // @[Rob.scala 1235:28]
  wire  difftest_1_io_clock; // @[Rob.scala 1235:28]
  wire [7:0] difftest_1_io_coreid; // @[Rob.scala 1235:28]
  wire [7:0] difftest_1_io_index; // @[Rob.scala 1235:28]
  wire  difftest_1_io_valid; // @[Rob.scala 1235:28]
  wire [7:0] difftest_1_io_special; // @[Rob.scala 1235:28]
  wire  difftest_1_io_skip; // @[Rob.scala 1235:28]
  wire  difftest_1_io_isRVC; // @[Rob.scala 1235:28]
  wire  difftest_1_io_rfwen; // @[Rob.scala 1235:28]
  wire  difftest_1_io_fpwen; // @[Rob.scala 1235:28]
  wire [31:0] difftest_1_io_wpdest; // @[Rob.scala 1235:28]
  wire [7:0] difftest_1_io_wdest; // @[Rob.scala 1235:28]
  reg  dt_isXSTrap [0:31]; // @[Rob.scala 1290:26]
  wire  dt_isXSTrap_trapVec_MPORT_en; // @[Rob.scala 1290:26]
  wire [4:0] dt_isXSTrap_trapVec_MPORT_addr; // @[Rob.scala 1290:26]
  wire  dt_isXSTrap_trapVec_MPORT_data; // @[Rob.scala 1290:26]
  wire  dt_isXSTrap_trapVec_MPORT_1_en; // @[Rob.scala 1290:26]
  wire [4:0] dt_isXSTrap_trapVec_MPORT_1_addr; // @[Rob.scala 1290:26]
  wire  dt_isXSTrap_trapVec_MPORT_1_data; // @[Rob.scala 1290:26]
  wire  dt_isXSTrap_MPORT_309_data; // @[Rob.scala 1290:26]
  wire [4:0] dt_isXSTrap_MPORT_309_addr; // @[Rob.scala 1290:26]
  wire  dt_isXSTrap_MPORT_309_mask; // @[Rob.scala 1290:26]
  wire  dt_isXSTrap_MPORT_309_en; // @[Rob.scala 1290:26]
  wire  dt_isXSTrap_MPORT_310_data; // @[Rob.scala 1290:26]
  wire [4:0] dt_isXSTrap_MPORT_310_addr; // @[Rob.scala 1290:26]
  wire  dt_isXSTrap_MPORT_310_mask; // @[Rob.scala 1290:26]
  wire  dt_isXSTrap_MPORT_310_en; // @[Rob.scala 1290:26]
  wire  difftest_2_io_clock; // @[Rob.scala 1298:26]
  wire [7:0] difftest_2_io_coreid; // @[Rob.scala 1298:26]
  wire  difftest_2_io_valid; // @[Rob.scala 1298:26]
  wire [63:0] difftest_2_io_cycleCnt; // @[Rob.scala 1298:26]
  wire [63:0] difftest_2_io_instrCnt; // @[Rob.scala 1298:26]
  wire  difftest_2_io_hasWFI; // @[Rob.scala 1298:26]
  reg  valid_0; // @[Rob.scala 426:22]
  reg  valid_1; // @[Rob.scala 426:22]
  reg  valid_2; // @[Rob.scala 426:22]
  reg  valid_3; // @[Rob.scala 426:22]
  reg  valid_4; // @[Rob.scala 426:22]
  reg  valid_5; // @[Rob.scala 426:22]
  reg  valid_6; // @[Rob.scala 426:22]
  reg  valid_7; // @[Rob.scala 426:22]
  reg  valid_8; // @[Rob.scala 426:22]
  reg  valid_9; // @[Rob.scala 426:22]
  reg  valid_10; // @[Rob.scala 426:22]
  reg  valid_11; // @[Rob.scala 426:22]
  reg  valid_12; // @[Rob.scala 426:22]
  reg  valid_13; // @[Rob.scala 426:22]
  reg  valid_14; // @[Rob.scala 426:22]
  reg  valid_15; // @[Rob.scala 426:22]
  reg  valid_16; // @[Rob.scala 426:22]
  reg  valid_17; // @[Rob.scala 426:22]
  reg  valid_18; // @[Rob.scala 426:22]
  reg  valid_19; // @[Rob.scala 426:22]
  reg  valid_20; // @[Rob.scala 426:22]
  reg  valid_21; // @[Rob.scala 426:22]
  reg  valid_22; // @[Rob.scala 426:22]
  reg  valid_23; // @[Rob.scala 426:22]
  reg  valid_24; // @[Rob.scala 426:22]
  reg  valid_25; // @[Rob.scala 426:22]
  reg  valid_26; // @[Rob.scala 426:22]
  reg  valid_27; // @[Rob.scala 426:22]
  reg  valid_28; // @[Rob.scala 426:22]
  reg  valid_29; // @[Rob.scala 426:22]
  reg  valid_30; // @[Rob.scala 426:22]
  reg  valid_31; // @[Rob.scala 426:22]
  reg  mmio_0; // @[Rob.scala 431:21]
  reg  mmio_1; // @[Rob.scala 431:21]
  reg  mmio_2; // @[Rob.scala 431:21]
  reg  mmio_3; // @[Rob.scala 431:21]
  reg  mmio_4; // @[Rob.scala 431:21]
  reg  mmio_5; // @[Rob.scala 431:21]
  reg  mmio_6; // @[Rob.scala 431:21]
  reg  mmio_7; // @[Rob.scala 431:21]
  reg  mmio_8; // @[Rob.scala 431:21]
  reg  mmio_9; // @[Rob.scala 431:21]
  reg  mmio_10; // @[Rob.scala 431:21]
  reg  mmio_11; // @[Rob.scala 431:21]
  reg  mmio_12; // @[Rob.scala 431:21]
  reg  mmio_13; // @[Rob.scala 431:21]
  reg  mmio_14; // @[Rob.scala 431:21]
  reg  mmio_15; // @[Rob.scala 431:21]
  reg  mmio_16; // @[Rob.scala 431:21]
  reg  mmio_17; // @[Rob.scala 431:21]
  reg  mmio_18; // @[Rob.scala 431:21]
  reg  mmio_19; // @[Rob.scala 431:21]
  reg  mmio_20; // @[Rob.scala 431:21]
  reg  mmio_21; // @[Rob.scala 431:21]
  reg  mmio_22; // @[Rob.scala 431:21]
  reg  mmio_23; // @[Rob.scala 431:21]
  reg  mmio_24; // @[Rob.scala 431:21]
  reg  mmio_25; // @[Rob.scala 431:21]
  reg  mmio_26; // @[Rob.scala 431:21]
  reg  mmio_27; // @[Rob.scala 431:21]
  reg  mmio_28; // @[Rob.scala 431:21]
  reg  mmio_29; // @[Rob.scala 431:21]
  reg  mmio_30; // @[Rob.scala 431:21]
  reg  mmio_31; // @[Rob.scala 431:21]
  reg  walkPtrVec_0_flag; // @[Rob.scala 450:23]
  reg [4:0] walkPtrVec_0_value; // @[Rob.scala 450:23]
  reg  walkPtrVec_1_flag; // @[Rob.scala 450:23]
  reg [4:0] walkPtrVec_1_value; // @[Rob.scala 450:23]
  reg  allowEnqueue; // @[Rob.scala 451:29]
  wire  enqPtrVec_0_flag = enqPtrGenModule_io_out_0_flag; // @[Rob.scala 447:23 791:13]
  wire [4:0] enqPtrVec_0_value = enqPtrGenModule_io_out_0_value; // @[Rob.scala 447:23 791:13]
  wire [5:0] _isEmpty_T = {enqPtrVec_0_flag,enqPtrVec_0_value}; // @[CircularQueuePtr.scala 61:50]
  wire  deqPtrVec_0_flag = deqPtrGenModule_io_out_0_flag; // @[Rob.scala 448:23 783:13]
  wire [4:0] deqPtrVec_0_value = deqPtrGenModule_io_out_0_value; // @[Rob.scala 448:23 783:13]
  wire [5:0] _isEmpty_T_1 = {deqPtrVec_0_flag,deqPtrVec_0_value}; // @[CircularQueuePtr.scala 61:70]
  wire  isEmpty = _isEmpty_T == _isEmpty_T_1; // @[CircularQueuePtr.scala 61:52]
  wire  isReplaying = io_redirect_valid & io_redirect_bits_level; // @[Rob.scala 458:39]
  reg  state; // @[Rob.scala 464:22]
  reg  hasBlockBackward; // @[Rob.scala 490:33]
  reg  hasNoSpecExec; // @[Rob.scala 491:30]
  wire  _GEN_0 = isEmpty ? 1'h0 : hasBlockBackward; // @[Rob.scala 495:18 490:33 495:36]
  wire [1:0] _T = {io_commits_walkValid_1,io_commits_walkValid_0}; // @[Bundle.scala 390:48]
  wire  _T_2 = io_commits_isWalk & |_T; // @[Bundle.scala 390:35]
  wire [1:0] _T_3 = {io_commits_commitValid_1,io_commits_commitValid_0}; // @[Bundle.scala 391:54]
  wire  _T_5 = io_commits_isCommit & |_T_3; // @[Bundle.scala 391:39]
  wire  _GEN_1 = _T_2 | _T_5 ? 1'h0 : hasNoSpecExec; // @[Rob.scala 491:30 497:{63,78}]
  reg  hasWFI; // @[Rob.scala 502:23]
  reg [19:0] wfi_cycles; // @[Rob.scala 505:27]
  wire [19:0] _wfi_cycles_T_1 = wfi_cycles + 20'h1; // @[Rob.scala 507:30]
  reg  REG; // @[Rob.scala 508:33]
  wire  wfi_timeout = &wfi_cycles; // @[Rob.scala 511:32]
  reg  REG_1; // @[Rob.scala 512:24]
  reg  REG_2; // @[Rob.scala 512:16]
  wire  _GEN_4 = REG_2 | io_flushOut_valid | wfi_timeout ? 1'h0 : hasWFI; // @[Rob.scala 512:80 513:12 502:23]
  wire [4:0] enqPtrVec_1_value = enqPtrGenModule_io_out_1_value; // @[Rob.scala 447:23 791:13]
  wire [4:0] allocatePtrVec_1_value = io_enq_needAlloc_0 ? enqPtrVec_1_value : enqPtrVec_0_value; // @[Rob.scala 516:{31,31}]
  wire  canEnqueue_0 = io_enq_req_0_valid & io_enq_canAccept; // @[Rob.scala 519:51]
  wire  canEnqueue_1 = io_enq_req_1_valid & io_enq_canAccept; // @[Rob.scala 519:51]
  reg [63:0] timer; // @[GTimer.scala 23:20]
  wire  _GEN_329 = io_enq_req_0_bits_ctrl_blockBackward | _GEN_0; // @[Rob.scala 536:40 537:26]
  wire  _GEN_330 = io_enq_req_0_bits_ctrl_noSpecExec | _GEN_1; // @[Rob.scala 539:37 540:23]
  wire  enqHasTriggerHit = io_enq_req_0_bits_cf_trigger_frontendHit_0 | io_enq_req_0_bits_cf_trigger_frontendHit_1 |
    io_enq_req_0_bits_cf_trigger_frontendHit_2 | io_enq_req_0_bits_cf_trigger_frontendHit_3; // @[Bundle.scala 628:45]
  wire [15:0] _enqHasException_T = {2'h0,1'h0,io_enq_req_0_bits_cf_exceptionVec_12,4'h0,4'h0,1'h0,
    io_enq_req_0_bits_cf_exceptionVec_2,io_enq_req_0_bits_cf_exceptionVec_1,1'h0}; // @[Rob.scala 543:80]
  wire  enqHasException = |_enqHasException_T; // @[Rob.scala 543:87]
  wire  _T_11 = ~enqHasTriggerHit; // @[Rob.scala 545:12]
  wire  _T_12 = ~enqHasException; // @[Rob.scala 545:33]
  wire  _T_45 = io_enq_req_0_bits_ctrl_fuType == 4'h2 & io_enq_req_0_bits_ctrl_fuOpType == 7'h4; // @[Bundle.scala 192:43]
  wire  _GEN_333 = _T_45 & _T_12 & _T_11 | _GEN_4; // @[Rob.scala 557:73 558:16]
  wire  _GEN_334 = 5'h0 == enqPtrVec_0_value ? 1'h0 : mmio_0; // @[Rob.scala 431:21 562:{22,22}]
  wire  _GEN_335 = 5'h1 == enqPtrVec_0_value ? 1'h0 : mmio_1; // @[Rob.scala 431:21 562:{22,22}]
  wire  _GEN_336 = 5'h2 == enqPtrVec_0_value ? 1'h0 : mmio_2; // @[Rob.scala 431:21 562:{22,22}]
  wire  _GEN_337 = 5'h3 == enqPtrVec_0_value ? 1'h0 : mmio_3; // @[Rob.scala 431:21 562:{22,22}]
  wire  _GEN_338 = 5'h4 == enqPtrVec_0_value ? 1'h0 : mmio_4; // @[Rob.scala 431:21 562:{22,22}]
  wire  _GEN_339 = 5'h5 == enqPtrVec_0_value ? 1'h0 : mmio_5; // @[Rob.scala 431:21 562:{22,22}]
  wire  _GEN_340 = 5'h6 == enqPtrVec_0_value ? 1'h0 : mmio_6; // @[Rob.scala 431:21 562:{22,22}]
  wire  _GEN_341 = 5'h7 == enqPtrVec_0_value ? 1'h0 : mmio_7; // @[Rob.scala 431:21 562:{22,22}]
  wire  _GEN_342 = 5'h8 == enqPtrVec_0_value ? 1'h0 : mmio_8; // @[Rob.scala 431:21 562:{22,22}]
  wire  _GEN_343 = 5'h9 == enqPtrVec_0_value ? 1'h0 : mmio_9; // @[Rob.scala 431:21 562:{22,22}]
  wire  _GEN_344 = 5'ha == enqPtrVec_0_value ? 1'h0 : mmio_10; // @[Rob.scala 431:21 562:{22,22}]
  wire  _GEN_345 = 5'hb == enqPtrVec_0_value ? 1'h0 : mmio_11; // @[Rob.scala 431:21 562:{22,22}]
  wire  _GEN_346 = 5'hc == enqPtrVec_0_value ? 1'h0 : mmio_12; // @[Rob.scala 431:21 562:{22,22}]
  wire  _GEN_347 = 5'hd == enqPtrVec_0_value ? 1'h0 : mmio_13; // @[Rob.scala 431:21 562:{22,22}]
  wire  _GEN_348 = 5'he == enqPtrVec_0_value ? 1'h0 : mmio_14; // @[Rob.scala 431:21 562:{22,22}]
  wire  _GEN_349 = 5'hf == enqPtrVec_0_value ? 1'h0 : mmio_15; // @[Rob.scala 431:21 562:{22,22}]
  wire  _GEN_350 = 5'h10 == enqPtrVec_0_value ? 1'h0 : mmio_16; // @[Rob.scala 431:21 562:{22,22}]
  wire  _GEN_351 = 5'h11 == enqPtrVec_0_value ? 1'h0 : mmio_17; // @[Rob.scala 431:21 562:{22,22}]
  wire  _GEN_352 = 5'h12 == enqPtrVec_0_value ? 1'h0 : mmio_18; // @[Rob.scala 431:21 562:{22,22}]
  wire  _GEN_353 = 5'h13 == enqPtrVec_0_value ? 1'h0 : mmio_19; // @[Rob.scala 431:21 562:{22,22}]
  wire  _GEN_354 = 5'h14 == enqPtrVec_0_value ? 1'h0 : mmio_20; // @[Rob.scala 431:21 562:{22,22}]
  wire  _GEN_355 = 5'h15 == enqPtrVec_0_value ? 1'h0 : mmio_21; // @[Rob.scala 431:21 562:{22,22}]
  wire  _GEN_356 = 5'h16 == enqPtrVec_0_value ? 1'h0 : mmio_22; // @[Rob.scala 431:21 562:{22,22}]
  wire  _GEN_357 = 5'h17 == enqPtrVec_0_value ? 1'h0 : mmio_23; // @[Rob.scala 431:21 562:{22,22}]
  wire  _GEN_358 = 5'h18 == enqPtrVec_0_value ? 1'h0 : mmio_24; // @[Rob.scala 431:21 562:{22,22}]
  wire  _GEN_359 = 5'h19 == enqPtrVec_0_value ? 1'h0 : mmio_25; // @[Rob.scala 431:21 562:{22,22}]
  wire  _GEN_360 = 5'h1a == enqPtrVec_0_value ? 1'h0 : mmio_26; // @[Rob.scala 431:21 562:{22,22}]
  wire  _GEN_361 = 5'h1b == enqPtrVec_0_value ? 1'h0 : mmio_27; // @[Rob.scala 431:21 562:{22,22}]
  wire  _GEN_362 = 5'h1c == enqPtrVec_0_value ? 1'h0 : mmio_28; // @[Rob.scala 431:21 562:{22,22}]
  wire  _GEN_363 = 5'h1d == enqPtrVec_0_value ? 1'h0 : mmio_29; // @[Rob.scala 431:21 562:{22,22}]
  wire  _GEN_364 = 5'h1e == enqPtrVec_0_value ? 1'h0 : mmio_30; // @[Rob.scala 431:21 562:{22,22}]
  wire  _GEN_365 = 5'h1f == enqPtrVec_0_value ? 1'h0 : mmio_31; // @[Rob.scala 431:21 562:{22,22}]
  wire  _GEN_800 = canEnqueue_0 ? _GEN_329 : _GEN_0; // @[Rob.scala 523:26]
  wire  _GEN_801 = canEnqueue_0 ? _GEN_330 : _GEN_1; // @[Rob.scala 523:26]
  wire  _GEN_803 = canEnqueue_0 ? _GEN_333 : _GEN_4; // @[Rob.scala 523:26]
  wire  _GEN_804 = canEnqueue_0 ? _GEN_334 : mmio_0; // @[Rob.scala 431:21 523:26]
  wire  _GEN_805 = canEnqueue_0 ? _GEN_335 : mmio_1; // @[Rob.scala 431:21 523:26]
  wire  _GEN_806 = canEnqueue_0 ? _GEN_336 : mmio_2; // @[Rob.scala 431:21 523:26]
  wire  _GEN_807 = canEnqueue_0 ? _GEN_337 : mmio_3; // @[Rob.scala 431:21 523:26]
  wire  _GEN_808 = canEnqueue_0 ? _GEN_338 : mmio_4; // @[Rob.scala 431:21 523:26]
  wire  _GEN_809 = canEnqueue_0 ? _GEN_339 : mmio_5; // @[Rob.scala 431:21 523:26]
  wire  _GEN_810 = canEnqueue_0 ? _GEN_340 : mmio_6; // @[Rob.scala 431:21 523:26]
  wire  _GEN_811 = canEnqueue_0 ? _GEN_341 : mmio_7; // @[Rob.scala 431:21 523:26]
  wire  _GEN_812 = canEnqueue_0 ? _GEN_342 : mmio_8; // @[Rob.scala 431:21 523:26]
  wire  _GEN_813 = canEnqueue_0 ? _GEN_343 : mmio_9; // @[Rob.scala 431:21 523:26]
  wire  _GEN_814 = canEnqueue_0 ? _GEN_344 : mmio_10; // @[Rob.scala 431:21 523:26]
  wire  _GEN_815 = canEnqueue_0 ? _GEN_345 : mmio_11; // @[Rob.scala 431:21 523:26]
  wire  _GEN_816 = canEnqueue_0 ? _GEN_346 : mmio_12; // @[Rob.scala 431:21 523:26]
  wire  _GEN_817 = canEnqueue_0 ? _GEN_347 : mmio_13; // @[Rob.scala 431:21 523:26]
  wire  _GEN_818 = canEnqueue_0 ? _GEN_348 : mmio_14; // @[Rob.scala 431:21 523:26]
  wire  _GEN_819 = canEnqueue_0 ? _GEN_349 : mmio_15; // @[Rob.scala 431:21 523:26]
  wire  _GEN_820 = canEnqueue_0 ? _GEN_350 : mmio_16; // @[Rob.scala 431:21 523:26]
  wire  _GEN_821 = canEnqueue_0 ? _GEN_351 : mmio_17; // @[Rob.scala 431:21 523:26]
  wire  _GEN_822 = canEnqueue_0 ? _GEN_352 : mmio_18; // @[Rob.scala 431:21 523:26]
  wire  _GEN_823 = canEnqueue_0 ? _GEN_353 : mmio_19; // @[Rob.scala 431:21 523:26]
  wire  _GEN_824 = canEnqueue_0 ? _GEN_354 : mmio_20; // @[Rob.scala 431:21 523:26]
  wire  _GEN_825 = canEnqueue_0 ? _GEN_355 : mmio_21; // @[Rob.scala 431:21 523:26]
  wire  _GEN_826 = canEnqueue_0 ? _GEN_356 : mmio_22; // @[Rob.scala 431:21 523:26]
  wire  _GEN_827 = canEnqueue_0 ? _GEN_357 : mmio_23; // @[Rob.scala 431:21 523:26]
  wire  _GEN_828 = canEnqueue_0 ? _GEN_358 : mmio_24; // @[Rob.scala 431:21 523:26]
  wire  _GEN_829 = canEnqueue_0 ? _GEN_359 : mmio_25; // @[Rob.scala 431:21 523:26]
  wire  _GEN_830 = canEnqueue_0 ? _GEN_360 : mmio_26; // @[Rob.scala 431:21 523:26]
  wire  _GEN_831 = canEnqueue_0 ? _GEN_361 : mmio_27; // @[Rob.scala 431:21 523:26]
  wire  _GEN_832 = canEnqueue_0 ? _GEN_362 : mmio_28; // @[Rob.scala 431:21 523:26]
  wire  _GEN_833 = canEnqueue_0 ? _GEN_363 : mmio_29; // @[Rob.scala 431:21 523:26]
  wire  _GEN_834 = canEnqueue_0 ? _GEN_364 : mmio_30; // @[Rob.scala 431:21 523:26]
  wire  _GEN_835 = canEnqueue_0 ? _GEN_365 : mmio_31; // @[Rob.scala 431:21 523:26]
  wire  _GEN_1156 = io_enq_req_1_bits_ctrl_blockBackward | _GEN_800; // @[Rob.scala 536:40 537:26]
  wire  _GEN_1157 = io_enq_req_1_bits_ctrl_noSpecExec | _GEN_801; // @[Rob.scala 539:37 540:23]
  wire  enqHasTriggerHit_1 = io_enq_req_1_bits_cf_trigger_frontendHit_0 | io_enq_req_1_bits_cf_trigger_frontendHit_1 |
    io_enq_req_1_bits_cf_trigger_frontendHit_2 | io_enq_req_1_bits_cf_trigger_frontendHit_3; // @[Bundle.scala 628:45]
  wire [15:0] _enqHasException_T_1 = {2'h0,1'h0,io_enq_req_1_bits_cf_exceptionVec_12,4'h0,4'h0,1'h0,
    io_enq_req_1_bits_cf_exceptionVec_2,io_enq_req_1_bits_cf_exceptionVec_1,1'h0}; // @[Rob.scala 543:80]
  wire  enqHasException_1 = |_enqHasException_T_1; // @[Rob.scala 543:87]
  wire  _T_50 = ~enqHasTriggerHit_1; // @[Rob.scala 545:12]
  wire  _T_51 = ~enqHasException_1; // @[Rob.scala 545:33]
  wire  _T_84 = io_enq_req_1_bits_ctrl_fuType == 4'h2 & io_enq_req_1_bits_ctrl_fuOpType == 7'h4; // @[Bundle.scala 192:43]
  wire  _GEN_1160 = _T_84 & _T_51 & _T_50 | _GEN_803; // @[Rob.scala 557:73 558:16]
  wire  _GEN_1161 = 5'h0 == allocatePtrVec_1_value ? 1'h0 : _GEN_804; // @[Rob.scala 562:{22,22}]
  wire  _GEN_1162 = 5'h1 == allocatePtrVec_1_value ? 1'h0 : _GEN_805; // @[Rob.scala 562:{22,22}]
  wire  _GEN_1163 = 5'h2 == allocatePtrVec_1_value ? 1'h0 : _GEN_806; // @[Rob.scala 562:{22,22}]
  wire  _GEN_1164 = 5'h3 == allocatePtrVec_1_value ? 1'h0 : _GEN_807; // @[Rob.scala 562:{22,22}]
  wire  _GEN_1165 = 5'h4 == allocatePtrVec_1_value ? 1'h0 : _GEN_808; // @[Rob.scala 562:{22,22}]
  wire  _GEN_1166 = 5'h5 == allocatePtrVec_1_value ? 1'h0 : _GEN_809; // @[Rob.scala 562:{22,22}]
  wire  _GEN_1167 = 5'h6 == allocatePtrVec_1_value ? 1'h0 : _GEN_810; // @[Rob.scala 562:{22,22}]
  wire  _GEN_1168 = 5'h7 == allocatePtrVec_1_value ? 1'h0 : _GEN_811; // @[Rob.scala 562:{22,22}]
  wire  _GEN_1169 = 5'h8 == allocatePtrVec_1_value ? 1'h0 : _GEN_812; // @[Rob.scala 562:{22,22}]
  wire  _GEN_1170 = 5'h9 == allocatePtrVec_1_value ? 1'h0 : _GEN_813; // @[Rob.scala 562:{22,22}]
  wire  _GEN_1171 = 5'ha == allocatePtrVec_1_value ? 1'h0 : _GEN_814; // @[Rob.scala 562:{22,22}]
  wire  _GEN_1172 = 5'hb == allocatePtrVec_1_value ? 1'h0 : _GEN_815; // @[Rob.scala 562:{22,22}]
  wire  _GEN_1173 = 5'hc == allocatePtrVec_1_value ? 1'h0 : _GEN_816; // @[Rob.scala 562:{22,22}]
  wire  _GEN_1174 = 5'hd == allocatePtrVec_1_value ? 1'h0 : _GEN_817; // @[Rob.scala 562:{22,22}]
  wire  _GEN_1175 = 5'he == allocatePtrVec_1_value ? 1'h0 : _GEN_818; // @[Rob.scala 562:{22,22}]
  wire  _GEN_1176 = 5'hf == allocatePtrVec_1_value ? 1'h0 : _GEN_819; // @[Rob.scala 562:{22,22}]
  wire  _GEN_1177 = 5'h10 == allocatePtrVec_1_value ? 1'h0 : _GEN_820; // @[Rob.scala 562:{22,22}]
  wire  _GEN_1178 = 5'h11 == allocatePtrVec_1_value ? 1'h0 : _GEN_821; // @[Rob.scala 562:{22,22}]
  wire  _GEN_1179 = 5'h12 == allocatePtrVec_1_value ? 1'h0 : _GEN_822; // @[Rob.scala 562:{22,22}]
  wire  _GEN_1180 = 5'h13 == allocatePtrVec_1_value ? 1'h0 : _GEN_823; // @[Rob.scala 562:{22,22}]
  wire  _GEN_1181 = 5'h14 == allocatePtrVec_1_value ? 1'h0 : _GEN_824; // @[Rob.scala 562:{22,22}]
  wire  _GEN_1182 = 5'h15 == allocatePtrVec_1_value ? 1'h0 : _GEN_825; // @[Rob.scala 562:{22,22}]
  wire  _GEN_1183 = 5'h16 == allocatePtrVec_1_value ? 1'h0 : _GEN_826; // @[Rob.scala 562:{22,22}]
  wire  _GEN_1184 = 5'h17 == allocatePtrVec_1_value ? 1'h0 : _GEN_827; // @[Rob.scala 562:{22,22}]
  wire  _GEN_1185 = 5'h18 == allocatePtrVec_1_value ? 1'h0 : _GEN_828; // @[Rob.scala 562:{22,22}]
  wire  _GEN_1186 = 5'h19 == allocatePtrVec_1_value ? 1'h0 : _GEN_829; // @[Rob.scala 562:{22,22}]
  wire  _GEN_1187 = 5'h1a == allocatePtrVec_1_value ? 1'h0 : _GEN_830; // @[Rob.scala 562:{22,22}]
  wire  _GEN_1188 = 5'h1b == allocatePtrVec_1_value ? 1'h0 : _GEN_831; // @[Rob.scala 562:{22,22}]
  wire  _GEN_1189 = 5'h1c == allocatePtrVec_1_value ? 1'h0 : _GEN_832; // @[Rob.scala 562:{22,22}]
  wire  _GEN_1190 = 5'h1d == allocatePtrVec_1_value ? 1'h0 : _GEN_833; // @[Rob.scala 562:{22,22}]
  wire  _GEN_1191 = 5'h1e == allocatePtrVec_1_value ? 1'h0 : _GEN_834; // @[Rob.scala 562:{22,22}]
  wire  _GEN_1192 = 5'h1f == allocatePtrVec_1_value ? 1'h0 : _GEN_835; // @[Rob.scala 562:{22,22}]
  wire  _GEN_1631 = canEnqueue_1 ? _GEN_1161 : _GEN_804; // @[Rob.scala 523:26]
  wire  _GEN_1632 = canEnqueue_1 ? _GEN_1162 : _GEN_805; // @[Rob.scala 523:26]
  wire  _GEN_1633 = canEnqueue_1 ? _GEN_1163 : _GEN_806; // @[Rob.scala 523:26]
  wire  _GEN_1634 = canEnqueue_1 ? _GEN_1164 : _GEN_807; // @[Rob.scala 523:26]
  wire  _GEN_1635 = canEnqueue_1 ? _GEN_1165 : _GEN_808; // @[Rob.scala 523:26]
  wire  _GEN_1636 = canEnqueue_1 ? _GEN_1166 : _GEN_809; // @[Rob.scala 523:26]
  wire  _GEN_1637 = canEnqueue_1 ? _GEN_1167 : _GEN_810; // @[Rob.scala 523:26]
  wire  _GEN_1638 = canEnqueue_1 ? _GEN_1168 : _GEN_811; // @[Rob.scala 523:26]
  wire  _GEN_1639 = canEnqueue_1 ? _GEN_1169 : _GEN_812; // @[Rob.scala 523:26]
  wire  _GEN_1640 = canEnqueue_1 ? _GEN_1170 : _GEN_813; // @[Rob.scala 523:26]
  wire  _GEN_1641 = canEnqueue_1 ? _GEN_1171 : _GEN_814; // @[Rob.scala 523:26]
  wire  _GEN_1642 = canEnqueue_1 ? _GEN_1172 : _GEN_815; // @[Rob.scala 523:26]
  wire  _GEN_1643 = canEnqueue_1 ? _GEN_1173 : _GEN_816; // @[Rob.scala 523:26]
  wire  _GEN_1644 = canEnqueue_1 ? _GEN_1174 : _GEN_817; // @[Rob.scala 523:26]
  wire  _GEN_1645 = canEnqueue_1 ? _GEN_1175 : _GEN_818; // @[Rob.scala 523:26]
  wire  _GEN_1646 = canEnqueue_1 ? _GEN_1176 : _GEN_819; // @[Rob.scala 523:26]
  wire  _GEN_1647 = canEnqueue_1 ? _GEN_1177 : _GEN_820; // @[Rob.scala 523:26]
  wire  _GEN_1648 = canEnqueue_1 ? _GEN_1178 : _GEN_821; // @[Rob.scala 523:26]
  wire  _GEN_1649 = canEnqueue_1 ? _GEN_1179 : _GEN_822; // @[Rob.scala 523:26]
  wire  _GEN_1650 = canEnqueue_1 ? _GEN_1180 : _GEN_823; // @[Rob.scala 523:26]
  wire  _GEN_1651 = canEnqueue_1 ? _GEN_1181 : _GEN_824; // @[Rob.scala 523:26]
  wire  _GEN_1652 = canEnqueue_1 ? _GEN_1182 : _GEN_825; // @[Rob.scala 523:26]
  wire  _GEN_1653 = canEnqueue_1 ? _GEN_1183 : _GEN_826; // @[Rob.scala 523:26]
  wire  _GEN_1654 = canEnqueue_1 ? _GEN_1184 : _GEN_827; // @[Rob.scala 523:26]
  wire  _GEN_1655 = canEnqueue_1 ? _GEN_1185 : _GEN_828; // @[Rob.scala 523:26]
  wire  _GEN_1656 = canEnqueue_1 ? _GEN_1186 : _GEN_829; // @[Rob.scala 523:26]
  wire  _GEN_1657 = canEnqueue_1 ? _GEN_1187 : _GEN_830; // @[Rob.scala 523:26]
  wire  _GEN_1658 = canEnqueue_1 ? _GEN_1188 : _GEN_831; // @[Rob.scala 523:26]
  wire  _GEN_1659 = canEnqueue_1 ? _GEN_1189 : _GEN_832; // @[Rob.scala 523:26]
  wire  _GEN_1660 = canEnqueue_1 ? _GEN_1190 : _GEN_833; // @[Rob.scala 523:26]
  wire  _GEN_1661 = canEnqueue_1 ? _GEN_1191 : _GEN_834; // @[Rob.scala 523:26]
  wire  _GEN_1662 = canEnqueue_1 ? _GEN_1192 : _GEN_835; // @[Rob.scala 523:26]
  wire [1:0] _dispatchNum_T = io_enq_req_0_valid + io_enq_req_1_valid; // @[Bitwise.scala 48:55]
  wire [1:0] dispatchNum = io_enq_canAccept ? _dispatchNum_T : 2'h0; // @[Rob.scala 565:24]
  wire [1:0] _io_enq_isEmpty_T = {io_enq_req_1_valid,io_enq_req_0_valid}; // @[Rob.scala 566:76]
  reg  io_enq_isEmpty_REG; // @[Rob.scala 566:30]
  reg  REG_3; // @[Rob.scala 606:18]
  reg [4:0] REG_4; // @[Rob.scala 607:19]
  wire  _GEN_4679 = 5'h0 == REG_4 | _GEN_1631; // @[Rob.scala 607:{49,49}]
  wire  _GEN_4680 = 5'h1 == REG_4 | _GEN_1632; // @[Rob.scala 607:{49,49}]
  wire  _GEN_4681 = 5'h2 == REG_4 | _GEN_1633; // @[Rob.scala 607:{49,49}]
  wire  _GEN_4682 = 5'h3 == REG_4 | _GEN_1634; // @[Rob.scala 607:{49,49}]
  wire  _GEN_4683 = 5'h4 == REG_4 | _GEN_1635; // @[Rob.scala 607:{49,49}]
  wire  _GEN_4684 = 5'h5 == REG_4 | _GEN_1636; // @[Rob.scala 607:{49,49}]
  wire  _GEN_4685 = 5'h6 == REG_4 | _GEN_1637; // @[Rob.scala 607:{49,49}]
  wire  _GEN_4686 = 5'h7 == REG_4 | _GEN_1638; // @[Rob.scala 607:{49,49}]
  wire  _GEN_4687 = 5'h8 == REG_4 | _GEN_1639; // @[Rob.scala 607:{49,49}]
  wire  _GEN_4688 = 5'h9 == REG_4 | _GEN_1640; // @[Rob.scala 607:{49,49}]
  wire  _GEN_4689 = 5'ha == REG_4 | _GEN_1641; // @[Rob.scala 607:{49,49}]
  wire  _GEN_4690 = 5'hb == REG_4 | _GEN_1642; // @[Rob.scala 607:{49,49}]
  wire  _GEN_4691 = 5'hc == REG_4 | _GEN_1643; // @[Rob.scala 607:{49,49}]
  wire  _GEN_4692 = 5'hd == REG_4 | _GEN_1644; // @[Rob.scala 607:{49,49}]
  wire  _GEN_4693 = 5'he == REG_4 | _GEN_1645; // @[Rob.scala 607:{49,49}]
  wire  _GEN_4694 = 5'hf == REG_4 | _GEN_1646; // @[Rob.scala 607:{49,49}]
  wire  _GEN_4695 = 5'h10 == REG_4 | _GEN_1647; // @[Rob.scala 607:{49,49}]
  wire  _GEN_4696 = 5'h11 == REG_4 | _GEN_1648; // @[Rob.scala 607:{49,49}]
  wire  _GEN_4697 = 5'h12 == REG_4 | _GEN_1649; // @[Rob.scala 607:{49,49}]
  wire  _GEN_4698 = 5'h13 == REG_4 | _GEN_1650; // @[Rob.scala 607:{49,49}]
  wire  _GEN_4699 = 5'h14 == REG_4 | _GEN_1651; // @[Rob.scala 607:{49,49}]
  wire  _GEN_4700 = 5'h15 == REG_4 | _GEN_1652; // @[Rob.scala 607:{49,49}]
  wire  _GEN_4701 = 5'h16 == REG_4 | _GEN_1653; // @[Rob.scala 607:{49,49}]
  wire  _GEN_4702 = 5'h17 == REG_4 | _GEN_1654; // @[Rob.scala 607:{49,49}]
  wire  _GEN_4703 = 5'h18 == REG_4 | _GEN_1655; // @[Rob.scala 607:{49,49}]
  wire  _GEN_4704 = 5'h19 == REG_4 | _GEN_1656; // @[Rob.scala 607:{49,49}]
  wire  _GEN_4705 = 5'h1a == REG_4 | _GEN_1657; // @[Rob.scala 607:{49,49}]
  wire  _GEN_4706 = 5'h1b == REG_4 | _GEN_1658; // @[Rob.scala 607:{49,49}]
  wire  _GEN_4707 = 5'h1c == REG_4 | _GEN_1659; // @[Rob.scala 607:{49,49}]
  wire  _GEN_4708 = 5'h1d == REG_4 | _GEN_1660; // @[Rob.scala 607:{49,49}]
  wire  _GEN_4709 = 5'h1e == REG_4 | _GEN_1661; // @[Rob.scala 607:{49,49}]
  wire  _GEN_4710 = 5'h1f == REG_4 | _GEN_1662; // @[Rob.scala 607:{49,49}]
  wire  _GEN_4711 = REG_3 ? _GEN_4679 : _GEN_1631; // @[Rob.scala 606:38]
  wire  _GEN_4712 = REG_3 ? _GEN_4680 : _GEN_1632; // @[Rob.scala 606:38]
  wire  _GEN_4713 = REG_3 ? _GEN_4681 : _GEN_1633; // @[Rob.scala 606:38]
  wire  _GEN_4714 = REG_3 ? _GEN_4682 : _GEN_1634; // @[Rob.scala 606:38]
  wire  _GEN_4715 = REG_3 ? _GEN_4683 : _GEN_1635; // @[Rob.scala 606:38]
  wire  _GEN_4716 = REG_3 ? _GEN_4684 : _GEN_1636; // @[Rob.scala 606:38]
  wire  _GEN_4717 = REG_3 ? _GEN_4685 : _GEN_1637; // @[Rob.scala 606:38]
  wire  _GEN_4718 = REG_3 ? _GEN_4686 : _GEN_1638; // @[Rob.scala 606:38]
  wire  _GEN_4719 = REG_3 ? _GEN_4687 : _GEN_1639; // @[Rob.scala 606:38]
  wire  _GEN_4720 = REG_3 ? _GEN_4688 : _GEN_1640; // @[Rob.scala 606:38]
  wire  _GEN_4721 = REG_3 ? _GEN_4689 : _GEN_1641; // @[Rob.scala 606:38]
  wire  _GEN_4722 = REG_3 ? _GEN_4690 : _GEN_1642; // @[Rob.scala 606:38]
  wire  _GEN_4723 = REG_3 ? _GEN_4691 : _GEN_1643; // @[Rob.scala 606:38]
  wire  _GEN_4724 = REG_3 ? _GEN_4692 : _GEN_1644; // @[Rob.scala 606:38]
  wire  _GEN_4725 = REG_3 ? _GEN_4693 : _GEN_1645; // @[Rob.scala 606:38]
  wire  _GEN_4726 = REG_3 ? _GEN_4694 : _GEN_1646; // @[Rob.scala 606:38]
  wire  _GEN_4727 = REG_3 ? _GEN_4695 : _GEN_1647; // @[Rob.scala 606:38]
  wire  _GEN_4728 = REG_3 ? _GEN_4696 : _GEN_1648; // @[Rob.scala 606:38]
  wire  _GEN_4729 = REG_3 ? _GEN_4697 : _GEN_1649; // @[Rob.scala 606:38]
  wire  _GEN_4730 = REG_3 ? _GEN_4698 : _GEN_1650; // @[Rob.scala 606:38]
  wire  _GEN_4731 = REG_3 ? _GEN_4699 : _GEN_1651; // @[Rob.scala 606:38]
  wire  _GEN_4732 = REG_3 ? _GEN_4700 : _GEN_1652; // @[Rob.scala 606:38]
  wire  _GEN_4733 = REG_3 ? _GEN_4701 : _GEN_1653; // @[Rob.scala 606:38]
  wire  _GEN_4734 = REG_3 ? _GEN_4702 : _GEN_1654; // @[Rob.scala 606:38]
  wire  _GEN_4735 = REG_3 ? _GEN_4703 : _GEN_1655; // @[Rob.scala 606:38]
  wire  _GEN_4736 = REG_3 ? _GEN_4704 : _GEN_1656; // @[Rob.scala 606:38]
  wire  _GEN_4737 = REG_3 ? _GEN_4705 : _GEN_1657; // @[Rob.scala 606:38]
  wire  _GEN_4738 = REG_3 ? _GEN_4706 : _GEN_1658; // @[Rob.scala 606:38]
  wire  _GEN_4739 = REG_3 ? _GEN_4707 : _GEN_1659; // @[Rob.scala 606:38]
  wire  _GEN_4740 = REG_3 ? _GEN_4708 : _GEN_1660; // @[Rob.scala 606:38]
  wire  _GEN_4741 = REG_3 ? _GEN_4709 : _GEN_1661; // @[Rob.scala 606:38]
  wire  _GEN_4742 = REG_3 ? _GEN_4710 : _GEN_1662; // @[Rob.scala 606:38]
  reg  REG_5; // @[Rob.scala 606:18]
  reg [4:0] REG_6; // @[Rob.scala 607:19]
  wire  _GEN_4743 = 5'h0 == REG_6 | _GEN_4711; // @[Rob.scala 607:{49,49}]
  wire  _GEN_4744 = 5'h1 == REG_6 | _GEN_4712; // @[Rob.scala 607:{49,49}]
  wire  _GEN_4745 = 5'h2 == REG_6 | _GEN_4713; // @[Rob.scala 607:{49,49}]
  wire  _GEN_4746 = 5'h3 == REG_6 | _GEN_4714; // @[Rob.scala 607:{49,49}]
  wire  _GEN_4747 = 5'h4 == REG_6 | _GEN_4715; // @[Rob.scala 607:{49,49}]
  wire  _GEN_4748 = 5'h5 == REG_6 | _GEN_4716; // @[Rob.scala 607:{49,49}]
  wire  _GEN_4749 = 5'h6 == REG_6 | _GEN_4717; // @[Rob.scala 607:{49,49}]
  wire  _GEN_4750 = 5'h7 == REG_6 | _GEN_4718; // @[Rob.scala 607:{49,49}]
  wire  _GEN_4751 = 5'h8 == REG_6 | _GEN_4719; // @[Rob.scala 607:{49,49}]
  wire  _GEN_4752 = 5'h9 == REG_6 | _GEN_4720; // @[Rob.scala 607:{49,49}]
  wire  _GEN_4753 = 5'ha == REG_6 | _GEN_4721; // @[Rob.scala 607:{49,49}]
  wire  _GEN_4754 = 5'hb == REG_6 | _GEN_4722; // @[Rob.scala 607:{49,49}]
  wire  _GEN_4755 = 5'hc == REG_6 | _GEN_4723; // @[Rob.scala 607:{49,49}]
  wire  _GEN_4756 = 5'hd == REG_6 | _GEN_4724; // @[Rob.scala 607:{49,49}]
  wire  _GEN_4757 = 5'he == REG_6 | _GEN_4725; // @[Rob.scala 607:{49,49}]
  wire  _GEN_4758 = 5'hf == REG_6 | _GEN_4726; // @[Rob.scala 607:{49,49}]
  wire  _GEN_4759 = 5'h10 == REG_6 | _GEN_4727; // @[Rob.scala 607:{49,49}]
  wire  _GEN_4760 = 5'h11 == REG_6 | _GEN_4728; // @[Rob.scala 607:{49,49}]
  wire  _GEN_4761 = 5'h12 == REG_6 | _GEN_4729; // @[Rob.scala 607:{49,49}]
  wire  _GEN_4762 = 5'h13 == REG_6 | _GEN_4730; // @[Rob.scala 607:{49,49}]
  wire  _GEN_4763 = 5'h14 == REG_6 | _GEN_4731; // @[Rob.scala 607:{49,49}]
  wire  _GEN_4764 = 5'h15 == REG_6 | _GEN_4732; // @[Rob.scala 607:{49,49}]
  wire  _GEN_4765 = 5'h16 == REG_6 | _GEN_4733; // @[Rob.scala 607:{49,49}]
  wire  _GEN_4766 = 5'h17 == REG_6 | _GEN_4734; // @[Rob.scala 607:{49,49}]
  wire  _GEN_4767 = 5'h18 == REG_6 | _GEN_4735; // @[Rob.scala 607:{49,49}]
  wire  _GEN_4768 = 5'h19 == REG_6 | _GEN_4736; // @[Rob.scala 607:{49,49}]
  wire  _GEN_4769 = 5'h1a == REG_6 | _GEN_4737; // @[Rob.scala 607:{49,49}]
  wire  _GEN_4770 = 5'h1b == REG_6 | _GEN_4738; // @[Rob.scala 607:{49,49}]
  wire  _GEN_4771 = 5'h1c == REG_6 | _GEN_4739; // @[Rob.scala 607:{49,49}]
  wire  _GEN_4772 = 5'h1d == REG_6 | _GEN_4740; // @[Rob.scala 607:{49,49}]
  wire  _GEN_4773 = 5'h1e == REG_6 | _GEN_4741; // @[Rob.scala 607:{49,49}]
  wire  _GEN_4774 = 5'h1f == REG_6 | _GEN_4742; // @[Rob.scala 607:{49,49}]
  reg  intrBitSetReg; // @[Rob.scala 617:30]
  wire  intrEnable = intrBitSetReg & ~hasNoSpecExec & interrupt_safe_intrEnable_MPORT_data; // @[Rob.scala 618:52]
  wire [5:0] _deqHasExceptionOrFlush_T = {exceptionGen_io_state_bits_robIdx_flag,exceptionGen_io_state_bits_robIdx_value
    }; // @[CircularQueuePtr.scala 61:50]
  wire  _deqHasExceptionOrFlush_T_2 = _deqHasExceptionOrFlush_T == _isEmpty_T_1; // @[CircularQueuePtr.scala 61:52]
  wire  deqHasExceptionOrFlush = exceptionGen_io_state_valid & _deqHasExceptionOrFlush_T_2; // @[Rob.scala 619:56]
  wire [7:0] deqHasException_lo = {exceptionGen_io_state_bits_exceptionVec_7,exceptionGen_io_state_bits_exceptionVec_6,
    exceptionGen_io_state_bits_exceptionVec_5,exceptionGen_io_state_bits_exceptionVec_4,
    exceptionGen_io_state_bits_exceptionVec_3,exceptionGen_io_state_bits_exceptionVec_2,
    exceptionGen_io_state_bits_exceptionVec_1,exceptionGen_io_state_bits_exceptionVec_0}; // @[Rob.scala 620:88]
  wire [15:0] _deqHasException_T = {exceptionGen_io_state_bits_exceptionVec_15,
    exceptionGen_io_state_bits_exceptionVec_14,exceptionGen_io_state_bits_exceptionVec_13,
    exceptionGen_io_state_bits_exceptionVec_12,exceptionGen_io_state_bits_exceptionVec_11,
    exceptionGen_io_state_bits_exceptionVec_10,exceptionGen_io_state_bits_exceptionVec_9,
    exceptionGen_io_state_bits_exceptionVec_8,deqHasException_lo}; // @[Rob.scala 620:88]
  wire  _deqHasException_T_2 = |_deqHasException_T | exceptionGen_io_state_bits_singleStep; // @[Rob.scala 620:99]
  wire  _deqHasException_T_5 = exceptionGen_io_state_bits_trigger_frontendHit_0 |
    exceptionGen_io_state_bits_trigger_frontendHit_1 | exceptionGen_io_state_bits_trigger_frontendHit_2 |
    exceptionGen_io_state_bits_trigger_frontendHit_3; // @[Bundle.scala 628:45]
  wire  _deqHasException_T_10 = exceptionGen_io_state_bits_trigger_backendHit_0 |
    exceptionGen_io_state_bits_trigger_backendHit_1 | exceptionGen_io_state_bits_trigger_backendHit_2 |
    exceptionGen_io_state_bits_trigger_backendHit_3 | exceptionGen_io_state_bits_trigger_backendHit_4 |
    exceptionGen_io_state_bits_trigger_backendHit_5; // @[Bundle.scala 629:43]
  wire  _deqHasException_T_11 = _deqHasException_T_5 | _deqHasException_T_10; // @[Bundle.scala 630:28]
  wire  _deqHasException_T_12 = _deqHasException_T_2 | _deqHasException_T_11; // @[Rob.scala 621:39]
  wire  deqHasException = deqHasExceptionOrFlush & _deqHasException_T_12; // @[Rob.scala 620:48]
  wire  deqHasFlushPipe = deqHasExceptionOrFlush & exceptionGen_io_state_bits_flushPipe; // @[Rob.scala 622:48]
  wire  deqHasReplayInst = deqHasExceptionOrFlush & exceptionGen_io_state_bits_replayInst; // @[Rob.scala 623:49]
  wire  exceptionEnable = writebacked_exceptionEnable_MPORT_data & deqHasException; // @[Rob.scala 624:51]
  wire  isFlushPipe = writebacked_isFlushPipe_MPORT_data & (deqHasFlushPipe | deqHasReplayInst); // @[Rob.scala 630:47]
  reg  lastCycleFlush; // @[Rob.scala 634:31]
  wire  _io_flushOut_valid_T = ~state; // @[Rob.scala 636:31]
  wire  _GEN_4808 = 5'h1 == deqPtrVec_0_value ? valid_1 : valid_0; // @[Rob.scala 636:{43,43}]
  wire  _GEN_4809 = 5'h2 == deqPtrVec_0_value ? valid_2 : _GEN_4808; // @[Rob.scala 636:{43,43}]
  wire  _GEN_4810 = 5'h3 == deqPtrVec_0_value ? valid_3 : _GEN_4809; // @[Rob.scala 636:{43,43}]
  wire  _GEN_4811 = 5'h4 == deqPtrVec_0_value ? valid_4 : _GEN_4810; // @[Rob.scala 636:{43,43}]
  wire  _GEN_4812 = 5'h5 == deqPtrVec_0_value ? valid_5 : _GEN_4811; // @[Rob.scala 636:{43,43}]
  wire  _GEN_4813 = 5'h6 == deqPtrVec_0_value ? valid_6 : _GEN_4812; // @[Rob.scala 636:{43,43}]
  wire  _GEN_4814 = 5'h7 == deqPtrVec_0_value ? valid_7 : _GEN_4813; // @[Rob.scala 636:{43,43}]
  wire  _GEN_4815 = 5'h8 == deqPtrVec_0_value ? valid_8 : _GEN_4814; // @[Rob.scala 636:{43,43}]
  wire  _GEN_4816 = 5'h9 == deqPtrVec_0_value ? valid_9 : _GEN_4815; // @[Rob.scala 636:{43,43}]
  wire  _GEN_4817 = 5'ha == deqPtrVec_0_value ? valid_10 : _GEN_4816; // @[Rob.scala 636:{43,43}]
  wire  _GEN_4818 = 5'hb == deqPtrVec_0_value ? valid_11 : _GEN_4817; // @[Rob.scala 636:{43,43}]
  wire  _GEN_4819 = 5'hc == deqPtrVec_0_value ? valid_12 : _GEN_4818; // @[Rob.scala 636:{43,43}]
  wire  _GEN_4820 = 5'hd == deqPtrVec_0_value ? valid_13 : _GEN_4819; // @[Rob.scala 636:{43,43}]
  wire  _GEN_4821 = 5'he == deqPtrVec_0_value ? valid_14 : _GEN_4820; // @[Rob.scala 636:{43,43}]
  wire  _GEN_4822 = 5'hf == deqPtrVec_0_value ? valid_15 : _GEN_4821; // @[Rob.scala 636:{43,43}]
  wire  _GEN_4823 = 5'h10 == deqPtrVec_0_value ? valid_16 : _GEN_4822; // @[Rob.scala 636:{43,43}]
  wire  _GEN_4824 = 5'h11 == deqPtrVec_0_value ? valid_17 : _GEN_4823; // @[Rob.scala 636:{43,43}]
  wire  _GEN_4825 = 5'h12 == deqPtrVec_0_value ? valid_18 : _GEN_4824; // @[Rob.scala 636:{43,43}]
  wire  _GEN_4826 = 5'h13 == deqPtrVec_0_value ? valid_19 : _GEN_4825; // @[Rob.scala 636:{43,43}]
  wire  _GEN_4827 = 5'h14 == deqPtrVec_0_value ? valid_20 : _GEN_4826; // @[Rob.scala 636:{43,43}]
  wire  _GEN_4828 = 5'h15 == deqPtrVec_0_value ? valid_21 : _GEN_4827; // @[Rob.scala 636:{43,43}]
  wire  _GEN_4829 = 5'h16 == deqPtrVec_0_value ? valid_22 : _GEN_4828; // @[Rob.scala 636:{43,43}]
  wire  _GEN_4830 = 5'h17 == deqPtrVec_0_value ? valid_23 : _GEN_4829; // @[Rob.scala 636:{43,43}]
  wire  _GEN_4831 = 5'h18 == deqPtrVec_0_value ? valid_24 : _GEN_4830; // @[Rob.scala 636:{43,43}]
  wire  _GEN_4832 = 5'h19 == deqPtrVec_0_value ? valid_25 : _GEN_4831; // @[Rob.scala 636:{43,43}]
  wire  _GEN_4833 = 5'h1a == deqPtrVec_0_value ? valid_26 : _GEN_4832; // @[Rob.scala 636:{43,43}]
  wire  _GEN_4834 = 5'h1b == deqPtrVec_0_value ? valid_27 : _GEN_4833; // @[Rob.scala 636:{43,43}]
  wire  _GEN_4835 = 5'h1c == deqPtrVec_0_value ? valid_28 : _GEN_4834; // @[Rob.scala 636:{43,43}]
  wire  _GEN_4836 = 5'h1d == deqPtrVec_0_value ? valid_29 : _GEN_4835; // @[Rob.scala 636:{43,43}]
  wire  _GEN_4837 = 5'h1e == deqPtrVec_0_value ? valid_30 : _GEN_4836; // @[Rob.scala 636:{43,43}]
  wire  commit_v_0 = 5'h1f == deqPtrVec_0_value ? valid_31 : _GEN_4837; // @[Rob.scala 636:{43,43}]
  wire  _io_flushOut_valid_T_1 = ~state & commit_v_0; // @[Rob.scala 636:43]
  wire  _io_flushOut_valid_T_2 = intrEnable | exceptionEnable; // @[Rob.scala 636:81]
  wire  _io_flushOut_valid_T_5 = ~lastCycleFlush; // @[Rob.scala 636:119]
  wire  _T_108 = io_flushOut_valid & isFlushPipe; // @[Rob.scala 645:56]
  wire  exceptionHappen = _io_flushOut_valid_T_1 & _io_flushOut_valid_T_2 & _io_flushOut_valid_T_5; // @[Rob.scala 648:102]
  reg  io_exception_valid_REG; // @[Rob.scala 649:32]
  reg [2:0] io_exception_bits_uop_ctrl_commitType_r; // @[Reg.scala 16:16]
  reg  r_0; // @[Reg.scala 16:16]
  reg  r_1; // @[Reg.scala 16:16]
  reg  r_2; // @[Reg.scala 16:16]
  reg  r_3; // @[Reg.scala 16:16]
  reg  r_4; // @[Reg.scala 16:16]
  reg  r_5; // @[Reg.scala 16:16]
  reg  r_6; // @[Reg.scala 16:16]
  reg  r_7; // @[Reg.scala 16:16]
  reg  r_8; // @[Reg.scala 16:16]
  reg  r_9; // @[Reg.scala 16:16]
  reg  r_11; // @[Reg.scala 16:16]
  reg  r_12; // @[Reg.scala 16:16]
  reg  r_13; // @[Reg.scala 16:16]
  reg  r_15; // @[Reg.scala 16:16]
  reg  io_exception_bits_uop_ctrl_singleStep_r; // @[Reg.scala 16:16]
  reg  io_exception_bits_uop_cf_crossPageIPFFix_r; // @[Reg.scala 16:16]
  reg  io_exception_bits_isInterrupt_r; // @[Reg.scala 16:16]
  reg  io_exception_bits_uop_cf_trigger_rfrontendHit_0; // @[Reg.scala 16:16]
  reg  io_exception_bits_uop_cf_trigger_rfrontendHit_1; // @[Reg.scala 16:16]
  reg  io_exception_bits_uop_cf_trigger_rfrontendHit_2; // @[Reg.scala 16:16]
  reg  io_exception_bits_uop_cf_trigger_rfrontendHit_3; // @[Reg.scala 16:16]
  reg  io_exception_bits_uop_cf_trigger_rbackendHit_0; // @[Reg.scala 16:16]
  reg  io_exception_bits_uop_cf_trigger_rbackendHit_1; // @[Reg.scala 16:16]
  reg  io_exception_bits_uop_cf_trigger_rbackendHit_2; // @[Reg.scala 16:16]
  reg  io_exception_bits_uop_cf_trigger_rbackendHit_3; // @[Reg.scala 16:16]
  reg  io_exception_bits_uop_cf_trigger_rbackendHit_4; // @[Reg.scala 16:16]
  reg  io_exception_bits_uop_cf_trigger_rbackendHit_5; // @[Reg.scala 16:16]
  reg [5:0] walkCounter; // @[Rob.scala 668:24]
  wire  walkFinished = walkCounter <= 6'h2; // @[Rob.scala 670:34]
  wire  wflags_0 = io_commits_commitValid_0 & io_commits_info_0_wflags; // @[Rob.scala 678:8]
  wire  fpWen_0 = io_commits_commitValid_0 & io_commits_info_0_fpWen; // @[Rob.scala 678:25]
  wire  wflags_1 = io_commits_commitValid_1 & io_commits_info_1_wflags; // @[Rob.scala 678:8]
  wire  fpWen_1 = io_commits_commitValid_1 & io_commits_info_1_fpWen; // @[Rob.scala 678:25]
  wire [1:0] _fflags_valid_T = {wflags_1,wflags_0}; // @[Rob.scala 681:58]
  wire [4:0] fflagsDataRead_0 = fflagsDataModule_io_rdata_0; // @[Rob.scala 1016:18 482:28]
  wire [4:0] _fflags_bits_T = wflags_0 ? fflagsDataRead_0 : 5'h0; // @[Rob.scala 683:23]
  wire [4:0] fflagsDataRead_1 = fflagsDataModule_io_rdata_1; // @[Rob.scala 1016:18 482:28]
  wire [4:0] _fflags_bits_T_1 = wflags_1 ? fflagsDataRead_1 : 5'h0; // @[Rob.scala 683:23]
  wire [1:0] _dirty_fs_T = {fpWen_1,fpWen_0}; // @[Rob.scala 685:56]
  wire  _misPredWb_T = io_writeback_1_0_bits_redirect_cfiUpdate_isMisPred & io_writeback_1_0_bits_redirectValid; // @[Rob.scala 690:42]
  wire  _misPredWb_T_1 = io_writeback_1_1_bits_redirect_cfiUpdate_isMisPred & io_writeback_1_1_bits_redirectValid; // @[Rob.scala 690:42]
  wire  _misPredWb_T_4 = io_writeback_1_4_bits_redirect_cfiUpdate_isMisPred & io_writeback_1_4_bits_redirectValid; // @[Rob.scala 690:42]
  wire  _misPredWb_T_6 = io_writeback_1_6_bits_redirect_cfiUpdate_isMisPred & io_writeback_1_6_bits_redirectValid; // @[Rob.scala 690:42]
  wire  _misPredWb_T_7 = io_writeback_1_7_bits_redirect_cfiUpdate_isMisPred & io_writeback_1_7_bits_redirectValid; // @[Rob.scala 690:42]
  wire  _misPredWb_T_8 = io_writeback_1_8_bits_redirect_cfiUpdate_isMisPred & io_writeback_1_8_bits_redirectValid; // @[Rob.scala 690:42]
  wire [8:0] _misPredWb_T_9 = {_misPredWb_T,_misPredWb_T_1,1'h0,1'h0,_misPredWb_T_4,1'h0,_misPredWb_T_6,_misPredWb_T_7,
    _misPredWb_T_8}; // @[Cat.scala 31:58]
  wire  misPredWb = |_misPredWb_T_9; // @[Rob.scala 691:7]
  reg [2:0] misPredBlockCounter; // @[Rob.scala 692:32]
  wire [2:0] _misPredBlockCounter_T = {{1'd0}, misPredBlockCounter[2:1]}; // @[Rob.scala 695:25]
  wire  misPredBlock = misPredBlockCounter[0]; // @[Rob.scala 697:41]
  wire  blockCommit = misPredBlock | isReplaying | lastCycleFlush | hasWFI; // @[Rob.scala 698:67]
  wire [4:0] deqPtrVec_1_value = deqPtrGenModule_io_out_1_value; // @[Rob.scala 448:23 783:13]
  wire  _GEN_5044 = 5'h1 == deqPtrVec_1_value ? valid_1 : valid_0; // @[Rob.scala 703:{25,25}]
  wire  _GEN_5045 = 5'h2 == deqPtrVec_1_value ? valid_2 : _GEN_5044; // @[Rob.scala 703:{25,25}]
  wire  _GEN_5046 = 5'h3 == deqPtrVec_1_value ? valid_3 : _GEN_5045; // @[Rob.scala 703:{25,25}]
  wire  _GEN_5047 = 5'h4 == deqPtrVec_1_value ? valid_4 : _GEN_5046; // @[Rob.scala 703:{25,25}]
  wire  _GEN_5048 = 5'h5 == deqPtrVec_1_value ? valid_5 : _GEN_5047; // @[Rob.scala 703:{25,25}]
  wire  _GEN_5049 = 5'h6 == deqPtrVec_1_value ? valid_6 : _GEN_5048; // @[Rob.scala 703:{25,25}]
  wire  _GEN_5050 = 5'h7 == deqPtrVec_1_value ? valid_7 : _GEN_5049; // @[Rob.scala 703:{25,25}]
  wire  _GEN_5051 = 5'h8 == deqPtrVec_1_value ? valid_8 : _GEN_5050; // @[Rob.scala 703:{25,25}]
  wire  _GEN_5052 = 5'h9 == deqPtrVec_1_value ? valid_9 : _GEN_5051; // @[Rob.scala 703:{25,25}]
  wire  _GEN_5053 = 5'ha == deqPtrVec_1_value ? valid_10 : _GEN_5052; // @[Rob.scala 703:{25,25}]
  wire  _GEN_5054 = 5'hb == deqPtrVec_1_value ? valid_11 : _GEN_5053; // @[Rob.scala 703:{25,25}]
  wire  _GEN_5055 = 5'hc == deqPtrVec_1_value ? valid_12 : _GEN_5054; // @[Rob.scala 703:{25,25}]
  wire  _GEN_5056 = 5'hd == deqPtrVec_1_value ? valid_13 : _GEN_5055; // @[Rob.scala 703:{25,25}]
  wire  _GEN_5057 = 5'he == deqPtrVec_1_value ? valid_14 : _GEN_5056; // @[Rob.scala 703:{25,25}]
  wire  _GEN_5058 = 5'hf == deqPtrVec_1_value ? valid_15 : _GEN_5057; // @[Rob.scala 703:{25,25}]
  wire  _GEN_5059 = 5'h10 == deqPtrVec_1_value ? valid_16 : _GEN_5058; // @[Rob.scala 703:{25,25}]
  wire  _GEN_5060 = 5'h11 == deqPtrVec_1_value ? valid_17 : _GEN_5059; // @[Rob.scala 703:{25,25}]
  wire  _GEN_5061 = 5'h12 == deqPtrVec_1_value ? valid_18 : _GEN_5060; // @[Rob.scala 703:{25,25}]
  wire  _GEN_5062 = 5'h13 == deqPtrVec_1_value ? valid_19 : _GEN_5061; // @[Rob.scala 703:{25,25}]
  wire  _GEN_5063 = 5'h14 == deqPtrVec_1_value ? valid_20 : _GEN_5062; // @[Rob.scala 703:{25,25}]
  wire  _GEN_5064 = 5'h15 == deqPtrVec_1_value ? valid_21 : _GEN_5063; // @[Rob.scala 703:{25,25}]
  wire  _GEN_5065 = 5'h16 == deqPtrVec_1_value ? valid_22 : _GEN_5064; // @[Rob.scala 703:{25,25}]
  wire  _GEN_5066 = 5'h17 == deqPtrVec_1_value ? valid_23 : _GEN_5065; // @[Rob.scala 703:{25,25}]
  wire  _GEN_5067 = 5'h18 == deqPtrVec_1_value ? valid_24 : _GEN_5066; // @[Rob.scala 703:{25,25}]
  wire  _GEN_5068 = 5'h19 == deqPtrVec_1_value ? valid_25 : _GEN_5067; // @[Rob.scala 703:{25,25}]
  wire  _GEN_5069 = 5'h1a == deqPtrVec_1_value ? valid_26 : _GEN_5068; // @[Rob.scala 703:{25,25}]
  wire  _GEN_5070 = 5'h1b == deqPtrVec_1_value ? valid_27 : _GEN_5069; // @[Rob.scala 703:{25,25}]
  wire  _GEN_5071 = 5'h1c == deqPtrVec_1_value ? valid_28 : _GEN_5070; // @[Rob.scala 703:{25,25}]
  wire  _GEN_5072 = 5'h1d == deqPtrVec_1_value ? valid_29 : _GEN_5071; // @[Rob.scala 703:{25,25}]
  wire  _GEN_5073 = 5'h1e == deqPtrVec_1_value ? valid_30 : _GEN_5072; // @[Rob.scala 703:{25,25}]
  wire  commit_v_1 = 5'h1f == deqPtrVec_1_value ? valid_31 : _GEN_5073; // @[Rob.scala 703:{25,25}]
  wire  commit_w0 = writebacked_commit_wMPORT_data & store_data_writebacked_commit_wMPORT_1_data; // @[Rob.scala 705:70]
  wire  commit_w1 = writebacked_commit_wMPORT_2_data & store_data_writebacked_commit_wMPORT_3_data; // @[Rob.scala 705:70]
  wire  deqPtrVec_1_flag = deqPtrGenModule_io_out_1_flag; // @[Rob.scala 448:23 783:13]
  wire  commit_exception_differentFlag = exceptionGen_io_state_bits_robIdx_flag ^ deqPtrVec_1_flag; // @[CircularQueuePtr.scala 86:35]
  wire  commit_exception_compare = exceptionGen_io_state_bits_robIdx_value > deqPtrVec_1_value; // @[CircularQueuePtr.scala 87:30]
  wire  _commit_exception_T = commit_exception_differentFlag ^ commit_exception_compare; // @[CircularQueuePtr.scala 88:19]
  wire  commit_exception = exceptionGen_io_state_valid & ~_commit_exception_T; // @[Rob.scala 706:50]
  wire  commit_block_0 = ~commit_w0; // @[Rob.scala 707:61]
  wire  allowOnlyOneCommit = commit_exception | intrBitSetReg; // @[Rob.scala 708:45]
  wire  isBlocked = intrEnable | deqHasException | deqHasReplayInst; // @[Rob.scala 713:120]
  wire  _T_117 = io_commits_isCommit & io_commits_commitValid_0; // @[Rob.scala 724:32]
  wire  isBlocked_1 = |commit_block_0 | allowOnlyOneCommit; // @[Rob.scala 713:63]
  wire  _T_125 = io_commits_isCommit & io_commits_commitValid_1; // @[Rob.scala 724:32]
  reg  io_csr_fflags_REG_valid; // @[Rob.scala 746:27]
  reg [4:0] io_csr_fflags_REG_bits; // @[Rob.scala 746:27]
  reg  io_csr_dirty_fs_REG; // @[Rob.scala 747:29]
  wire  _ldCommitVec_T = io_commits_info_0_commitType == 3'h2; // @[Rob.scala 750:119]
  wire  ldCommitVec_0 = io_commits_commitValid_0 & io_commits_info_0_commitType == 3'h2; // @[Rob.scala 750:86]
  wire  _ldCommitVec_T_2 = io_commits_info_1_commitType == 3'h2; // @[Rob.scala 750:119]
  wire  ldCommitVec_1 = io_commits_commitValid_1 & io_commits_info_1_commitType == 3'h2; // @[Rob.scala 750:86]
  wire  _stCommitVec_T = io_commits_info_0_commitType == 3'h3; // @[Rob.scala 751:119]
  wire  stCommitVec_0 = io_commits_commitValid_0 & io_commits_info_0_commitType == 3'h3; // @[Rob.scala 751:86]
  wire  _stCommitVec_T_2 = io_commits_info_1_commitType == 3'h3; // @[Rob.scala 751:119]
  wire  stCommitVec_1 = io_commits_commitValid_1 & io_commits_info_1_commitType == 3'h3; // @[Rob.scala 751:86]
  wire [1:0] _io_lsq_scommit_T = stCommitVec_0 + stCommitVec_1; // @[Bitwise.scala 48:55]
  reg [1:0] io_lsq_scommit_REG; // @[Rob.scala 753:28]
  wire  _GEN_5078 = 5'h1 == deqPtrVec_0_value ? mmio_1 : mmio_0; // @[Rob.scala 755:{127,127}]
  wire  _GEN_5079 = 5'h2 == deqPtrVec_0_value ? mmio_2 : _GEN_5078; // @[Rob.scala 755:{127,127}]
  wire  _GEN_5080 = 5'h3 == deqPtrVec_0_value ? mmio_3 : _GEN_5079; // @[Rob.scala 755:{127,127}]
  wire  _GEN_5081 = 5'h4 == deqPtrVec_0_value ? mmio_4 : _GEN_5080; // @[Rob.scala 755:{127,127}]
  wire  _GEN_5082 = 5'h5 == deqPtrVec_0_value ? mmio_5 : _GEN_5081; // @[Rob.scala 755:{127,127}]
  wire  _GEN_5083 = 5'h6 == deqPtrVec_0_value ? mmio_6 : _GEN_5082; // @[Rob.scala 755:{127,127}]
  wire  _GEN_5084 = 5'h7 == deqPtrVec_0_value ? mmio_7 : _GEN_5083; // @[Rob.scala 755:{127,127}]
  wire  _GEN_5085 = 5'h8 == deqPtrVec_0_value ? mmio_8 : _GEN_5084; // @[Rob.scala 755:{127,127}]
  wire  _GEN_5086 = 5'h9 == deqPtrVec_0_value ? mmio_9 : _GEN_5085; // @[Rob.scala 755:{127,127}]
  wire  _GEN_5087 = 5'ha == deqPtrVec_0_value ? mmio_10 : _GEN_5086; // @[Rob.scala 755:{127,127}]
  wire  _GEN_5088 = 5'hb == deqPtrVec_0_value ? mmio_11 : _GEN_5087; // @[Rob.scala 755:{127,127}]
  wire  _GEN_5089 = 5'hc == deqPtrVec_0_value ? mmio_12 : _GEN_5088; // @[Rob.scala 755:{127,127}]
  wire  _GEN_5090 = 5'hd == deqPtrVec_0_value ? mmio_13 : _GEN_5089; // @[Rob.scala 755:{127,127}]
  wire  _GEN_5091 = 5'he == deqPtrVec_0_value ? mmio_14 : _GEN_5090; // @[Rob.scala 755:{127,127}]
  wire  _GEN_5092 = 5'hf == deqPtrVec_0_value ? mmio_15 : _GEN_5091; // @[Rob.scala 755:{127,127}]
  wire  _GEN_5093 = 5'h10 == deqPtrVec_0_value ? mmio_16 : _GEN_5092; // @[Rob.scala 755:{127,127}]
  wire  _GEN_5094 = 5'h11 == deqPtrVec_0_value ? mmio_17 : _GEN_5093; // @[Rob.scala 755:{127,127}]
  wire  _GEN_5095 = 5'h12 == deqPtrVec_0_value ? mmio_18 : _GEN_5094; // @[Rob.scala 755:{127,127}]
  wire  _GEN_5096 = 5'h13 == deqPtrVec_0_value ? mmio_19 : _GEN_5095; // @[Rob.scala 755:{127,127}]
  wire  _GEN_5097 = 5'h14 == deqPtrVec_0_value ? mmio_20 : _GEN_5096; // @[Rob.scala 755:{127,127}]
  wire  _GEN_5098 = 5'h15 == deqPtrVec_0_value ? mmio_21 : _GEN_5097; // @[Rob.scala 755:{127,127}]
  wire  _GEN_5099 = 5'h16 == deqPtrVec_0_value ? mmio_22 : _GEN_5098; // @[Rob.scala 755:{127,127}]
  wire  _GEN_5100 = 5'h17 == deqPtrVec_0_value ? mmio_23 : _GEN_5099; // @[Rob.scala 755:{127,127}]
  wire  _GEN_5101 = 5'h18 == deqPtrVec_0_value ? mmio_24 : _GEN_5100; // @[Rob.scala 755:{127,127}]
  wire  _GEN_5102 = 5'h19 == deqPtrVec_0_value ? mmio_25 : _GEN_5101; // @[Rob.scala 755:{127,127}]
  wire  _GEN_5103 = 5'h1a == deqPtrVec_0_value ? mmio_26 : _GEN_5102; // @[Rob.scala 755:{127,127}]
  wire  _GEN_5104 = 5'h1b == deqPtrVec_0_value ? mmio_27 : _GEN_5103; // @[Rob.scala 755:{127,127}]
  wire  _GEN_5105 = 5'h1c == deqPtrVec_0_value ? mmio_28 : _GEN_5104; // @[Rob.scala 755:{127,127}]
  wire  _GEN_5106 = 5'h1d == deqPtrVec_0_value ? mmio_29 : _GEN_5105; // @[Rob.scala 755:{127,127}]
  wire  _GEN_5107 = 5'h1e == deqPtrVec_0_value ? mmio_30 : _GEN_5106; // @[Rob.scala 755:{127,127}]
  wire  _GEN_5108 = 5'h1f == deqPtrVec_0_value ? mmio_31 : _GEN_5107; // @[Rob.scala 755:{127,127}]
  reg  io_lsq_pendingld_REG; // @[Rob.scala 755:30]
  reg  io_lsq_pendingst_REG; // @[Rob.scala 756:30]
  reg  io_lsq_commit_REG; // @[Rob.scala 757:27]
  wire  _state_next_T_2 = state & walkFinished ? 1'h0 : state; // @[Rob.scala 764:54]
  wire  state_next = io_redirect_valid | _state_next_T_2; // @[Rob.scala 764:23]
  wire  _T_129 = ~state_next; // @[Rob.scala 765:80]
  wire [5:0] thisCycleWalkCount = walkFinished ? walkCounter : 6'h2; // @[Rob.scala 793:31]
  wire [5:0] _walkPtrVec_next_new_ptr_T = {walkPtrVec_0_flag,walkPtrVec_0_value}; // @[Cat.scala 31:58]
  wire [5:0] _walkPtrVec_next_new_ptr_T_2 = _walkPtrVec_next_new_ptr_T + 6'h2; // @[CircularQueuePtr.scala 39:46]
  wire [4:0] walkPtrVec_next_new_ptr_value = _walkPtrVec_next_new_ptr_T_2[4:0]; // @[CircularQueuePtr.scala 39:59]
  wire  walkPtrVec_next_new_ptr_flag = _walkPtrVec_next_new_ptr_T_2[5]; // @[CircularQueuePtr.scala 39:59]
  wire [5:0] _walkPtrVec_next_new_ptr_T_5 = {walkPtrVec_1_flag,walkPtrVec_1_value}; // @[Cat.scala 31:58]
  wire [5:0] _walkPtrVec_next_new_ptr_T_7 = _walkPtrVec_next_new_ptr_T_5 + 6'h2; // @[CircularQueuePtr.scala 39:46]
  wire [4:0] walkPtrVec_next_new_ptr_1_value = _walkPtrVec_next_new_ptr_T_7[4:0]; // @[CircularQueuePtr.scala 39:59]
  wire  walkPtrVec_next_new_ptr_1_flag = _walkPtrVec_next_new_ptr_T_7[5]; // @[CircularQueuePtr.scala 39:59]
  wire [4:0] _walkPtrVec_next_T_1_0_value = state ? walkPtrVec_next_new_ptr_value : walkPtrVec_0_value; // @[Rob.scala 799:8]
  wire [4:0] _walkPtrVec_next_T_1_1_value = state ? walkPtrVec_next_new_ptr_1_value : walkPtrVec_1_value; // @[Rob.scala 799:8]
  wire [4:0] walkPtrVec_next_0_value = io_redirect_valid ? deqPtrGenModule_io_next_out_0_value :
    _walkPtrVec_next_T_1_0_value; // @[Rob.scala 797:28]
  wire [4:0] walkPtrVec_next_1_value = io_redirect_valid ? deqPtrGenModule_io_next_out_1_value :
    _walkPtrVec_next_T_1_1_value; // @[Rob.scala 797:28]
  wire [4:0] _numValidEntries_T_2 = enqPtrVec_0_value - deqPtrVec_0_value; // @[CircularQueuePtr.scala 81:21]
  wire [5:0] _GEN_11213 = {{1'd0}, enqPtrVec_0_value}; // @[CircularQueuePtr.scala 82:25]
  wire [5:0] _numValidEntries_T_4 = 6'h20 + _GEN_11213; // @[CircularQueuePtr.scala 82:25]
  wire [5:0] _GEN_11214 = {{1'd0}, deqPtrVec_0_value}; // @[CircularQueuePtr.scala 82:41]
  wire [5:0] _numValidEntries_T_6 = _numValidEntries_T_4 - _GEN_11214; // @[CircularQueuePtr.scala 82:41]
  wire [5:0] numValidEntries = enqPtrVec_0_flag == deqPtrVec_0_flag ? {{1'd0}, _numValidEntries_T_2} :
    _numValidEntries_T_6; // @[CircularQueuePtr.scala 80:8]
  wire [1:0] commitCnt = io_commits_commitValid_0 + io_commits_commitValid_1; // @[Bitwise.scala 48:55]
  wire [5:0] _GEN_11215 = {{4'd0}, dispatchNum}; // @[Rob.scala 806:35]
  wire [5:0] _allowEnqueue_T_1 = numValidEntries + _GEN_11215; // @[Rob.scala 806:35]
  wire [4:0] _redirectWalkDistance_T_2 = io_redirect_bits_robIdx_value - deqPtrGenModule_io_next_out_0_value; // @[CircularQueuePtr.scala 81:21]
  wire [5:0] _GEN_11216 = {{1'd0}, io_redirect_bits_robIdx_value}; // @[CircularQueuePtr.scala 82:25]
  wire [5:0] _redirectWalkDistance_T_4 = 6'h20 + _GEN_11216; // @[CircularQueuePtr.scala 82:25]
  wire [5:0] _GEN_11217 = {{1'd0}, deqPtrGenModule_io_next_out_0_value}; // @[CircularQueuePtr.scala 82:41]
  wire [5:0] _redirectWalkDistance_T_6 = _redirectWalkDistance_T_4 - _GEN_11217; // @[CircularQueuePtr.scala 82:41]
  wire [5:0] redirectWalkDistance = io_redirect_bits_robIdx_flag == deqPtrGenModule_io_next_out_0_flag ? {{1'd0},
    _redirectWalkDistance_T_2} : _redirectWalkDistance_T_6; // @[CircularQueuePtr.scala 80:8]
  wire  walkCounter_differentFlag = io_redirect_bits_robIdx_flag ^ deqPtrGenModule_io_next_out_0_flag; // @[CircularQueuePtr.scala 92:35]
  wire  walkCounter_compare = io_redirect_bits_robIdx_value < deqPtrGenModule_io_next_out_0_value; // @[CircularQueuePtr.scala 93:30]
  wire  _walkCounter_T = walkCounter_differentFlag ^ walkCounter_compare; // @[CircularQueuePtr.scala 94:19]
  wire  _walkCounter_T_2 = ~io_redirect_bits_level; // @[Rob.scala 825:48]
  wire [5:0] _GEN_11218 = {{5'd0}, _walkCounter_T_2}; // @[Rob.scala 825:45]
  wire [6:0] _walkCounter_T_3 = redirectWalkDistance + _GEN_11218; // @[Rob.scala 825:45]
  wire [6:0] _walkCounter_T_4 = _walkCounter_T ? 7'h0 : _walkCounter_T_3; // @[Rob.scala 824:23]
  wire [5:0] _walkCounter_T_6 = walkCounter - thisCycleWalkCount; // @[Rob.scala 827:32]
  wire [5:0] _GEN_5109 = state ? _walkCounter_T_6 : walkCounter; // @[Rob.scala 826:33 827:17 668:24]
  wire [6:0] _GEN_5110 = io_redirect_valid ? _walkCounter_T_4 : {{1'd0}, _GEN_5109}; // @[Rob.scala 810:28 824:17]
  wire [4:0] commitReadAddr_0 = _io_flushOut_valid_T ? deqPtrVec_0_value : walkPtrVec_0_value; // @[Rob.scala 839:27]
  wire [4:0] commitReadAddr_1 = _io_flushOut_valid_T ? deqPtrVec_1_value : walkPtrVec_1_value; // @[Rob.scala 839:27]
  reg  redirectHeadVec_0_flag; // @[Rob.scala 842:28]
  reg [4:0] redirectHeadVec_0_value; // @[Rob.scala 842:28]
  reg  redirectHeadVec_1_flag; // @[Rob.scala 842:28]
  reg [4:0] redirectHeadVec_1_value; // @[Rob.scala 842:28]
  reg  redirectTail_flag; // @[Rob.scala 843:25]
  reg [4:0] redirectTail_value; // @[Rob.scala 843:25]
  reg  redirectState; // @[Rob.scala 845:30]
  wire  invMask_differentFlag = redirectHeadVec_0_flag ^ redirectTail_flag; // @[CircularQueuePtr.scala 92:35]
  wire  invMask_compare = redirectHeadVec_0_value < redirectTail_value; // @[CircularQueuePtr.scala 93:30]
  wire  invMask_0 = invMask_differentFlag ^ invMask_compare; // @[CircularQueuePtr.scala 94:19]
  wire  invMask_differentFlag_1 = redirectHeadVec_1_flag ^ redirectTail_flag; // @[CircularQueuePtr.scala 92:35]
  wire  invMask_compare_1 = redirectHeadVec_1_value < redirectTail_value; // @[CircularQueuePtr.scala 93:30]
  wire  invMask_1 = invMask_differentFlag_1 ^ invMask_compare_1; // @[CircularQueuePtr.scala 94:19]
  wire [5:0] _redirectHeadVec_0_new_ptr_T = {redirectHeadVec_0_flag,redirectHeadVec_0_value}; // @[Cat.scala 31:58]
  wire [5:0] _redirectHeadVec_0_new_ptr_T_2 = _redirectHeadVec_0_new_ptr_T + 6'h2; // @[CircularQueuePtr.scala 39:46]
  wire [4:0] redirectHeadVec_0_new_ptr_value = _redirectHeadVec_0_new_ptr_T_2[4:0]; // @[CircularQueuePtr.scala 39:59]
  wire  redirectHeadVec_0_new_ptr_flag = _redirectHeadVec_0_new_ptr_T_2[5]; // @[CircularQueuePtr.scala 39:59]
  wire [5:0] _redirectHeadVec_1_new_ptr_T = {redirectHeadVec_1_flag,redirectHeadVec_1_value}; // @[Cat.scala 31:58]
  wire [5:0] _redirectHeadVec_1_new_ptr_T_2 = _redirectHeadVec_1_new_ptr_T + 6'h2; // @[CircularQueuePtr.scala 39:46]
  wire [4:0] redirectHeadVec_1_new_ptr_value = _redirectHeadVec_1_new_ptr_T_2[4:0]; // @[CircularQueuePtr.scala 39:59]
  wire  redirectHeadVec_1_new_ptr_flag = _redirectHeadVec_1_new_ptr_T_2[5]; // @[CircularQueuePtr.scala 39:59]
  wire  _GEN_5111 = 5'h0 == redirectHeadVec_0_value ? 1'h0 : valid_0; // @[Rob.scala 426:22 851:{35,35}]
  wire  _GEN_5112 = 5'h1 == redirectHeadVec_0_value ? 1'h0 : valid_1; // @[Rob.scala 426:22 851:{35,35}]
  wire  _GEN_5113 = 5'h2 == redirectHeadVec_0_value ? 1'h0 : valid_2; // @[Rob.scala 426:22 851:{35,35}]
  wire  _GEN_5114 = 5'h3 == redirectHeadVec_0_value ? 1'h0 : valid_3; // @[Rob.scala 426:22 851:{35,35}]
  wire  _GEN_5115 = 5'h4 == redirectHeadVec_0_value ? 1'h0 : valid_4; // @[Rob.scala 426:22 851:{35,35}]
  wire  _GEN_5116 = 5'h5 == redirectHeadVec_0_value ? 1'h0 : valid_5; // @[Rob.scala 426:22 851:{35,35}]
  wire  _GEN_5117 = 5'h6 == redirectHeadVec_0_value ? 1'h0 : valid_6; // @[Rob.scala 426:22 851:{35,35}]
  wire  _GEN_5118 = 5'h7 == redirectHeadVec_0_value ? 1'h0 : valid_7; // @[Rob.scala 426:22 851:{35,35}]
  wire  _GEN_5119 = 5'h8 == redirectHeadVec_0_value ? 1'h0 : valid_8; // @[Rob.scala 426:22 851:{35,35}]
  wire  _GEN_5120 = 5'h9 == redirectHeadVec_0_value ? 1'h0 : valid_9; // @[Rob.scala 426:22 851:{35,35}]
  wire  _GEN_5121 = 5'ha == redirectHeadVec_0_value ? 1'h0 : valid_10; // @[Rob.scala 426:22 851:{35,35}]
  wire  _GEN_5122 = 5'hb == redirectHeadVec_0_value ? 1'h0 : valid_11; // @[Rob.scala 426:22 851:{35,35}]
  wire  _GEN_5123 = 5'hc == redirectHeadVec_0_value ? 1'h0 : valid_12; // @[Rob.scala 426:22 851:{35,35}]
  wire  _GEN_5124 = 5'hd == redirectHeadVec_0_value ? 1'h0 : valid_13; // @[Rob.scala 426:22 851:{35,35}]
  wire  _GEN_5125 = 5'he == redirectHeadVec_0_value ? 1'h0 : valid_14; // @[Rob.scala 426:22 851:{35,35}]
  wire  _GEN_5126 = 5'hf == redirectHeadVec_0_value ? 1'h0 : valid_15; // @[Rob.scala 426:22 851:{35,35}]
  wire  _GEN_5127 = 5'h10 == redirectHeadVec_0_value ? 1'h0 : valid_16; // @[Rob.scala 426:22 851:{35,35}]
  wire  _GEN_5128 = 5'h11 == redirectHeadVec_0_value ? 1'h0 : valid_17; // @[Rob.scala 426:22 851:{35,35}]
  wire  _GEN_5129 = 5'h12 == redirectHeadVec_0_value ? 1'h0 : valid_18; // @[Rob.scala 426:22 851:{35,35}]
  wire  _GEN_5130 = 5'h13 == redirectHeadVec_0_value ? 1'h0 : valid_19; // @[Rob.scala 426:22 851:{35,35}]
  wire  _GEN_5131 = 5'h14 == redirectHeadVec_0_value ? 1'h0 : valid_20; // @[Rob.scala 426:22 851:{35,35}]
  wire  _GEN_5132 = 5'h15 == redirectHeadVec_0_value ? 1'h0 : valid_21; // @[Rob.scala 426:22 851:{35,35}]
  wire  _GEN_5133 = 5'h16 == redirectHeadVec_0_value ? 1'h0 : valid_22; // @[Rob.scala 426:22 851:{35,35}]
  wire  _GEN_5134 = 5'h17 == redirectHeadVec_0_value ? 1'h0 : valid_23; // @[Rob.scala 426:22 851:{35,35}]
  wire  _GEN_5135 = 5'h18 == redirectHeadVec_0_value ? 1'h0 : valid_24; // @[Rob.scala 426:22 851:{35,35}]
  wire  _GEN_5136 = 5'h19 == redirectHeadVec_0_value ? 1'h0 : valid_25; // @[Rob.scala 426:22 851:{35,35}]
  wire  _GEN_5137 = 5'h1a == redirectHeadVec_0_value ? 1'h0 : valid_26; // @[Rob.scala 426:22 851:{35,35}]
  wire  _GEN_5138 = 5'h1b == redirectHeadVec_0_value ? 1'h0 : valid_27; // @[Rob.scala 426:22 851:{35,35}]
  wire  _GEN_5139 = 5'h1c == redirectHeadVec_0_value ? 1'h0 : valid_28; // @[Rob.scala 426:22 851:{35,35}]
  wire  _GEN_5140 = 5'h1d == redirectHeadVec_0_value ? 1'h0 : valid_29; // @[Rob.scala 426:22 851:{35,35}]
  wire  _GEN_5141 = 5'h1e == redirectHeadVec_0_value ? 1'h0 : valid_30; // @[Rob.scala 426:22 851:{35,35}]
  wire  _GEN_5142 = 5'h1f == redirectHeadVec_0_value ? 1'h0 : valid_31; // @[Rob.scala 426:22 851:{35,35}]
  wire  _GEN_5143 = invMask_0 ? _GEN_5111 : valid_0; // @[Rob.scala 426:22 850:45]
  wire  _GEN_5144 = invMask_0 ? _GEN_5112 : valid_1; // @[Rob.scala 426:22 850:45]
  wire  _GEN_5145 = invMask_0 ? _GEN_5113 : valid_2; // @[Rob.scala 426:22 850:45]
  wire  _GEN_5146 = invMask_0 ? _GEN_5114 : valid_3; // @[Rob.scala 426:22 850:45]
  wire  _GEN_5147 = invMask_0 ? _GEN_5115 : valid_4; // @[Rob.scala 426:22 850:45]
  wire  _GEN_5148 = invMask_0 ? _GEN_5116 : valid_5; // @[Rob.scala 426:22 850:45]
  wire  _GEN_5149 = invMask_0 ? _GEN_5117 : valid_6; // @[Rob.scala 426:22 850:45]
  wire  _GEN_5150 = invMask_0 ? _GEN_5118 : valid_7; // @[Rob.scala 426:22 850:45]
  wire  _GEN_5151 = invMask_0 ? _GEN_5119 : valid_8; // @[Rob.scala 426:22 850:45]
  wire  _GEN_5152 = invMask_0 ? _GEN_5120 : valid_9; // @[Rob.scala 426:22 850:45]
  wire  _GEN_5153 = invMask_0 ? _GEN_5121 : valid_10; // @[Rob.scala 426:22 850:45]
  wire  _GEN_5154 = invMask_0 ? _GEN_5122 : valid_11; // @[Rob.scala 426:22 850:45]
  wire  _GEN_5155 = invMask_0 ? _GEN_5123 : valid_12; // @[Rob.scala 426:22 850:45]
  wire  _GEN_5156 = invMask_0 ? _GEN_5124 : valid_13; // @[Rob.scala 426:22 850:45]
  wire  _GEN_5157 = invMask_0 ? _GEN_5125 : valid_14; // @[Rob.scala 426:22 850:45]
  wire  _GEN_5158 = invMask_0 ? _GEN_5126 : valid_15; // @[Rob.scala 426:22 850:45]
  wire  _GEN_5159 = invMask_0 ? _GEN_5127 : valid_16; // @[Rob.scala 426:22 850:45]
  wire  _GEN_5160 = invMask_0 ? _GEN_5128 : valid_17; // @[Rob.scala 426:22 850:45]
  wire  _GEN_5161 = invMask_0 ? _GEN_5129 : valid_18; // @[Rob.scala 426:22 850:45]
  wire  _GEN_5162 = invMask_0 ? _GEN_5130 : valid_19; // @[Rob.scala 426:22 850:45]
  wire  _GEN_5163 = invMask_0 ? _GEN_5131 : valid_20; // @[Rob.scala 426:22 850:45]
  wire  _GEN_5164 = invMask_0 ? _GEN_5132 : valid_21; // @[Rob.scala 426:22 850:45]
  wire  _GEN_5165 = invMask_0 ? _GEN_5133 : valid_22; // @[Rob.scala 426:22 850:45]
  wire  _GEN_5166 = invMask_0 ? _GEN_5134 : valid_23; // @[Rob.scala 426:22 850:45]
  wire  _GEN_5167 = invMask_0 ? _GEN_5135 : valid_24; // @[Rob.scala 426:22 850:45]
  wire  _GEN_5168 = invMask_0 ? _GEN_5136 : valid_25; // @[Rob.scala 426:22 850:45]
  wire  _GEN_5169 = invMask_0 ? _GEN_5137 : valid_26; // @[Rob.scala 426:22 850:45]
  wire  _GEN_5170 = invMask_0 ? _GEN_5138 : valid_27; // @[Rob.scala 426:22 850:45]
  wire  _GEN_5171 = invMask_0 ? _GEN_5139 : valid_28; // @[Rob.scala 426:22 850:45]
  wire  _GEN_5172 = invMask_0 ? _GEN_5140 : valid_29; // @[Rob.scala 426:22 850:45]
  wire  _GEN_5173 = invMask_0 ? _GEN_5141 : valid_30; // @[Rob.scala 426:22 850:45]
  wire  _GEN_5174 = invMask_0 ? _GEN_5142 : valid_31; // @[Rob.scala 426:22 850:45]
  wire  _GEN_5175 = 5'h0 == redirectHeadVec_1_value ? 1'h0 : _GEN_5143; // @[Rob.scala 851:{35,35}]
  wire  _GEN_5176 = 5'h1 == redirectHeadVec_1_value ? 1'h0 : _GEN_5144; // @[Rob.scala 851:{35,35}]
  wire  _GEN_5177 = 5'h2 == redirectHeadVec_1_value ? 1'h0 : _GEN_5145; // @[Rob.scala 851:{35,35}]
  wire  _GEN_5178 = 5'h3 == redirectHeadVec_1_value ? 1'h0 : _GEN_5146; // @[Rob.scala 851:{35,35}]
  wire  _GEN_5179 = 5'h4 == redirectHeadVec_1_value ? 1'h0 : _GEN_5147; // @[Rob.scala 851:{35,35}]
  wire  _GEN_5180 = 5'h5 == redirectHeadVec_1_value ? 1'h0 : _GEN_5148; // @[Rob.scala 851:{35,35}]
  wire  _GEN_5181 = 5'h6 == redirectHeadVec_1_value ? 1'h0 : _GEN_5149; // @[Rob.scala 851:{35,35}]
  wire  _GEN_5182 = 5'h7 == redirectHeadVec_1_value ? 1'h0 : _GEN_5150; // @[Rob.scala 851:{35,35}]
  wire  _GEN_5183 = 5'h8 == redirectHeadVec_1_value ? 1'h0 : _GEN_5151; // @[Rob.scala 851:{35,35}]
  wire  _GEN_5184 = 5'h9 == redirectHeadVec_1_value ? 1'h0 : _GEN_5152; // @[Rob.scala 851:{35,35}]
  wire  _GEN_5185 = 5'ha == redirectHeadVec_1_value ? 1'h0 : _GEN_5153; // @[Rob.scala 851:{35,35}]
  wire  _GEN_5186 = 5'hb == redirectHeadVec_1_value ? 1'h0 : _GEN_5154; // @[Rob.scala 851:{35,35}]
  wire  _GEN_5187 = 5'hc == redirectHeadVec_1_value ? 1'h0 : _GEN_5155; // @[Rob.scala 851:{35,35}]
  wire  _GEN_5188 = 5'hd == redirectHeadVec_1_value ? 1'h0 : _GEN_5156; // @[Rob.scala 851:{35,35}]
  wire  _GEN_5189 = 5'he == redirectHeadVec_1_value ? 1'h0 : _GEN_5157; // @[Rob.scala 851:{35,35}]
  wire  _GEN_5190 = 5'hf == redirectHeadVec_1_value ? 1'h0 : _GEN_5158; // @[Rob.scala 851:{35,35}]
  wire  _GEN_5191 = 5'h10 == redirectHeadVec_1_value ? 1'h0 : _GEN_5159; // @[Rob.scala 851:{35,35}]
  wire  _GEN_5192 = 5'h11 == redirectHeadVec_1_value ? 1'h0 : _GEN_5160; // @[Rob.scala 851:{35,35}]
  wire  _GEN_5193 = 5'h12 == redirectHeadVec_1_value ? 1'h0 : _GEN_5161; // @[Rob.scala 851:{35,35}]
  wire  _GEN_5194 = 5'h13 == redirectHeadVec_1_value ? 1'h0 : _GEN_5162; // @[Rob.scala 851:{35,35}]
  wire  _GEN_5195 = 5'h14 == redirectHeadVec_1_value ? 1'h0 : _GEN_5163; // @[Rob.scala 851:{35,35}]
  wire  _GEN_5196 = 5'h15 == redirectHeadVec_1_value ? 1'h0 : _GEN_5164; // @[Rob.scala 851:{35,35}]
  wire  _GEN_5197 = 5'h16 == redirectHeadVec_1_value ? 1'h0 : _GEN_5165; // @[Rob.scala 851:{35,35}]
  wire  _GEN_5198 = 5'h17 == redirectHeadVec_1_value ? 1'h0 : _GEN_5166; // @[Rob.scala 851:{35,35}]
  wire  _GEN_5199 = 5'h18 == redirectHeadVec_1_value ? 1'h0 : _GEN_5167; // @[Rob.scala 851:{35,35}]
  wire  _GEN_5200 = 5'h19 == redirectHeadVec_1_value ? 1'h0 : _GEN_5168; // @[Rob.scala 851:{35,35}]
  wire  _GEN_5201 = 5'h1a == redirectHeadVec_1_value ? 1'h0 : _GEN_5169; // @[Rob.scala 851:{35,35}]
  wire  _GEN_5202 = 5'h1b == redirectHeadVec_1_value ? 1'h0 : _GEN_5170; // @[Rob.scala 851:{35,35}]
  wire  _GEN_5203 = 5'h1c == redirectHeadVec_1_value ? 1'h0 : _GEN_5171; // @[Rob.scala 851:{35,35}]
  wire  _GEN_5204 = 5'h1d == redirectHeadVec_1_value ? 1'h0 : _GEN_5172; // @[Rob.scala 851:{35,35}]
  wire  _GEN_5205 = 5'h1e == redirectHeadVec_1_value ? 1'h0 : _GEN_5173; // @[Rob.scala 851:{35,35}]
  wire  _GEN_5206 = 5'h1f == redirectHeadVec_1_value ? 1'h0 : _GEN_5174; // @[Rob.scala 851:{35,35}]
  wire  _GEN_5207 = invMask_1 ? _GEN_5175 : _GEN_5143; // @[Rob.scala 850:45]
  wire  _GEN_5208 = invMask_1 ? _GEN_5176 : _GEN_5144; // @[Rob.scala 850:45]
  wire  _GEN_5209 = invMask_1 ? _GEN_5177 : _GEN_5145; // @[Rob.scala 850:45]
  wire  _GEN_5210 = invMask_1 ? _GEN_5178 : _GEN_5146; // @[Rob.scala 850:45]
  wire  _GEN_5211 = invMask_1 ? _GEN_5179 : _GEN_5147; // @[Rob.scala 850:45]
  wire  _GEN_5212 = invMask_1 ? _GEN_5180 : _GEN_5148; // @[Rob.scala 850:45]
  wire  _GEN_5213 = invMask_1 ? _GEN_5181 : _GEN_5149; // @[Rob.scala 850:45]
  wire  _GEN_5214 = invMask_1 ? _GEN_5182 : _GEN_5150; // @[Rob.scala 850:45]
  wire  _GEN_5215 = invMask_1 ? _GEN_5183 : _GEN_5151; // @[Rob.scala 850:45]
  wire  _GEN_5216 = invMask_1 ? _GEN_5184 : _GEN_5152; // @[Rob.scala 850:45]
  wire  _GEN_5217 = invMask_1 ? _GEN_5185 : _GEN_5153; // @[Rob.scala 850:45]
  wire  _GEN_5218 = invMask_1 ? _GEN_5186 : _GEN_5154; // @[Rob.scala 850:45]
  wire  _GEN_5219 = invMask_1 ? _GEN_5187 : _GEN_5155; // @[Rob.scala 850:45]
  wire  _GEN_5220 = invMask_1 ? _GEN_5188 : _GEN_5156; // @[Rob.scala 850:45]
  wire  _GEN_5221 = invMask_1 ? _GEN_5189 : _GEN_5157; // @[Rob.scala 850:45]
  wire  _GEN_5222 = invMask_1 ? _GEN_5190 : _GEN_5158; // @[Rob.scala 850:45]
  wire  _GEN_5223 = invMask_1 ? _GEN_5191 : _GEN_5159; // @[Rob.scala 850:45]
  wire  _GEN_5224 = invMask_1 ? _GEN_5192 : _GEN_5160; // @[Rob.scala 850:45]
  wire  _GEN_5225 = invMask_1 ? _GEN_5193 : _GEN_5161; // @[Rob.scala 850:45]
  wire  _GEN_5226 = invMask_1 ? _GEN_5194 : _GEN_5162; // @[Rob.scala 850:45]
  wire  _GEN_5227 = invMask_1 ? _GEN_5195 : _GEN_5163; // @[Rob.scala 850:45]
  wire  _GEN_5228 = invMask_1 ? _GEN_5196 : _GEN_5164; // @[Rob.scala 850:45]
  wire  _GEN_5229 = invMask_1 ? _GEN_5197 : _GEN_5165; // @[Rob.scala 850:45]
  wire  _GEN_5230 = invMask_1 ? _GEN_5198 : _GEN_5166; // @[Rob.scala 850:45]
  wire  _GEN_5231 = invMask_1 ? _GEN_5199 : _GEN_5167; // @[Rob.scala 850:45]
  wire  _GEN_5232 = invMask_1 ? _GEN_5200 : _GEN_5168; // @[Rob.scala 850:45]
  wire  _GEN_5233 = invMask_1 ? _GEN_5201 : _GEN_5169; // @[Rob.scala 850:45]
  wire  _GEN_5234 = invMask_1 ? _GEN_5202 : _GEN_5170; // @[Rob.scala 850:45]
  wire  _GEN_5235 = invMask_1 ? _GEN_5203 : _GEN_5171; // @[Rob.scala 850:45]
  wire  _GEN_5236 = invMask_1 ? _GEN_5204 : _GEN_5172; // @[Rob.scala 850:45]
  wire  _GEN_5237 = invMask_1 ? _GEN_5205 : _GEN_5173; // @[Rob.scala 850:45]
  wire  _GEN_5238 = invMask_1 ? _GEN_5206 : _GEN_5174; // @[Rob.scala 850:45]
  wire  _GEN_5239 = ~invMask_1 ? 1'h0 : redirectState; // @[Rob.scala 854:25 855:21 845:30]
  wire  _GEN_5244 = redirectState ? _GEN_5207 : valid_0; // @[Rob.scala 426:22 847:40]
  wire  _GEN_5245 = redirectState ? _GEN_5208 : valid_1; // @[Rob.scala 426:22 847:40]
  wire  _GEN_5246 = redirectState ? _GEN_5209 : valid_2; // @[Rob.scala 426:22 847:40]
  wire  _GEN_5247 = redirectState ? _GEN_5210 : valid_3; // @[Rob.scala 426:22 847:40]
  wire  _GEN_5248 = redirectState ? _GEN_5211 : valid_4; // @[Rob.scala 426:22 847:40]
  wire  _GEN_5249 = redirectState ? _GEN_5212 : valid_5; // @[Rob.scala 426:22 847:40]
  wire  _GEN_5250 = redirectState ? _GEN_5213 : valid_6; // @[Rob.scala 426:22 847:40]
  wire  _GEN_5251 = redirectState ? _GEN_5214 : valid_7; // @[Rob.scala 426:22 847:40]
  wire  _GEN_5252 = redirectState ? _GEN_5215 : valid_8; // @[Rob.scala 426:22 847:40]
  wire  _GEN_5253 = redirectState ? _GEN_5216 : valid_9; // @[Rob.scala 426:22 847:40]
  wire  _GEN_5254 = redirectState ? _GEN_5217 : valid_10; // @[Rob.scala 426:22 847:40]
  wire  _GEN_5255 = redirectState ? _GEN_5218 : valid_11; // @[Rob.scala 426:22 847:40]
  wire  _GEN_5256 = redirectState ? _GEN_5219 : valid_12; // @[Rob.scala 426:22 847:40]
  wire  _GEN_5257 = redirectState ? _GEN_5220 : valid_13; // @[Rob.scala 426:22 847:40]
  wire  _GEN_5258 = redirectState ? _GEN_5221 : valid_14; // @[Rob.scala 426:22 847:40]
  wire  _GEN_5259 = redirectState ? _GEN_5222 : valid_15; // @[Rob.scala 426:22 847:40]
  wire  _GEN_5260 = redirectState ? _GEN_5223 : valid_16; // @[Rob.scala 426:22 847:40]
  wire  _GEN_5261 = redirectState ? _GEN_5224 : valid_17; // @[Rob.scala 426:22 847:40]
  wire  _GEN_5262 = redirectState ? _GEN_5225 : valid_18; // @[Rob.scala 426:22 847:40]
  wire  _GEN_5263 = redirectState ? _GEN_5226 : valid_19; // @[Rob.scala 426:22 847:40]
  wire  _GEN_5264 = redirectState ? _GEN_5227 : valid_20; // @[Rob.scala 426:22 847:40]
  wire  _GEN_5265 = redirectState ? _GEN_5228 : valid_21; // @[Rob.scala 426:22 847:40]
  wire  _GEN_5266 = redirectState ? _GEN_5229 : valid_22; // @[Rob.scala 426:22 847:40]
  wire  _GEN_5267 = redirectState ? _GEN_5230 : valid_23; // @[Rob.scala 426:22 847:40]
  wire  _GEN_5268 = redirectState ? _GEN_5231 : valid_24; // @[Rob.scala 426:22 847:40]
  wire  _GEN_5269 = redirectState ? _GEN_5232 : valid_25; // @[Rob.scala 426:22 847:40]
  wire  _GEN_5270 = redirectState ? _GEN_5233 : valid_26; // @[Rob.scala 426:22 847:40]
  wire  _GEN_5271 = redirectState ? _GEN_5234 : valid_27; // @[Rob.scala 426:22 847:40]
  wire  _GEN_5272 = redirectState ? _GEN_5235 : valid_28; // @[Rob.scala 426:22 847:40]
  wire  _GEN_5273 = redirectState ? _GEN_5236 : valid_29; // @[Rob.scala 426:22 847:40]
  wire  _GEN_5274 = redirectState ? _GEN_5237 : valid_30; // @[Rob.scala 426:22 847:40]
  wire  _GEN_5275 = redirectState ? _GEN_5238 : valid_31; // @[Rob.scala 426:22 847:40]
  wire  _GEN_5276 = redirectState ? _GEN_5239 : redirectState; // @[Rob.scala 845:30 847:40]
  wire [5:0] _redirectHeadVec_0_new_ptr_T_5 = {io_redirect_bits_robIdx_flag,io_redirect_bits_robIdx_value}; // @[Cat.scala 31:58]
  wire [6:0] _redirectHeadVec_0_new_ptr_T_6 = {{1'd0}, _redirectHeadVec_0_new_ptr_T_5}; // @[CircularQueuePtr.scala 39:46]
  wire [4:0] redirectHeadVec_0_new_ptr_1_value = _redirectHeadVec_0_new_ptr_T_6[4:0]; // @[CircularQueuePtr.scala 39:59]
  wire  redirectHeadVec_0_new_ptr_1_flag = _redirectHeadVec_0_new_ptr_T_6[5]; // @[CircularQueuePtr.scala 39:59]
  wire [5:0] _redirectHeadVec_0_new_ptr_T_12 = _redirectHeadVec_0_new_ptr_T_5 + 6'h1; // @[CircularQueuePtr.scala 39:46]
  wire [4:0] redirectHeadVec_0_new_ptr_2_value = _redirectHeadVec_0_new_ptr_T_12[4:0]; // @[CircularQueuePtr.scala 39:59]
  wire  redirectHeadVec_0_new_ptr_2_flag = _redirectHeadVec_0_new_ptr_T_12[5]; // @[CircularQueuePtr.scala 39:59]
  wire [5:0] _redirectHeadVec_1_new_ptr_T_12 = _redirectHeadVec_0_new_ptr_T_5 + 6'h2; // @[CircularQueuePtr.scala 39:46]
  wire [4:0] redirectHeadVec_1_new_ptr_2_value = _redirectHeadVec_1_new_ptr_T_12[4:0]; // @[CircularQueuePtr.scala 39:59]
  wire  redirectHeadVec_1_new_ptr_2_flag = _redirectHeadVec_1_new_ptr_T_12[5]; // @[CircularQueuePtr.scala 39:59]
  wire  _GEN_5286 = 5'h0 == enqPtrVec_0_value | _GEN_5244; // @[Rob.scala 870:{38,38}]
  wire  _GEN_5287 = 5'h1 == enqPtrVec_0_value | _GEN_5245; // @[Rob.scala 870:{38,38}]
  wire  _GEN_5288 = 5'h2 == enqPtrVec_0_value | _GEN_5246; // @[Rob.scala 870:{38,38}]
  wire  _GEN_5289 = 5'h3 == enqPtrVec_0_value | _GEN_5247; // @[Rob.scala 870:{38,38}]
  wire  _GEN_5290 = 5'h4 == enqPtrVec_0_value | _GEN_5248; // @[Rob.scala 870:{38,38}]
  wire  _GEN_5291 = 5'h5 == enqPtrVec_0_value | _GEN_5249; // @[Rob.scala 870:{38,38}]
  wire  _GEN_5292 = 5'h6 == enqPtrVec_0_value | _GEN_5250; // @[Rob.scala 870:{38,38}]
  wire  _GEN_5293 = 5'h7 == enqPtrVec_0_value | _GEN_5251; // @[Rob.scala 870:{38,38}]
  wire  _GEN_5294 = 5'h8 == enqPtrVec_0_value | _GEN_5252; // @[Rob.scala 870:{38,38}]
  wire  _GEN_5295 = 5'h9 == enqPtrVec_0_value | _GEN_5253; // @[Rob.scala 870:{38,38}]
  wire  _GEN_5296 = 5'ha == enqPtrVec_0_value | _GEN_5254; // @[Rob.scala 870:{38,38}]
  wire  _GEN_5297 = 5'hb == enqPtrVec_0_value | _GEN_5255; // @[Rob.scala 870:{38,38}]
  wire  _GEN_5298 = 5'hc == enqPtrVec_0_value | _GEN_5256; // @[Rob.scala 870:{38,38}]
  wire  _GEN_5299 = 5'hd == enqPtrVec_0_value | _GEN_5257; // @[Rob.scala 870:{38,38}]
  wire  _GEN_5300 = 5'he == enqPtrVec_0_value | _GEN_5258; // @[Rob.scala 870:{38,38}]
  wire  _GEN_5301 = 5'hf == enqPtrVec_0_value | _GEN_5259; // @[Rob.scala 870:{38,38}]
  wire  _GEN_5302 = 5'h10 == enqPtrVec_0_value | _GEN_5260; // @[Rob.scala 870:{38,38}]
  wire  _GEN_5303 = 5'h11 == enqPtrVec_0_value | _GEN_5261; // @[Rob.scala 870:{38,38}]
  wire  _GEN_5304 = 5'h12 == enqPtrVec_0_value | _GEN_5262; // @[Rob.scala 870:{38,38}]
  wire  _GEN_5305 = 5'h13 == enqPtrVec_0_value | _GEN_5263; // @[Rob.scala 870:{38,38}]
  wire  _GEN_5306 = 5'h14 == enqPtrVec_0_value | _GEN_5264; // @[Rob.scala 870:{38,38}]
  wire  _GEN_5307 = 5'h15 == enqPtrVec_0_value | _GEN_5265; // @[Rob.scala 870:{38,38}]
  wire  _GEN_5308 = 5'h16 == enqPtrVec_0_value | _GEN_5266; // @[Rob.scala 870:{38,38}]
  wire  _GEN_5309 = 5'h17 == enqPtrVec_0_value | _GEN_5267; // @[Rob.scala 870:{38,38}]
  wire  _GEN_5310 = 5'h18 == enqPtrVec_0_value | _GEN_5268; // @[Rob.scala 870:{38,38}]
  wire  _GEN_5311 = 5'h19 == enqPtrVec_0_value | _GEN_5269; // @[Rob.scala 870:{38,38}]
  wire  _GEN_5312 = 5'h1a == enqPtrVec_0_value | _GEN_5270; // @[Rob.scala 870:{38,38}]
  wire  _GEN_5313 = 5'h1b == enqPtrVec_0_value | _GEN_5271; // @[Rob.scala 870:{38,38}]
  wire  _GEN_5314 = 5'h1c == enqPtrVec_0_value | _GEN_5272; // @[Rob.scala 870:{38,38}]
  wire  _GEN_5315 = 5'h1d == enqPtrVec_0_value | _GEN_5273; // @[Rob.scala 870:{38,38}]
  wire  _GEN_5316 = 5'h1e == enqPtrVec_0_value | _GEN_5274; // @[Rob.scala 870:{38,38}]
  wire  _GEN_5317 = 5'h1f == enqPtrVec_0_value | _GEN_5275; // @[Rob.scala 870:{38,38}]
  wire  _GEN_5318 = canEnqueue_0 & ~io_redirect_valid ? _GEN_5286 : _GEN_5244; // @[Rob.scala 869:48]
  wire  _GEN_5319 = canEnqueue_0 & ~io_redirect_valid ? _GEN_5287 : _GEN_5245; // @[Rob.scala 869:48]
  wire  _GEN_5320 = canEnqueue_0 & ~io_redirect_valid ? _GEN_5288 : _GEN_5246; // @[Rob.scala 869:48]
  wire  _GEN_5321 = canEnqueue_0 & ~io_redirect_valid ? _GEN_5289 : _GEN_5247; // @[Rob.scala 869:48]
  wire  _GEN_5322 = canEnqueue_0 & ~io_redirect_valid ? _GEN_5290 : _GEN_5248; // @[Rob.scala 869:48]
  wire  _GEN_5323 = canEnqueue_0 & ~io_redirect_valid ? _GEN_5291 : _GEN_5249; // @[Rob.scala 869:48]
  wire  _GEN_5324 = canEnqueue_0 & ~io_redirect_valid ? _GEN_5292 : _GEN_5250; // @[Rob.scala 869:48]
  wire  _GEN_5325 = canEnqueue_0 & ~io_redirect_valid ? _GEN_5293 : _GEN_5251; // @[Rob.scala 869:48]
  wire  _GEN_5326 = canEnqueue_0 & ~io_redirect_valid ? _GEN_5294 : _GEN_5252; // @[Rob.scala 869:48]
  wire  _GEN_5327 = canEnqueue_0 & ~io_redirect_valid ? _GEN_5295 : _GEN_5253; // @[Rob.scala 869:48]
  wire  _GEN_5328 = canEnqueue_0 & ~io_redirect_valid ? _GEN_5296 : _GEN_5254; // @[Rob.scala 869:48]
  wire  _GEN_5329 = canEnqueue_0 & ~io_redirect_valid ? _GEN_5297 : _GEN_5255; // @[Rob.scala 869:48]
  wire  _GEN_5330 = canEnqueue_0 & ~io_redirect_valid ? _GEN_5298 : _GEN_5256; // @[Rob.scala 869:48]
  wire  _GEN_5331 = canEnqueue_0 & ~io_redirect_valid ? _GEN_5299 : _GEN_5257; // @[Rob.scala 869:48]
  wire  _GEN_5332 = canEnqueue_0 & ~io_redirect_valid ? _GEN_5300 : _GEN_5258; // @[Rob.scala 869:48]
  wire  _GEN_5333 = canEnqueue_0 & ~io_redirect_valid ? _GEN_5301 : _GEN_5259; // @[Rob.scala 869:48]
  wire  _GEN_5334 = canEnqueue_0 & ~io_redirect_valid ? _GEN_5302 : _GEN_5260; // @[Rob.scala 869:48]
  wire  _GEN_5335 = canEnqueue_0 & ~io_redirect_valid ? _GEN_5303 : _GEN_5261; // @[Rob.scala 869:48]
  wire  _GEN_5336 = canEnqueue_0 & ~io_redirect_valid ? _GEN_5304 : _GEN_5262; // @[Rob.scala 869:48]
  wire  _GEN_5337 = canEnqueue_0 & ~io_redirect_valid ? _GEN_5305 : _GEN_5263; // @[Rob.scala 869:48]
  wire  _GEN_5338 = canEnqueue_0 & ~io_redirect_valid ? _GEN_5306 : _GEN_5264; // @[Rob.scala 869:48]
  wire  _GEN_5339 = canEnqueue_0 & ~io_redirect_valid ? _GEN_5307 : _GEN_5265; // @[Rob.scala 869:48]
  wire  _GEN_5340 = canEnqueue_0 & ~io_redirect_valid ? _GEN_5308 : _GEN_5266; // @[Rob.scala 869:48]
  wire  _GEN_5341 = canEnqueue_0 & ~io_redirect_valid ? _GEN_5309 : _GEN_5267; // @[Rob.scala 869:48]
  wire  _GEN_5342 = canEnqueue_0 & ~io_redirect_valid ? _GEN_5310 : _GEN_5268; // @[Rob.scala 869:48]
  wire  _GEN_5343 = canEnqueue_0 & ~io_redirect_valid ? _GEN_5311 : _GEN_5269; // @[Rob.scala 869:48]
  wire  _GEN_5344 = canEnqueue_0 & ~io_redirect_valid ? _GEN_5312 : _GEN_5270; // @[Rob.scala 869:48]
  wire  _GEN_5345 = canEnqueue_0 & ~io_redirect_valid ? _GEN_5313 : _GEN_5271; // @[Rob.scala 869:48]
  wire  _GEN_5346 = canEnqueue_0 & ~io_redirect_valid ? _GEN_5314 : _GEN_5272; // @[Rob.scala 869:48]
  wire  _GEN_5347 = canEnqueue_0 & ~io_redirect_valid ? _GEN_5315 : _GEN_5273; // @[Rob.scala 869:48]
  wire  _GEN_5348 = canEnqueue_0 & ~io_redirect_valid ? _GEN_5316 : _GEN_5274; // @[Rob.scala 869:48]
  wire  _GEN_5349 = canEnqueue_0 & ~io_redirect_valid ? _GEN_5317 : _GEN_5275; // @[Rob.scala 869:48]
  wire  _GEN_5350 = 5'h0 == allocatePtrVec_1_value | _GEN_5318; // @[Rob.scala 870:{38,38}]
  wire  _GEN_5351 = 5'h1 == allocatePtrVec_1_value | _GEN_5319; // @[Rob.scala 870:{38,38}]
  wire  _GEN_5352 = 5'h2 == allocatePtrVec_1_value | _GEN_5320; // @[Rob.scala 870:{38,38}]
  wire  _GEN_5353 = 5'h3 == allocatePtrVec_1_value | _GEN_5321; // @[Rob.scala 870:{38,38}]
  wire  _GEN_5354 = 5'h4 == allocatePtrVec_1_value | _GEN_5322; // @[Rob.scala 870:{38,38}]
  wire  _GEN_5355 = 5'h5 == allocatePtrVec_1_value | _GEN_5323; // @[Rob.scala 870:{38,38}]
  wire  _GEN_5356 = 5'h6 == allocatePtrVec_1_value | _GEN_5324; // @[Rob.scala 870:{38,38}]
  wire  _GEN_5357 = 5'h7 == allocatePtrVec_1_value | _GEN_5325; // @[Rob.scala 870:{38,38}]
  wire  _GEN_5358 = 5'h8 == allocatePtrVec_1_value | _GEN_5326; // @[Rob.scala 870:{38,38}]
  wire  _GEN_5359 = 5'h9 == allocatePtrVec_1_value | _GEN_5327; // @[Rob.scala 870:{38,38}]
  wire  _GEN_5360 = 5'ha == allocatePtrVec_1_value | _GEN_5328; // @[Rob.scala 870:{38,38}]
  wire  _GEN_5361 = 5'hb == allocatePtrVec_1_value | _GEN_5329; // @[Rob.scala 870:{38,38}]
  wire  _GEN_5362 = 5'hc == allocatePtrVec_1_value | _GEN_5330; // @[Rob.scala 870:{38,38}]
  wire  _GEN_5363 = 5'hd == allocatePtrVec_1_value | _GEN_5331; // @[Rob.scala 870:{38,38}]
  wire  _GEN_5364 = 5'he == allocatePtrVec_1_value | _GEN_5332; // @[Rob.scala 870:{38,38}]
  wire  _GEN_5365 = 5'hf == allocatePtrVec_1_value | _GEN_5333; // @[Rob.scala 870:{38,38}]
  wire  _GEN_5366 = 5'h10 == allocatePtrVec_1_value | _GEN_5334; // @[Rob.scala 870:{38,38}]
  wire  _GEN_5367 = 5'h11 == allocatePtrVec_1_value | _GEN_5335; // @[Rob.scala 870:{38,38}]
  wire  _GEN_5368 = 5'h12 == allocatePtrVec_1_value | _GEN_5336; // @[Rob.scala 870:{38,38}]
  wire  _GEN_5369 = 5'h13 == allocatePtrVec_1_value | _GEN_5337; // @[Rob.scala 870:{38,38}]
  wire  _GEN_5370 = 5'h14 == allocatePtrVec_1_value | _GEN_5338; // @[Rob.scala 870:{38,38}]
  wire  _GEN_5371 = 5'h15 == allocatePtrVec_1_value | _GEN_5339; // @[Rob.scala 870:{38,38}]
  wire  _GEN_5372 = 5'h16 == allocatePtrVec_1_value | _GEN_5340; // @[Rob.scala 870:{38,38}]
  wire  _GEN_5373 = 5'h17 == allocatePtrVec_1_value | _GEN_5341; // @[Rob.scala 870:{38,38}]
  wire  _GEN_5374 = 5'h18 == allocatePtrVec_1_value | _GEN_5342; // @[Rob.scala 870:{38,38}]
  wire  _GEN_5375 = 5'h19 == allocatePtrVec_1_value | _GEN_5343; // @[Rob.scala 870:{38,38}]
  wire  _GEN_5376 = 5'h1a == allocatePtrVec_1_value | _GEN_5344; // @[Rob.scala 870:{38,38}]
  wire  _GEN_5377 = 5'h1b == allocatePtrVec_1_value | _GEN_5345; // @[Rob.scala 870:{38,38}]
  wire  _GEN_5378 = 5'h1c == allocatePtrVec_1_value | _GEN_5346; // @[Rob.scala 870:{38,38}]
  wire  _GEN_5379 = 5'h1d == allocatePtrVec_1_value | _GEN_5347; // @[Rob.scala 870:{38,38}]
  wire  _GEN_5380 = 5'h1e == allocatePtrVec_1_value | _GEN_5348; // @[Rob.scala 870:{38,38}]
  wire  _GEN_5381 = 5'h1f == allocatePtrVec_1_value | _GEN_5349; // @[Rob.scala 870:{38,38}]
  wire  _GEN_5382 = canEnqueue_1 & ~io_redirect_valid ? _GEN_5350 : _GEN_5318; // @[Rob.scala 869:48]
  wire  _GEN_5383 = canEnqueue_1 & ~io_redirect_valid ? _GEN_5351 : _GEN_5319; // @[Rob.scala 869:48]
  wire  _GEN_5384 = canEnqueue_1 & ~io_redirect_valid ? _GEN_5352 : _GEN_5320; // @[Rob.scala 869:48]
  wire  _GEN_5385 = canEnqueue_1 & ~io_redirect_valid ? _GEN_5353 : _GEN_5321; // @[Rob.scala 869:48]
  wire  _GEN_5386 = canEnqueue_1 & ~io_redirect_valid ? _GEN_5354 : _GEN_5322; // @[Rob.scala 869:48]
  wire  _GEN_5387 = canEnqueue_1 & ~io_redirect_valid ? _GEN_5355 : _GEN_5323; // @[Rob.scala 869:48]
  wire  _GEN_5388 = canEnqueue_1 & ~io_redirect_valid ? _GEN_5356 : _GEN_5324; // @[Rob.scala 869:48]
  wire  _GEN_5389 = canEnqueue_1 & ~io_redirect_valid ? _GEN_5357 : _GEN_5325; // @[Rob.scala 869:48]
  wire  _GEN_5390 = canEnqueue_1 & ~io_redirect_valid ? _GEN_5358 : _GEN_5326; // @[Rob.scala 869:48]
  wire  _GEN_5391 = canEnqueue_1 & ~io_redirect_valid ? _GEN_5359 : _GEN_5327; // @[Rob.scala 869:48]
  wire  _GEN_5392 = canEnqueue_1 & ~io_redirect_valid ? _GEN_5360 : _GEN_5328; // @[Rob.scala 869:48]
  wire  _GEN_5393 = canEnqueue_1 & ~io_redirect_valid ? _GEN_5361 : _GEN_5329; // @[Rob.scala 869:48]
  wire  _GEN_5394 = canEnqueue_1 & ~io_redirect_valid ? _GEN_5362 : _GEN_5330; // @[Rob.scala 869:48]
  wire  _GEN_5395 = canEnqueue_1 & ~io_redirect_valid ? _GEN_5363 : _GEN_5331; // @[Rob.scala 869:48]
  wire  _GEN_5396 = canEnqueue_1 & ~io_redirect_valid ? _GEN_5364 : _GEN_5332; // @[Rob.scala 869:48]
  wire  _GEN_5397 = canEnqueue_1 & ~io_redirect_valid ? _GEN_5365 : _GEN_5333; // @[Rob.scala 869:48]
  wire  _GEN_5398 = canEnqueue_1 & ~io_redirect_valid ? _GEN_5366 : _GEN_5334; // @[Rob.scala 869:48]
  wire  _GEN_5399 = canEnqueue_1 & ~io_redirect_valid ? _GEN_5367 : _GEN_5335; // @[Rob.scala 869:48]
  wire  _GEN_5400 = canEnqueue_1 & ~io_redirect_valid ? _GEN_5368 : _GEN_5336; // @[Rob.scala 869:48]
  wire  _GEN_5401 = canEnqueue_1 & ~io_redirect_valid ? _GEN_5369 : _GEN_5337; // @[Rob.scala 869:48]
  wire  _GEN_5402 = canEnqueue_1 & ~io_redirect_valid ? _GEN_5370 : _GEN_5338; // @[Rob.scala 869:48]
  wire  _GEN_5403 = canEnqueue_1 & ~io_redirect_valid ? _GEN_5371 : _GEN_5339; // @[Rob.scala 869:48]
  wire  _GEN_5404 = canEnqueue_1 & ~io_redirect_valid ? _GEN_5372 : _GEN_5340; // @[Rob.scala 869:48]
  wire  _GEN_5405 = canEnqueue_1 & ~io_redirect_valid ? _GEN_5373 : _GEN_5341; // @[Rob.scala 869:48]
  wire  _GEN_5406 = canEnqueue_1 & ~io_redirect_valid ? _GEN_5374 : _GEN_5342; // @[Rob.scala 869:48]
  wire  _GEN_5407 = canEnqueue_1 & ~io_redirect_valid ? _GEN_5375 : _GEN_5343; // @[Rob.scala 869:48]
  wire  _GEN_5408 = canEnqueue_1 & ~io_redirect_valid ? _GEN_5376 : _GEN_5344; // @[Rob.scala 869:48]
  wire  _GEN_5409 = canEnqueue_1 & ~io_redirect_valid ? _GEN_5377 : _GEN_5345; // @[Rob.scala 869:48]
  wire  _GEN_5410 = canEnqueue_1 & ~io_redirect_valid ? _GEN_5378 : _GEN_5346; // @[Rob.scala 869:48]
  wire  _GEN_5411 = canEnqueue_1 & ~io_redirect_valid ? _GEN_5379 : _GEN_5347; // @[Rob.scala 869:48]
  wire  _GEN_5412 = canEnqueue_1 & ~io_redirect_valid ? _GEN_5380 : _GEN_5348; // @[Rob.scala 869:48]
  wire  _GEN_5413 = canEnqueue_1 & ~io_redirect_valid ? _GEN_5381 : _GEN_5349; // @[Rob.scala 869:48]
  wire  _GEN_5414 = 5'h0 == commitReadAddr_0 ? 1'h0 : _GEN_5382; // @[Rob.scala 877:{32,32}]
  wire  _GEN_5415 = 5'h1 == commitReadAddr_0 ? 1'h0 : _GEN_5383; // @[Rob.scala 877:{32,32}]
  wire  _GEN_5416 = 5'h2 == commitReadAddr_0 ? 1'h0 : _GEN_5384; // @[Rob.scala 877:{32,32}]
  wire  _GEN_5417 = 5'h3 == commitReadAddr_0 ? 1'h0 : _GEN_5385; // @[Rob.scala 877:{32,32}]
  wire  _GEN_5418 = 5'h4 == commitReadAddr_0 ? 1'h0 : _GEN_5386; // @[Rob.scala 877:{32,32}]
  wire  _GEN_5419 = 5'h5 == commitReadAddr_0 ? 1'h0 : _GEN_5387; // @[Rob.scala 877:{32,32}]
  wire  _GEN_5420 = 5'h6 == commitReadAddr_0 ? 1'h0 : _GEN_5388; // @[Rob.scala 877:{32,32}]
  wire  _GEN_5421 = 5'h7 == commitReadAddr_0 ? 1'h0 : _GEN_5389; // @[Rob.scala 877:{32,32}]
  wire  _GEN_5422 = 5'h8 == commitReadAddr_0 ? 1'h0 : _GEN_5390; // @[Rob.scala 877:{32,32}]
  wire  _GEN_5423 = 5'h9 == commitReadAddr_0 ? 1'h0 : _GEN_5391; // @[Rob.scala 877:{32,32}]
  wire  _GEN_5424 = 5'ha == commitReadAddr_0 ? 1'h0 : _GEN_5392; // @[Rob.scala 877:{32,32}]
  wire  _GEN_5425 = 5'hb == commitReadAddr_0 ? 1'h0 : _GEN_5393; // @[Rob.scala 877:{32,32}]
  wire  _GEN_5426 = 5'hc == commitReadAddr_0 ? 1'h0 : _GEN_5394; // @[Rob.scala 877:{32,32}]
  wire  _GEN_5427 = 5'hd == commitReadAddr_0 ? 1'h0 : _GEN_5395; // @[Rob.scala 877:{32,32}]
  wire  _GEN_5428 = 5'he == commitReadAddr_0 ? 1'h0 : _GEN_5396; // @[Rob.scala 877:{32,32}]
  wire  _GEN_5429 = 5'hf == commitReadAddr_0 ? 1'h0 : _GEN_5397; // @[Rob.scala 877:{32,32}]
  wire  _GEN_5430 = 5'h10 == commitReadAddr_0 ? 1'h0 : _GEN_5398; // @[Rob.scala 877:{32,32}]
  wire  _GEN_5431 = 5'h11 == commitReadAddr_0 ? 1'h0 : _GEN_5399; // @[Rob.scala 877:{32,32}]
  wire  _GEN_5432 = 5'h12 == commitReadAddr_0 ? 1'h0 : _GEN_5400; // @[Rob.scala 877:{32,32}]
  wire  _GEN_5433 = 5'h13 == commitReadAddr_0 ? 1'h0 : _GEN_5401; // @[Rob.scala 877:{32,32}]
  wire  _GEN_5434 = 5'h14 == commitReadAddr_0 ? 1'h0 : _GEN_5402; // @[Rob.scala 877:{32,32}]
  wire  _GEN_5435 = 5'h15 == commitReadAddr_0 ? 1'h0 : _GEN_5403; // @[Rob.scala 877:{32,32}]
  wire  _GEN_5436 = 5'h16 == commitReadAddr_0 ? 1'h0 : _GEN_5404; // @[Rob.scala 877:{32,32}]
  wire  _GEN_5437 = 5'h17 == commitReadAddr_0 ? 1'h0 : _GEN_5405; // @[Rob.scala 877:{32,32}]
  wire  _GEN_5438 = 5'h18 == commitReadAddr_0 ? 1'h0 : _GEN_5406; // @[Rob.scala 877:{32,32}]
  wire  _GEN_5439 = 5'h19 == commitReadAddr_0 ? 1'h0 : _GEN_5407; // @[Rob.scala 877:{32,32}]
  wire  _GEN_5440 = 5'h1a == commitReadAddr_0 ? 1'h0 : _GEN_5408; // @[Rob.scala 877:{32,32}]
  wire  _GEN_5441 = 5'h1b == commitReadAddr_0 ? 1'h0 : _GEN_5409; // @[Rob.scala 877:{32,32}]
  wire  _GEN_5442 = 5'h1c == commitReadAddr_0 ? 1'h0 : _GEN_5410; // @[Rob.scala 877:{32,32}]
  wire  _GEN_5443 = 5'h1d == commitReadAddr_0 ? 1'h0 : _GEN_5411; // @[Rob.scala 877:{32,32}]
  wire  _GEN_5444 = 5'h1e == commitReadAddr_0 ? 1'h0 : _GEN_5412; // @[Rob.scala 877:{32,32}]
  wire  _GEN_5445 = 5'h1f == commitReadAddr_0 ? 1'h0 : _GEN_5413; // @[Rob.scala 877:{32,32}]
  wire  _GEN_5446 = _T_117 ? _GEN_5414 : _GEN_5382; // @[Rob.scala 876:24]
  wire  _GEN_5447 = _T_117 ? _GEN_5415 : _GEN_5383; // @[Rob.scala 876:24]
  wire  _GEN_5448 = _T_117 ? _GEN_5416 : _GEN_5384; // @[Rob.scala 876:24]
  wire  _GEN_5449 = _T_117 ? _GEN_5417 : _GEN_5385; // @[Rob.scala 876:24]
  wire  _GEN_5450 = _T_117 ? _GEN_5418 : _GEN_5386; // @[Rob.scala 876:24]
  wire  _GEN_5451 = _T_117 ? _GEN_5419 : _GEN_5387; // @[Rob.scala 876:24]
  wire  _GEN_5452 = _T_117 ? _GEN_5420 : _GEN_5388; // @[Rob.scala 876:24]
  wire  _GEN_5453 = _T_117 ? _GEN_5421 : _GEN_5389; // @[Rob.scala 876:24]
  wire  _GEN_5454 = _T_117 ? _GEN_5422 : _GEN_5390; // @[Rob.scala 876:24]
  wire  _GEN_5455 = _T_117 ? _GEN_5423 : _GEN_5391; // @[Rob.scala 876:24]
  wire  _GEN_5456 = _T_117 ? _GEN_5424 : _GEN_5392; // @[Rob.scala 876:24]
  wire  _GEN_5457 = _T_117 ? _GEN_5425 : _GEN_5393; // @[Rob.scala 876:24]
  wire  _GEN_5458 = _T_117 ? _GEN_5426 : _GEN_5394; // @[Rob.scala 876:24]
  wire  _GEN_5459 = _T_117 ? _GEN_5427 : _GEN_5395; // @[Rob.scala 876:24]
  wire  _GEN_5460 = _T_117 ? _GEN_5428 : _GEN_5396; // @[Rob.scala 876:24]
  wire  _GEN_5461 = _T_117 ? _GEN_5429 : _GEN_5397; // @[Rob.scala 876:24]
  wire  _GEN_5462 = _T_117 ? _GEN_5430 : _GEN_5398; // @[Rob.scala 876:24]
  wire  _GEN_5463 = _T_117 ? _GEN_5431 : _GEN_5399; // @[Rob.scala 876:24]
  wire  _GEN_5464 = _T_117 ? _GEN_5432 : _GEN_5400; // @[Rob.scala 876:24]
  wire  _GEN_5465 = _T_117 ? _GEN_5433 : _GEN_5401; // @[Rob.scala 876:24]
  wire  _GEN_5466 = _T_117 ? _GEN_5434 : _GEN_5402; // @[Rob.scala 876:24]
  wire  _GEN_5467 = _T_117 ? _GEN_5435 : _GEN_5403; // @[Rob.scala 876:24]
  wire  _GEN_5468 = _T_117 ? _GEN_5436 : _GEN_5404; // @[Rob.scala 876:24]
  wire  _GEN_5469 = _T_117 ? _GEN_5437 : _GEN_5405; // @[Rob.scala 876:24]
  wire  _GEN_5470 = _T_117 ? _GEN_5438 : _GEN_5406; // @[Rob.scala 876:24]
  wire  _GEN_5471 = _T_117 ? _GEN_5439 : _GEN_5407; // @[Rob.scala 876:24]
  wire  _GEN_5472 = _T_117 ? _GEN_5440 : _GEN_5408; // @[Rob.scala 876:24]
  wire  _GEN_5473 = _T_117 ? _GEN_5441 : _GEN_5409; // @[Rob.scala 876:24]
  wire  _GEN_5474 = _T_117 ? _GEN_5442 : _GEN_5410; // @[Rob.scala 876:24]
  wire  _GEN_5475 = _T_117 ? _GEN_5443 : _GEN_5411; // @[Rob.scala 876:24]
  wire  _GEN_5476 = _T_117 ? _GEN_5444 : _GEN_5412; // @[Rob.scala 876:24]
  wire  _GEN_5477 = _T_117 ? _GEN_5445 : _GEN_5413; // @[Rob.scala 876:24]
  wire  _T_149 = io_enq_req_0_bits_eliminatedMove & _T_12; // @[Rob.scala 894:64]
  wire  isStu = io_enq_req_0_bits_ctrl_fuType == 4'hd; // @[Rob.scala 895:50]
  wire  _T_154 = io_enq_req_1_bits_eliminatedMove & _T_51; // @[Rob.scala 894:64]
  wire  isStu_1 = io_enq_req_1_bits_ctrl_fuType == 4'hd; // @[Rob.scala 895:50]
  wire [15:0] _wbHasException_T_2 = {2'h0,io_writeback_1_2_bits_uop_cf_exceptionVec_13,1'h0,4'h0,2'h0,
    io_writeback_1_2_bits_uop_cf_exceptionVec_5,io_writeback_1_2_bits_uop_cf_exceptionVec_4,4'h0}; // @[Rob.scala 908:87]
  wire  wbHasException_2 = |_wbHasException_T_2; // @[Rob.scala 908:94]
  wire  wbHasTriggerHit_2 = io_writeback_1_2_bits_uop_cf_trigger_backendHit_0 |
    io_writeback_1_2_bits_uop_cf_trigger_backendHit_1 | io_writeback_1_2_bits_uop_cf_trigger_backendHit_2 |
    io_writeback_1_2_bits_uop_cf_trigger_backendHit_3 | io_writeback_1_2_bits_uop_cf_trigger_backendHit_4 |
    io_writeback_1_2_bits_uop_cf_trigger_backendHit_5; // @[Bundle.scala 629:43]
  wire  block_wb_2 = wbHasException_2 | io_writeback_1_2_bits_uop_ctrl_flushPipe |
    io_writeback_1_2_bits_uop_ctrl_replayInst | wbHasTriggerHit_2; // @[Rob.scala 912:74]
  wire [15:0] _wbHasException_T_3 = {2'h0,io_writeback_1_3_bits_uop_cf_exceptionVec_13,1'h0,4'h0,2'h0,
    io_writeback_1_3_bits_uop_cf_exceptionVec_5,io_writeback_1_3_bits_uop_cf_exceptionVec_4,4'h0}; // @[Rob.scala 908:87]
  wire  wbHasException_3 = |_wbHasException_T_3; // @[Rob.scala 908:94]
  wire  wbHasTriggerHit_3 = io_writeback_1_3_bits_uop_cf_trigger_backendHit_0 |
    io_writeback_1_3_bits_uop_cf_trigger_backendHit_1 | io_writeback_1_3_bits_uop_cf_trigger_backendHit_2 |
    io_writeback_1_3_bits_uop_cf_trigger_backendHit_3 | io_writeback_1_3_bits_uop_cf_trigger_backendHit_4 |
    io_writeback_1_3_bits_uop_cf_trigger_backendHit_5; // @[Bundle.scala 629:43]
  wire  block_wb_3 = wbHasException_3 | io_writeback_1_3_bits_uop_ctrl_flushPipe |
    io_writeback_1_3_bits_uop_ctrl_replayInst | wbHasTriggerHit_3; // @[Rob.scala 912:74]
  wire [15:0] _wbHasException_T_4 = {4'h0,io_writeback_1_4_bits_uop_cf_exceptionVec_11,1'h0,
    io_writeback_1_4_bits_uop_cf_exceptionVec_9,io_writeback_1_4_bits_uop_cf_exceptionVec_8,4'h0,
    io_writeback_1_4_bits_uop_cf_exceptionVec_3,io_writeback_1_4_bits_uop_cf_exceptionVec_2,2'h0}; // @[Rob.scala 908:87]
  wire  wbHasException_4 = |_wbHasException_T_4; // @[Rob.scala 908:94]
  wire  block_wb_4 = wbHasException_4 | io_writeback_1_4_bits_uop_ctrl_flushPipe; // @[Rob.scala 912:37]
  wire  wbHasTriggerHit_5 = io_writeback_1_5_bits_uop_cf_trigger_backendHit_0 |
    io_writeback_1_5_bits_uop_cf_trigger_backendHit_1 | io_writeback_1_5_bits_uop_cf_trigger_backendHit_2 |
    io_writeback_1_5_bits_uop_cf_trigger_backendHit_3 | io_writeback_1_5_bits_uop_cf_trigger_backendHit_4 |
    io_writeback_1_5_bits_uop_cf_trigger_backendHit_5; // @[Bundle.scala 629:43]
  wire [15:0] _wbHasException_T_6 = {4'h0,io_writeback_1_6_bits_uop_cf_exceptionVec_11,1'h0,
    io_writeback_1_6_bits_uop_cf_exceptionVec_9,io_writeback_1_6_bits_uop_cf_exceptionVec_8,4'h0,
    io_writeback_1_6_bits_uop_cf_exceptionVec_3,io_writeback_1_6_bits_uop_cf_exceptionVec_2,2'h0}; // @[Rob.scala 908:87]
  wire  wbHasException_6 = |_wbHasException_T_6; // @[Rob.scala 908:94]
  wire  block_wb_6 = wbHasException_6 | io_writeback_1_6_bits_uop_ctrl_flushPipe; // @[Rob.scala 912:37]
  wire [15:0] _wbHasException_T_7 = {io_writeback_1_7_bits_uop_cf_exceptionVec_15,1'h0,
    io_writeback_1_7_bits_uop_cf_exceptionVec_13,1'h0,4'h0,io_writeback_1_7_bits_uop_cf_exceptionVec_7,
    io_writeback_1_7_bits_uop_cf_exceptionVec_6,io_writeback_1_7_bits_uop_cf_exceptionVec_5,
    io_writeback_1_7_bits_uop_cf_exceptionVec_4,4'h0}; // @[Rob.scala 908:87]
  wire  wbHasException_7 = |_wbHasException_T_7; // @[Rob.scala 908:94]
  wire  wbHasTriggerHit_7 = io_writeback_1_7_bits_uop_cf_trigger_backendHit_0 |
    io_writeback_1_7_bits_uop_cf_trigger_backendHit_1 | io_writeback_1_7_bits_uop_cf_trigger_backendHit_2 |
    io_writeback_1_7_bits_uop_cf_trigger_backendHit_3 | io_writeback_1_7_bits_uop_cf_trigger_backendHit_4 |
    io_writeback_1_7_bits_uop_cf_trigger_backendHit_5; // @[Bundle.scala 629:43]
  wire  block_wb_7 = wbHasException_7 | wbHasTriggerHit_7; // @[Rob.scala 912:74]
  wire [15:0] _wbHasException_T_8 = {io_writeback_1_8_bits_uop_cf_exceptionVec_15,1'h0,
    io_writeback_1_8_bits_uop_cf_exceptionVec_13,1'h0,4'h0,io_writeback_1_8_bits_uop_cf_exceptionVec_7,
    io_writeback_1_8_bits_uop_cf_exceptionVec_6,io_writeback_1_8_bits_uop_cf_exceptionVec_5,
    io_writeback_1_8_bits_uop_cf_exceptionVec_4,4'h0}; // @[Rob.scala 908:87]
  wire  wbHasException_8 = |_wbHasException_T_8; // @[Rob.scala 908:94]
  wire  wbHasTriggerHit_8 = io_writeback_1_8_bits_uop_cf_trigger_backendHit_0 |
    io_writeback_1_8_bits_uop_cf_trigger_backendHit_1 | io_writeback_1_8_bits_uop_cf_trigger_backendHit_2 |
    io_writeback_1_8_bits_uop_cf_trigger_backendHit_3 | io_writeback_1_8_bits_uop_cf_trigger_backendHit_4 |
    io_writeback_1_8_bits_uop_cf_trigger_backendHit_5; // @[Bundle.scala 629:43]
  wire  block_wb_8 = wbHasException_8 | wbHasTriggerHit_8; // @[Rob.scala 912:74]
  reg  REG_7; // @[Rob.scala 918:17]
  reg [4:0] REG_8; // @[Rob.scala 919:37]
  reg  REG_9; // @[Rob.scala 918:17]
  reg [4:0] REG_10; // @[Rob.scala 919:37]
  reg  REG_11; // @[Rob.scala 935:18]
  wire  _allow_interrupts_T_3 = ~io_enq_req_0_bits_ctrl_commitType[2] & io_enq_req_0_bits_ctrl_commitType[1]; // @[package.scala 135:68]
  reg [4:0] REG_12; // @[Rob.scala 943:29]
  reg  REG_13; // @[Rob.scala 943:66]
  reg  REG_14; // @[Rob.scala 935:18]
  wire  _allow_interrupts_T_7 = ~io_enq_req_1_bits_ctrl_commitType[2] & io_enq_req_1_bits_ctrl_commitType[1]; // @[package.scala 135:68]
  reg [4:0] REG_15; // @[Rob.scala 943:29]
  reg  REG_16; // @[Rob.scala 943:66]
  wire [4:0] _commitReadAddr_next_WIRE__0 = deqPtrGenModule_io_next_out_0_value; // @[Rob.scala 951:{12,12}]
  wire [4:0] _commitReadAddr_next_WIRE__1 = deqPtrGenModule_io_next_out_1_value; // @[Rob.scala 951:{12,12}]
  reg [63:0] instrCntReg; // @[Rob.scala 1018:28]
  reg  fuseCommitCnt_REG; // @[Rob.scala 1019:103]
  reg  fuseCommitCnt_REG_1; // @[Rob.scala 1019:103]
  wire [1:0] fuseCommitCnt = fuseCommitCnt_REG + fuseCommitCnt_REG_1; // @[Bitwise.scala 48:55]
  reg [1:0] trueCommitCnt_REG; // @[Rob.scala 1020:30]
  wire [2:0] trueCommitCnt = trueCommitCnt_REG + fuseCommitCnt; // @[Rob.scala 1020:42]
  reg  retireCounter_REG; // @[Rob.scala 1021:34]
  wire [2:0] retireCounter = retireCounter_REG ? trueCommitCnt : 3'h0; // @[Rob.scala 1021:26]
  wire [63:0] _GEN_11347 = {{61'd0}, retireCounter}; // @[Rob.scala 1022:30]
  wire [1:0] _T_433 = valid_0 + valid_1; // @[Bitwise.scala 48:55]
  wire [1:0] _T_435 = valid_2 + valid_3; // @[Bitwise.scala 48:55]
  wire [2:0] _T_437 = _T_433 + _T_435; // @[Bitwise.scala 48:55]
  wire [1:0] _T_439 = valid_4 + valid_5; // @[Bitwise.scala 48:55]
  wire [1:0] _T_441 = valid_6 + valid_7; // @[Bitwise.scala 48:55]
  wire [2:0] _T_443 = _T_439 + _T_441; // @[Bitwise.scala 48:55]
  wire [3:0] _T_445 = _T_437 + _T_443; // @[Bitwise.scala 48:55]
  wire [1:0] _T_447 = valid_8 + valid_9; // @[Bitwise.scala 48:55]
  wire [1:0] _T_449 = valid_10 + valid_11; // @[Bitwise.scala 48:55]
  wire [2:0] _T_451 = _T_447 + _T_449; // @[Bitwise.scala 48:55]
  wire [1:0] _T_453 = valid_12 + valid_13; // @[Bitwise.scala 48:55]
  wire [1:0] _T_455 = valid_14 + valid_15; // @[Bitwise.scala 48:55]
  wire [2:0] _T_457 = _T_453 + _T_455; // @[Bitwise.scala 48:55]
  wire [3:0] _T_459 = _T_451 + _T_457; // @[Bitwise.scala 48:55]
  wire [4:0] _T_461 = _T_445 + _T_459; // @[Bitwise.scala 48:55]
  wire [1:0] _T_463 = valid_16 + valid_17; // @[Bitwise.scala 48:55]
  wire [1:0] _T_465 = valid_18 + valid_19; // @[Bitwise.scala 48:55]
  wire [2:0] _T_467 = _T_463 + _T_465; // @[Bitwise.scala 48:55]
  wire [1:0] _T_469 = valid_20 + valid_21; // @[Bitwise.scala 48:55]
  wire [1:0] _T_471 = valid_22 + valid_23; // @[Bitwise.scala 48:55]
  wire [2:0] _T_473 = _T_469 + _T_471; // @[Bitwise.scala 48:55]
  wire [3:0] _T_475 = _T_467 + _T_473; // @[Bitwise.scala 48:55]
  wire [1:0] _T_477 = valid_24 + valid_25; // @[Bitwise.scala 48:55]
  wire [1:0] _T_479 = valid_26 + valid_27; // @[Bitwise.scala 48:55]
  wire [2:0] _T_481 = _T_477 + _T_479; // @[Bitwise.scala 48:55]
  wire [1:0] _T_483 = valid_28 + valid_29; // @[Bitwise.scala 48:55]
  wire [1:0] _T_485 = valid_30 + valid_31; // @[Bitwise.scala 48:55]
  wire [2:0] _T_487 = _T_483 + _T_485; // @[Bitwise.scala 48:55]
  wire [3:0] _T_489 = _T_481 + _T_487; // @[Bitwise.scala 48:55]
  wire [4:0] _T_491 = _T_475 + _T_489; // @[Bitwise.scala 48:55]
  wire  commitIsBranch_0 = io_commits_info_0_commitType == 3'h1; // @[Rob.scala 1066:64]
  wire  commitIsBranch_1 = io_commits_info_1_commitType == 3'h1; // @[Rob.scala 1066:64]
  wire [1:0] _T_619 = io_commits_walkValid_0 + io_commits_walkValid_1; // @[Bitwise.scala 48:55]
  reg  dt_exuDebug_0_isMMIO; // @[Rob.scala 1214:26]
  reg  dt_exuDebug_0_isPerfCnt; // @[Rob.scala 1214:26]
  reg  dt_exuDebug_1_isMMIO; // @[Rob.scala 1214:26]
  reg  dt_exuDebug_1_isPerfCnt; // @[Rob.scala 1214:26]
  reg  dt_exuDebug_2_isMMIO; // @[Rob.scala 1214:26]
  reg  dt_exuDebug_2_isPerfCnt; // @[Rob.scala 1214:26]
  reg  dt_exuDebug_3_isMMIO; // @[Rob.scala 1214:26]
  reg  dt_exuDebug_3_isPerfCnt; // @[Rob.scala 1214:26]
  reg  dt_exuDebug_4_isMMIO; // @[Rob.scala 1214:26]
  reg  dt_exuDebug_4_isPerfCnt; // @[Rob.scala 1214:26]
  reg  dt_exuDebug_5_isMMIO; // @[Rob.scala 1214:26]
  reg  dt_exuDebug_5_isPerfCnt; // @[Rob.scala 1214:26]
  reg  dt_exuDebug_6_isMMIO; // @[Rob.scala 1214:26]
  reg  dt_exuDebug_6_isPerfCnt; // @[Rob.scala 1214:26]
  reg  dt_exuDebug_7_isMMIO; // @[Rob.scala 1214:26]
  reg  dt_exuDebug_7_isPerfCnt; // @[Rob.scala 1214:26]
  reg  dt_exuDebug_8_isMMIO; // @[Rob.scala 1214:26]
  reg  dt_exuDebug_8_isPerfCnt; // @[Rob.scala 1214:26]
  reg  dt_exuDebug_9_isMMIO; // @[Rob.scala 1214:26]
  reg  dt_exuDebug_9_isPerfCnt; // @[Rob.scala 1214:26]
  reg  dt_exuDebug_10_isMMIO; // @[Rob.scala 1214:26]
  reg  dt_exuDebug_10_isPerfCnt; // @[Rob.scala 1214:26]
  reg  dt_exuDebug_11_isMMIO; // @[Rob.scala 1214:26]
  reg  dt_exuDebug_11_isPerfCnt; // @[Rob.scala 1214:26]
  reg  dt_exuDebug_12_isMMIO; // @[Rob.scala 1214:26]
  reg  dt_exuDebug_12_isPerfCnt; // @[Rob.scala 1214:26]
  reg  dt_exuDebug_13_isMMIO; // @[Rob.scala 1214:26]
  reg  dt_exuDebug_13_isPerfCnt; // @[Rob.scala 1214:26]
  reg  dt_exuDebug_14_isMMIO; // @[Rob.scala 1214:26]
  reg  dt_exuDebug_14_isPerfCnt; // @[Rob.scala 1214:26]
  reg  dt_exuDebug_15_isMMIO; // @[Rob.scala 1214:26]
  reg  dt_exuDebug_15_isPerfCnt; // @[Rob.scala 1214:26]
  reg  dt_exuDebug_16_isMMIO; // @[Rob.scala 1214:26]
  reg  dt_exuDebug_16_isPerfCnt; // @[Rob.scala 1214:26]
  reg  dt_exuDebug_17_isMMIO; // @[Rob.scala 1214:26]
  reg  dt_exuDebug_17_isPerfCnt; // @[Rob.scala 1214:26]
  reg  dt_exuDebug_18_isMMIO; // @[Rob.scala 1214:26]
  reg  dt_exuDebug_18_isPerfCnt; // @[Rob.scala 1214:26]
  reg  dt_exuDebug_19_isMMIO; // @[Rob.scala 1214:26]
  reg  dt_exuDebug_19_isPerfCnt; // @[Rob.scala 1214:26]
  reg  dt_exuDebug_20_isMMIO; // @[Rob.scala 1214:26]
  reg  dt_exuDebug_20_isPerfCnt; // @[Rob.scala 1214:26]
  reg  dt_exuDebug_21_isMMIO; // @[Rob.scala 1214:26]
  reg  dt_exuDebug_21_isPerfCnt; // @[Rob.scala 1214:26]
  reg  dt_exuDebug_22_isMMIO; // @[Rob.scala 1214:26]
  reg  dt_exuDebug_22_isPerfCnt; // @[Rob.scala 1214:26]
  reg  dt_exuDebug_23_isMMIO; // @[Rob.scala 1214:26]
  reg  dt_exuDebug_23_isPerfCnt; // @[Rob.scala 1214:26]
  reg  dt_exuDebug_24_isMMIO; // @[Rob.scala 1214:26]
  reg  dt_exuDebug_24_isPerfCnt; // @[Rob.scala 1214:26]
  reg  dt_exuDebug_25_isMMIO; // @[Rob.scala 1214:26]
  reg  dt_exuDebug_25_isPerfCnt; // @[Rob.scala 1214:26]
  reg  dt_exuDebug_26_isMMIO; // @[Rob.scala 1214:26]
  reg  dt_exuDebug_26_isPerfCnt; // @[Rob.scala 1214:26]
  reg  dt_exuDebug_27_isMMIO; // @[Rob.scala 1214:26]
  reg  dt_exuDebug_27_isPerfCnt; // @[Rob.scala 1214:26]
  reg  dt_exuDebug_28_isMMIO; // @[Rob.scala 1214:26]
  reg  dt_exuDebug_28_isPerfCnt; // @[Rob.scala 1214:26]
  reg  dt_exuDebug_29_isMMIO; // @[Rob.scala 1214:26]
  reg  dt_exuDebug_29_isPerfCnt; // @[Rob.scala 1214:26]
  reg  dt_exuDebug_30_isMMIO; // @[Rob.scala 1214:26]
  reg  dt_exuDebug_30_isPerfCnt; // @[Rob.scala 1214:26]
  reg  dt_exuDebug_31_isMMIO; // @[Rob.scala 1214:26]
  reg  dt_exuDebug_31_isPerfCnt; // @[Rob.scala 1214:26]
  wire  _GEN_8715 = 5'h0 == io_writeback_1_0_bits_uop_robIdx_value ? 1'h0 : dt_exuDebug_0_isMMIO; // @[Rob.scala 1214:26 1224:{28,28}]
  wire  _GEN_8716 = 5'h1 == io_writeback_1_0_bits_uop_robIdx_value ? 1'h0 : dt_exuDebug_1_isMMIO; // @[Rob.scala 1214:26 1224:{28,28}]
  wire  _GEN_8717 = 5'h2 == io_writeback_1_0_bits_uop_robIdx_value ? 1'h0 : dt_exuDebug_2_isMMIO; // @[Rob.scala 1214:26 1224:{28,28}]
  wire  _GEN_8718 = 5'h3 == io_writeback_1_0_bits_uop_robIdx_value ? 1'h0 : dt_exuDebug_3_isMMIO; // @[Rob.scala 1214:26 1224:{28,28}]
  wire  _GEN_8719 = 5'h4 == io_writeback_1_0_bits_uop_robIdx_value ? 1'h0 : dt_exuDebug_4_isMMIO; // @[Rob.scala 1214:26 1224:{28,28}]
  wire  _GEN_8720 = 5'h5 == io_writeback_1_0_bits_uop_robIdx_value ? 1'h0 : dt_exuDebug_5_isMMIO; // @[Rob.scala 1214:26 1224:{28,28}]
  wire  _GEN_8721 = 5'h6 == io_writeback_1_0_bits_uop_robIdx_value ? 1'h0 : dt_exuDebug_6_isMMIO; // @[Rob.scala 1214:26 1224:{28,28}]
  wire  _GEN_8722 = 5'h7 == io_writeback_1_0_bits_uop_robIdx_value ? 1'h0 : dt_exuDebug_7_isMMIO; // @[Rob.scala 1214:26 1224:{28,28}]
  wire  _GEN_8723 = 5'h8 == io_writeback_1_0_bits_uop_robIdx_value ? 1'h0 : dt_exuDebug_8_isMMIO; // @[Rob.scala 1214:26 1224:{28,28}]
  wire  _GEN_8724 = 5'h9 == io_writeback_1_0_bits_uop_robIdx_value ? 1'h0 : dt_exuDebug_9_isMMIO; // @[Rob.scala 1214:26 1224:{28,28}]
  wire  _GEN_8725 = 5'ha == io_writeback_1_0_bits_uop_robIdx_value ? 1'h0 : dt_exuDebug_10_isMMIO; // @[Rob.scala 1214:26 1224:{28,28}]
  wire  _GEN_8726 = 5'hb == io_writeback_1_0_bits_uop_robIdx_value ? 1'h0 : dt_exuDebug_11_isMMIO; // @[Rob.scala 1214:26 1224:{28,28}]
  wire  _GEN_8727 = 5'hc == io_writeback_1_0_bits_uop_robIdx_value ? 1'h0 : dt_exuDebug_12_isMMIO; // @[Rob.scala 1214:26 1224:{28,28}]
  wire  _GEN_8728 = 5'hd == io_writeback_1_0_bits_uop_robIdx_value ? 1'h0 : dt_exuDebug_13_isMMIO; // @[Rob.scala 1214:26 1224:{28,28}]
  wire  _GEN_8729 = 5'he == io_writeback_1_0_bits_uop_robIdx_value ? 1'h0 : dt_exuDebug_14_isMMIO; // @[Rob.scala 1214:26 1224:{28,28}]
  wire  _GEN_8730 = 5'hf == io_writeback_1_0_bits_uop_robIdx_value ? 1'h0 : dt_exuDebug_15_isMMIO; // @[Rob.scala 1214:26 1224:{28,28}]
  wire  _GEN_8731 = 5'h10 == io_writeback_1_0_bits_uop_robIdx_value ? 1'h0 : dt_exuDebug_16_isMMIO; // @[Rob.scala 1214:26 1224:{28,28}]
  wire  _GEN_8732 = 5'h11 == io_writeback_1_0_bits_uop_robIdx_value ? 1'h0 : dt_exuDebug_17_isMMIO; // @[Rob.scala 1214:26 1224:{28,28}]
  wire  _GEN_8733 = 5'h12 == io_writeback_1_0_bits_uop_robIdx_value ? 1'h0 : dt_exuDebug_18_isMMIO; // @[Rob.scala 1214:26 1224:{28,28}]
  wire  _GEN_8734 = 5'h13 == io_writeback_1_0_bits_uop_robIdx_value ? 1'h0 : dt_exuDebug_19_isMMIO; // @[Rob.scala 1214:26 1224:{28,28}]
  wire  _GEN_8735 = 5'h14 == io_writeback_1_0_bits_uop_robIdx_value ? 1'h0 : dt_exuDebug_20_isMMIO; // @[Rob.scala 1214:26 1224:{28,28}]
  wire  _GEN_8736 = 5'h15 == io_writeback_1_0_bits_uop_robIdx_value ? 1'h0 : dt_exuDebug_21_isMMIO; // @[Rob.scala 1214:26 1224:{28,28}]
  wire  _GEN_8737 = 5'h16 == io_writeback_1_0_bits_uop_robIdx_value ? 1'h0 : dt_exuDebug_22_isMMIO; // @[Rob.scala 1214:26 1224:{28,28}]
  wire  _GEN_8738 = 5'h17 == io_writeback_1_0_bits_uop_robIdx_value ? 1'h0 : dt_exuDebug_23_isMMIO; // @[Rob.scala 1214:26 1224:{28,28}]
  wire  _GEN_8739 = 5'h18 == io_writeback_1_0_bits_uop_robIdx_value ? 1'h0 : dt_exuDebug_24_isMMIO; // @[Rob.scala 1214:26 1224:{28,28}]
  wire  _GEN_8740 = 5'h19 == io_writeback_1_0_bits_uop_robIdx_value ? 1'h0 : dt_exuDebug_25_isMMIO; // @[Rob.scala 1214:26 1224:{28,28}]
  wire  _GEN_8741 = 5'h1a == io_writeback_1_0_bits_uop_robIdx_value ? 1'h0 : dt_exuDebug_26_isMMIO; // @[Rob.scala 1214:26 1224:{28,28}]
  wire  _GEN_8742 = 5'h1b == io_writeback_1_0_bits_uop_robIdx_value ? 1'h0 : dt_exuDebug_27_isMMIO; // @[Rob.scala 1214:26 1224:{28,28}]
  wire  _GEN_8743 = 5'h1c == io_writeback_1_0_bits_uop_robIdx_value ? 1'h0 : dt_exuDebug_28_isMMIO; // @[Rob.scala 1214:26 1224:{28,28}]
  wire  _GEN_8744 = 5'h1d == io_writeback_1_0_bits_uop_robIdx_value ? 1'h0 : dt_exuDebug_29_isMMIO; // @[Rob.scala 1214:26 1224:{28,28}]
  wire  _GEN_8745 = 5'h1e == io_writeback_1_0_bits_uop_robIdx_value ? 1'h0 : dt_exuDebug_30_isMMIO; // @[Rob.scala 1214:26 1224:{28,28}]
  wire  _GEN_8746 = 5'h1f == io_writeback_1_0_bits_uop_robIdx_value ? 1'h0 : dt_exuDebug_31_isMMIO; // @[Rob.scala 1214:26 1224:{28,28}]
  wire  _GEN_8747 = 5'h0 == io_writeback_1_0_bits_uop_robIdx_value ? 1'h0 : dt_exuDebug_0_isPerfCnt; // @[Rob.scala 1214:26 1224:{28,28}]
  wire  _GEN_8748 = 5'h1 == io_writeback_1_0_bits_uop_robIdx_value ? 1'h0 : dt_exuDebug_1_isPerfCnt; // @[Rob.scala 1214:26 1224:{28,28}]
  wire  _GEN_8749 = 5'h2 == io_writeback_1_0_bits_uop_robIdx_value ? 1'h0 : dt_exuDebug_2_isPerfCnt; // @[Rob.scala 1214:26 1224:{28,28}]
  wire  _GEN_8750 = 5'h3 == io_writeback_1_0_bits_uop_robIdx_value ? 1'h0 : dt_exuDebug_3_isPerfCnt; // @[Rob.scala 1214:26 1224:{28,28}]
  wire  _GEN_8751 = 5'h4 == io_writeback_1_0_bits_uop_robIdx_value ? 1'h0 : dt_exuDebug_4_isPerfCnt; // @[Rob.scala 1214:26 1224:{28,28}]
  wire  _GEN_8752 = 5'h5 == io_writeback_1_0_bits_uop_robIdx_value ? 1'h0 : dt_exuDebug_5_isPerfCnt; // @[Rob.scala 1214:26 1224:{28,28}]
  wire  _GEN_8753 = 5'h6 == io_writeback_1_0_bits_uop_robIdx_value ? 1'h0 : dt_exuDebug_6_isPerfCnt; // @[Rob.scala 1214:26 1224:{28,28}]
  wire  _GEN_8754 = 5'h7 == io_writeback_1_0_bits_uop_robIdx_value ? 1'h0 : dt_exuDebug_7_isPerfCnt; // @[Rob.scala 1214:26 1224:{28,28}]
  wire  _GEN_8755 = 5'h8 == io_writeback_1_0_bits_uop_robIdx_value ? 1'h0 : dt_exuDebug_8_isPerfCnt; // @[Rob.scala 1214:26 1224:{28,28}]
  wire  _GEN_8756 = 5'h9 == io_writeback_1_0_bits_uop_robIdx_value ? 1'h0 : dt_exuDebug_9_isPerfCnt; // @[Rob.scala 1214:26 1224:{28,28}]
  wire  _GEN_8757 = 5'ha == io_writeback_1_0_bits_uop_robIdx_value ? 1'h0 : dt_exuDebug_10_isPerfCnt; // @[Rob.scala 1214:26 1224:{28,28}]
  wire  _GEN_8758 = 5'hb == io_writeback_1_0_bits_uop_robIdx_value ? 1'h0 : dt_exuDebug_11_isPerfCnt; // @[Rob.scala 1214:26 1224:{28,28}]
  wire  _GEN_8759 = 5'hc == io_writeback_1_0_bits_uop_robIdx_value ? 1'h0 : dt_exuDebug_12_isPerfCnt; // @[Rob.scala 1214:26 1224:{28,28}]
  wire  _GEN_8760 = 5'hd == io_writeback_1_0_bits_uop_robIdx_value ? 1'h0 : dt_exuDebug_13_isPerfCnt; // @[Rob.scala 1214:26 1224:{28,28}]
  wire  _GEN_8761 = 5'he == io_writeback_1_0_bits_uop_robIdx_value ? 1'h0 : dt_exuDebug_14_isPerfCnt; // @[Rob.scala 1214:26 1224:{28,28}]
  wire  _GEN_8762 = 5'hf == io_writeback_1_0_bits_uop_robIdx_value ? 1'h0 : dt_exuDebug_15_isPerfCnt; // @[Rob.scala 1214:26 1224:{28,28}]
  wire  _GEN_8763 = 5'h10 == io_writeback_1_0_bits_uop_robIdx_value ? 1'h0 : dt_exuDebug_16_isPerfCnt; // @[Rob.scala 1214:26 1224:{28,28}]
  wire  _GEN_8764 = 5'h11 == io_writeback_1_0_bits_uop_robIdx_value ? 1'h0 : dt_exuDebug_17_isPerfCnt; // @[Rob.scala 1214:26 1224:{28,28}]
  wire  _GEN_8765 = 5'h12 == io_writeback_1_0_bits_uop_robIdx_value ? 1'h0 : dt_exuDebug_18_isPerfCnt; // @[Rob.scala 1214:26 1224:{28,28}]
  wire  _GEN_8766 = 5'h13 == io_writeback_1_0_bits_uop_robIdx_value ? 1'h0 : dt_exuDebug_19_isPerfCnt; // @[Rob.scala 1214:26 1224:{28,28}]
  wire  _GEN_8767 = 5'h14 == io_writeback_1_0_bits_uop_robIdx_value ? 1'h0 : dt_exuDebug_20_isPerfCnt; // @[Rob.scala 1214:26 1224:{28,28}]
  wire  _GEN_8768 = 5'h15 == io_writeback_1_0_bits_uop_robIdx_value ? 1'h0 : dt_exuDebug_21_isPerfCnt; // @[Rob.scala 1214:26 1224:{28,28}]
  wire  _GEN_8769 = 5'h16 == io_writeback_1_0_bits_uop_robIdx_value ? 1'h0 : dt_exuDebug_22_isPerfCnt; // @[Rob.scala 1214:26 1224:{28,28}]
  wire  _GEN_8770 = 5'h17 == io_writeback_1_0_bits_uop_robIdx_value ? 1'h0 : dt_exuDebug_23_isPerfCnt; // @[Rob.scala 1214:26 1224:{28,28}]
  wire  _GEN_8771 = 5'h18 == io_writeback_1_0_bits_uop_robIdx_value ? 1'h0 : dt_exuDebug_24_isPerfCnt; // @[Rob.scala 1214:26 1224:{28,28}]
  wire  _GEN_8772 = 5'h19 == io_writeback_1_0_bits_uop_robIdx_value ? 1'h0 : dt_exuDebug_25_isPerfCnt; // @[Rob.scala 1214:26 1224:{28,28}]
  wire  _GEN_8773 = 5'h1a == io_writeback_1_0_bits_uop_robIdx_value ? 1'h0 : dt_exuDebug_26_isPerfCnt; // @[Rob.scala 1214:26 1224:{28,28}]
  wire  _GEN_8774 = 5'h1b == io_writeback_1_0_bits_uop_robIdx_value ? 1'h0 : dt_exuDebug_27_isPerfCnt; // @[Rob.scala 1214:26 1224:{28,28}]
  wire  _GEN_8775 = 5'h1c == io_writeback_1_0_bits_uop_robIdx_value ? 1'h0 : dt_exuDebug_28_isPerfCnt; // @[Rob.scala 1214:26 1224:{28,28}]
  wire  _GEN_8776 = 5'h1d == io_writeback_1_0_bits_uop_robIdx_value ? 1'h0 : dt_exuDebug_29_isPerfCnt; // @[Rob.scala 1214:26 1224:{28,28}]
  wire  _GEN_8777 = 5'h1e == io_writeback_1_0_bits_uop_robIdx_value ? 1'h0 : dt_exuDebug_30_isPerfCnt; // @[Rob.scala 1214:26 1224:{28,28}]
  wire  _GEN_8778 = 5'h1f == io_writeback_1_0_bits_uop_robIdx_value ? 1'h0 : dt_exuDebug_31_isPerfCnt; // @[Rob.scala 1214:26 1224:{28,28}]
  wire  _GEN_8843 = io_writeback_1_0_valid ? _GEN_8715 : dt_exuDebug_0_isMMIO; // @[Rob.scala 1222:23 1214:26]
  wire  _GEN_8844 = io_writeback_1_0_valid ? _GEN_8716 : dt_exuDebug_1_isMMIO; // @[Rob.scala 1222:23 1214:26]
  wire  _GEN_8845 = io_writeback_1_0_valid ? _GEN_8717 : dt_exuDebug_2_isMMIO; // @[Rob.scala 1222:23 1214:26]
  wire  _GEN_8846 = io_writeback_1_0_valid ? _GEN_8718 : dt_exuDebug_3_isMMIO; // @[Rob.scala 1222:23 1214:26]
  wire  _GEN_8847 = io_writeback_1_0_valid ? _GEN_8719 : dt_exuDebug_4_isMMIO; // @[Rob.scala 1222:23 1214:26]
  wire  _GEN_8848 = io_writeback_1_0_valid ? _GEN_8720 : dt_exuDebug_5_isMMIO; // @[Rob.scala 1222:23 1214:26]
  wire  _GEN_8849 = io_writeback_1_0_valid ? _GEN_8721 : dt_exuDebug_6_isMMIO; // @[Rob.scala 1222:23 1214:26]
  wire  _GEN_8850 = io_writeback_1_0_valid ? _GEN_8722 : dt_exuDebug_7_isMMIO; // @[Rob.scala 1222:23 1214:26]
  wire  _GEN_8851 = io_writeback_1_0_valid ? _GEN_8723 : dt_exuDebug_8_isMMIO; // @[Rob.scala 1222:23 1214:26]
  wire  _GEN_8852 = io_writeback_1_0_valid ? _GEN_8724 : dt_exuDebug_9_isMMIO; // @[Rob.scala 1222:23 1214:26]
  wire  _GEN_8853 = io_writeback_1_0_valid ? _GEN_8725 : dt_exuDebug_10_isMMIO; // @[Rob.scala 1222:23 1214:26]
  wire  _GEN_8854 = io_writeback_1_0_valid ? _GEN_8726 : dt_exuDebug_11_isMMIO; // @[Rob.scala 1222:23 1214:26]
  wire  _GEN_8855 = io_writeback_1_0_valid ? _GEN_8727 : dt_exuDebug_12_isMMIO; // @[Rob.scala 1222:23 1214:26]
  wire  _GEN_8856 = io_writeback_1_0_valid ? _GEN_8728 : dt_exuDebug_13_isMMIO; // @[Rob.scala 1222:23 1214:26]
  wire  _GEN_8857 = io_writeback_1_0_valid ? _GEN_8729 : dt_exuDebug_14_isMMIO; // @[Rob.scala 1222:23 1214:26]
  wire  _GEN_8858 = io_writeback_1_0_valid ? _GEN_8730 : dt_exuDebug_15_isMMIO; // @[Rob.scala 1222:23 1214:26]
  wire  _GEN_8859 = io_writeback_1_0_valid ? _GEN_8731 : dt_exuDebug_16_isMMIO; // @[Rob.scala 1222:23 1214:26]
  wire  _GEN_8860 = io_writeback_1_0_valid ? _GEN_8732 : dt_exuDebug_17_isMMIO; // @[Rob.scala 1222:23 1214:26]
  wire  _GEN_8861 = io_writeback_1_0_valid ? _GEN_8733 : dt_exuDebug_18_isMMIO; // @[Rob.scala 1222:23 1214:26]
  wire  _GEN_8862 = io_writeback_1_0_valid ? _GEN_8734 : dt_exuDebug_19_isMMIO; // @[Rob.scala 1222:23 1214:26]
  wire  _GEN_8863 = io_writeback_1_0_valid ? _GEN_8735 : dt_exuDebug_20_isMMIO; // @[Rob.scala 1222:23 1214:26]
  wire  _GEN_8864 = io_writeback_1_0_valid ? _GEN_8736 : dt_exuDebug_21_isMMIO; // @[Rob.scala 1222:23 1214:26]
  wire  _GEN_8865 = io_writeback_1_0_valid ? _GEN_8737 : dt_exuDebug_22_isMMIO; // @[Rob.scala 1222:23 1214:26]
  wire  _GEN_8866 = io_writeback_1_0_valid ? _GEN_8738 : dt_exuDebug_23_isMMIO; // @[Rob.scala 1222:23 1214:26]
  wire  _GEN_8867 = io_writeback_1_0_valid ? _GEN_8739 : dt_exuDebug_24_isMMIO; // @[Rob.scala 1222:23 1214:26]
  wire  _GEN_8868 = io_writeback_1_0_valid ? _GEN_8740 : dt_exuDebug_25_isMMIO; // @[Rob.scala 1222:23 1214:26]
  wire  _GEN_8869 = io_writeback_1_0_valid ? _GEN_8741 : dt_exuDebug_26_isMMIO; // @[Rob.scala 1222:23 1214:26]
  wire  _GEN_8870 = io_writeback_1_0_valid ? _GEN_8742 : dt_exuDebug_27_isMMIO; // @[Rob.scala 1222:23 1214:26]
  wire  _GEN_8871 = io_writeback_1_0_valid ? _GEN_8743 : dt_exuDebug_28_isMMIO; // @[Rob.scala 1222:23 1214:26]
  wire  _GEN_8872 = io_writeback_1_0_valid ? _GEN_8744 : dt_exuDebug_29_isMMIO; // @[Rob.scala 1222:23 1214:26]
  wire  _GEN_8873 = io_writeback_1_0_valid ? _GEN_8745 : dt_exuDebug_30_isMMIO; // @[Rob.scala 1222:23 1214:26]
  wire  _GEN_8874 = io_writeback_1_0_valid ? _GEN_8746 : dt_exuDebug_31_isMMIO; // @[Rob.scala 1222:23 1214:26]
  wire  _GEN_8875 = io_writeback_1_0_valid ? _GEN_8747 : dt_exuDebug_0_isPerfCnt; // @[Rob.scala 1222:23 1214:26]
  wire  _GEN_8876 = io_writeback_1_0_valid ? _GEN_8748 : dt_exuDebug_1_isPerfCnt; // @[Rob.scala 1222:23 1214:26]
  wire  _GEN_8877 = io_writeback_1_0_valid ? _GEN_8749 : dt_exuDebug_2_isPerfCnt; // @[Rob.scala 1222:23 1214:26]
  wire  _GEN_8878 = io_writeback_1_0_valid ? _GEN_8750 : dt_exuDebug_3_isPerfCnt; // @[Rob.scala 1222:23 1214:26]
  wire  _GEN_8879 = io_writeback_1_0_valid ? _GEN_8751 : dt_exuDebug_4_isPerfCnt; // @[Rob.scala 1222:23 1214:26]
  wire  _GEN_8880 = io_writeback_1_0_valid ? _GEN_8752 : dt_exuDebug_5_isPerfCnt; // @[Rob.scala 1222:23 1214:26]
  wire  _GEN_8881 = io_writeback_1_0_valid ? _GEN_8753 : dt_exuDebug_6_isPerfCnt; // @[Rob.scala 1222:23 1214:26]
  wire  _GEN_8882 = io_writeback_1_0_valid ? _GEN_8754 : dt_exuDebug_7_isPerfCnt; // @[Rob.scala 1222:23 1214:26]
  wire  _GEN_8883 = io_writeback_1_0_valid ? _GEN_8755 : dt_exuDebug_8_isPerfCnt; // @[Rob.scala 1222:23 1214:26]
  wire  _GEN_8884 = io_writeback_1_0_valid ? _GEN_8756 : dt_exuDebug_9_isPerfCnt; // @[Rob.scala 1222:23 1214:26]
  wire  _GEN_8885 = io_writeback_1_0_valid ? _GEN_8757 : dt_exuDebug_10_isPerfCnt; // @[Rob.scala 1222:23 1214:26]
  wire  _GEN_8886 = io_writeback_1_0_valid ? _GEN_8758 : dt_exuDebug_11_isPerfCnt; // @[Rob.scala 1222:23 1214:26]
  wire  _GEN_8887 = io_writeback_1_0_valid ? _GEN_8759 : dt_exuDebug_12_isPerfCnt; // @[Rob.scala 1222:23 1214:26]
  wire  _GEN_8888 = io_writeback_1_0_valid ? _GEN_8760 : dt_exuDebug_13_isPerfCnt; // @[Rob.scala 1222:23 1214:26]
  wire  _GEN_8889 = io_writeback_1_0_valid ? _GEN_8761 : dt_exuDebug_14_isPerfCnt; // @[Rob.scala 1222:23 1214:26]
  wire  _GEN_8890 = io_writeback_1_0_valid ? _GEN_8762 : dt_exuDebug_15_isPerfCnt; // @[Rob.scala 1222:23 1214:26]
  wire  _GEN_8891 = io_writeback_1_0_valid ? _GEN_8763 : dt_exuDebug_16_isPerfCnt; // @[Rob.scala 1222:23 1214:26]
  wire  _GEN_8892 = io_writeback_1_0_valid ? _GEN_8764 : dt_exuDebug_17_isPerfCnt; // @[Rob.scala 1222:23 1214:26]
  wire  _GEN_8893 = io_writeback_1_0_valid ? _GEN_8765 : dt_exuDebug_18_isPerfCnt; // @[Rob.scala 1222:23 1214:26]
  wire  _GEN_8894 = io_writeback_1_0_valid ? _GEN_8766 : dt_exuDebug_19_isPerfCnt; // @[Rob.scala 1222:23 1214:26]
  wire  _GEN_8895 = io_writeback_1_0_valid ? _GEN_8767 : dt_exuDebug_20_isPerfCnt; // @[Rob.scala 1222:23 1214:26]
  wire  _GEN_8896 = io_writeback_1_0_valid ? _GEN_8768 : dt_exuDebug_21_isPerfCnt; // @[Rob.scala 1222:23 1214:26]
  wire  _GEN_8897 = io_writeback_1_0_valid ? _GEN_8769 : dt_exuDebug_22_isPerfCnt; // @[Rob.scala 1222:23 1214:26]
  wire  _GEN_8898 = io_writeback_1_0_valid ? _GEN_8770 : dt_exuDebug_23_isPerfCnt; // @[Rob.scala 1222:23 1214:26]
  wire  _GEN_8899 = io_writeback_1_0_valid ? _GEN_8771 : dt_exuDebug_24_isPerfCnt; // @[Rob.scala 1222:23 1214:26]
  wire  _GEN_8900 = io_writeback_1_0_valid ? _GEN_8772 : dt_exuDebug_25_isPerfCnt; // @[Rob.scala 1222:23 1214:26]
  wire  _GEN_8901 = io_writeback_1_0_valid ? _GEN_8773 : dt_exuDebug_26_isPerfCnt; // @[Rob.scala 1222:23 1214:26]
  wire  _GEN_8902 = io_writeback_1_0_valid ? _GEN_8774 : dt_exuDebug_27_isPerfCnt; // @[Rob.scala 1222:23 1214:26]
  wire  _GEN_8903 = io_writeback_1_0_valid ? _GEN_8775 : dt_exuDebug_28_isPerfCnt; // @[Rob.scala 1222:23 1214:26]
  wire  _GEN_8904 = io_writeback_1_0_valid ? _GEN_8776 : dt_exuDebug_29_isPerfCnt; // @[Rob.scala 1222:23 1214:26]
  wire  _GEN_8905 = io_writeback_1_0_valid ? _GEN_8777 : dt_exuDebug_30_isPerfCnt; // @[Rob.scala 1222:23 1214:26]
  wire  _GEN_8906 = io_writeback_1_0_valid ? _GEN_8778 : dt_exuDebug_31_isPerfCnt; // @[Rob.scala 1222:23 1214:26]
  wire  _GEN_8971 = 5'h0 == io_writeback_1_1_bits_uop_robIdx_value ? 1'h0 : _GEN_8843; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_8972 = 5'h1 == io_writeback_1_1_bits_uop_robIdx_value ? 1'h0 : _GEN_8844; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_8973 = 5'h2 == io_writeback_1_1_bits_uop_robIdx_value ? 1'h0 : _GEN_8845; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_8974 = 5'h3 == io_writeback_1_1_bits_uop_robIdx_value ? 1'h0 : _GEN_8846; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_8975 = 5'h4 == io_writeback_1_1_bits_uop_robIdx_value ? 1'h0 : _GEN_8847; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_8976 = 5'h5 == io_writeback_1_1_bits_uop_robIdx_value ? 1'h0 : _GEN_8848; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_8977 = 5'h6 == io_writeback_1_1_bits_uop_robIdx_value ? 1'h0 : _GEN_8849; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_8978 = 5'h7 == io_writeback_1_1_bits_uop_robIdx_value ? 1'h0 : _GEN_8850; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_8979 = 5'h8 == io_writeback_1_1_bits_uop_robIdx_value ? 1'h0 : _GEN_8851; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_8980 = 5'h9 == io_writeback_1_1_bits_uop_robIdx_value ? 1'h0 : _GEN_8852; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_8981 = 5'ha == io_writeback_1_1_bits_uop_robIdx_value ? 1'h0 : _GEN_8853; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_8982 = 5'hb == io_writeback_1_1_bits_uop_robIdx_value ? 1'h0 : _GEN_8854; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_8983 = 5'hc == io_writeback_1_1_bits_uop_robIdx_value ? 1'h0 : _GEN_8855; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_8984 = 5'hd == io_writeback_1_1_bits_uop_robIdx_value ? 1'h0 : _GEN_8856; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_8985 = 5'he == io_writeback_1_1_bits_uop_robIdx_value ? 1'h0 : _GEN_8857; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_8986 = 5'hf == io_writeback_1_1_bits_uop_robIdx_value ? 1'h0 : _GEN_8858; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_8987 = 5'h10 == io_writeback_1_1_bits_uop_robIdx_value ? 1'h0 : _GEN_8859; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_8988 = 5'h11 == io_writeback_1_1_bits_uop_robIdx_value ? 1'h0 : _GEN_8860; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_8989 = 5'h12 == io_writeback_1_1_bits_uop_robIdx_value ? 1'h0 : _GEN_8861; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_8990 = 5'h13 == io_writeback_1_1_bits_uop_robIdx_value ? 1'h0 : _GEN_8862; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_8991 = 5'h14 == io_writeback_1_1_bits_uop_robIdx_value ? 1'h0 : _GEN_8863; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_8992 = 5'h15 == io_writeback_1_1_bits_uop_robIdx_value ? 1'h0 : _GEN_8864; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_8993 = 5'h16 == io_writeback_1_1_bits_uop_robIdx_value ? 1'h0 : _GEN_8865; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_8994 = 5'h17 == io_writeback_1_1_bits_uop_robIdx_value ? 1'h0 : _GEN_8866; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_8995 = 5'h18 == io_writeback_1_1_bits_uop_robIdx_value ? 1'h0 : _GEN_8867; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_8996 = 5'h19 == io_writeback_1_1_bits_uop_robIdx_value ? 1'h0 : _GEN_8868; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_8997 = 5'h1a == io_writeback_1_1_bits_uop_robIdx_value ? 1'h0 : _GEN_8869; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_8998 = 5'h1b == io_writeback_1_1_bits_uop_robIdx_value ? 1'h0 : _GEN_8870; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_8999 = 5'h1c == io_writeback_1_1_bits_uop_robIdx_value ? 1'h0 : _GEN_8871; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9000 = 5'h1d == io_writeback_1_1_bits_uop_robIdx_value ? 1'h0 : _GEN_8872; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9001 = 5'h1e == io_writeback_1_1_bits_uop_robIdx_value ? 1'h0 : _GEN_8873; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9002 = 5'h1f == io_writeback_1_1_bits_uop_robIdx_value ? 1'h0 : _GEN_8874; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9003 = 5'h0 == io_writeback_1_1_bits_uop_robIdx_value ? 1'h0 : _GEN_8875; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9004 = 5'h1 == io_writeback_1_1_bits_uop_robIdx_value ? 1'h0 : _GEN_8876; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9005 = 5'h2 == io_writeback_1_1_bits_uop_robIdx_value ? 1'h0 : _GEN_8877; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9006 = 5'h3 == io_writeback_1_1_bits_uop_robIdx_value ? 1'h0 : _GEN_8878; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9007 = 5'h4 == io_writeback_1_1_bits_uop_robIdx_value ? 1'h0 : _GEN_8879; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9008 = 5'h5 == io_writeback_1_1_bits_uop_robIdx_value ? 1'h0 : _GEN_8880; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9009 = 5'h6 == io_writeback_1_1_bits_uop_robIdx_value ? 1'h0 : _GEN_8881; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9010 = 5'h7 == io_writeback_1_1_bits_uop_robIdx_value ? 1'h0 : _GEN_8882; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9011 = 5'h8 == io_writeback_1_1_bits_uop_robIdx_value ? 1'h0 : _GEN_8883; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9012 = 5'h9 == io_writeback_1_1_bits_uop_robIdx_value ? 1'h0 : _GEN_8884; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9013 = 5'ha == io_writeback_1_1_bits_uop_robIdx_value ? 1'h0 : _GEN_8885; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9014 = 5'hb == io_writeback_1_1_bits_uop_robIdx_value ? 1'h0 : _GEN_8886; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9015 = 5'hc == io_writeback_1_1_bits_uop_robIdx_value ? 1'h0 : _GEN_8887; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9016 = 5'hd == io_writeback_1_1_bits_uop_robIdx_value ? 1'h0 : _GEN_8888; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9017 = 5'he == io_writeback_1_1_bits_uop_robIdx_value ? 1'h0 : _GEN_8889; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9018 = 5'hf == io_writeback_1_1_bits_uop_robIdx_value ? 1'h0 : _GEN_8890; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9019 = 5'h10 == io_writeback_1_1_bits_uop_robIdx_value ? 1'h0 : _GEN_8891; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9020 = 5'h11 == io_writeback_1_1_bits_uop_robIdx_value ? 1'h0 : _GEN_8892; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9021 = 5'h12 == io_writeback_1_1_bits_uop_robIdx_value ? 1'h0 : _GEN_8893; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9022 = 5'h13 == io_writeback_1_1_bits_uop_robIdx_value ? 1'h0 : _GEN_8894; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9023 = 5'h14 == io_writeback_1_1_bits_uop_robIdx_value ? 1'h0 : _GEN_8895; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9024 = 5'h15 == io_writeback_1_1_bits_uop_robIdx_value ? 1'h0 : _GEN_8896; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9025 = 5'h16 == io_writeback_1_1_bits_uop_robIdx_value ? 1'h0 : _GEN_8897; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9026 = 5'h17 == io_writeback_1_1_bits_uop_robIdx_value ? 1'h0 : _GEN_8898; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9027 = 5'h18 == io_writeback_1_1_bits_uop_robIdx_value ? 1'h0 : _GEN_8899; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9028 = 5'h19 == io_writeback_1_1_bits_uop_robIdx_value ? 1'h0 : _GEN_8900; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9029 = 5'h1a == io_writeback_1_1_bits_uop_robIdx_value ? 1'h0 : _GEN_8901; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9030 = 5'h1b == io_writeback_1_1_bits_uop_robIdx_value ? 1'h0 : _GEN_8902; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9031 = 5'h1c == io_writeback_1_1_bits_uop_robIdx_value ? 1'h0 : _GEN_8903; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9032 = 5'h1d == io_writeback_1_1_bits_uop_robIdx_value ? 1'h0 : _GEN_8904; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9033 = 5'h1e == io_writeback_1_1_bits_uop_robIdx_value ? 1'h0 : _GEN_8905; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9034 = 5'h1f == io_writeback_1_1_bits_uop_robIdx_value ? 1'h0 : _GEN_8906; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9099 = io_writeback_1_1_valid ? _GEN_8971 : _GEN_8843; // @[Rob.scala 1222:23]
  wire  _GEN_9100 = io_writeback_1_1_valid ? _GEN_8972 : _GEN_8844; // @[Rob.scala 1222:23]
  wire  _GEN_9101 = io_writeback_1_1_valid ? _GEN_8973 : _GEN_8845; // @[Rob.scala 1222:23]
  wire  _GEN_9102 = io_writeback_1_1_valid ? _GEN_8974 : _GEN_8846; // @[Rob.scala 1222:23]
  wire  _GEN_9103 = io_writeback_1_1_valid ? _GEN_8975 : _GEN_8847; // @[Rob.scala 1222:23]
  wire  _GEN_9104 = io_writeback_1_1_valid ? _GEN_8976 : _GEN_8848; // @[Rob.scala 1222:23]
  wire  _GEN_9105 = io_writeback_1_1_valid ? _GEN_8977 : _GEN_8849; // @[Rob.scala 1222:23]
  wire  _GEN_9106 = io_writeback_1_1_valid ? _GEN_8978 : _GEN_8850; // @[Rob.scala 1222:23]
  wire  _GEN_9107 = io_writeback_1_1_valid ? _GEN_8979 : _GEN_8851; // @[Rob.scala 1222:23]
  wire  _GEN_9108 = io_writeback_1_1_valid ? _GEN_8980 : _GEN_8852; // @[Rob.scala 1222:23]
  wire  _GEN_9109 = io_writeback_1_1_valid ? _GEN_8981 : _GEN_8853; // @[Rob.scala 1222:23]
  wire  _GEN_9110 = io_writeback_1_1_valid ? _GEN_8982 : _GEN_8854; // @[Rob.scala 1222:23]
  wire  _GEN_9111 = io_writeback_1_1_valid ? _GEN_8983 : _GEN_8855; // @[Rob.scala 1222:23]
  wire  _GEN_9112 = io_writeback_1_1_valid ? _GEN_8984 : _GEN_8856; // @[Rob.scala 1222:23]
  wire  _GEN_9113 = io_writeback_1_1_valid ? _GEN_8985 : _GEN_8857; // @[Rob.scala 1222:23]
  wire  _GEN_9114 = io_writeback_1_1_valid ? _GEN_8986 : _GEN_8858; // @[Rob.scala 1222:23]
  wire  _GEN_9115 = io_writeback_1_1_valid ? _GEN_8987 : _GEN_8859; // @[Rob.scala 1222:23]
  wire  _GEN_9116 = io_writeback_1_1_valid ? _GEN_8988 : _GEN_8860; // @[Rob.scala 1222:23]
  wire  _GEN_9117 = io_writeback_1_1_valid ? _GEN_8989 : _GEN_8861; // @[Rob.scala 1222:23]
  wire  _GEN_9118 = io_writeback_1_1_valid ? _GEN_8990 : _GEN_8862; // @[Rob.scala 1222:23]
  wire  _GEN_9119 = io_writeback_1_1_valid ? _GEN_8991 : _GEN_8863; // @[Rob.scala 1222:23]
  wire  _GEN_9120 = io_writeback_1_1_valid ? _GEN_8992 : _GEN_8864; // @[Rob.scala 1222:23]
  wire  _GEN_9121 = io_writeback_1_1_valid ? _GEN_8993 : _GEN_8865; // @[Rob.scala 1222:23]
  wire  _GEN_9122 = io_writeback_1_1_valid ? _GEN_8994 : _GEN_8866; // @[Rob.scala 1222:23]
  wire  _GEN_9123 = io_writeback_1_1_valid ? _GEN_8995 : _GEN_8867; // @[Rob.scala 1222:23]
  wire  _GEN_9124 = io_writeback_1_1_valid ? _GEN_8996 : _GEN_8868; // @[Rob.scala 1222:23]
  wire  _GEN_9125 = io_writeback_1_1_valid ? _GEN_8997 : _GEN_8869; // @[Rob.scala 1222:23]
  wire  _GEN_9126 = io_writeback_1_1_valid ? _GEN_8998 : _GEN_8870; // @[Rob.scala 1222:23]
  wire  _GEN_9127 = io_writeback_1_1_valid ? _GEN_8999 : _GEN_8871; // @[Rob.scala 1222:23]
  wire  _GEN_9128 = io_writeback_1_1_valid ? _GEN_9000 : _GEN_8872; // @[Rob.scala 1222:23]
  wire  _GEN_9129 = io_writeback_1_1_valid ? _GEN_9001 : _GEN_8873; // @[Rob.scala 1222:23]
  wire  _GEN_9130 = io_writeback_1_1_valid ? _GEN_9002 : _GEN_8874; // @[Rob.scala 1222:23]
  wire  _GEN_9131 = io_writeback_1_1_valid ? _GEN_9003 : _GEN_8875; // @[Rob.scala 1222:23]
  wire  _GEN_9132 = io_writeback_1_1_valid ? _GEN_9004 : _GEN_8876; // @[Rob.scala 1222:23]
  wire  _GEN_9133 = io_writeback_1_1_valid ? _GEN_9005 : _GEN_8877; // @[Rob.scala 1222:23]
  wire  _GEN_9134 = io_writeback_1_1_valid ? _GEN_9006 : _GEN_8878; // @[Rob.scala 1222:23]
  wire  _GEN_9135 = io_writeback_1_1_valid ? _GEN_9007 : _GEN_8879; // @[Rob.scala 1222:23]
  wire  _GEN_9136 = io_writeback_1_1_valid ? _GEN_9008 : _GEN_8880; // @[Rob.scala 1222:23]
  wire  _GEN_9137 = io_writeback_1_1_valid ? _GEN_9009 : _GEN_8881; // @[Rob.scala 1222:23]
  wire  _GEN_9138 = io_writeback_1_1_valid ? _GEN_9010 : _GEN_8882; // @[Rob.scala 1222:23]
  wire  _GEN_9139 = io_writeback_1_1_valid ? _GEN_9011 : _GEN_8883; // @[Rob.scala 1222:23]
  wire  _GEN_9140 = io_writeback_1_1_valid ? _GEN_9012 : _GEN_8884; // @[Rob.scala 1222:23]
  wire  _GEN_9141 = io_writeback_1_1_valid ? _GEN_9013 : _GEN_8885; // @[Rob.scala 1222:23]
  wire  _GEN_9142 = io_writeback_1_1_valid ? _GEN_9014 : _GEN_8886; // @[Rob.scala 1222:23]
  wire  _GEN_9143 = io_writeback_1_1_valid ? _GEN_9015 : _GEN_8887; // @[Rob.scala 1222:23]
  wire  _GEN_9144 = io_writeback_1_1_valid ? _GEN_9016 : _GEN_8888; // @[Rob.scala 1222:23]
  wire  _GEN_9145 = io_writeback_1_1_valid ? _GEN_9017 : _GEN_8889; // @[Rob.scala 1222:23]
  wire  _GEN_9146 = io_writeback_1_1_valid ? _GEN_9018 : _GEN_8890; // @[Rob.scala 1222:23]
  wire  _GEN_9147 = io_writeback_1_1_valid ? _GEN_9019 : _GEN_8891; // @[Rob.scala 1222:23]
  wire  _GEN_9148 = io_writeback_1_1_valid ? _GEN_9020 : _GEN_8892; // @[Rob.scala 1222:23]
  wire  _GEN_9149 = io_writeback_1_1_valid ? _GEN_9021 : _GEN_8893; // @[Rob.scala 1222:23]
  wire  _GEN_9150 = io_writeback_1_1_valid ? _GEN_9022 : _GEN_8894; // @[Rob.scala 1222:23]
  wire  _GEN_9151 = io_writeback_1_1_valid ? _GEN_9023 : _GEN_8895; // @[Rob.scala 1222:23]
  wire  _GEN_9152 = io_writeback_1_1_valid ? _GEN_9024 : _GEN_8896; // @[Rob.scala 1222:23]
  wire  _GEN_9153 = io_writeback_1_1_valid ? _GEN_9025 : _GEN_8897; // @[Rob.scala 1222:23]
  wire  _GEN_9154 = io_writeback_1_1_valid ? _GEN_9026 : _GEN_8898; // @[Rob.scala 1222:23]
  wire  _GEN_9155 = io_writeback_1_1_valid ? _GEN_9027 : _GEN_8899; // @[Rob.scala 1222:23]
  wire  _GEN_9156 = io_writeback_1_1_valid ? _GEN_9028 : _GEN_8900; // @[Rob.scala 1222:23]
  wire  _GEN_9157 = io_writeback_1_1_valid ? _GEN_9029 : _GEN_8901; // @[Rob.scala 1222:23]
  wire  _GEN_9158 = io_writeback_1_1_valid ? _GEN_9030 : _GEN_8902; // @[Rob.scala 1222:23]
  wire  _GEN_9159 = io_writeback_1_1_valid ? _GEN_9031 : _GEN_8903; // @[Rob.scala 1222:23]
  wire  _GEN_9160 = io_writeback_1_1_valid ? _GEN_9032 : _GEN_8904; // @[Rob.scala 1222:23]
  wire  _GEN_9161 = io_writeback_1_1_valid ? _GEN_9033 : _GEN_8905; // @[Rob.scala 1222:23]
  wire  _GEN_9162 = io_writeback_1_1_valid ? _GEN_9034 : _GEN_8906; // @[Rob.scala 1222:23]
  wire  _GEN_9227 = 5'h0 == io_writeback_1_2_bits_uop_robIdx_value ? io_writeback_1_2_bits_debug_isMMIO : _GEN_9099; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9228 = 5'h1 == io_writeback_1_2_bits_uop_robIdx_value ? io_writeback_1_2_bits_debug_isMMIO : _GEN_9100; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9229 = 5'h2 == io_writeback_1_2_bits_uop_robIdx_value ? io_writeback_1_2_bits_debug_isMMIO : _GEN_9101; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9230 = 5'h3 == io_writeback_1_2_bits_uop_robIdx_value ? io_writeback_1_2_bits_debug_isMMIO : _GEN_9102; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9231 = 5'h4 == io_writeback_1_2_bits_uop_robIdx_value ? io_writeback_1_2_bits_debug_isMMIO : _GEN_9103; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9232 = 5'h5 == io_writeback_1_2_bits_uop_robIdx_value ? io_writeback_1_2_bits_debug_isMMIO : _GEN_9104; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9233 = 5'h6 == io_writeback_1_2_bits_uop_robIdx_value ? io_writeback_1_2_bits_debug_isMMIO : _GEN_9105; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9234 = 5'h7 == io_writeback_1_2_bits_uop_robIdx_value ? io_writeback_1_2_bits_debug_isMMIO : _GEN_9106; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9235 = 5'h8 == io_writeback_1_2_bits_uop_robIdx_value ? io_writeback_1_2_bits_debug_isMMIO : _GEN_9107; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9236 = 5'h9 == io_writeback_1_2_bits_uop_robIdx_value ? io_writeback_1_2_bits_debug_isMMIO : _GEN_9108; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9237 = 5'ha == io_writeback_1_2_bits_uop_robIdx_value ? io_writeback_1_2_bits_debug_isMMIO : _GEN_9109; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9238 = 5'hb == io_writeback_1_2_bits_uop_robIdx_value ? io_writeback_1_2_bits_debug_isMMIO : _GEN_9110; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9239 = 5'hc == io_writeback_1_2_bits_uop_robIdx_value ? io_writeback_1_2_bits_debug_isMMIO : _GEN_9111; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9240 = 5'hd == io_writeback_1_2_bits_uop_robIdx_value ? io_writeback_1_2_bits_debug_isMMIO : _GEN_9112; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9241 = 5'he == io_writeback_1_2_bits_uop_robIdx_value ? io_writeback_1_2_bits_debug_isMMIO : _GEN_9113; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9242 = 5'hf == io_writeback_1_2_bits_uop_robIdx_value ? io_writeback_1_2_bits_debug_isMMIO : _GEN_9114; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9243 = 5'h10 == io_writeback_1_2_bits_uop_robIdx_value ? io_writeback_1_2_bits_debug_isMMIO : _GEN_9115; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9244 = 5'h11 == io_writeback_1_2_bits_uop_robIdx_value ? io_writeback_1_2_bits_debug_isMMIO : _GEN_9116; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9245 = 5'h12 == io_writeback_1_2_bits_uop_robIdx_value ? io_writeback_1_2_bits_debug_isMMIO : _GEN_9117; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9246 = 5'h13 == io_writeback_1_2_bits_uop_robIdx_value ? io_writeback_1_2_bits_debug_isMMIO : _GEN_9118; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9247 = 5'h14 == io_writeback_1_2_bits_uop_robIdx_value ? io_writeback_1_2_bits_debug_isMMIO : _GEN_9119; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9248 = 5'h15 == io_writeback_1_2_bits_uop_robIdx_value ? io_writeback_1_2_bits_debug_isMMIO : _GEN_9120; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9249 = 5'h16 == io_writeback_1_2_bits_uop_robIdx_value ? io_writeback_1_2_bits_debug_isMMIO : _GEN_9121; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9250 = 5'h17 == io_writeback_1_2_bits_uop_robIdx_value ? io_writeback_1_2_bits_debug_isMMIO : _GEN_9122; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9251 = 5'h18 == io_writeback_1_2_bits_uop_robIdx_value ? io_writeback_1_2_bits_debug_isMMIO : _GEN_9123; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9252 = 5'h19 == io_writeback_1_2_bits_uop_robIdx_value ? io_writeback_1_2_bits_debug_isMMIO : _GEN_9124; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9253 = 5'h1a == io_writeback_1_2_bits_uop_robIdx_value ? io_writeback_1_2_bits_debug_isMMIO : _GEN_9125; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9254 = 5'h1b == io_writeback_1_2_bits_uop_robIdx_value ? io_writeback_1_2_bits_debug_isMMIO : _GEN_9126; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9255 = 5'h1c == io_writeback_1_2_bits_uop_robIdx_value ? io_writeback_1_2_bits_debug_isMMIO : _GEN_9127; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9256 = 5'h1d == io_writeback_1_2_bits_uop_robIdx_value ? io_writeback_1_2_bits_debug_isMMIO : _GEN_9128; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9257 = 5'h1e == io_writeback_1_2_bits_uop_robIdx_value ? io_writeback_1_2_bits_debug_isMMIO : _GEN_9129; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9258 = 5'h1f == io_writeback_1_2_bits_uop_robIdx_value ? io_writeback_1_2_bits_debug_isMMIO : _GEN_9130; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9259 = 5'h0 == io_writeback_1_2_bits_uop_robIdx_value ? 1'h0 : _GEN_9131; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9260 = 5'h1 == io_writeback_1_2_bits_uop_robIdx_value ? 1'h0 : _GEN_9132; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9261 = 5'h2 == io_writeback_1_2_bits_uop_robIdx_value ? 1'h0 : _GEN_9133; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9262 = 5'h3 == io_writeback_1_2_bits_uop_robIdx_value ? 1'h0 : _GEN_9134; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9263 = 5'h4 == io_writeback_1_2_bits_uop_robIdx_value ? 1'h0 : _GEN_9135; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9264 = 5'h5 == io_writeback_1_2_bits_uop_robIdx_value ? 1'h0 : _GEN_9136; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9265 = 5'h6 == io_writeback_1_2_bits_uop_robIdx_value ? 1'h0 : _GEN_9137; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9266 = 5'h7 == io_writeback_1_2_bits_uop_robIdx_value ? 1'h0 : _GEN_9138; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9267 = 5'h8 == io_writeback_1_2_bits_uop_robIdx_value ? 1'h0 : _GEN_9139; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9268 = 5'h9 == io_writeback_1_2_bits_uop_robIdx_value ? 1'h0 : _GEN_9140; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9269 = 5'ha == io_writeback_1_2_bits_uop_robIdx_value ? 1'h0 : _GEN_9141; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9270 = 5'hb == io_writeback_1_2_bits_uop_robIdx_value ? 1'h0 : _GEN_9142; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9271 = 5'hc == io_writeback_1_2_bits_uop_robIdx_value ? 1'h0 : _GEN_9143; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9272 = 5'hd == io_writeback_1_2_bits_uop_robIdx_value ? 1'h0 : _GEN_9144; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9273 = 5'he == io_writeback_1_2_bits_uop_robIdx_value ? 1'h0 : _GEN_9145; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9274 = 5'hf == io_writeback_1_2_bits_uop_robIdx_value ? 1'h0 : _GEN_9146; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9275 = 5'h10 == io_writeback_1_2_bits_uop_robIdx_value ? 1'h0 : _GEN_9147; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9276 = 5'h11 == io_writeback_1_2_bits_uop_robIdx_value ? 1'h0 : _GEN_9148; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9277 = 5'h12 == io_writeback_1_2_bits_uop_robIdx_value ? 1'h0 : _GEN_9149; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9278 = 5'h13 == io_writeback_1_2_bits_uop_robIdx_value ? 1'h0 : _GEN_9150; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9279 = 5'h14 == io_writeback_1_2_bits_uop_robIdx_value ? 1'h0 : _GEN_9151; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9280 = 5'h15 == io_writeback_1_2_bits_uop_robIdx_value ? 1'h0 : _GEN_9152; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9281 = 5'h16 == io_writeback_1_2_bits_uop_robIdx_value ? 1'h0 : _GEN_9153; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9282 = 5'h17 == io_writeback_1_2_bits_uop_robIdx_value ? 1'h0 : _GEN_9154; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9283 = 5'h18 == io_writeback_1_2_bits_uop_robIdx_value ? 1'h0 : _GEN_9155; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9284 = 5'h19 == io_writeback_1_2_bits_uop_robIdx_value ? 1'h0 : _GEN_9156; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9285 = 5'h1a == io_writeback_1_2_bits_uop_robIdx_value ? 1'h0 : _GEN_9157; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9286 = 5'h1b == io_writeback_1_2_bits_uop_robIdx_value ? 1'h0 : _GEN_9158; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9287 = 5'h1c == io_writeback_1_2_bits_uop_robIdx_value ? 1'h0 : _GEN_9159; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9288 = 5'h1d == io_writeback_1_2_bits_uop_robIdx_value ? 1'h0 : _GEN_9160; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9289 = 5'h1e == io_writeback_1_2_bits_uop_robIdx_value ? 1'h0 : _GEN_9161; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9290 = 5'h1f == io_writeback_1_2_bits_uop_robIdx_value ? 1'h0 : _GEN_9162; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9355 = io_writeback_1_2_valid ? _GEN_9227 : _GEN_9099; // @[Rob.scala 1222:23]
  wire  _GEN_9356 = io_writeback_1_2_valid ? _GEN_9228 : _GEN_9100; // @[Rob.scala 1222:23]
  wire  _GEN_9357 = io_writeback_1_2_valid ? _GEN_9229 : _GEN_9101; // @[Rob.scala 1222:23]
  wire  _GEN_9358 = io_writeback_1_2_valid ? _GEN_9230 : _GEN_9102; // @[Rob.scala 1222:23]
  wire  _GEN_9359 = io_writeback_1_2_valid ? _GEN_9231 : _GEN_9103; // @[Rob.scala 1222:23]
  wire  _GEN_9360 = io_writeback_1_2_valid ? _GEN_9232 : _GEN_9104; // @[Rob.scala 1222:23]
  wire  _GEN_9361 = io_writeback_1_2_valid ? _GEN_9233 : _GEN_9105; // @[Rob.scala 1222:23]
  wire  _GEN_9362 = io_writeback_1_2_valid ? _GEN_9234 : _GEN_9106; // @[Rob.scala 1222:23]
  wire  _GEN_9363 = io_writeback_1_2_valid ? _GEN_9235 : _GEN_9107; // @[Rob.scala 1222:23]
  wire  _GEN_9364 = io_writeback_1_2_valid ? _GEN_9236 : _GEN_9108; // @[Rob.scala 1222:23]
  wire  _GEN_9365 = io_writeback_1_2_valid ? _GEN_9237 : _GEN_9109; // @[Rob.scala 1222:23]
  wire  _GEN_9366 = io_writeback_1_2_valid ? _GEN_9238 : _GEN_9110; // @[Rob.scala 1222:23]
  wire  _GEN_9367 = io_writeback_1_2_valid ? _GEN_9239 : _GEN_9111; // @[Rob.scala 1222:23]
  wire  _GEN_9368 = io_writeback_1_2_valid ? _GEN_9240 : _GEN_9112; // @[Rob.scala 1222:23]
  wire  _GEN_9369 = io_writeback_1_2_valid ? _GEN_9241 : _GEN_9113; // @[Rob.scala 1222:23]
  wire  _GEN_9370 = io_writeback_1_2_valid ? _GEN_9242 : _GEN_9114; // @[Rob.scala 1222:23]
  wire  _GEN_9371 = io_writeback_1_2_valid ? _GEN_9243 : _GEN_9115; // @[Rob.scala 1222:23]
  wire  _GEN_9372 = io_writeback_1_2_valid ? _GEN_9244 : _GEN_9116; // @[Rob.scala 1222:23]
  wire  _GEN_9373 = io_writeback_1_2_valid ? _GEN_9245 : _GEN_9117; // @[Rob.scala 1222:23]
  wire  _GEN_9374 = io_writeback_1_2_valid ? _GEN_9246 : _GEN_9118; // @[Rob.scala 1222:23]
  wire  _GEN_9375 = io_writeback_1_2_valid ? _GEN_9247 : _GEN_9119; // @[Rob.scala 1222:23]
  wire  _GEN_9376 = io_writeback_1_2_valid ? _GEN_9248 : _GEN_9120; // @[Rob.scala 1222:23]
  wire  _GEN_9377 = io_writeback_1_2_valid ? _GEN_9249 : _GEN_9121; // @[Rob.scala 1222:23]
  wire  _GEN_9378 = io_writeback_1_2_valid ? _GEN_9250 : _GEN_9122; // @[Rob.scala 1222:23]
  wire  _GEN_9379 = io_writeback_1_2_valid ? _GEN_9251 : _GEN_9123; // @[Rob.scala 1222:23]
  wire  _GEN_9380 = io_writeback_1_2_valid ? _GEN_9252 : _GEN_9124; // @[Rob.scala 1222:23]
  wire  _GEN_9381 = io_writeback_1_2_valid ? _GEN_9253 : _GEN_9125; // @[Rob.scala 1222:23]
  wire  _GEN_9382 = io_writeback_1_2_valid ? _GEN_9254 : _GEN_9126; // @[Rob.scala 1222:23]
  wire  _GEN_9383 = io_writeback_1_2_valid ? _GEN_9255 : _GEN_9127; // @[Rob.scala 1222:23]
  wire  _GEN_9384 = io_writeback_1_2_valid ? _GEN_9256 : _GEN_9128; // @[Rob.scala 1222:23]
  wire  _GEN_9385 = io_writeback_1_2_valid ? _GEN_9257 : _GEN_9129; // @[Rob.scala 1222:23]
  wire  _GEN_9386 = io_writeback_1_2_valid ? _GEN_9258 : _GEN_9130; // @[Rob.scala 1222:23]
  wire  _GEN_9387 = io_writeback_1_2_valid ? _GEN_9259 : _GEN_9131; // @[Rob.scala 1222:23]
  wire  _GEN_9388 = io_writeback_1_2_valid ? _GEN_9260 : _GEN_9132; // @[Rob.scala 1222:23]
  wire  _GEN_9389 = io_writeback_1_2_valid ? _GEN_9261 : _GEN_9133; // @[Rob.scala 1222:23]
  wire  _GEN_9390 = io_writeback_1_2_valid ? _GEN_9262 : _GEN_9134; // @[Rob.scala 1222:23]
  wire  _GEN_9391 = io_writeback_1_2_valid ? _GEN_9263 : _GEN_9135; // @[Rob.scala 1222:23]
  wire  _GEN_9392 = io_writeback_1_2_valid ? _GEN_9264 : _GEN_9136; // @[Rob.scala 1222:23]
  wire  _GEN_9393 = io_writeback_1_2_valid ? _GEN_9265 : _GEN_9137; // @[Rob.scala 1222:23]
  wire  _GEN_9394 = io_writeback_1_2_valid ? _GEN_9266 : _GEN_9138; // @[Rob.scala 1222:23]
  wire  _GEN_9395 = io_writeback_1_2_valid ? _GEN_9267 : _GEN_9139; // @[Rob.scala 1222:23]
  wire  _GEN_9396 = io_writeback_1_2_valid ? _GEN_9268 : _GEN_9140; // @[Rob.scala 1222:23]
  wire  _GEN_9397 = io_writeback_1_2_valid ? _GEN_9269 : _GEN_9141; // @[Rob.scala 1222:23]
  wire  _GEN_9398 = io_writeback_1_2_valid ? _GEN_9270 : _GEN_9142; // @[Rob.scala 1222:23]
  wire  _GEN_9399 = io_writeback_1_2_valid ? _GEN_9271 : _GEN_9143; // @[Rob.scala 1222:23]
  wire  _GEN_9400 = io_writeback_1_2_valid ? _GEN_9272 : _GEN_9144; // @[Rob.scala 1222:23]
  wire  _GEN_9401 = io_writeback_1_2_valid ? _GEN_9273 : _GEN_9145; // @[Rob.scala 1222:23]
  wire  _GEN_9402 = io_writeback_1_2_valid ? _GEN_9274 : _GEN_9146; // @[Rob.scala 1222:23]
  wire  _GEN_9403 = io_writeback_1_2_valid ? _GEN_9275 : _GEN_9147; // @[Rob.scala 1222:23]
  wire  _GEN_9404 = io_writeback_1_2_valid ? _GEN_9276 : _GEN_9148; // @[Rob.scala 1222:23]
  wire  _GEN_9405 = io_writeback_1_2_valid ? _GEN_9277 : _GEN_9149; // @[Rob.scala 1222:23]
  wire  _GEN_9406 = io_writeback_1_2_valid ? _GEN_9278 : _GEN_9150; // @[Rob.scala 1222:23]
  wire  _GEN_9407 = io_writeback_1_2_valid ? _GEN_9279 : _GEN_9151; // @[Rob.scala 1222:23]
  wire  _GEN_9408 = io_writeback_1_2_valid ? _GEN_9280 : _GEN_9152; // @[Rob.scala 1222:23]
  wire  _GEN_9409 = io_writeback_1_2_valid ? _GEN_9281 : _GEN_9153; // @[Rob.scala 1222:23]
  wire  _GEN_9410 = io_writeback_1_2_valid ? _GEN_9282 : _GEN_9154; // @[Rob.scala 1222:23]
  wire  _GEN_9411 = io_writeback_1_2_valid ? _GEN_9283 : _GEN_9155; // @[Rob.scala 1222:23]
  wire  _GEN_9412 = io_writeback_1_2_valid ? _GEN_9284 : _GEN_9156; // @[Rob.scala 1222:23]
  wire  _GEN_9413 = io_writeback_1_2_valid ? _GEN_9285 : _GEN_9157; // @[Rob.scala 1222:23]
  wire  _GEN_9414 = io_writeback_1_2_valid ? _GEN_9286 : _GEN_9158; // @[Rob.scala 1222:23]
  wire  _GEN_9415 = io_writeback_1_2_valid ? _GEN_9287 : _GEN_9159; // @[Rob.scala 1222:23]
  wire  _GEN_9416 = io_writeback_1_2_valid ? _GEN_9288 : _GEN_9160; // @[Rob.scala 1222:23]
  wire  _GEN_9417 = io_writeback_1_2_valid ? _GEN_9289 : _GEN_9161; // @[Rob.scala 1222:23]
  wire  _GEN_9418 = io_writeback_1_2_valid ? _GEN_9290 : _GEN_9162; // @[Rob.scala 1222:23]
  wire  _GEN_9483 = 5'h0 == io_writeback_1_3_bits_uop_robIdx_value ? io_writeback_1_3_bits_debug_isMMIO : _GEN_9355; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9484 = 5'h1 == io_writeback_1_3_bits_uop_robIdx_value ? io_writeback_1_3_bits_debug_isMMIO : _GEN_9356; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9485 = 5'h2 == io_writeback_1_3_bits_uop_robIdx_value ? io_writeback_1_3_bits_debug_isMMIO : _GEN_9357; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9486 = 5'h3 == io_writeback_1_3_bits_uop_robIdx_value ? io_writeback_1_3_bits_debug_isMMIO : _GEN_9358; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9487 = 5'h4 == io_writeback_1_3_bits_uop_robIdx_value ? io_writeback_1_3_bits_debug_isMMIO : _GEN_9359; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9488 = 5'h5 == io_writeback_1_3_bits_uop_robIdx_value ? io_writeback_1_3_bits_debug_isMMIO : _GEN_9360; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9489 = 5'h6 == io_writeback_1_3_bits_uop_robIdx_value ? io_writeback_1_3_bits_debug_isMMIO : _GEN_9361; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9490 = 5'h7 == io_writeback_1_3_bits_uop_robIdx_value ? io_writeback_1_3_bits_debug_isMMIO : _GEN_9362; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9491 = 5'h8 == io_writeback_1_3_bits_uop_robIdx_value ? io_writeback_1_3_bits_debug_isMMIO : _GEN_9363; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9492 = 5'h9 == io_writeback_1_3_bits_uop_robIdx_value ? io_writeback_1_3_bits_debug_isMMIO : _GEN_9364; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9493 = 5'ha == io_writeback_1_3_bits_uop_robIdx_value ? io_writeback_1_3_bits_debug_isMMIO : _GEN_9365; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9494 = 5'hb == io_writeback_1_3_bits_uop_robIdx_value ? io_writeback_1_3_bits_debug_isMMIO : _GEN_9366; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9495 = 5'hc == io_writeback_1_3_bits_uop_robIdx_value ? io_writeback_1_3_bits_debug_isMMIO : _GEN_9367; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9496 = 5'hd == io_writeback_1_3_bits_uop_robIdx_value ? io_writeback_1_3_bits_debug_isMMIO : _GEN_9368; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9497 = 5'he == io_writeback_1_3_bits_uop_robIdx_value ? io_writeback_1_3_bits_debug_isMMIO : _GEN_9369; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9498 = 5'hf == io_writeback_1_3_bits_uop_robIdx_value ? io_writeback_1_3_bits_debug_isMMIO : _GEN_9370; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9499 = 5'h10 == io_writeback_1_3_bits_uop_robIdx_value ? io_writeback_1_3_bits_debug_isMMIO : _GEN_9371; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9500 = 5'h11 == io_writeback_1_3_bits_uop_robIdx_value ? io_writeback_1_3_bits_debug_isMMIO : _GEN_9372; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9501 = 5'h12 == io_writeback_1_3_bits_uop_robIdx_value ? io_writeback_1_3_bits_debug_isMMIO : _GEN_9373; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9502 = 5'h13 == io_writeback_1_3_bits_uop_robIdx_value ? io_writeback_1_3_bits_debug_isMMIO : _GEN_9374; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9503 = 5'h14 == io_writeback_1_3_bits_uop_robIdx_value ? io_writeback_1_3_bits_debug_isMMIO : _GEN_9375; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9504 = 5'h15 == io_writeback_1_3_bits_uop_robIdx_value ? io_writeback_1_3_bits_debug_isMMIO : _GEN_9376; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9505 = 5'h16 == io_writeback_1_3_bits_uop_robIdx_value ? io_writeback_1_3_bits_debug_isMMIO : _GEN_9377; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9506 = 5'h17 == io_writeback_1_3_bits_uop_robIdx_value ? io_writeback_1_3_bits_debug_isMMIO : _GEN_9378; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9507 = 5'h18 == io_writeback_1_3_bits_uop_robIdx_value ? io_writeback_1_3_bits_debug_isMMIO : _GEN_9379; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9508 = 5'h19 == io_writeback_1_3_bits_uop_robIdx_value ? io_writeback_1_3_bits_debug_isMMIO : _GEN_9380; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9509 = 5'h1a == io_writeback_1_3_bits_uop_robIdx_value ? io_writeback_1_3_bits_debug_isMMIO : _GEN_9381; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9510 = 5'h1b == io_writeback_1_3_bits_uop_robIdx_value ? io_writeback_1_3_bits_debug_isMMIO : _GEN_9382; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9511 = 5'h1c == io_writeback_1_3_bits_uop_robIdx_value ? io_writeback_1_3_bits_debug_isMMIO : _GEN_9383; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9512 = 5'h1d == io_writeback_1_3_bits_uop_robIdx_value ? io_writeback_1_3_bits_debug_isMMIO : _GEN_9384; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9513 = 5'h1e == io_writeback_1_3_bits_uop_robIdx_value ? io_writeback_1_3_bits_debug_isMMIO : _GEN_9385; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9514 = 5'h1f == io_writeback_1_3_bits_uop_robIdx_value ? io_writeback_1_3_bits_debug_isMMIO : _GEN_9386; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9515 = 5'h0 == io_writeback_1_3_bits_uop_robIdx_value ? 1'h0 : _GEN_9387; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9516 = 5'h1 == io_writeback_1_3_bits_uop_robIdx_value ? 1'h0 : _GEN_9388; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9517 = 5'h2 == io_writeback_1_3_bits_uop_robIdx_value ? 1'h0 : _GEN_9389; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9518 = 5'h3 == io_writeback_1_3_bits_uop_robIdx_value ? 1'h0 : _GEN_9390; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9519 = 5'h4 == io_writeback_1_3_bits_uop_robIdx_value ? 1'h0 : _GEN_9391; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9520 = 5'h5 == io_writeback_1_3_bits_uop_robIdx_value ? 1'h0 : _GEN_9392; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9521 = 5'h6 == io_writeback_1_3_bits_uop_robIdx_value ? 1'h0 : _GEN_9393; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9522 = 5'h7 == io_writeback_1_3_bits_uop_robIdx_value ? 1'h0 : _GEN_9394; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9523 = 5'h8 == io_writeback_1_3_bits_uop_robIdx_value ? 1'h0 : _GEN_9395; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9524 = 5'h9 == io_writeback_1_3_bits_uop_robIdx_value ? 1'h0 : _GEN_9396; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9525 = 5'ha == io_writeback_1_3_bits_uop_robIdx_value ? 1'h0 : _GEN_9397; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9526 = 5'hb == io_writeback_1_3_bits_uop_robIdx_value ? 1'h0 : _GEN_9398; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9527 = 5'hc == io_writeback_1_3_bits_uop_robIdx_value ? 1'h0 : _GEN_9399; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9528 = 5'hd == io_writeback_1_3_bits_uop_robIdx_value ? 1'h0 : _GEN_9400; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9529 = 5'he == io_writeback_1_3_bits_uop_robIdx_value ? 1'h0 : _GEN_9401; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9530 = 5'hf == io_writeback_1_3_bits_uop_robIdx_value ? 1'h0 : _GEN_9402; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9531 = 5'h10 == io_writeback_1_3_bits_uop_robIdx_value ? 1'h0 : _GEN_9403; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9532 = 5'h11 == io_writeback_1_3_bits_uop_robIdx_value ? 1'h0 : _GEN_9404; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9533 = 5'h12 == io_writeback_1_3_bits_uop_robIdx_value ? 1'h0 : _GEN_9405; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9534 = 5'h13 == io_writeback_1_3_bits_uop_robIdx_value ? 1'h0 : _GEN_9406; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9535 = 5'h14 == io_writeback_1_3_bits_uop_robIdx_value ? 1'h0 : _GEN_9407; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9536 = 5'h15 == io_writeback_1_3_bits_uop_robIdx_value ? 1'h0 : _GEN_9408; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9537 = 5'h16 == io_writeback_1_3_bits_uop_robIdx_value ? 1'h0 : _GEN_9409; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9538 = 5'h17 == io_writeback_1_3_bits_uop_robIdx_value ? 1'h0 : _GEN_9410; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9539 = 5'h18 == io_writeback_1_3_bits_uop_robIdx_value ? 1'h0 : _GEN_9411; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9540 = 5'h19 == io_writeback_1_3_bits_uop_robIdx_value ? 1'h0 : _GEN_9412; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9541 = 5'h1a == io_writeback_1_3_bits_uop_robIdx_value ? 1'h0 : _GEN_9413; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9542 = 5'h1b == io_writeback_1_3_bits_uop_robIdx_value ? 1'h0 : _GEN_9414; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9543 = 5'h1c == io_writeback_1_3_bits_uop_robIdx_value ? 1'h0 : _GEN_9415; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9544 = 5'h1d == io_writeback_1_3_bits_uop_robIdx_value ? 1'h0 : _GEN_9416; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9545 = 5'h1e == io_writeback_1_3_bits_uop_robIdx_value ? 1'h0 : _GEN_9417; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9546 = 5'h1f == io_writeback_1_3_bits_uop_robIdx_value ? 1'h0 : _GEN_9418; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9611 = io_writeback_1_3_valid ? _GEN_9483 : _GEN_9355; // @[Rob.scala 1222:23]
  wire  _GEN_9612 = io_writeback_1_3_valid ? _GEN_9484 : _GEN_9356; // @[Rob.scala 1222:23]
  wire  _GEN_9613 = io_writeback_1_3_valid ? _GEN_9485 : _GEN_9357; // @[Rob.scala 1222:23]
  wire  _GEN_9614 = io_writeback_1_3_valid ? _GEN_9486 : _GEN_9358; // @[Rob.scala 1222:23]
  wire  _GEN_9615 = io_writeback_1_3_valid ? _GEN_9487 : _GEN_9359; // @[Rob.scala 1222:23]
  wire  _GEN_9616 = io_writeback_1_3_valid ? _GEN_9488 : _GEN_9360; // @[Rob.scala 1222:23]
  wire  _GEN_9617 = io_writeback_1_3_valid ? _GEN_9489 : _GEN_9361; // @[Rob.scala 1222:23]
  wire  _GEN_9618 = io_writeback_1_3_valid ? _GEN_9490 : _GEN_9362; // @[Rob.scala 1222:23]
  wire  _GEN_9619 = io_writeback_1_3_valid ? _GEN_9491 : _GEN_9363; // @[Rob.scala 1222:23]
  wire  _GEN_9620 = io_writeback_1_3_valid ? _GEN_9492 : _GEN_9364; // @[Rob.scala 1222:23]
  wire  _GEN_9621 = io_writeback_1_3_valid ? _GEN_9493 : _GEN_9365; // @[Rob.scala 1222:23]
  wire  _GEN_9622 = io_writeback_1_3_valid ? _GEN_9494 : _GEN_9366; // @[Rob.scala 1222:23]
  wire  _GEN_9623 = io_writeback_1_3_valid ? _GEN_9495 : _GEN_9367; // @[Rob.scala 1222:23]
  wire  _GEN_9624 = io_writeback_1_3_valid ? _GEN_9496 : _GEN_9368; // @[Rob.scala 1222:23]
  wire  _GEN_9625 = io_writeback_1_3_valid ? _GEN_9497 : _GEN_9369; // @[Rob.scala 1222:23]
  wire  _GEN_9626 = io_writeback_1_3_valid ? _GEN_9498 : _GEN_9370; // @[Rob.scala 1222:23]
  wire  _GEN_9627 = io_writeback_1_3_valid ? _GEN_9499 : _GEN_9371; // @[Rob.scala 1222:23]
  wire  _GEN_9628 = io_writeback_1_3_valid ? _GEN_9500 : _GEN_9372; // @[Rob.scala 1222:23]
  wire  _GEN_9629 = io_writeback_1_3_valid ? _GEN_9501 : _GEN_9373; // @[Rob.scala 1222:23]
  wire  _GEN_9630 = io_writeback_1_3_valid ? _GEN_9502 : _GEN_9374; // @[Rob.scala 1222:23]
  wire  _GEN_9631 = io_writeback_1_3_valid ? _GEN_9503 : _GEN_9375; // @[Rob.scala 1222:23]
  wire  _GEN_9632 = io_writeback_1_3_valid ? _GEN_9504 : _GEN_9376; // @[Rob.scala 1222:23]
  wire  _GEN_9633 = io_writeback_1_3_valid ? _GEN_9505 : _GEN_9377; // @[Rob.scala 1222:23]
  wire  _GEN_9634 = io_writeback_1_3_valid ? _GEN_9506 : _GEN_9378; // @[Rob.scala 1222:23]
  wire  _GEN_9635 = io_writeback_1_3_valid ? _GEN_9507 : _GEN_9379; // @[Rob.scala 1222:23]
  wire  _GEN_9636 = io_writeback_1_3_valid ? _GEN_9508 : _GEN_9380; // @[Rob.scala 1222:23]
  wire  _GEN_9637 = io_writeback_1_3_valid ? _GEN_9509 : _GEN_9381; // @[Rob.scala 1222:23]
  wire  _GEN_9638 = io_writeback_1_3_valid ? _GEN_9510 : _GEN_9382; // @[Rob.scala 1222:23]
  wire  _GEN_9639 = io_writeback_1_3_valid ? _GEN_9511 : _GEN_9383; // @[Rob.scala 1222:23]
  wire  _GEN_9640 = io_writeback_1_3_valid ? _GEN_9512 : _GEN_9384; // @[Rob.scala 1222:23]
  wire  _GEN_9641 = io_writeback_1_3_valid ? _GEN_9513 : _GEN_9385; // @[Rob.scala 1222:23]
  wire  _GEN_9642 = io_writeback_1_3_valid ? _GEN_9514 : _GEN_9386; // @[Rob.scala 1222:23]
  wire  _GEN_9643 = io_writeback_1_3_valid ? _GEN_9515 : _GEN_9387; // @[Rob.scala 1222:23]
  wire  _GEN_9644 = io_writeback_1_3_valid ? _GEN_9516 : _GEN_9388; // @[Rob.scala 1222:23]
  wire  _GEN_9645 = io_writeback_1_3_valid ? _GEN_9517 : _GEN_9389; // @[Rob.scala 1222:23]
  wire  _GEN_9646 = io_writeback_1_3_valid ? _GEN_9518 : _GEN_9390; // @[Rob.scala 1222:23]
  wire  _GEN_9647 = io_writeback_1_3_valid ? _GEN_9519 : _GEN_9391; // @[Rob.scala 1222:23]
  wire  _GEN_9648 = io_writeback_1_3_valid ? _GEN_9520 : _GEN_9392; // @[Rob.scala 1222:23]
  wire  _GEN_9649 = io_writeback_1_3_valid ? _GEN_9521 : _GEN_9393; // @[Rob.scala 1222:23]
  wire  _GEN_9650 = io_writeback_1_3_valid ? _GEN_9522 : _GEN_9394; // @[Rob.scala 1222:23]
  wire  _GEN_9651 = io_writeback_1_3_valid ? _GEN_9523 : _GEN_9395; // @[Rob.scala 1222:23]
  wire  _GEN_9652 = io_writeback_1_3_valid ? _GEN_9524 : _GEN_9396; // @[Rob.scala 1222:23]
  wire  _GEN_9653 = io_writeback_1_3_valid ? _GEN_9525 : _GEN_9397; // @[Rob.scala 1222:23]
  wire  _GEN_9654 = io_writeback_1_3_valid ? _GEN_9526 : _GEN_9398; // @[Rob.scala 1222:23]
  wire  _GEN_9655 = io_writeback_1_3_valid ? _GEN_9527 : _GEN_9399; // @[Rob.scala 1222:23]
  wire  _GEN_9656 = io_writeback_1_3_valid ? _GEN_9528 : _GEN_9400; // @[Rob.scala 1222:23]
  wire  _GEN_9657 = io_writeback_1_3_valid ? _GEN_9529 : _GEN_9401; // @[Rob.scala 1222:23]
  wire  _GEN_9658 = io_writeback_1_3_valid ? _GEN_9530 : _GEN_9402; // @[Rob.scala 1222:23]
  wire  _GEN_9659 = io_writeback_1_3_valid ? _GEN_9531 : _GEN_9403; // @[Rob.scala 1222:23]
  wire  _GEN_9660 = io_writeback_1_3_valid ? _GEN_9532 : _GEN_9404; // @[Rob.scala 1222:23]
  wire  _GEN_9661 = io_writeback_1_3_valid ? _GEN_9533 : _GEN_9405; // @[Rob.scala 1222:23]
  wire  _GEN_9662 = io_writeback_1_3_valid ? _GEN_9534 : _GEN_9406; // @[Rob.scala 1222:23]
  wire  _GEN_9663 = io_writeback_1_3_valid ? _GEN_9535 : _GEN_9407; // @[Rob.scala 1222:23]
  wire  _GEN_9664 = io_writeback_1_3_valid ? _GEN_9536 : _GEN_9408; // @[Rob.scala 1222:23]
  wire  _GEN_9665 = io_writeback_1_3_valid ? _GEN_9537 : _GEN_9409; // @[Rob.scala 1222:23]
  wire  _GEN_9666 = io_writeback_1_3_valid ? _GEN_9538 : _GEN_9410; // @[Rob.scala 1222:23]
  wire  _GEN_9667 = io_writeback_1_3_valid ? _GEN_9539 : _GEN_9411; // @[Rob.scala 1222:23]
  wire  _GEN_9668 = io_writeback_1_3_valid ? _GEN_9540 : _GEN_9412; // @[Rob.scala 1222:23]
  wire  _GEN_9669 = io_writeback_1_3_valid ? _GEN_9541 : _GEN_9413; // @[Rob.scala 1222:23]
  wire  _GEN_9670 = io_writeback_1_3_valid ? _GEN_9542 : _GEN_9414; // @[Rob.scala 1222:23]
  wire  _GEN_9671 = io_writeback_1_3_valid ? _GEN_9543 : _GEN_9415; // @[Rob.scala 1222:23]
  wire  _GEN_9672 = io_writeback_1_3_valid ? _GEN_9544 : _GEN_9416; // @[Rob.scala 1222:23]
  wire  _GEN_9673 = io_writeback_1_3_valid ? _GEN_9545 : _GEN_9417; // @[Rob.scala 1222:23]
  wire  _GEN_9674 = io_writeback_1_3_valid ? _GEN_9546 : _GEN_9418; // @[Rob.scala 1222:23]
  wire  _GEN_9739 = 5'h0 == io_writeback_1_4_bits_uop_robIdx_value ? 1'h0 : _GEN_9611; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9740 = 5'h1 == io_writeback_1_4_bits_uop_robIdx_value ? 1'h0 : _GEN_9612; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9741 = 5'h2 == io_writeback_1_4_bits_uop_robIdx_value ? 1'h0 : _GEN_9613; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9742 = 5'h3 == io_writeback_1_4_bits_uop_robIdx_value ? 1'h0 : _GEN_9614; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9743 = 5'h4 == io_writeback_1_4_bits_uop_robIdx_value ? 1'h0 : _GEN_9615; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9744 = 5'h5 == io_writeback_1_4_bits_uop_robIdx_value ? 1'h0 : _GEN_9616; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9745 = 5'h6 == io_writeback_1_4_bits_uop_robIdx_value ? 1'h0 : _GEN_9617; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9746 = 5'h7 == io_writeback_1_4_bits_uop_robIdx_value ? 1'h0 : _GEN_9618; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9747 = 5'h8 == io_writeback_1_4_bits_uop_robIdx_value ? 1'h0 : _GEN_9619; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9748 = 5'h9 == io_writeback_1_4_bits_uop_robIdx_value ? 1'h0 : _GEN_9620; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9749 = 5'ha == io_writeback_1_4_bits_uop_robIdx_value ? 1'h0 : _GEN_9621; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9750 = 5'hb == io_writeback_1_4_bits_uop_robIdx_value ? 1'h0 : _GEN_9622; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9751 = 5'hc == io_writeback_1_4_bits_uop_robIdx_value ? 1'h0 : _GEN_9623; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9752 = 5'hd == io_writeback_1_4_bits_uop_robIdx_value ? 1'h0 : _GEN_9624; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9753 = 5'he == io_writeback_1_4_bits_uop_robIdx_value ? 1'h0 : _GEN_9625; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9754 = 5'hf == io_writeback_1_4_bits_uop_robIdx_value ? 1'h0 : _GEN_9626; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9755 = 5'h10 == io_writeback_1_4_bits_uop_robIdx_value ? 1'h0 : _GEN_9627; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9756 = 5'h11 == io_writeback_1_4_bits_uop_robIdx_value ? 1'h0 : _GEN_9628; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9757 = 5'h12 == io_writeback_1_4_bits_uop_robIdx_value ? 1'h0 : _GEN_9629; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9758 = 5'h13 == io_writeback_1_4_bits_uop_robIdx_value ? 1'h0 : _GEN_9630; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9759 = 5'h14 == io_writeback_1_4_bits_uop_robIdx_value ? 1'h0 : _GEN_9631; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9760 = 5'h15 == io_writeback_1_4_bits_uop_robIdx_value ? 1'h0 : _GEN_9632; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9761 = 5'h16 == io_writeback_1_4_bits_uop_robIdx_value ? 1'h0 : _GEN_9633; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9762 = 5'h17 == io_writeback_1_4_bits_uop_robIdx_value ? 1'h0 : _GEN_9634; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9763 = 5'h18 == io_writeback_1_4_bits_uop_robIdx_value ? 1'h0 : _GEN_9635; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9764 = 5'h19 == io_writeback_1_4_bits_uop_robIdx_value ? 1'h0 : _GEN_9636; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9765 = 5'h1a == io_writeback_1_4_bits_uop_robIdx_value ? 1'h0 : _GEN_9637; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9766 = 5'h1b == io_writeback_1_4_bits_uop_robIdx_value ? 1'h0 : _GEN_9638; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9767 = 5'h1c == io_writeback_1_4_bits_uop_robIdx_value ? 1'h0 : _GEN_9639; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9768 = 5'h1d == io_writeback_1_4_bits_uop_robIdx_value ? 1'h0 : _GEN_9640; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9769 = 5'h1e == io_writeback_1_4_bits_uop_robIdx_value ? 1'h0 : _GEN_9641; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9770 = 5'h1f == io_writeback_1_4_bits_uop_robIdx_value ? 1'h0 : _GEN_9642; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9771 = 5'h0 == io_writeback_1_4_bits_uop_robIdx_value ? io_writeback_1_4_bits_debug_isPerfCnt : _GEN_9643; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9772 = 5'h1 == io_writeback_1_4_bits_uop_robIdx_value ? io_writeback_1_4_bits_debug_isPerfCnt : _GEN_9644; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9773 = 5'h2 == io_writeback_1_4_bits_uop_robIdx_value ? io_writeback_1_4_bits_debug_isPerfCnt : _GEN_9645; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9774 = 5'h3 == io_writeback_1_4_bits_uop_robIdx_value ? io_writeback_1_4_bits_debug_isPerfCnt : _GEN_9646; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9775 = 5'h4 == io_writeback_1_4_bits_uop_robIdx_value ? io_writeback_1_4_bits_debug_isPerfCnt : _GEN_9647; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9776 = 5'h5 == io_writeback_1_4_bits_uop_robIdx_value ? io_writeback_1_4_bits_debug_isPerfCnt : _GEN_9648; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9777 = 5'h6 == io_writeback_1_4_bits_uop_robIdx_value ? io_writeback_1_4_bits_debug_isPerfCnt : _GEN_9649; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9778 = 5'h7 == io_writeback_1_4_bits_uop_robIdx_value ? io_writeback_1_4_bits_debug_isPerfCnt : _GEN_9650; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9779 = 5'h8 == io_writeback_1_4_bits_uop_robIdx_value ? io_writeback_1_4_bits_debug_isPerfCnt : _GEN_9651; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9780 = 5'h9 == io_writeback_1_4_bits_uop_robIdx_value ? io_writeback_1_4_bits_debug_isPerfCnt : _GEN_9652; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9781 = 5'ha == io_writeback_1_4_bits_uop_robIdx_value ? io_writeback_1_4_bits_debug_isPerfCnt : _GEN_9653; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9782 = 5'hb == io_writeback_1_4_bits_uop_robIdx_value ? io_writeback_1_4_bits_debug_isPerfCnt : _GEN_9654; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9783 = 5'hc == io_writeback_1_4_bits_uop_robIdx_value ? io_writeback_1_4_bits_debug_isPerfCnt : _GEN_9655; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9784 = 5'hd == io_writeback_1_4_bits_uop_robIdx_value ? io_writeback_1_4_bits_debug_isPerfCnt : _GEN_9656; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9785 = 5'he == io_writeback_1_4_bits_uop_robIdx_value ? io_writeback_1_4_bits_debug_isPerfCnt : _GEN_9657; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9786 = 5'hf == io_writeback_1_4_bits_uop_robIdx_value ? io_writeback_1_4_bits_debug_isPerfCnt : _GEN_9658; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9787 = 5'h10 == io_writeback_1_4_bits_uop_robIdx_value ? io_writeback_1_4_bits_debug_isPerfCnt : _GEN_9659; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9788 = 5'h11 == io_writeback_1_4_bits_uop_robIdx_value ? io_writeback_1_4_bits_debug_isPerfCnt : _GEN_9660; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9789 = 5'h12 == io_writeback_1_4_bits_uop_robIdx_value ? io_writeback_1_4_bits_debug_isPerfCnt : _GEN_9661; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9790 = 5'h13 == io_writeback_1_4_bits_uop_robIdx_value ? io_writeback_1_4_bits_debug_isPerfCnt : _GEN_9662; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9791 = 5'h14 == io_writeback_1_4_bits_uop_robIdx_value ? io_writeback_1_4_bits_debug_isPerfCnt : _GEN_9663; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9792 = 5'h15 == io_writeback_1_4_bits_uop_robIdx_value ? io_writeback_1_4_bits_debug_isPerfCnt : _GEN_9664; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9793 = 5'h16 == io_writeback_1_4_bits_uop_robIdx_value ? io_writeback_1_4_bits_debug_isPerfCnt : _GEN_9665; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9794 = 5'h17 == io_writeback_1_4_bits_uop_robIdx_value ? io_writeback_1_4_bits_debug_isPerfCnt : _GEN_9666; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9795 = 5'h18 == io_writeback_1_4_bits_uop_robIdx_value ? io_writeback_1_4_bits_debug_isPerfCnt : _GEN_9667; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9796 = 5'h19 == io_writeback_1_4_bits_uop_robIdx_value ? io_writeback_1_4_bits_debug_isPerfCnt : _GEN_9668; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9797 = 5'h1a == io_writeback_1_4_bits_uop_robIdx_value ? io_writeback_1_4_bits_debug_isPerfCnt : _GEN_9669; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9798 = 5'h1b == io_writeback_1_4_bits_uop_robIdx_value ? io_writeback_1_4_bits_debug_isPerfCnt : _GEN_9670; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9799 = 5'h1c == io_writeback_1_4_bits_uop_robIdx_value ? io_writeback_1_4_bits_debug_isPerfCnt : _GEN_9671; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9800 = 5'h1d == io_writeback_1_4_bits_uop_robIdx_value ? io_writeback_1_4_bits_debug_isPerfCnt : _GEN_9672; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9801 = 5'h1e == io_writeback_1_4_bits_uop_robIdx_value ? io_writeback_1_4_bits_debug_isPerfCnt : _GEN_9673; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9802 = 5'h1f == io_writeback_1_4_bits_uop_robIdx_value ? io_writeback_1_4_bits_debug_isPerfCnt : _GEN_9674; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9867 = io_writeback_1_4_valid ? _GEN_9739 : _GEN_9611; // @[Rob.scala 1222:23]
  wire  _GEN_9868 = io_writeback_1_4_valid ? _GEN_9740 : _GEN_9612; // @[Rob.scala 1222:23]
  wire  _GEN_9869 = io_writeback_1_4_valid ? _GEN_9741 : _GEN_9613; // @[Rob.scala 1222:23]
  wire  _GEN_9870 = io_writeback_1_4_valid ? _GEN_9742 : _GEN_9614; // @[Rob.scala 1222:23]
  wire  _GEN_9871 = io_writeback_1_4_valid ? _GEN_9743 : _GEN_9615; // @[Rob.scala 1222:23]
  wire  _GEN_9872 = io_writeback_1_4_valid ? _GEN_9744 : _GEN_9616; // @[Rob.scala 1222:23]
  wire  _GEN_9873 = io_writeback_1_4_valid ? _GEN_9745 : _GEN_9617; // @[Rob.scala 1222:23]
  wire  _GEN_9874 = io_writeback_1_4_valid ? _GEN_9746 : _GEN_9618; // @[Rob.scala 1222:23]
  wire  _GEN_9875 = io_writeback_1_4_valid ? _GEN_9747 : _GEN_9619; // @[Rob.scala 1222:23]
  wire  _GEN_9876 = io_writeback_1_4_valid ? _GEN_9748 : _GEN_9620; // @[Rob.scala 1222:23]
  wire  _GEN_9877 = io_writeback_1_4_valid ? _GEN_9749 : _GEN_9621; // @[Rob.scala 1222:23]
  wire  _GEN_9878 = io_writeback_1_4_valid ? _GEN_9750 : _GEN_9622; // @[Rob.scala 1222:23]
  wire  _GEN_9879 = io_writeback_1_4_valid ? _GEN_9751 : _GEN_9623; // @[Rob.scala 1222:23]
  wire  _GEN_9880 = io_writeback_1_4_valid ? _GEN_9752 : _GEN_9624; // @[Rob.scala 1222:23]
  wire  _GEN_9881 = io_writeback_1_4_valid ? _GEN_9753 : _GEN_9625; // @[Rob.scala 1222:23]
  wire  _GEN_9882 = io_writeback_1_4_valid ? _GEN_9754 : _GEN_9626; // @[Rob.scala 1222:23]
  wire  _GEN_9883 = io_writeback_1_4_valid ? _GEN_9755 : _GEN_9627; // @[Rob.scala 1222:23]
  wire  _GEN_9884 = io_writeback_1_4_valid ? _GEN_9756 : _GEN_9628; // @[Rob.scala 1222:23]
  wire  _GEN_9885 = io_writeback_1_4_valid ? _GEN_9757 : _GEN_9629; // @[Rob.scala 1222:23]
  wire  _GEN_9886 = io_writeback_1_4_valid ? _GEN_9758 : _GEN_9630; // @[Rob.scala 1222:23]
  wire  _GEN_9887 = io_writeback_1_4_valid ? _GEN_9759 : _GEN_9631; // @[Rob.scala 1222:23]
  wire  _GEN_9888 = io_writeback_1_4_valid ? _GEN_9760 : _GEN_9632; // @[Rob.scala 1222:23]
  wire  _GEN_9889 = io_writeback_1_4_valid ? _GEN_9761 : _GEN_9633; // @[Rob.scala 1222:23]
  wire  _GEN_9890 = io_writeback_1_4_valid ? _GEN_9762 : _GEN_9634; // @[Rob.scala 1222:23]
  wire  _GEN_9891 = io_writeback_1_4_valid ? _GEN_9763 : _GEN_9635; // @[Rob.scala 1222:23]
  wire  _GEN_9892 = io_writeback_1_4_valid ? _GEN_9764 : _GEN_9636; // @[Rob.scala 1222:23]
  wire  _GEN_9893 = io_writeback_1_4_valid ? _GEN_9765 : _GEN_9637; // @[Rob.scala 1222:23]
  wire  _GEN_9894 = io_writeback_1_4_valid ? _GEN_9766 : _GEN_9638; // @[Rob.scala 1222:23]
  wire  _GEN_9895 = io_writeback_1_4_valid ? _GEN_9767 : _GEN_9639; // @[Rob.scala 1222:23]
  wire  _GEN_9896 = io_writeback_1_4_valid ? _GEN_9768 : _GEN_9640; // @[Rob.scala 1222:23]
  wire  _GEN_9897 = io_writeback_1_4_valid ? _GEN_9769 : _GEN_9641; // @[Rob.scala 1222:23]
  wire  _GEN_9898 = io_writeback_1_4_valid ? _GEN_9770 : _GEN_9642; // @[Rob.scala 1222:23]
  wire  _GEN_9899 = io_writeback_1_4_valid ? _GEN_9771 : _GEN_9643; // @[Rob.scala 1222:23]
  wire  _GEN_9900 = io_writeback_1_4_valid ? _GEN_9772 : _GEN_9644; // @[Rob.scala 1222:23]
  wire  _GEN_9901 = io_writeback_1_4_valid ? _GEN_9773 : _GEN_9645; // @[Rob.scala 1222:23]
  wire  _GEN_9902 = io_writeback_1_4_valid ? _GEN_9774 : _GEN_9646; // @[Rob.scala 1222:23]
  wire  _GEN_9903 = io_writeback_1_4_valid ? _GEN_9775 : _GEN_9647; // @[Rob.scala 1222:23]
  wire  _GEN_9904 = io_writeback_1_4_valid ? _GEN_9776 : _GEN_9648; // @[Rob.scala 1222:23]
  wire  _GEN_9905 = io_writeback_1_4_valid ? _GEN_9777 : _GEN_9649; // @[Rob.scala 1222:23]
  wire  _GEN_9906 = io_writeback_1_4_valid ? _GEN_9778 : _GEN_9650; // @[Rob.scala 1222:23]
  wire  _GEN_9907 = io_writeback_1_4_valid ? _GEN_9779 : _GEN_9651; // @[Rob.scala 1222:23]
  wire  _GEN_9908 = io_writeback_1_4_valid ? _GEN_9780 : _GEN_9652; // @[Rob.scala 1222:23]
  wire  _GEN_9909 = io_writeback_1_4_valid ? _GEN_9781 : _GEN_9653; // @[Rob.scala 1222:23]
  wire  _GEN_9910 = io_writeback_1_4_valid ? _GEN_9782 : _GEN_9654; // @[Rob.scala 1222:23]
  wire  _GEN_9911 = io_writeback_1_4_valid ? _GEN_9783 : _GEN_9655; // @[Rob.scala 1222:23]
  wire  _GEN_9912 = io_writeback_1_4_valid ? _GEN_9784 : _GEN_9656; // @[Rob.scala 1222:23]
  wire  _GEN_9913 = io_writeback_1_4_valid ? _GEN_9785 : _GEN_9657; // @[Rob.scala 1222:23]
  wire  _GEN_9914 = io_writeback_1_4_valid ? _GEN_9786 : _GEN_9658; // @[Rob.scala 1222:23]
  wire  _GEN_9915 = io_writeback_1_4_valid ? _GEN_9787 : _GEN_9659; // @[Rob.scala 1222:23]
  wire  _GEN_9916 = io_writeback_1_4_valid ? _GEN_9788 : _GEN_9660; // @[Rob.scala 1222:23]
  wire  _GEN_9917 = io_writeback_1_4_valid ? _GEN_9789 : _GEN_9661; // @[Rob.scala 1222:23]
  wire  _GEN_9918 = io_writeback_1_4_valid ? _GEN_9790 : _GEN_9662; // @[Rob.scala 1222:23]
  wire  _GEN_9919 = io_writeback_1_4_valid ? _GEN_9791 : _GEN_9663; // @[Rob.scala 1222:23]
  wire  _GEN_9920 = io_writeback_1_4_valid ? _GEN_9792 : _GEN_9664; // @[Rob.scala 1222:23]
  wire  _GEN_9921 = io_writeback_1_4_valid ? _GEN_9793 : _GEN_9665; // @[Rob.scala 1222:23]
  wire  _GEN_9922 = io_writeback_1_4_valid ? _GEN_9794 : _GEN_9666; // @[Rob.scala 1222:23]
  wire  _GEN_9923 = io_writeback_1_4_valid ? _GEN_9795 : _GEN_9667; // @[Rob.scala 1222:23]
  wire  _GEN_9924 = io_writeback_1_4_valid ? _GEN_9796 : _GEN_9668; // @[Rob.scala 1222:23]
  wire  _GEN_9925 = io_writeback_1_4_valid ? _GEN_9797 : _GEN_9669; // @[Rob.scala 1222:23]
  wire  _GEN_9926 = io_writeback_1_4_valid ? _GEN_9798 : _GEN_9670; // @[Rob.scala 1222:23]
  wire  _GEN_9927 = io_writeback_1_4_valid ? _GEN_9799 : _GEN_9671; // @[Rob.scala 1222:23]
  wire  _GEN_9928 = io_writeback_1_4_valid ? _GEN_9800 : _GEN_9672; // @[Rob.scala 1222:23]
  wire  _GEN_9929 = io_writeback_1_4_valid ? _GEN_9801 : _GEN_9673; // @[Rob.scala 1222:23]
  wire  _GEN_9930 = io_writeback_1_4_valid ? _GEN_9802 : _GEN_9674; // @[Rob.scala 1222:23]
  wire  _GEN_9995 = 5'h0 == io_writeback_1_5_bits_uop_robIdx_value ? 1'h0 : _GEN_9867; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9996 = 5'h1 == io_writeback_1_5_bits_uop_robIdx_value ? 1'h0 : _GEN_9868; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9997 = 5'h2 == io_writeback_1_5_bits_uop_robIdx_value ? 1'h0 : _GEN_9869; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9998 = 5'h3 == io_writeback_1_5_bits_uop_robIdx_value ? 1'h0 : _GEN_9870; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_9999 = 5'h4 == io_writeback_1_5_bits_uop_robIdx_value ? 1'h0 : _GEN_9871; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10000 = 5'h5 == io_writeback_1_5_bits_uop_robIdx_value ? 1'h0 : _GEN_9872; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10001 = 5'h6 == io_writeback_1_5_bits_uop_robIdx_value ? 1'h0 : _GEN_9873; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10002 = 5'h7 == io_writeback_1_5_bits_uop_robIdx_value ? 1'h0 : _GEN_9874; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10003 = 5'h8 == io_writeback_1_5_bits_uop_robIdx_value ? 1'h0 : _GEN_9875; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10004 = 5'h9 == io_writeback_1_5_bits_uop_robIdx_value ? 1'h0 : _GEN_9876; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10005 = 5'ha == io_writeback_1_5_bits_uop_robIdx_value ? 1'h0 : _GEN_9877; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10006 = 5'hb == io_writeback_1_5_bits_uop_robIdx_value ? 1'h0 : _GEN_9878; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10007 = 5'hc == io_writeback_1_5_bits_uop_robIdx_value ? 1'h0 : _GEN_9879; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10008 = 5'hd == io_writeback_1_5_bits_uop_robIdx_value ? 1'h0 : _GEN_9880; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10009 = 5'he == io_writeback_1_5_bits_uop_robIdx_value ? 1'h0 : _GEN_9881; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10010 = 5'hf == io_writeback_1_5_bits_uop_robIdx_value ? 1'h0 : _GEN_9882; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10011 = 5'h10 == io_writeback_1_5_bits_uop_robIdx_value ? 1'h0 : _GEN_9883; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10012 = 5'h11 == io_writeback_1_5_bits_uop_robIdx_value ? 1'h0 : _GEN_9884; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10013 = 5'h12 == io_writeback_1_5_bits_uop_robIdx_value ? 1'h0 : _GEN_9885; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10014 = 5'h13 == io_writeback_1_5_bits_uop_robIdx_value ? 1'h0 : _GEN_9886; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10015 = 5'h14 == io_writeback_1_5_bits_uop_robIdx_value ? 1'h0 : _GEN_9887; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10016 = 5'h15 == io_writeback_1_5_bits_uop_robIdx_value ? 1'h0 : _GEN_9888; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10017 = 5'h16 == io_writeback_1_5_bits_uop_robIdx_value ? 1'h0 : _GEN_9889; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10018 = 5'h17 == io_writeback_1_5_bits_uop_robIdx_value ? 1'h0 : _GEN_9890; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10019 = 5'h18 == io_writeback_1_5_bits_uop_robIdx_value ? 1'h0 : _GEN_9891; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10020 = 5'h19 == io_writeback_1_5_bits_uop_robIdx_value ? 1'h0 : _GEN_9892; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10021 = 5'h1a == io_writeback_1_5_bits_uop_robIdx_value ? 1'h0 : _GEN_9893; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10022 = 5'h1b == io_writeback_1_5_bits_uop_robIdx_value ? 1'h0 : _GEN_9894; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10023 = 5'h1c == io_writeback_1_5_bits_uop_robIdx_value ? 1'h0 : _GEN_9895; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10024 = 5'h1d == io_writeback_1_5_bits_uop_robIdx_value ? 1'h0 : _GEN_9896; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10025 = 5'h1e == io_writeback_1_5_bits_uop_robIdx_value ? 1'h0 : _GEN_9897; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10026 = 5'h1f == io_writeback_1_5_bits_uop_robIdx_value ? 1'h0 : _GEN_9898; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10027 = 5'h0 == io_writeback_1_5_bits_uop_robIdx_value ? 1'h0 : _GEN_9899; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10028 = 5'h1 == io_writeback_1_5_bits_uop_robIdx_value ? 1'h0 : _GEN_9900; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10029 = 5'h2 == io_writeback_1_5_bits_uop_robIdx_value ? 1'h0 : _GEN_9901; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10030 = 5'h3 == io_writeback_1_5_bits_uop_robIdx_value ? 1'h0 : _GEN_9902; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10031 = 5'h4 == io_writeback_1_5_bits_uop_robIdx_value ? 1'h0 : _GEN_9903; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10032 = 5'h5 == io_writeback_1_5_bits_uop_robIdx_value ? 1'h0 : _GEN_9904; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10033 = 5'h6 == io_writeback_1_5_bits_uop_robIdx_value ? 1'h0 : _GEN_9905; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10034 = 5'h7 == io_writeback_1_5_bits_uop_robIdx_value ? 1'h0 : _GEN_9906; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10035 = 5'h8 == io_writeback_1_5_bits_uop_robIdx_value ? 1'h0 : _GEN_9907; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10036 = 5'h9 == io_writeback_1_5_bits_uop_robIdx_value ? 1'h0 : _GEN_9908; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10037 = 5'ha == io_writeback_1_5_bits_uop_robIdx_value ? 1'h0 : _GEN_9909; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10038 = 5'hb == io_writeback_1_5_bits_uop_robIdx_value ? 1'h0 : _GEN_9910; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10039 = 5'hc == io_writeback_1_5_bits_uop_robIdx_value ? 1'h0 : _GEN_9911; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10040 = 5'hd == io_writeback_1_5_bits_uop_robIdx_value ? 1'h0 : _GEN_9912; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10041 = 5'he == io_writeback_1_5_bits_uop_robIdx_value ? 1'h0 : _GEN_9913; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10042 = 5'hf == io_writeback_1_5_bits_uop_robIdx_value ? 1'h0 : _GEN_9914; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10043 = 5'h10 == io_writeback_1_5_bits_uop_robIdx_value ? 1'h0 : _GEN_9915; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10044 = 5'h11 == io_writeback_1_5_bits_uop_robIdx_value ? 1'h0 : _GEN_9916; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10045 = 5'h12 == io_writeback_1_5_bits_uop_robIdx_value ? 1'h0 : _GEN_9917; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10046 = 5'h13 == io_writeback_1_5_bits_uop_robIdx_value ? 1'h0 : _GEN_9918; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10047 = 5'h14 == io_writeback_1_5_bits_uop_robIdx_value ? 1'h0 : _GEN_9919; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10048 = 5'h15 == io_writeback_1_5_bits_uop_robIdx_value ? 1'h0 : _GEN_9920; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10049 = 5'h16 == io_writeback_1_5_bits_uop_robIdx_value ? 1'h0 : _GEN_9921; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10050 = 5'h17 == io_writeback_1_5_bits_uop_robIdx_value ? 1'h0 : _GEN_9922; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10051 = 5'h18 == io_writeback_1_5_bits_uop_robIdx_value ? 1'h0 : _GEN_9923; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10052 = 5'h19 == io_writeback_1_5_bits_uop_robIdx_value ? 1'h0 : _GEN_9924; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10053 = 5'h1a == io_writeback_1_5_bits_uop_robIdx_value ? 1'h0 : _GEN_9925; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10054 = 5'h1b == io_writeback_1_5_bits_uop_robIdx_value ? 1'h0 : _GEN_9926; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10055 = 5'h1c == io_writeback_1_5_bits_uop_robIdx_value ? 1'h0 : _GEN_9927; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10056 = 5'h1d == io_writeback_1_5_bits_uop_robIdx_value ? 1'h0 : _GEN_9928; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10057 = 5'h1e == io_writeback_1_5_bits_uop_robIdx_value ? 1'h0 : _GEN_9929; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10058 = 5'h1f == io_writeback_1_5_bits_uop_robIdx_value ? 1'h0 : _GEN_9930; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10123 = io_writeback_1_5_valid ? _GEN_9995 : _GEN_9867; // @[Rob.scala 1222:23]
  wire  _GEN_10124 = io_writeback_1_5_valid ? _GEN_9996 : _GEN_9868; // @[Rob.scala 1222:23]
  wire  _GEN_10125 = io_writeback_1_5_valid ? _GEN_9997 : _GEN_9869; // @[Rob.scala 1222:23]
  wire  _GEN_10126 = io_writeback_1_5_valid ? _GEN_9998 : _GEN_9870; // @[Rob.scala 1222:23]
  wire  _GEN_10127 = io_writeback_1_5_valid ? _GEN_9999 : _GEN_9871; // @[Rob.scala 1222:23]
  wire  _GEN_10128 = io_writeback_1_5_valid ? _GEN_10000 : _GEN_9872; // @[Rob.scala 1222:23]
  wire  _GEN_10129 = io_writeback_1_5_valid ? _GEN_10001 : _GEN_9873; // @[Rob.scala 1222:23]
  wire  _GEN_10130 = io_writeback_1_5_valid ? _GEN_10002 : _GEN_9874; // @[Rob.scala 1222:23]
  wire  _GEN_10131 = io_writeback_1_5_valid ? _GEN_10003 : _GEN_9875; // @[Rob.scala 1222:23]
  wire  _GEN_10132 = io_writeback_1_5_valid ? _GEN_10004 : _GEN_9876; // @[Rob.scala 1222:23]
  wire  _GEN_10133 = io_writeback_1_5_valid ? _GEN_10005 : _GEN_9877; // @[Rob.scala 1222:23]
  wire  _GEN_10134 = io_writeback_1_5_valid ? _GEN_10006 : _GEN_9878; // @[Rob.scala 1222:23]
  wire  _GEN_10135 = io_writeback_1_5_valid ? _GEN_10007 : _GEN_9879; // @[Rob.scala 1222:23]
  wire  _GEN_10136 = io_writeback_1_5_valid ? _GEN_10008 : _GEN_9880; // @[Rob.scala 1222:23]
  wire  _GEN_10137 = io_writeback_1_5_valid ? _GEN_10009 : _GEN_9881; // @[Rob.scala 1222:23]
  wire  _GEN_10138 = io_writeback_1_5_valid ? _GEN_10010 : _GEN_9882; // @[Rob.scala 1222:23]
  wire  _GEN_10139 = io_writeback_1_5_valid ? _GEN_10011 : _GEN_9883; // @[Rob.scala 1222:23]
  wire  _GEN_10140 = io_writeback_1_5_valid ? _GEN_10012 : _GEN_9884; // @[Rob.scala 1222:23]
  wire  _GEN_10141 = io_writeback_1_5_valid ? _GEN_10013 : _GEN_9885; // @[Rob.scala 1222:23]
  wire  _GEN_10142 = io_writeback_1_5_valid ? _GEN_10014 : _GEN_9886; // @[Rob.scala 1222:23]
  wire  _GEN_10143 = io_writeback_1_5_valid ? _GEN_10015 : _GEN_9887; // @[Rob.scala 1222:23]
  wire  _GEN_10144 = io_writeback_1_5_valid ? _GEN_10016 : _GEN_9888; // @[Rob.scala 1222:23]
  wire  _GEN_10145 = io_writeback_1_5_valid ? _GEN_10017 : _GEN_9889; // @[Rob.scala 1222:23]
  wire  _GEN_10146 = io_writeback_1_5_valid ? _GEN_10018 : _GEN_9890; // @[Rob.scala 1222:23]
  wire  _GEN_10147 = io_writeback_1_5_valid ? _GEN_10019 : _GEN_9891; // @[Rob.scala 1222:23]
  wire  _GEN_10148 = io_writeback_1_5_valid ? _GEN_10020 : _GEN_9892; // @[Rob.scala 1222:23]
  wire  _GEN_10149 = io_writeback_1_5_valid ? _GEN_10021 : _GEN_9893; // @[Rob.scala 1222:23]
  wire  _GEN_10150 = io_writeback_1_5_valid ? _GEN_10022 : _GEN_9894; // @[Rob.scala 1222:23]
  wire  _GEN_10151 = io_writeback_1_5_valid ? _GEN_10023 : _GEN_9895; // @[Rob.scala 1222:23]
  wire  _GEN_10152 = io_writeback_1_5_valid ? _GEN_10024 : _GEN_9896; // @[Rob.scala 1222:23]
  wire  _GEN_10153 = io_writeback_1_5_valid ? _GEN_10025 : _GEN_9897; // @[Rob.scala 1222:23]
  wire  _GEN_10154 = io_writeback_1_5_valid ? _GEN_10026 : _GEN_9898; // @[Rob.scala 1222:23]
  wire  _GEN_10155 = io_writeback_1_5_valid ? _GEN_10027 : _GEN_9899; // @[Rob.scala 1222:23]
  wire  _GEN_10156 = io_writeback_1_5_valid ? _GEN_10028 : _GEN_9900; // @[Rob.scala 1222:23]
  wire  _GEN_10157 = io_writeback_1_5_valid ? _GEN_10029 : _GEN_9901; // @[Rob.scala 1222:23]
  wire  _GEN_10158 = io_writeback_1_5_valid ? _GEN_10030 : _GEN_9902; // @[Rob.scala 1222:23]
  wire  _GEN_10159 = io_writeback_1_5_valid ? _GEN_10031 : _GEN_9903; // @[Rob.scala 1222:23]
  wire  _GEN_10160 = io_writeback_1_5_valid ? _GEN_10032 : _GEN_9904; // @[Rob.scala 1222:23]
  wire  _GEN_10161 = io_writeback_1_5_valid ? _GEN_10033 : _GEN_9905; // @[Rob.scala 1222:23]
  wire  _GEN_10162 = io_writeback_1_5_valid ? _GEN_10034 : _GEN_9906; // @[Rob.scala 1222:23]
  wire  _GEN_10163 = io_writeback_1_5_valid ? _GEN_10035 : _GEN_9907; // @[Rob.scala 1222:23]
  wire  _GEN_10164 = io_writeback_1_5_valid ? _GEN_10036 : _GEN_9908; // @[Rob.scala 1222:23]
  wire  _GEN_10165 = io_writeback_1_5_valid ? _GEN_10037 : _GEN_9909; // @[Rob.scala 1222:23]
  wire  _GEN_10166 = io_writeback_1_5_valid ? _GEN_10038 : _GEN_9910; // @[Rob.scala 1222:23]
  wire  _GEN_10167 = io_writeback_1_5_valid ? _GEN_10039 : _GEN_9911; // @[Rob.scala 1222:23]
  wire  _GEN_10168 = io_writeback_1_5_valid ? _GEN_10040 : _GEN_9912; // @[Rob.scala 1222:23]
  wire  _GEN_10169 = io_writeback_1_5_valid ? _GEN_10041 : _GEN_9913; // @[Rob.scala 1222:23]
  wire  _GEN_10170 = io_writeback_1_5_valid ? _GEN_10042 : _GEN_9914; // @[Rob.scala 1222:23]
  wire  _GEN_10171 = io_writeback_1_5_valid ? _GEN_10043 : _GEN_9915; // @[Rob.scala 1222:23]
  wire  _GEN_10172 = io_writeback_1_5_valid ? _GEN_10044 : _GEN_9916; // @[Rob.scala 1222:23]
  wire  _GEN_10173 = io_writeback_1_5_valid ? _GEN_10045 : _GEN_9917; // @[Rob.scala 1222:23]
  wire  _GEN_10174 = io_writeback_1_5_valid ? _GEN_10046 : _GEN_9918; // @[Rob.scala 1222:23]
  wire  _GEN_10175 = io_writeback_1_5_valid ? _GEN_10047 : _GEN_9919; // @[Rob.scala 1222:23]
  wire  _GEN_10176 = io_writeback_1_5_valid ? _GEN_10048 : _GEN_9920; // @[Rob.scala 1222:23]
  wire  _GEN_10177 = io_writeback_1_5_valid ? _GEN_10049 : _GEN_9921; // @[Rob.scala 1222:23]
  wire  _GEN_10178 = io_writeback_1_5_valid ? _GEN_10050 : _GEN_9922; // @[Rob.scala 1222:23]
  wire  _GEN_10179 = io_writeback_1_5_valid ? _GEN_10051 : _GEN_9923; // @[Rob.scala 1222:23]
  wire  _GEN_10180 = io_writeback_1_5_valid ? _GEN_10052 : _GEN_9924; // @[Rob.scala 1222:23]
  wire  _GEN_10181 = io_writeback_1_5_valid ? _GEN_10053 : _GEN_9925; // @[Rob.scala 1222:23]
  wire  _GEN_10182 = io_writeback_1_5_valid ? _GEN_10054 : _GEN_9926; // @[Rob.scala 1222:23]
  wire  _GEN_10183 = io_writeback_1_5_valid ? _GEN_10055 : _GEN_9927; // @[Rob.scala 1222:23]
  wire  _GEN_10184 = io_writeback_1_5_valid ? _GEN_10056 : _GEN_9928; // @[Rob.scala 1222:23]
  wire  _GEN_10185 = io_writeback_1_5_valid ? _GEN_10057 : _GEN_9929; // @[Rob.scala 1222:23]
  wire  _GEN_10186 = io_writeback_1_5_valid ? _GEN_10058 : _GEN_9930; // @[Rob.scala 1222:23]
  wire  _GEN_10251 = 5'h0 == io_writeback_1_6_bits_uop_robIdx_value ? 1'h0 : _GEN_10123; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10252 = 5'h1 == io_writeback_1_6_bits_uop_robIdx_value ? 1'h0 : _GEN_10124; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10253 = 5'h2 == io_writeback_1_6_bits_uop_robIdx_value ? 1'h0 : _GEN_10125; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10254 = 5'h3 == io_writeback_1_6_bits_uop_robIdx_value ? 1'h0 : _GEN_10126; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10255 = 5'h4 == io_writeback_1_6_bits_uop_robIdx_value ? 1'h0 : _GEN_10127; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10256 = 5'h5 == io_writeback_1_6_bits_uop_robIdx_value ? 1'h0 : _GEN_10128; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10257 = 5'h6 == io_writeback_1_6_bits_uop_robIdx_value ? 1'h0 : _GEN_10129; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10258 = 5'h7 == io_writeback_1_6_bits_uop_robIdx_value ? 1'h0 : _GEN_10130; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10259 = 5'h8 == io_writeback_1_6_bits_uop_robIdx_value ? 1'h0 : _GEN_10131; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10260 = 5'h9 == io_writeback_1_6_bits_uop_robIdx_value ? 1'h0 : _GEN_10132; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10261 = 5'ha == io_writeback_1_6_bits_uop_robIdx_value ? 1'h0 : _GEN_10133; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10262 = 5'hb == io_writeback_1_6_bits_uop_robIdx_value ? 1'h0 : _GEN_10134; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10263 = 5'hc == io_writeback_1_6_bits_uop_robIdx_value ? 1'h0 : _GEN_10135; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10264 = 5'hd == io_writeback_1_6_bits_uop_robIdx_value ? 1'h0 : _GEN_10136; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10265 = 5'he == io_writeback_1_6_bits_uop_robIdx_value ? 1'h0 : _GEN_10137; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10266 = 5'hf == io_writeback_1_6_bits_uop_robIdx_value ? 1'h0 : _GEN_10138; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10267 = 5'h10 == io_writeback_1_6_bits_uop_robIdx_value ? 1'h0 : _GEN_10139; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10268 = 5'h11 == io_writeback_1_6_bits_uop_robIdx_value ? 1'h0 : _GEN_10140; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10269 = 5'h12 == io_writeback_1_6_bits_uop_robIdx_value ? 1'h0 : _GEN_10141; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10270 = 5'h13 == io_writeback_1_6_bits_uop_robIdx_value ? 1'h0 : _GEN_10142; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10271 = 5'h14 == io_writeback_1_6_bits_uop_robIdx_value ? 1'h0 : _GEN_10143; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10272 = 5'h15 == io_writeback_1_6_bits_uop_robIdx_value ? 1'h0 : _GEN_10144; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10273 = 5'h16 == io_writeback_1_6_bits_uop_robIdx_value ? 1'h0 : _GEN_10145; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10274 = 5'h17 == io_writeback_1_6_bits_uop_robIdx_value ? 1'h0 : _GEN_10146; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10275 = 5'h18 == io_writeback_1_6_bits_uop_robIdx_value ? 1'h0 : _GEN_10147; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10276 = 5'h19 == io_writeback_1_6_bits_uop_robIdx_value ? 1'h0 : _GEN_10148; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10277 = 5'h1a == io_writeback_1_6_bits_uop_robIdx_value ? 1'h0 : _GEN_10149; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10278 = 5'h1b == io_writeback_1_6_bits_uop_robIdx_value ? 1'h0 : _GEN_10150; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10279 = 5'h1c == io_writeback_1_6_bits_uop_robIdx_value ? 1'h0 : _GEN_10151; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10280 = 5'h1d == io_writeback_1_6_bits_uop_robIdx_value ? 1'h0 : _GEN_10152; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10281 = 5'h1e == io_writeback_1_6_bits_uop_robIdx_value ? 1'h0 : _GEN_10153; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10282 = 5'h1f == io_writeback_1_6_bits_uop_robIdx_value ? 1'h0 : _GEN_10154; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10283 = 5'h0 == io_writeback_1_6_bits_uop_robIdx_value ? io_writeback_1_6_bits_debug_isPerfCnt : _GEN_10155
    ; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10284 = 5'h1 == io_writeback_1_6_bits_uop_robIdx_value ? io_writeback_1_6_bits_debug_isPerfCnt : _GEN_10156
    ; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10285 = 5'h2 == io_writeback_1_6_bits_uop_robIdx_value ? io_writeback_1_6_bits_debug_isPerfCnt : _GEN_10157
    ; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10286 = 5'h3 == io_writeback_1_6_bits_uop_robIdx_value ? io_writeback_1_6_bits_debug_isPerfCnt : _GEN_10158
    ; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10287 = 5'h4 == io_writeback_1_6_bits_uop_robIdx_value ? io_writeback_1_6_bits_debug_isPerfCnt : _GEN_10159
    ; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10288 = 5'h5 == io_writeback_1_6_bits_uop_robIdx_value ? io_writeback_1_6_bits_debug_isPerfCnt : _GEN_10160
    ; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10289 = 5'h6 == io_writeback_1_6_bits_uop_robIdx_value ? io_writeback_1_6_bits_debug_isPerfCnt : _GEN_10161
    ; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10290 = 5'h7 == io_writeback_1_6_bits_uop_robIdx_value ? io_writeback_1_6_bits_debug_isPerfCnt : _GEN_10162
    ; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10291 = 5'h8 == io_writeback_1_6_bits_uop_robIdx_value ? io_writeback_1_6_bits_debug_isPerfCnt : _GEN_10163
    ; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10292 = 5'h9 == io_writeback_1_6_bits_uop_robIdx_value ? io_writeback_1_6_bits_debug_isPerfCnt : _GEN_10164
    ; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10293 = 5'ha == io_writeback_1_6_bits_uop_robIdx_value ? io_writeback_1_6_bits_debug_isPerfCnt : _GEN_10165
    ; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10294 = 5'hb == io_writeback_1_6_bits_uop_robIdx_value ? io_writeback_1_6_bits_debug_isPerfCnt : _GEN_10166
    ; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10295 = 5'hc == io_writeback_1_6_bits_uop_robIdx_value ? io_writeback_1_6_bits_debug_isPerfCnt : _GEN_10167
    ; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10296 = 5'hd == io_writeback_1_6_bits_uop_robIdx_value ? io_writeback_1_6_bits_debug_isPerfCnt : _GEN_10168
    ; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10297 = 5'he == io_writeback_1_6_bits_uop_robIdx_value ? io_writeback_1_6_bits_debug_isPerfCnt : _GEN_10169
    ; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10298 = 5'hf == io_writeback_1_6_bits_uop_robIdx_value ? io_writeback_1_6_bits_debug_isPerfCnt : _GEN_10170
    ; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10299 = 5'h10 == io_writeback_1_6_bits_uop_robIdx_value ? io_writeback_1_6_bits_debug_isPerfCnt :
    _GEN_10171; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10300 = 5'h11 == io_writeback_1_6_bits_uop_robIdx_value ? io_writeback_1_6_bits_debug_isPerfCnt :
    _GEN_10172; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10301 = 5'h12 == io_writeback_1_6_bits_uop_robIdx_value ? io_writeback_1_6_bits_debug_isPerfCnt :
    _GEN_10173; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10302 = 5'h13 == io_writeback_1_6_bits_uop_robIdx_value ? io_writeback_1_6_bits_debug_isPerfCnt :
    _GEN_10174; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10303 = 5'h14 == io_writeback_1_6_bits_uop_robIdx_value ? io_writeback_1_6_bits_debug_isPerfCnt :
    _GEN_10175; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10304 = 5'h15 == io_writeback_1_6_bits_uop_robIdx_value ? io_writeback_1_6_bits_debug_isPerfCnt :
    _GEN_10176; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10305 = 5'h16 == io_writeback_1_6_bits_uop_robIdx_value ? io_writeback_1_6_bits_debug_isPerfCnt :
    _GEN_10177; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10306 = 5'h17 == io_writeback_1_6_bits_uop_robIdx_value ? io_writeback_1_6_bits_debug_isPerfCnt :
    _GEN_10178; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10307 = 5'h18 == io_writeback_1_6_bits_uop_robIdx_value ? io_writeback_1_6_bits_debug_isPerfCnt :
    _GEN_10179; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10308 = 5'h19 == io_writeback_1_6_bits_uop_robIdx_value ? io_writeback_1_6_bits_debug_isPerfCnt :
    _GEN_10180; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10309 = 5'h1a == io_writeback_1_6_bits_uop_robIdx_value ? io_writeback_1_6_bits_debug_isPerfCnt :
    _GEN_10181; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10310 = 5'h1b == io_writeback_1_6_bits_uop_robIdx_value ? io_writeback_1_6_bits_debug_isPerfCnt :
    _GEN_10182; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10311 = 5'h1c == io_writeback_1_6_bits_uop_robIdx_value ? io_writeback_1_6_bits_debug_isPerfCnt :
    _GEN_10183; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10312 = 5'h1d == io_writeback_1_6_bits_uop_robIdx_value ? io_writeback_1_6_bits_debug_isPerfCnt :
    _GEN_10184; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10313 = 5'h1e == io_writeback_1_6_bits_uop_robIdx_value ? io_writeback_1_6_bits_debug_isPerfCnt :
    _GEN_10185; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10314 = 5'h1f == io_writeback_1_6_bits_uop_robIdx_value ? io_writeback_1_6_bits_debug_isPerfCnt :
    _GEN_10186; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10379 = io_writeback_1_6_valid ? _GEN_10251 : _GEN_10123; // @[Rob.scala 1222:23]
  wire  _GEN_10380 = io_writeback_1_6_valid ? _GEN_10252 : _GEN_10124; // @[Rob.scala 1222:23]
  wire  _GEN_10381 = io_writeback_1_6_valid ? _GEN_10253 : _GEN_10125; // @[Rob.scala 1222:23]
  wire  _GEN_10382 = io_writeback_1_6_valid ? _GEN_10254 : _GEN_10126; // @[Rob.scala 1222:23]
  wire  _GEN_10383 = io_writeback_1_6_valid ? _GEN_10255 : _GEN_10127; // @[Rob.scala 1222:23]
  wire  _GEN_10384 = io_writeback_1_6_valid ? _GEN_10256 : _GEN_10128; // @[Rob.scala 1222:23]
  wire  _GEN_10385 = io_writeback_1_6_valid ? _GEN_10257 : _GEN_10129; // @[Rob.scala 1222:23]
  wire  _GEN_10386 = io_writeback_1_6_valid ? _GEN_10258 : _GEN_10130; // @[Rob.scala 1222:23]
  wire  _GEN_10387 = io_writeback_1_6_valid ? _GEN_10259 : _GEN_10131; // @[Rob.scala 1222:23]
  wire  _GEN_10388 = io_writeback_1_6_valid ? _GEN_10260 : _GEN_10132; // @[Rob.scala 1222:23]
  wire  _GEN_10389 = io_writeback_1_6_valid ? _GEN_10261 : _GEN_10133; // @[Rob.scala 1222:23]
  wire  _GEN_10390 = io_writeback_1_6_valid ? _GEN_10262 : _GEN_10134; // @[Rob.scala 1222:23]
  wire  _GEN_10391 = io_writeback_1_6_valid ? _GEN_10263 : _GEN_10135; // @[Rob.scala 1222:23]
  wire  _GEN_10392 = io_writeback_1_6_valid ? _GEN_10264 : _GEN_10136; // @[Rob.scala 1222:23]
  wire  _GEN_10393 = io_writeback_1_6_valid ? _GEN_10265 : _GEN_10137; // @[Rob.scala 1222:23]
  wire  _GEN_10394 = io_writeback_1_6_valid ? _GEN_10266 : _GEN_10138; // @[Rob.scala 1222:23]
  wire  _GEN_10395 = io_writeback_1_6_valid ? _GEN_10267 : _GEN_10139; // @[Rob.scala 1222:23]
  wire  _GEN_10396 = io_writeback_1_6_valid ? _GEN_10268 : _GEN_10140; // @[Rob.scala 1222:23]
  wire  _GEN_10397 = io_writeback_1_6_valid ? _GEN_10269 : _GEN_10141; // @[Rob.scala 1222:23]
  wire  _GEN_10398 = io_writeback_1_6_valid ? _GEN_10270 : _GEN_10142; // @[Rob.scala 1222:23]
  wire  _GEN_10399 = io_writeback_1_6_valid ? _GEN_10271 : _GEN_10143; // @[Rob.scala 1222:23]
  wire  _GEN_10400 = io_writeback_1_6_valid ? _GEN_10272 : _GEN_10144; // @[Rob.scala 1222:23]
  wire  _GEN_10401 = io_writeback_1_6_valid ? _GEN_10273 : _GEN_10145; // @[Rob.scala 1222:23]
  wire  _GEN_10402 = io_writeback_1_6_valid ? _GEN_10274 : _GEN_10146; // @[Rob.scala 1222:23]
  wire  _GEN_10403 = io_writeback_1_6_valid ? _GEN_10275 : _GEN_10147; // @[Rob.scala 1222:23]
  wire  _GEN_10404 = io_writeback_1_6_valid ? _GEN_10276 : _GEN_10148; // @[Rob.scala 1222:23]
  wire  _GEN_10405 = io_writeback_1_6_valid ? _GEN_10277 : _GEN_10149; // @[Rob.scala 1222:23]
  wire  _GEN_10406 = io_writeback_1_6_valid ? _GEN_10278 : _GEN_10150; // @[Rob.scala 1222:23]
  wire  _GEN_10407 = io_writeback_1_6_valid ? _GEN_10279 : _GEN_10151; // @[Rob.scala 1222:23]
  wire  _GEN_10408 = io_writeback_1_6_valid ? _GEN_10280 : _GEN_10152; // @[Rob.scala 1222:23]
  wire  _GEN_10409 = io_writeback_1_6_valid ? _GEN_10281 : _GEN_10153; // @[Rob.scala 1222:23]
  wire  _GEN_10410 = io_writeback_1_6_valid ? _GEN_10282 : _GEN_10154; // @[Rob.scala 1222:23]
  wire  _GEN_10411 = io_writeback_1_6_valid ? _GEN_10283 : _GEN_10155; // @[Rob.scala 1222:23]
  wire  _GEN_10412 = io_writeback_1_6_valid ? _GEN_10284 : _GEN_10156; // @[Rob.scala 1222:23]
  wire  _GEN_10413 = io_writeback_1_6_valid ? _GEN_10285 : _GEN_10157; // @[Rob.scala 1222:23]
  wire  _GEN_10414 = io_writeback_1_6_valid ? _GEN_10286 : _GEN_10158; // @[Rob.scala 1222:23]
  wire  _GEN_10415 = io_writeback_1_6_valid ? _GEN_10287 : _GEN_10159; // @[Rob.scala 1222:23]
  wire  _GEN_10416 = io_writeback_1_6_valid ? _GEN_10288 : _GEN_10160; // @[Rob.scala 1222:23]
  wire  _GEN_10417 = io_writeback_1_6_valid ? _GEN_10289 : _GEN_10161; // @[Rob.scala 1222:23]
  wire  _GEN_10418 = io_writeback_1_6_valid ? _GEN_10290 : _GEN_10162; // @[Rob.scala 1222:23]
  wire  _GEN_10419 = io_writeback_1_6_valid ? _GEN_10291 : _GEN_10163; // @[Rob.scala 1222:23]
  wire  _GEN_10420 = io_writeback_1_6_valid ? _GEN_10292 : _GEN_10164; // @[Rob.scala 1222:23]
  wire  _GEN_10421 = io_writeback_1_6_valid ? _GEN_10293 : _GEN_10165; // @[Rob.scala 1222:23]
  wire  _GEN_10422 = io_writeback_1_6_valid ? _GEN_10294 : _GEN_10166; // @[Rob.scala 1222:23]
  wire  _GEN_10423 = io_writeback_1_6_valid ? _GEN_10295 : _GEN_10167; // @[Rob.scala 1222:23]
  wire  _GEN_10424 = io_writeback_1_6_valid ? _GEN_10296 : _GEN_10168; // @[Rob.scala 1222:23]
  wire  _GEN_10425 = io_writeback_1_6_valid ? _GEN_10297 : _GEN_10169; // @[Rob.scala 1222:23]
  wire  _GEN_10426 = io_writeback_1_6_valid ? _GEN_10298 : _GEN_10170; // @[Rob.scala 1222:23]
  wire  _GEN_10427 = io_writeback_1_6_valid ? _GEN_10299 : _GEN_10171; // @[Rob.scala 1222:23]
  wire  _GEN_10428 = io_writeback_1_6_valid ? _GEN_10300 : _GEN_10172; // @[Rob.scala 1222:23]
  wire  _GEN_10429 = io_writeback_1_6_valid ? _GEN_10301 : _GEN_10173; // @[Rob.scala 1222:23]
  wire  _GEN_10430 = io_writeback_1_6_valid ? _GEN_10302 : _GEN_10174; // @[Rob.scala 1222:23]
  wire  _GEN_10431 = io_writeback_1_6_valid ? _GEN_10303 : _GEN_10175; // @[Rob.scala 1222:23]
  wire  _GEN_10432 = io_writeback_1_6_valid ? _GEN_10304 : _GEN_10176; // @[Rob.scala 1222:23]
  wire  _GEN_10433 = io_writeback_1_6_valid ? _GEN_10305 : _GEN_10177; // @[Rob.scala 1222:23]
  wire  _GEN_10434 = io_writeback_1_6_valid ? _GEN_10306 : _GEN_10178; // @[Rob.scala 1222:23]
  wire  _GEN_10435 = io_writeback_1_6_valid ? _GEN_10307 : _GEN_10179; // @[Rob.scala 1222:23]
  wire  _GEN_10436 = io_writeback_1_6_valid ? _GEN_10308 : _GEN_10180; // @[Rob.scala 1222:23]
  wire  _GEN_10437 = io_writeback_1_6_valid ? _GEN_10309 : _GEN_10181; // @[Rob.scala 1222:23]
  wire  _GEN_10438 = io_writeback_1_6_valid ? _GEN_10310 : _GEN_10182; // @[Rob.scala 1222:23]
  wire  _GEN_10439 = io_writeback_1_6_valid ? _GEN_10311 : _GEN_10183; // @[Rob.scala 1222:23]
  wire  _GEN_10440 = io_writeback_1_6_valid ? _GEN_10312 : _GEN_10184; // @[Rob.scala 1222:23]
  wire  _GEN_10441 = io_writeback_1_6_valid ? _GEN_10313 : _GEN_10185; // @[Rob.scala 1222:23]
  wire  _GEN_10442 = io_writeback_1_6_valid ? _GEN_10314 : _GEN_10186; // @[Rob.scala 1222:23]
  wire  _GEN_10507 = 5'h0 == io_writeback_1_7_bits_uop_robIdx_value ? io_writeback_1_7_bits_debug_isMMIO : _GEN_10379; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10508 = 5'h1 == io_writeback_1_7_bits_uop_robIdx_value ? io_writeback_1_7_bits_debug_isMMIO : _GEN_10380; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10509 = 5'h2 == io_writeback_1_7_bits_uop_robIdx_value ? io_writeback_1_7_bits_debug_isMMIO : _GEN_10381; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10510 = 5'h3 == io_writeback_1_7_bits_uop_robIdx_value ? io_writeback_1_7_bits_debug_isMMIO : _GEN_10382; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10511 = 5'h4 == io_writeback_1_7_bits_uop_robIdx_value ? io_writeback_1_7_bits_debug_isMMIO : _GEN_10383; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10512 = 5'h5 == io_writeback_1_7_bits_uop_robIdx_value ? io_writeback_1_7_bits_debug_isMMIO : _GEN_10384; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10513 = 5'h6 == io_writeback_1_7_bits_uop_robIdx_value ? io_writeback_1_7_bits_debug_isMMIO : _GEN_10385; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10514 = 5'h7 == io_writeback_1_7_bits_uop_robIdx_value ? io_writeback_1_7_bits_debug_isMMIO : _GEN_10386; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10515 = 5'h8 == io_writeback_1_7_bits_uop_robIdx_value ? io_writeback_1_7_bits_debug_isMMIO : _GEN_10387; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10516 = 5'h9 == io_writeback_1_7_bits_uop_robIdx_value ? io_writeback_1_7_bits_debug_isMMIO : _GEN_10388; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10517 = 5'ha == io_writeback_1_7_bits_uop_robIdx_value ? io_writeback_1_7_bits_debug_isMMIO : _GEN_10389; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10518 = 5'hb == io_writeback_1_7_bits_uop_robIdx_value ? io_writeback_1_7_bits_debug_isMMIO : _GEN_10390; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10519 = 5'hc == io_writeback_1_7_bits_uop_robIdx_value ? io_writeback_1_7_bits_debug_isMMIO : _GEN_10391; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10520 = 5'hd == io_writeback_1_7_bits_uop_robIdx_value ? io_writeback_1_7_bits_debug_isMMIO : _GEN_10392; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10521 = 5'he == io_writeback_1_7_bits_uop_robIdx_value ? io_writeback_1_7_bits_debug_isMMIO : _GEN_10393; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10522 = 5'hf == io_writeback_1_7_bits_uop_robIdx_value ? io_writeback_1_7_bits_debug_isMMIO : _GEN_10394; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10523 = 5'h10 == io_writeback_1_7_bits_uop_robIdx_value ? io_writeback_1_7_bits_debug_isMMIO : _GEN_10395; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10524 = 5'h11 == io_writeback_1_7_bits_uop_robIdx_value ? io_writeback_1_7_bits_debug_isMMIO : _GEN_10396; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10525 = 5'h12 == io_writeback_1_7_bits_uop_robIdx_value ? io_writeback_1_7_bits_debug_isMMIO : _GEN_10397; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10526 = 5'h13 == io_writeback_1_7_bits_uop_robIdx_value ? io_writeback_1_7_bits_debug_isMMIO : _GEN_10398; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10527 = 5'h14 == io_writeback_1_7_bits_uop_robIdx_value ? io_writeback_1_7_bits_debug_isMMIO : _GEN_10399; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10528 = 5'h15 == io_writeback_1_7_bits_uop_robIdx_value ? io_writeback_1_7_bits_debug_isMMIO : _GEN_10400; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10529 = 5'h16 == io_writeback_1_7_bits_uop_robIdx_value ? io_writeback_1_7_bits_debug_isMMIO : _GEN_10401; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10530 = 5'h17 == io_writeback_1_7_bits_uop_robIdx_value ? io_writeback_1_7_bits_debug_isMMIO : _GEN_10402; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10531 = 5'h18 == io_writeback_1_7_bits_uop_robIdx_value ? io_writeback_1_7_bits_debug_isMMIO : _GEN_10403; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10532 = 5'h19 == io_writeback_1_7_bits_uop_robIdx_value ? io_writeback_1_7_bits_debug_isMMIO : _GEN_10404; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10533 = 5'h1a == io_writeback_1_7_bits_uop_robIdx_value ? io_writeback_1_7_bits_debug_isMMIO : _GEN_10405; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10534 = 5'h1b == io_writeback_1_7_bits_uop_robIdx_value ? io_writeback_1_7_bits_debug_isMMIO : _GEN_10406; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10535 = 5'h1c == io_writeback_1_7_bits_uop_robIdx_value ? io_writeback_1_7_bits_debug_isMMIO : _GEN_10407; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10536 = 5'h1d == io_writeback_1_7_bits_uop_robIdx_value ? io_writeback_1_7_bits_debug_isMMIO : _GEN_10408; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10537 = 5'h1e == io_writeback_1_7_bits_uop_robIdx_value ? io_writeback_1_7_bits_debug_isMMIO : _GEN_10409; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10538 = 5'h1f == io_writeback_1_7_bits_uop_robIdx_value ? io_writeback_1_7_bits_debug_isMMIO : _GEN_10410; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10539 = 5'h0 == io_writeback_1_7_bits_uop_robIdx_value ? io_writeback_1_7_bits_debug_isPerfCnt : _GEN_10411
    ; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10540 = 5'h1 == io_writeback_1_7_bits_uop_robIdx_value ? io_writeback_1_7_bits_debug_isPerfCnt : _GEN_10412
    ; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10541 = 5'h2 == io_writeback_1_7_bits_uop_robIdx_value ? io_writeback_1_7_bits_debug_isPerfCnt : _GEN_10413
    ; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10542 = 5'h3 == io_writeback_1_7_bits_uop_robIdx_value ? io_writeback_1_7_bits_debug_isPerfCnt : _GEN_10414
    ; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10543 = 5'h4 == io_writeback_1_7_bits_uop_robIdx_value ? io_writeback_1_7_bits_debug_isPerfCnt : _GEN_10415
    ; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10544 = 5'h5 == io_writeback_1_7_bits_uop_robIdx_value ? io_writeback_1_7_bits_debug_isPerfCnt : _GEN_10416
    ; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10545 = 5'h6 == io_writeback_1_7_bits_uop_robIdx_value ? io_writeback_1_7_bits_debug_isPerfCnt : _GEN_10417
    ; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10546 = 5'h7 == io_writeback_1_7_bits_uop_robIdx_value ? io_writeback_1_7_bits_debug_isPerfCnt : _GEN_10418
    ; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10547 = 5'h8 == io_writeback_1_7_bits_uop_robIdx_value ? io_writeback_1_7_bits_debug_isPerfCnt : _GEN_10419
    ; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10548 = 5'h9 == io_writeback_1_7_bits_uop_robIdx_value ? io_writeback_1_7_bits_debug_isPerfCnt : _GEN_10420
    ; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10549 = 5'ha == io_writeback_1_7_bits_uop_robIdx_value ? io_writeback_1_7_bits_debug_isPerfCnt : _GEN_10421
    ; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10550 = 5'hb == io_writeback_1_7_bits_uop_robIdx_value ? io_writeback_1_7_bits_debug_isPerfCnt : _GEN_10422
    ; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10551 = 5'hc == io_writeback_1_7_bits_uop_robIdx_value ? io_writeback_1_7_bits_debug_isPerfCnt : _GEN_10423
    ; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10552 = 5'hd == io_writeback_1_7_bits_uop_robIdx_value ? io_writeback_1_7_bits_debug_isPerfCnt : _GEN_10424
    ; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10553 = 5'he == io_writeback_1_7_bits_uop_robIdx_value ? io_writeback_1_7_bits_debug_isPerfCnt : _GEN_10425
    ; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10554 = 5'hf == io_writeback_1_7_bits_uop_robIdx_value ? io_writeback_1_7_bits_debug_isPerfCnt : _GEN_10426
    ; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10555 = 5'h10 == io_writeback_1_7_bits_uop_robIdx_value ? io_writeback_1_7_bits_debug_isPerfCnt :
    _GEN_10427; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10556 = 5'h11 == io_writeback_1_7_bits_uop_robIdx_value ? io_writeback_1_7_bits_debug_isPerfCnt :
    _GEN_10428; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10557 = 5'h12 == io_writeback_1_7_bits_uop_robIdx_value ? io_writeback_1_7_bits_debug_isPerfCnt :
    _GEN_10429; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10558 = 5'h13 == io_writeback_1_7_bits_uop_robIdx_value ? io_writeback_1_7_bits_debug_isPerfCnt :
    _GEN_10430; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10559 = 5'h14 == io_writeback_1_7_bits_uop_robIdx_value ? io_writeback_1_7_bits_debug_isPerfCnt :
    _GEN_10431; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10560 = 5'h15 == io_writeback_1_7_bits_uop_robIdx_value ? io_writeback_1_7_bits_debug_isPerfCnt :
    _GEN_10432; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10561 = 5'h16 == io_writeback_1_7_bits_uop_robIdx_value ? io_writeback_1_7_bits_debug_isPerfCnt :
    _GEN_10433; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10562 = 5'h17 == io_writeback_1_7_bits_uop_robIdx_value ? io_writeback_1_7_bits_debug_isPerfCnt :
    _GEN_10434; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10563 = 5'h18 == io_writeback_1_7_bits_uop_robIdx_value ? io_writeback_1_7_bits_debug_isPerfCnt :
    _GEN_10435; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10564 = 5'h19 == io_writeback_1_7_bits_uop_robIdx_value ? io_writeback_1_7_bits_debug_isPerfCnt :
    _GEN_10436; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10565 = 5'h1a == io_writeback_1_7_bits_uop_robIdx_value ? io_writeback_1_7_bits_debug_isPerfCnt :
    _GEN_10437; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10566 = 5'h1b == io_writeback_1_7_bits_uop_robIdx_value ? io_writeback_1_7_bits_debug_isPerfCnt :
    _GEN_10438; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10567 = 5'h1c == io_writeback_1_7_bits_uop_robIdx_value ? io_writeback_1_7_bits_debug_isPerfCnt :
    _GEN_10439; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10568 = 5'h1d == io_writeback_1_7_bits_uop_robIdx_value ? io_writeback_1_7_bits_debug_isPerfCnt :
    _GEN_10440; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10569 = 5'h1e == io_writeback_1_7_bits_uop_robIdx_value ? io_writeback_1_7_bits_debug_isPerfCnt :
    _GEN_10441; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10570 = 5'h1f == io_writeback_1_7_bits_uop_robIdx_value ? io_writeback_1_7_bits_debug_isPerfCnt :
    _GEN_10442; // @[Rob.scala 1224:{28,28}]
  wire  _GEN_10635 = io_writeback_1_7_valid ? _GEN_10507 : _GEN_10379; // @[Rob.scala 1222:23]
  wire  _GEN_10636 = io_writeback_1_7_valid ? _GEN_10508 : _GEN_10380; // @[Rob.scala 1222:23]
  wire  _GEN_10637 = io_writeback_1_7_valid ? _GEN_10509 : _GEN_10381; // @[Rob.scala 1222:23]
  wire  _GEN_10638 = io_writeback_1_7_valid ? _GEN_10510 : _GEN_10382; // @[Rob.scala 1222:23]
  wire  _GEN_10639 = io_writeback_1_7_valid ? _GEN_10511 : _GEN_10383; // @[Rob.scala 1222:23]
  wire  _GEN_10640 = io_writeback_1_7_valid ? _GEN_10512 : _GEN_10384; // @[Rob.scala 1222:23]
  wire  _GEN_10641 = io_writeback_1_7_valid ? _GEN_10513 : _GEN_10385; // @[Rob.scala 1222:23]
  wire  _GEN_10642 = io_writeback_1_7_valid ? _GEN_10514 : _GEN_10386; // @[Rob.scala 1222:23]
  wire  _GEN_10643 = io_writeback_1_7_valid ? _GEN_10515 : _GEN_10387; // @[Rob.scala 1222:23]
  wire  _GEN_10644 = io_writeback_1_7_valid ? _GEN_10516 : _GEN_10388; // @[Rob.scala 1222:23]
  wire  _GEN_10645 = io_writeback_1_7_valid ? _GEN_10517 : _GEN_10389; // @[Rob.scala 1222:23]
  wire  _GEN_10646 = io_writeback_1_7_valid ? _GEN_10518 : _GEN_10390; // @[Rob.scala 1222:23]
  wire  _GEN_10647 = io_writeback_1_7_valid ? _GEN_10519 : _GEN_10391; // @[Rob.scala 1222:23]
  wire  _GEN_10648 = io_writeback_1_7_valid ? _GEN_10520 : _GEN_10392; // @[Rob.scala 1222:23]
  wire  _GEN_10649 = io_writeback_1_7_valid ? _GEN_10521 : _GEN_10393; // @[Rob.scala 1222:23]
  wire  _GEN_10650 = io_writeback_1_7_valid ? _GEN_10522 : _GEN_10394; // @[Rob.scala 1222:23]
  wire  _GEN_10651 = io_writeback_1_7_valid ? _GEN_10523 : _GEN_10395; // @[Rob.scala 1222:23]
  wire  _GEN_10652 = io_writeback_1_7_valid ? _GEN_10524 : _GEN_10396; // @[Rob.scala 1222:23]
  wire  _GEN_10653 = io_writeback_1_7_valid ? _GEN_10525 : _GEN_10397; // @[Rob.scala 1222:23]
  wire  _GEN_10654 = io_writeback_1_7_valid ? _GEN_10526 : _GEN_10398; // @[Rob.scala 1222:23]
  wire  _GEN_10655 = io_writeback_1_7_valid ? _GEN_10527 : _GEN_10399; // @[Rob.scala 1222:23]
  wire  _GEN_10656 = io_writeback_1_7_valid ? _GEN_10528 : _GEN_10400; // @[Rob.scala 1222:23]
  wire  _GEN_10657 = io_writeback_1_7_valid ? _GEN_10529 : _GEN_10401; // @[Rob.scala 1222:23]
  wire  _GEN_10658 = io_writeback_1_7_valid ? _GEN_10530 : _GEN_10402; // @[Rob.scala 1222:23]
  wire  _GEN_10659 = io_writeback_1_7_valid ? _GEN_10531 : _GEN_10403; // @[Rob.scala 1222:23]
  wire  _GEN_10660 = io_writeback_1_7_valid ? _GEN_10532 : _GEN_10404; // @[Rob.scala 1222:23]
  wire  _GEN_10661 = io_writeback_1_7_valid ? _GEN_10533 : _GEN_10405; // @[Rob.scala 1222:23]
  wire  _GEN_10662 = io_writeback_1_7_valid ? _GEN_10534 : _GEN_10406; // @[Rob.scala 1222:23]
  wire  _GEN_10663 = io_writeback_1_7_valid ? _GEN_10535 : _GEN_10407; // @[Rob.scala 1222:23]
  wire  _GEN_10664 = io_writeback_1_7_valid ? _GEN_10536 : _GEN_10408; // @[Rob.scala 1222:23]
  wire  _GEN_10665 = io_writeback_1_7_valid ? _GEN_10537 : _GEN_10409; // @[Rob.scala 1222:23]
  wire  _GEN_10666 = io_writeback_1_7_valid ? _GEN_10538 : _GEN_10410; // @[Rob.scala 1222:23]
  wire  _GEN_10667 = io_writeback_1_7_valid ? _GEN_10539 : _GEN_10411; // @[Rob.scala 1222:23]
  wire  _GEN_10668 = io_writeback_1_7_valid ? _GEN_10540 : _GEN_10412; // @[Rob.scala 1222:23]
  wire  _GEN_10669 = io_writeback_1_7_valid ? _GEN_10541 : _GEN_10413; // @[Rob.scala 1222:23]
  wire  _GEN_10670 = io_writeback_1_7_valid ? _GEN_10542 : _GEN_10414; // @[Rob.scala 1222:23]
  wire  _GEN_10671 = io_writeback_1_7_valid ? _GEN_10543 : _GEN_10415; // @[Rob.scala 1222:23]
  wire  _GEN_10672 = io_writeback_1_7_valid ? _GEN_10544 : _GEN_10416; // @[Rob.scala 1222:23]
  wire  _GEN_10673 = io_writeback_1_7_valid ? _GEN_10545 : _GEN_10417; // @[Rob.scala 1222:23]
  wire  _GEN_10674 = io_writeback_1_7_valid ? _GEN_10546 : _GEN_10418; // @[Rob.scala 1222:23]
  wire  _GEN_10675 = io_writeback_1_7_valid ? _GEN_10547 : _GEN_10419; // @[Rob.scala 1222:23]
  wire  _GEN_10676 = io_writeback_1_7_valid ? _GEN_10548 : _GEN_10420; // @[Rob.scala 1222:23]
  wire  _GEN_10677 = io_writeback_1_7_valid ? _GEN_10549 : _GEN_10421; // @[Rob.scala 1222:23]
  wire  _GEN_10678 = io_writeback_1_7_valid ? _GEN_10550 : _GEN_10422; // @[Rob.scala 1222:23]
  wire  _GEN_10679 = io_writeback_1_7_valid ? _GEN_10551 : _GEN_10423; // @[Rob.scala 1222:23]
  wire  _GEN_10680 = io_writeback_1_7_valid ? _GEN_10552 : _GEN_10424; // @[Rob.scala 1222:23]
  wire  _GEN_10681 = io_writeback_1_7_valid ? _GEN_10553 : _GEN_10425; // @[Rob.scala 1222:23]
  wire  _GEN_10682 = io_writeback_1_7_valid ? _GEN_10554 : _GEN_10426; // @[Rob.scala 1222:23]
  wire  _GEN_10683 = io_writeback_1_7_valid ? _GEN_10555 : _GEN_10427; // @[Rob.scala 1222:23]
  wire  _GEN_10684 = io_writeback_1_7_valid ? _GEN_10556 : _GEN_10428; // @[Rob.scala 1222:23]
  wire  _GEN_10685 = io_writeback_1_7_valid ? _GEN_10557 : _GEN_10429; // @[Rob.scala 1222:23]
  wire  _GEN_10686 = io_writeback_1_7_valid ? _GEN_10558 : _GEN_10430; // @[Rob.scala 1222:23]
  wire  _GEN_10687 = io_writeback_1_7_valid ? _GEN_10559 : _GEN_10431; // @[Rob.scala 1222:23]
  wire  _GEN_10688 = io_writeback_1_7_valid ? _GEN_10560 : _GEN_10432; // @[Rob.scala 1222:23]
  wire  _GEN_10689 = io_writeback_1_7_valid ? _GEN_10561 : _GEN_10433; // @[Rob.scala 1222:23]
  wire  _GEN_10690 = io_writeback_1_7_valid ? _GEN_10562 : _GEN_10434; // @[Rob.scala 1222:23]
  wire  _GEN_10691 = io_writeback_1_7_valid ? _GEN_10563 : _GEN_10435; // @[Rob.scala 1222:23]
  wire  _GEN_10692 = io_writeback_1_7_valid ? _GEN_10564 : _GEN_10436; // @[Rob.scala 1222:23]
  wire  _GEN_10693 = io_writeback_1_7_valid ? _GEN_10565 : _GEN_10437; // @[Rob.scala 1222:23]
  wire  _GEN_10694 = io_writeback_1_7_valid ? _GEN_10566 : _GEN_10438; // @[Rob.scala 1222:23]
  wire  _GEN_10695 = io_writeback_1_7_valid ? _GEN_10567 : _GEN_10439; // @[Rob.scala 1222:23]
  wire  _GEN_10696 = io_writeback_1_7_valid ? _GEN_10568 : _GEN_10440; // @[Rob.scala 1222:23]
  wire  _GEN_10697 = io_writeback_1_7_valid ? _GEN_10569 : _GEN_10441; // @[Rob.scala 1222:23]
  wire  _GEN_10698 = io_writeback_1_7_valid ? _GEN_10570 : _GEN_10442; // @[Rob.scala 1222:23]
  reg  difftest_io_valid_REG; // @[Rob.scala 1239:53]
  reg  difftest_io_valid_REG_1; // @[Rob.scala 1239:45]
  reg  difftest_io_valid_REG_2; // @[Rob.scala 1239:37]
  reg  difftest_io_special_REG; // @[Rob.scala 1240:53]
  reg  difftest_io_special_REG_1; // @[Rob.scala 1240:45]
  reg  difftest_io_special_REG_2; // @[Rob.scala 1240:37]
  wire  _GEN_11020 = 5'h1 == deqPtrVec_0_value ? dt_exuDebug_1_isMMIO : dt_exuDebug_0_isMMIO; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11021 = 5'h2 == deqPtrVec_0_value ? dt_exuDebug_2_isMMIO : _GEN_11020; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11022 = 5'h3 == deqPtrVec_0_value ? dt_exuDebug_3_isMMIO : _GEN_11021; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11023 = 5'h4 == deqPtrVec_0_value ? dt_exuDebug_4_isMMIO : _GEN_11022; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11024 = 5'h5 == deqPtrVec_0_value ? dt_exuDebug_5_isMMIO : _GEN_11023; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11025 = 5'h6 == deqPtrVec_0_value ? dt_exuDebug_6_isMMIO : _GEN_11024; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11026 = 5'h7 == deqPtrVec_0_value ? dt_exuDebug_7_isMMIO : _GEN_11025; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11027 = 5'h8 == deqPtrVec_0_value ? dt_exuDebug_8_isMMIO : _GEN_11026; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11028 = 5'h9 == deqPtrVec_0_value ? dt_exuDebug_9_isMMIO : _GEN_11027; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11029 = 5'ha == deqPtrVec_0_value ? dt_exuDebug_10_isMMIO : _GEN_11028; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11030 = 5'hb == deqPtrVec_0_value ? dt_exuDebug_11_isMMIO : _GEN_11029; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11031 = 5'hc == deqPtrVec_0_value ? dt_exuDebug_12_isMMIO : _GEN_11030; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11032 = 5'hd == deqPtrVec_0_value ? dt_exuDebug_13_isMMIO : _GEN_11031; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11033 = 5'he == deqPtrVec_0_value ? dt_exuDebug_14_isMMIO : _GEN_11032; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11034 = 5'hf == deqPtrVec_0_value ? dt_exuDebug_15_isMMIO : _GEN_11033; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11035 = 5'h10 == deqPtrVec_0_value ? dt_exuDebug_16_isMMIO : _GEN_11034; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11036 = 5'h11 == deqPtrVec_0_value ? dt_exuDebug_17_isMMIO : _GEN_11035; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11037 = 5'h12 == deqPtrVec_0_value ? dt_exuDebug_18_isMMIO : _GEN_11036; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11038 = 5'h13 == deqPtrVec_0_value ? dt_exuDebug_19_isMMIO : _GEN_11037; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11039 = 5'h14 == deqPtrVec_0_value ? dt_exuDebug_20_isMMIO : _GEN_11038; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11040 = 5'h15 == deqPtrVec_0_value ? dt_exuDebug_21_isMMIO : _GEN_11039; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11041 = 5'h16 == deqPtrVec_0_value ? dt_exuDebug_22_isMMIO : _GEN_11040; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11042 = 5'h17 == deqPtrVec_0_value ? dt_exuDebug_23_isMMIO : _GEN_11041; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11043 = 5'h18 == deqPtrVec_0_value ? dt_exuDebug_24_isMMIO : _GEN_11042; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11044 = 5'h19 == deqPtrVec_0_value ? dt_exuDebug_25_isMMIO : _GEN_11043; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11045 = 5'h1a == deqPtrVec_0_value ? dt_exuDebug_26_isMMIO : _GEN_11044; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11046 = 5'h1b == deqPtrVec_0_value ? dt_exuDebug_27_isMMIO : _GEN_11045; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11047 = 5'h1c == deqPtrVec_0_value ? dt_exuDebug_28_isMMIO : _GEN_11046; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11048 = 5'h1d == deqPtrVec_0_value ? dt_exuDebug_29_isMMIO : _GEN_11047; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11049 = 5'h1e == deqPtrVec_0_value ? dt_exuDebug_30_isMMIO : _GEN_11048; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11050 = 5'h1f == deqPtrVec_0_value ? dt_exuDebug_31_isMMIO : _GEN_11049; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11052 = 5'h1 == deqPtrVec_0_value ? dt_exuDebug_1_isPerfCnt : dt_exuDebug_0_isPerfCnt; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11053 = 5'h2 == deqPtrVec_0_value ? dt_exuDebug_2_isPerfCnt : _GEN_11052; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11054 = 5'h3 == deqPtrVec_0_value ? dt_exuDebug_3_isPerfCnt : _GEN_11053; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11055 = 5'h4 == deqPtrVec_0_value ? dt_exuDebug_4_isPerfCnt : _GEN_11054; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11056 = 5'h5 == deqPtrVec_0_value ? dt_exuDebug_5_isPerfCnt : _GEN_11055; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11057 = 5'h6 == deqPtrVec_0_value ? dt_exuDebug_6_isPerfCnt : _GEN_11056; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11058 = 5'h7 == deqPtrVec_0_value ? dt_exuDebug_7_isPerfCnt : _GEN_11057; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11059 = 5'h8 == deqPtrVec_0_value ? dt_exuDebug_8_isPerfCnt : _GEN_11058; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11060 = 5'h9 == deqPtrVec_0_value ? dt_exuDebug_9_isPerfCnt : _GEN_11059; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11061 = 5'ha == deqPtrVec_0_value ? dt_exuDebug_10_isPerfCnt : _GEN_11060; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11062 = 5'hb == deqPtrVec_0_value ? dt_exuDebug_11_isPerfCnt : _GEN_11061; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11063 = 5'hc == deqPtrVec_0_value ? dt_exuDebug_12_isPerfCnt : _GEN_11062; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11064 = 5'hd == deqPtrVec_0_value ? dt_exuDebug_13_isPerfCnt : _GEN_11063; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11065 = 5'he == deqPtrVec_0_value ? dt_exuDebug_14_isPerfCnt : _GEN_11064; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11066 = 5'hf == deqPtrVec_0_value ? dt_exuDebug_15_isPerfCnt : _GEN_11065; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11067 = 5'h10 == deqPtrVec_0_value ? dt_exuDebug_16_isPerfCnt : _GEN_11066; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11068 = 5'h11 == deqPtrVec_0_value ? dt_exuDebug_17_isPerfCnt : _GEN_11067; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11069 = 5'h12 == deqPtrVec_0_value ? dt_exuDebug_18_isPerfCnt : _GEN_11068; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11070 = 5'h13 == deqPtrVec_0_value ? dt_exuDebug_19_isPerfCnt : _GEN_11069; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11071 = 5'h14 == deqPtrVec_0_value ? dt_exuDebug_20_isPerfCnt : _GEN_11070; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11072 = 5'h15 == deqPtrVec_0_value ? dt_exuDebug_21_isPerfCnt : _GEN_11071; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11073 = 5'h16 == deqPtrVec_0_value ? dt_exuDebug_22_isPerfCnt : _GEN_11072; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11074 = 5'h17 == deqPtrVec_0_value ? dt_exuDebug_23_isPerfCnt : _GEN_11073; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11075 = 5'h18 == deqPtrVec_0_value ? dt_exuDebug_24_isPerfCnt : _GEN_11074; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11076 = 5'h19 == deqPtrVec_0_value ? dt_exuDebug_25_isPerfCnt : _GEN_11075; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11077 = 5'h1a == deqPtrVec_0_value ? dt_exuDebug_26_isPerfCnt : _GEN_11076; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11078 = 5'h1b == deqPtrVec_0_value ? dt_exuDebug_27_isPerfCnt : _GEN_11077; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11079 = 5'h1c == deqPtrVec_0_value ? dt_exuDebug_28_isPerfCnt : _GEN_11078; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11080 = 5'h1d == deqPtrVec_0_value ? dt_exuDebug_29_isPerfCnt : _GEN_11079; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11081 = 5'h1e == deqPtrVec_0_value ? dt_exuDebug_30_isPerfCnt : _GEN_11080; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11082 = 5'h1f == deqPtrVec_0_value ? dt_exuDebug_31_isPerfCnt : _GEN_11081; // @[Rob.scala 1241:{97,97}]
  reg  difftest_io_skip_REG; // @[Rob.scala 1241:53]
  reg  difftest_io_skip_REG_1; // @[Rob.scala 1241:45]
  reg  difftest_io_skip_REG_2; // @[Rob.scala 1241:37]
  reg  difftest_io_isRVC_REG; // @[Rob.scala 1242:53]
  reg  difftest_io_isRVC_REG_1; // @[Rob.scala 1242:45]
  reg  difftest_io_isRVC_REG_2; // @[Rob.scala 1242:37]
  reg  difftest_io_rfwen_REG; // @[Rob.scala 1243:53]
  reg  difftest_io_rfwen_REG_1; // @[Rob.scala 1243:45]
  reg  difftest_io_rfwen_REG_2; // @[Rob.scala 1243:37]
  reg  difftest_io_fpwen_REG; // @[Rob.scala 1244:53]
  reg  difftest_io_fpwen_REG_1; // @[Rob.scala 1244:45]
  reg  difftest_io_fpwen_REG_2; // @[Rob.scala 1244:37]
  reg [5:0] difftest_io_wpdest_REG; // @[Rob.scala 1245:53]
  reg [5:0] difftest_io_wpdest_REG_1; // @[Rob.scala 1245:45]
  reg [5:0] difftest_io_wpdest_REG_2; // @[Rob.scala 1245:37]
  reg [4:0] difftest_io_wdest_REG; // @[Rob.scala 1246:53]
  reg [4:0] difftest_io_wdest_REG_1; // @[Rob.scala 1246:45]
  reg [4:0] difftest_io_wdest_REG_2; // @[Rob.scala 1246:37]
  reg  difftest_io_valid_REG_3; // @[Rob.scala 1239:53]
  reg  difftest_io_valid_REG_4; // @[Rob.scala 1239:45]
  reg  difftest_io_valid_REG_5; // @[Rob.scala 1239:37]
  reg  difftest_io_special_REG_3; // @[Rob.scala 1240:53]
  reg  difftest_io_special_REG_4; // @[Rob.scala 1240:45]
  reg  difftest_io_special_REG_5; // @[Rob.scala 1240:37]
  wire  _GEN_11084 = 5'h1 == deqPtrVec_1_value ? dt_exuDebug_1_isMMIO : dt_exuDebug_0_isMMIO; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11085 = 5'h2 == deqPtrVec_1_value ? dt_exuDebug_2_isMMIO : _GEN_11084; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11086 = 5'h3 == deqPtrVec_1_value ? dt_exuDebug_3_isMMIO : _GEN_11085; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11087 = 5'h4 == deqPtrVec_1_value ? dt_exuDebug_4_isMMIO : _GEN_11086; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11088 = 5'h5 == deqPtrVec_1_value ? dt_exuDebug_5_isMMIO : _GEN_11087; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11089 = 5'h6 == deqPtrVec_1_value ? dt_exuDebug_6_isMMIO : _GEN_11088; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11090 = 5'h7 == deqPtrVec_1_value ? dt_exuDebug_7_isMMIO : _GEN_11089; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11091 = 5'h8 == deqPtrVec_1_value ? dt_exuDebug_8_isMMIO : _GEN_11090; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11092 = 5'h9 == deqPtrVec_1_value ? dt_exuDebug_9_isMMIO : _GEN_11091; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11093 = 5'ha == deqPtrVec_1_value ? dt_exuDebug_10_isMMIO : _GEN_11092; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11094 = 5'hb == deqPtrVec_1_value ? dt_exuDebug_11_isMMIO : _GEN_11093; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11095 = 5'hc == deqPtrVec_1_value ? dt_exuDebug_12_isMMIO : _GEN_11094; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11096 = 5'hd == deqPtrVec_1_value ? dt_exuDebug_13_isMMIO : _GEN_11095; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11097 = 5'he == deqPtrVec_1_value ? dt_exuDebug_14_isMMIO : _GEN_11096; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11098 = 5'hf == deqPtrVec_1_value ? dt_exuDebug_15_isMMIO : _GEN_11097; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11099 = 5'h10 == deqPtrVec_1_value ? dt_exuDebug_16_isMMIO : _GEN_11098; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11100 = 5'h11 == deqPtrVec_1_value ? dt_exuDebug_17_isMMIO : _GEN_11099; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11101 = 5'h12 == deqPtrVec_1_value ? dt_exuDebug_18_isMMIO : _GEN_11100; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11102 = 5'h13 == deqPtrVec_1_value ? dt_exuDebug_19_isMMIO : _GEN_11101; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11103 = 5'h14 == deqPtrVec_1_value ? dt_exuDebug_20_isMMIO : _GEN_11102; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11104 = 5'h15 == deqPtrVec_1_value ? dt_exuDebug_21_isMMIO : _GEN_11103; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11105 = 5'h16 == deqPtrVec_1_value ? dt_exuDebug_22_isMMIO : _GEN_11104; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11106 = 5'h17 == deqPtrVec_1_value ? dt_exuDebug_23_isMMIO : _GEN_11105; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11107 = 5'h18 == deqPtrVec_1_value ? dt_exuDebug_24_isMMIO : _GEN_11106; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11108 = 5'h19 == deqPtrVec_1_value ? dt_exuDebug_25_isMMIO : _GEN_11107; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11109 = 5'h1a == deqPtrVec_1_value ? dt_exuDebug_26_isMMIO : _GEN_11108; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11110 = 5'h1b == deqPtrVec_1_value ? dt_exuDebug_27_isMMIO : _GEN_11109; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11111 = 5'h1c == deqPtrVec_1_value ? dt_exuDebug_28_isMMIO : _GEN_11110; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11112 = 5'h1d == deqPtrVec_1_value ? dt_exuDebug_29_isMMIO : _GEN_11111; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11113 = 5'h1e == deqPtrVec_1_value ? dt_exuDebug_30_isMMIO : _GEN_11112; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11114 = 5'h1f == deqPtrVec_1_value ? dt_exuDebug_31_isMMIO : _GEN_11113; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11116 = 5'h1 == deqPtrVec_1_value ? dt_exuDebug_1_isPerfCnt : dt_exuDebug_0_isPerfCnt; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11117 = 5'h2 == deqPtrVec_1_value ? dt_exuDebug_2_isPerfCnt : _GEN_11116; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11118 = 5'h3 == deqPtrVec_1_value ? dt_exuDebug_3_isPerfCnt : _GEN_11117; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11119 = 5'h4 == deqPtrVec_1_value ? dt_exuDebug_4_isPerfCnt : _GEN_11118; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11120 = 5'h5 == deqPtrVec_1_value ? dt_exuDebug_5_isPerfCnt : _GEN_11119; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11121 = 5'h6 == deqPtrVec_1_value ? dt_exuDebug_6_isPerfCnt : _GEN_11120; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11122 = 5'h7 == deqPtrVec_1_value ? dt_exuDebug_7_isPerfCnt : _GEN_11121; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11123 = 5'h8 == deqPtrVec_1_value ? dt_exuDebug_8_isPerfCnt : _GEN_11122; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11124 = 5'h9 == deqPtrVec_1_value ? dt_exuDebug_9_isPerfCnt : _GEN_11123; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11125 = 5'ha == deqPtrVec_1_value ? dt_exuDebug_10_isPerfCnt : _GEN_11124; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11126 = 5'hb == deqPtrVec_1_value ? dt_exuDebug_11_isPerfCnt : _GEN_11125; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11127 = 5'hc == deqPtrVec_1_value ? dt_exuDebug_12_isPerfCnt : _GEN_11126; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11128 = 5'hd == deqPtrVec_1_value ? dt_exuDebug_13_isPerfCnt : _GEN_11127; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11129 = 5'he == deqPtrVec_1_value ? dt_exuDebug_14_isPerfCnt : _GEN_11128; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11130 = 5'hf == deqPtrVec_1_value ? dt_exuDebug_15_isPerfCnt : _GEN_11129; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11131 = 5'h10 == deqPtrVec_1_value ? dt_exuDebug_16_isPerfCnt : _GEN_11130; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11132 = 5'h11 == deqPtrVec_1_value ? dt_exuDebug_17_isPerfCnt : _GEN_11131; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11133 = 5'h12 == deqPtrVec_1_value ? dt_exuDebug_18_isPerfCnt : _GEN_11132; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11134 = 5'h13 == deqPtrVec_1_value ? dt_exuDebug_19_isPerfCnt : _GEN_11133; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11135 = 5'h14 == deqPtrVec_1_value ? dt_exuDebug_20_isPerfCnt : _GEN_11134; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11136 = 5'h15 == deqPtrVec_1_value ? dt_exuDebug_21_isPerfCnt : _GEN_11135; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11137 = 5'h16 == deqPtrVec_1_value ? dt_exuDebug_22_isPerfCnt : _GEN_11136; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11138 = 5'h17 == deqPtrVec_1_value ? dt_exuDebug_23_isPerfCnt : _GEN_11137; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11139 = 5'h18 == deqPtrVec_1_value ? dt_exuDebug_24_isPerfCnt : _GEN_11138; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11140 = 5'h19 == deqPtrVec_1_value ? dt_exuDebug_25_isPerfCnt : _GEN_11139; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11141 = 5'h1a == deqPtrVec_1_value ? dt_exuDebug_26_isPerfCnt : _GEN_11140; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11142 = 5'h1b == deqPtrVec_1_value ? dt_exuDebug_27_isPerfCnt : _GEN_11141; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11143 = 5'h1c == deqPtrVec_1_value ? dt_exuDebug_28_isPerfCnt : _GEN_11142; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11144 = 5'h1d == deqPtrVec_1_value ? dt_exuDebug_29_isPerfCnt : _GEN_11143; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11145 = 5'h1e == deqPtrVec_1_value ? dt_exuDebug_30_isPerfCnt : _GEN_11144; // @[Rob.scala 1241:{97,97}]
  wire  _GEN_11146 = 5'h1f == deqPtrVec_1_value ? dt_exuDebug_31_isPerfCnt : _GEN_11145; // @[Rob.scala 1241:{97,97}]
  reg  difftest_io_skip_REG_3; // @[Rob.scala 1241:53]
  reg  difftest_io_skip_REG_4; // @[Rob.scala 1241:45]
  reg  difftest_io_skip_REG_5; // @[Rob.scala 1241:37]
  reg  difftest_io_isRVC_REG_3; // @[Rob.scala 1242:53]
  reg  difftest_io_isRVC_REG_4; // @[Rob.scala 1242:45]
  reg  difftest_io_isRVC_REG_5; // @[Rob.scala 1242:37]
  reg  difftest_io_rfwen_REG_3; // @[Rob.scala 1243:53]
  reg  difftest_io_rfwen_REG_4; // @[Rob.scala 1243:45]
  reg  difftest_io_rfwen_REG_5; // @[Rob.scala 1243:37]
  reg  difftest_io_fpwen_REG_3; // @[Rob.scala 1244:53]
  reg  difftest_io_fpwen_REG_4; // @[Rob.scala 1244:45]
  reg  difftest_io_fpwen_REG_5; // @[Rob.scala 1244:37]
  reg [5:0] difftest_io_wpdest_REG_3; // @[Rob.scala 1245:53]
  reg [5:0] difftest_io_wpdest_REG_4; // @[Rob.scala 1245:45]
  reg [5:0] difftest_io_wpdest_REG_5; // @[Rob.scala 1245:37]
  reg [4:0] difftest_io_wdest_REG_3; // @[Rob.scala 1246:53]
  reg [4:0] difftest_io_wdest_REG_4; // @[Rob.scala 1246:45]
  reg [4:0] difftest_io_wdest_REG_5; // @[Rob.scala 1246:37]
  wire  trapVec_0 = _T_117 & dt_isXSTrap_trapVec_MPORT_data; // @[Rob.scala 1296:102]
  wire  trapVec_1 = _T_125 & dt_isXSTrap_trapVec_MPORT_1_data; // @[Rob.scala 1296:102]
  reg [5:0] validEntriesBanks_0; // @[Rob.scala 1306:73]
  reg [5:0] validEntries; // @[Rob.scala 1307:29]
  reg  REG_19; // @[Rob.scala 1049:53]
  reg  REG_20_0; // @[Rob.scala 1320:61]
  reg  REG_20_1; // @[Rob.scala 1320:61]
  wire [1:0] _T_1083 = REG_20_0 + REG_20_1; // @[Bitwise.scala 48:55]
  reg  REG_21; // @[Rob.scala 1049:53]
  reg  REG_22; // @[Rob.scala 1049:53]
  reg  REG_23_0; // @[Rob.scala 1322:61]
  reg  REG_23_1; // @[Rob.scala 1322:61]
  wire [1:0] _T_1087 = REG_23_0 + REG_23_1; // @[Bitwise.scala 48:55]
  reg  REG_24; // @[Rob.scala 1049:53]
  reg  REG_25_0; // @[Rob.scala 1323:61]
  reg  REG_25_1; // @[Rob.scala 1323:61]
  wire [1:0] _T_1090 = REG_25_0 + REG_25_1; // @[Bitwise.scala 48:55]
  reg  REG_26; // @[Rob.scala 1049:53]
  reg  REG_27_0; // @[Rob.scala 1324:61]
  reg  REG_27_1; // @[Rob.scala 1324:61]
  wire [1:0] _T_1093 = REG_27_0 + REG_27_1; // @[Bitwise.scala 48:55]
  reg  REG_28; // @[Rob.scala 1049:53]
  reg  REG_29_0; // @[Rob.scala 1325:61]
  reg  REG_29_1; // @[Rob.scala 1325:61]
  wire [1:0] _T_1096 = REG_29_0 + REG_29_1; // @[Bitwise.scala 48:55]
  reg  REG_30; // @[Rob.scala 1049:53]
  reg  io_perf_0_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg  io_perf_0_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg  io_perf_1_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg  io_perf_1_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg  io_perf_2_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg  io_perf_2_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg  io_perf_3_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg  io_perf_3_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg [1:0] io_perf_4_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg [1:0] io_perf_4_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg [2:0] io_perf_5_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg [2:0] io_perf_5_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg [1:0] io_perf_6_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg [1:0] io_perf_6_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg [1:0] io_perf_7_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg [1:0] io_perf_7_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg [1:0] io_perf_8_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg [1:0] io_perf_8_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg [1:0] io_perf_9_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg [1:0] io_perf_9_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg [1:0] io_perf_10_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg [1:0] io_perf_10_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg [1:0] io_perf_11_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg [1:0] io_perf_11_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg [1:0] io_perf_12_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg [1:0] io_perf_12_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg  io_perf_13_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg  io_perf_13_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg  io_perf_14_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg  io_perf_14_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg  io_perf_15_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg  io_perf_15_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg  io_perf_16_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg  io_perf_16_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg  io_perf_17_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg  io_perf_17_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  SyncDataModuleTemplate__32entry dispatchData ( // @[Rob.scala 477:28]
    .clock(dispatchData_clock),
    .io_raddr_0(dispatchData_io_raddr_0),
    .io_raddr_1(dispatchData_io_raddr_1),
    .io_rdata_0_ldest(dispatchData_io_rdata_0_ldest),
    .io_rdata_0_rfWen(dispatchData_io_rdata_0_rfWen),
    .io_rdata_0_fpWen(dispatchData_io_rdata_0_fpWen),
    .io_rdata_0_wflags(dispatchData_io_rdata_0_wflags),
    .io_rdata_0_commitType(dispatchData_io_rdata_0_commitType),
    .io_rdata_0_pdest(dispatchData_io_rdata_0_pdest),
    .io_rdata_0_old_pdest(dispatchData_io_rdata_0_old_pdest),
    .io_rdata_0_ftqIdx_flag(dispatchData_io_rdata_0_ftqIdx_flag),
    .io_rdata_0_ftqIdx_value(dispatchData_io_rdata_0_ftqIdx_value),
    .io_rdata_0_ftqOffset(dispatchData_io_rdata_0_ftqOffset),
    .io_rdata_0_isMove(dispatchData_io_rdata_0_isMove),
    .io_rdata_1_ldest(dispatchData_io_rdata_1_ldest),
    .io_rdata_1_rfWen(dispatchData_io_rdata_1_rfWen),
    .io_rdata_1_fpWen(dispatchData_io_rdata_1_fpWen),
    .io_rdata_1_wflags(dispatchData_io_rdata_1_wflags),
    .io_rdata_1_commitType(dispatchData_io_rdata_1_commitType),
    .io_rdata_1_pdest(dispatchData_io_rdata_1_pdest),
    .io_rdata_1_old_pdest(dispatchData_io_rdata_1_old_pdest),
    .io_rdata_1_ftqIdx_flag(dispatchData_io_rdata_1_ftqIdx_flag),
    .io_rdata_1_ftqIdx_value(dispatchData_io_rdata_1_ftqIdx_value),
    .io_rdata_1_ftqOffset(dispatchData_io_rdata_1_ftqOffset),
    .io_rdata_1_isMove(dispatchData_io_rdata_1_isMove),
    .io_wen_0(dispatchData_io_wen_0),
    .io_wen_1(dispatchData_io_wen_1),
    .io_waddr_0(dispatchData_io_waddr_0),
    .io_waddr_1(dispatchData_io_waddr_1),
    .io_wdata_0_ldest(dispatchData_io_wdata_0_ldest),
    .io_wdata_0_rfWen(dispatchData_io_wdata_0_rfWen),
    .io_wdata_0_fpWen(dispatchData_io_wdata_0_fpWen),
    .io_wdata_0_wflags(dispatchData_io_wdata_0_wflags),
    .io_wdata_0_commitType(dispatchData_io_wdata_0_commitType),
    .io_wdata_0_pdest(dispatchData_io_wdata_0_pdest),
    .io_wdata_0_old_pdest(dispatchData_io_wdata_0_old_pdest),
    .io_wdata_0_ftqIdx_flag(dispatchData_io_wdata_0_ftqIdx_flag),
    .io_wdata_0_ftqIdx_value(dispatchData_io_wdata_0_ftqIdx_value),
    .io_wdata_0_ftqOffset(dispatchData_io_wdata_0_ftqOffset),
    .io_wdata_0_isMove(dispatchData_io_wdata_0_isMove),
    .io_wdata_1_ldest(dispatchData_io_wdata_1_ldest),
    .io_wdata_1_rfWen(dispatchData_io_wdata_1_rfWen),
    .io_wdata_1_fpWen(dispatchData_io_wdata_1_fpWen),
    .io_wdata_1_wflags(dispatchData_io_wdata_1_wflags),
    .io_wdata_1_commitType(dispatchData_io_wdata_1_commitType),
    .io_wdata_1_pdest(dispatchData_io_wdata_1_pdest),
    .io_wdata_1_old_pdest(dispatchData_io_wdata_1_old_pdest),
    .io_wdata_1_ftqIdx_flag(dispatchData_io_wdata_1_ftqIdx_flag),
    .io_wdata_1_ftqIdx_value(dispatchData_io_wdata_1_ftqIdx_value),
    .io_wdata_1_ftqOffset(dispatchData_io_wdata_1_ftqOffset),
    .io_wdata_1_isMove(dispatchData_io_wdata_1_isMove)
  );
  ExceptionGen exceptionGen ( // @[Rob.scala 480:28]
    .clock(exceptionGen_clock),
    .reset(exceptionGen_reset),
    .io_redirect_valid(exceptionGen_io_redirect_valid),
    .io_redirect_bits_robIdx_flag(exceptionGen_io_redirect_bits_robIdx_flag),
    .io_redirect_bits_robIdx_value(exceptionGen_io_redirect_bits_robIdx_value),
    .io_redirect_bits_level(exceptionGen_io_redirect_bits_level),
    .io_flush(exceptionGen_io_flush),
    .io_enq_0_valid(exceptionGen_io_enq_0_valid),
    .io_enq_0_bits_robIdx_flag(exceptionGen_io_enq_0_bits_robIdx_flag),
    .io_enq_0_bits_robIdx_value(exceptionGen_io_enq_0_bits_robIdx_value),
    .io_enq_0_bits_exceptionVec_1(exceptionGen_io_enq_0_bits_exceptionVec_1),
    .io_enq_0_bits_exceptionVec_2(exceptionGen_io_enq_0_bits_exceptionVec_2),
    .io_enq_0_bits_exceptionVec_12(exceptionGen_io_enq_0_bits_exceptionVec_12),
    .io_enq_0_bits_flushPipe(exceptionGen_io_enq_0_bits_flushPipe),
    .io_enq_0_bits_singleStep(exceptionGen_io_enq_0_bits_singleStep),
    .io_enq_0_bits_crossPageIPFFix(exceptionGen_io_enq_0_bits_crossPageIPFFix),
    .io_enq_0_bits_trigger_frontendHit_0(exceptionGen_io_enq_0_bits_trigger_frontendHit_0),
    .io_enq_0_bits_trigger_frontendHit_1(exceptionGen_io_enq_0_bits_trigger_frontendHit_1),
    .io_enq_0_bits_trigger_frontendHit_2(exceptionGen_io_enq_0_bits_trigger_frontendHit_2),
    .io_enq_0_bits_trigger_frontendHit_3(exceptionGen_io_enq_0_bits_trigger_frontendHit_3),
    .io_enq_1_valid(exceptionGen_io_enq_1_valid),
    .io_enq_1_bits_robIdx_flag(exceptionGen_io_enq_1_bits_robIdx_flag),
    .io_enq_1_bits_robIdx_value(exceptionGen_io_enq_1_bits_robIdx_value),
    .io_enq_1_bits_exceptionVec_1(exceptionGen_io_enq_1_bits_exceptionVec_1),
    .io_enq_1_bits_exceptionVec_2(exceptionGen_io_enq_1_bits_exceptionVec_2),
    .io_enq_1_bits_exceptionVec_12(exceptionGen_io_enq_1_bits_exceptionVec_12),
    .io_enq_1_bits_flushPipe(exceptionGen_io_enq_1_bits_flushPipe),
    .io_enq_1_bits_singleStep(exceptionGen_io_enq_1_bits_singleStep),
    .io_enq_1_bits_crossPageIPFFix(exceptionGen_io_enq_1_bits_crossPageIPFFix),
    .io_enq_1_bits_trigger_frontendHit_0(exceptionGen_io_enq_1_bits_trigger_frontendHit_0),
    .io_enq_1_bits_trigger_frontendHit_1(exceptionGen_io_enq_1_bits_trigger_frontendHit_1),
    .io_enq_1_bits_trigger_frontendHit_2(exceptionGen_io_enq_1_bits_trigger_frontendHit_2),
    .io_enq_1_bits_trigger_frontendHit_3(exceptionGen_io_enq_1_bits_trigger_frontendHit_3),
    .io_wb_0_valid(exceptionGen_io_wb_0_valid),
    .io_wb_0_bits_robIdx_flag(exceptionGen_io_wb_0_bits_robIdx_flag),
    .io_wb_0_bits_robIdx_value(exceptionGen_io_wb_0_bits_robIdx_value),
    .io_wb_0_bits_exceptionVec_2(exceptionGen_io_wb_0_bits_exceptionVec_2),
    .io_wb_0_bits_exceptionVec_3(exceptionGen_io_wb_0_bits_exceptionVec_3),
    .io_wb_0_bits_exceptionVec_8(exceptionGen_io_wb_0_bits_exceptionVec_8),
    .io_wb_0_bits_exceptionVec_9(exceptionGen_io_wb_0_bits_exceptionVec_9),
    .io_wb_0_bits_exceptionVec_11(exceptionGen_io_wb_0_bits_exceptionVec_11),
    .io_wb_0_bits_flushPipe(exceptionGen_io_wb_0_bits_flushPipe),
    .io_wb_1_valid(exceptionGen_io_wb_1_valid),
    .io_wb_1_bits_robIdx_flag(exceptionGen_io_wb_1_bits_robIdx_flag),
    .io_wb_1_bits_robIdx_value(exceptionGen_io_wb_1_bits_robIdx_value),
    .io_wb_1_bits_exceptionVec_4(exceptionGen_io_wb_1_bits_exceptionVec_4),
    .io_wb_1_bits_exceptionVec_5(exceptionGen_io_wb_1_bits_exceptionVec_5),
    .io_wb_1_bits_exceptionVec_13(exceptionGen_io_wb_1_bits_exceptionVec_13),
    .io_wb_1_bits_flushPipe(exceptionGen_io_wb_1_bits_flushPipe),
    .io_wb_1_bits_replayInst(exceptionGen_io_wb_1_bits_replayInst),
    .io_wb_1_bits_trigger_backendHit_0(exceptionGen_io_wb_1_bits_trigger_backendHit_0),
    .io_wb_1_bits_trigger_backendHit_1(exceptionGen_io_wb_1_bits_trigger_backendHit_1),
    .io_wb_1_bits_trigger_backendHit_2(exceptionGen_io_wb_1_bits_trigger_backendHit_2),
    .io_wb_1_bits_trigger_backendHit_3(exceptionGen_io_wb_1_bits_trigger_backendHit_3),
    .io_wb_1_bits_trigger_backendHit_4(exceptionGen_io_wb_1_bits_trigger_backendHit_4),
    .io_wb_1_bits_trigger_backendHit_5(exceptionGen_io_wb_1_bits_trigger_backendHit_5),
    .io_wb_2_valid(exceptionGen_io_wb_2_valid),
    .io_wb_2_bits_robIdx_flag(exceptionGen_io_wb_2_bits_robIdx_flag),
    .io_wb_2_bits_robIdx_value(exceptionGen_io_wb_2_bits_robIdx_value),
    .io_wb_2_bits_exceptionVec_4(exceptionGen_io_wb_2_bits_exceptionVec_4),
    .io_wb_2_bits_exceptionVec_5(exceptionGen_io_wb_2_bits_exceptionVec_5),
    .io_wb_2_bits_exceptionVec_13(exceptionGen_io_wb_2_bits_exceptionVec_13),
    .io_wb_2_bits_flushPipe(exceptionGen_io_wb_2_bits_flushPipe),
    .io_wb_2_bits_replayInst(exceptionGen_io_wb_2_bits_replayInst),
    .io_wb_2_bits_trigger_backendHit_0(exceptionGen_io_wb_2_bits_trigger_backendHit_0),
    .io_wb_2_bits_trigger_backendHit_1(exceptionGen_io_wb_2_bits_trigger_backendHit_1),
    .io_wb_2_bits_trigger_backendHit_2(exceptionGen_io_wb_2_bits_trigger_backendHit_2),
    .io_wb_2_bits_trigger_backendHit_3(exceptionGen_io_wb_2_bits_trigger_backendHit_3),
    .io_wb_2_bits_trigger_backendHit_4(exceptionGen_io_wb_2_bits_trigger_backendHit_4),
    .io_wb_2_bits_trigger_backendHit_5(exceptionGen_io_wb_2_bits_trigger_backendHit_5),
    .io_wb_3_valid(exceptionGen_io_wb_3_valid),
    .io_wb_3_bits_robIdx_flag(exceptionGen_io_wb_3_bits_robIdx_flag),
    .io_wb_3_bits_robIdx_value(exceptionGen_io_wb_3_bits_robIdx_value),
    .io_wb_3_bits_exceptionVec_4(exceptionGen_io_wb_3_bits_exceptionVec_4),
    .io_wb_3_bits_exceptionVec_5(exceptionGen_io_wb_3_bits_exceptionVec_5),
    .io_wb_3_bits_exceptionVec_6(exceptionGen_io_wb_3_bits_exceptionVec_6),
    .io_wb_3_bits_exceptionVec_7(exceptionGen_io_wb_3_bits_exceptionVec_7),
    .io_wb_3_bits_exceptionVec_13(exceptionGen_io_wb_3_bits_exceptionVec_13),
    .io_wb_3_bits_exceptionVec_15(exceptionGen_io_wb_3_bits_exceptionVec_15),
    .io_wb_3_bits_trigger_backendHit_0(exceptionGen_io_wb_3_bits_trigger_backendHit_0),
    .io_wb_3_bits_trigger_backendHit_1(exceptionGen_io_wb_3_bits_trigger_backendHit_1),
    .io_wb_3_bits_trigger_backendHit_2(exceptionGen_io_wb_3_bits_trigger_backendHit_2),
    .io_wb_3_bits_trigger_backendHit_3(exceptionGen_io_wb_3_bits_trigger_backendHit_3),
    .io_wb_3_bits_trigger_backendHit_4(exceptionGen_io_wb_3_bits_trigger_backendHit_4),
    .io_wb_3_bits_trigger_backendHit_5(exceptionGen_io_wb_3_bits_trigger_backendHit_5),
    .io_wb_4_valid(exceptionGen_io_wb_4_valid),
    .io_wb_4_bits_robIdx_flag(exceptionGen_io_wb_4_bits_robIdx_flag),
    .io_wb_4_bits_robIdx_value(exceptionGen_io_wb_4_bits_robIdx_value),
    .io_wb_4_bits_exceptionVec_6(exceptionGen_io_wb_4_bits_exceptionVec_6),
    .io_wb_4_bits_exceptionVec_7(exceptionGen_io_wb_4_bits_exceptionVec_7),
    .io_wb_4_bits_exceptionVec_15(exceptionGen_io_wb_4_bits_exceptionVec_15),
    .io_wb_4_bits_trigger_backendHit_0(exceptionGen_io_wb_4_bits_trigger_backendHit_0),
    .io_wb_4_bits_trigger_backendHit_1(exceptionGen_io_wb_4_bits_trigger_backendHit_1),
    .io_wb_4_bits_trigger_backendHit_4(exceptionGen_io_wb_4_bits_trigger_backendHit_4),
    .io_out_valid(exceptionGen_io_out_valid),
    .io_out_bits_robIdx_value(exceptionGen_io_out_bits_robIdx_value),
    .io_state_valid(exceptionGen_io_state_valid),
    .io_state_bits_robIdx_flag(exceptionGen_io_state_bits_robIdx_flag),
    .io_state_bits_robIdx_value(exceptionGen_io_state_bits_robIdx_value),
    .io_state_bits_exceptionVec_0(exceptionGen_io_state_bits_exceptionVec_0),
    .io_state_bits_exceptionVec_1(exceptionGen_io_state_bits_exceptionVec_1),
    .io_state_bits_exceptionVec_2(exceptionGen_io_state_bits_exceptionVec_2),
    .io_state_bits_exceptionVec_3(exceptionGen_io_state_bits_exceptionVec_3),
    .io_state_bits_exceptionVec_4(exceptionGen_io_state_bits_exceptionVec_4),
    .io_state_bits_exceptionVec_5(exceptionGen_io_state_bits_exceptionVec_5),
    .io_state_bits_exceptionVec_6(exceptionGen_io_state_bits_exceptionVec_6),
    .io_state_bits_exceptionVec_7(exceptionGen_io_state_bits_exceptionVec_7),
    .io_state_bits_exceptionVec_8(exceptionGen_io_state_bits_exceptionVec_8),
    .io_state_bits_exceptionVec_9(exceptionGen_io_state_bits_exceptionVec_9),
    .io_state_bits_exceptionVec_10(exceptionGen_io_state_bits_exceptionVec_10),
    .io_state_bits_exceptionVec_11(exceptionGen_io_state_bits_exceptionVec_11),
    .io_state_bits_exceptionVec_12(exceptionGen_io_state_bits_exceptionVec_12),
    .io_state_bits_exceptionVec_13(exceptionGen_io_state_bits_exceptionVec_13),
    .io_state_bits_exceptionVec_14(exceptionGen_io_state_bits_exceptionVec_14),
    .io_state_bits_exceptionVec_15(exceptionGen_io_state_bits_exceptionVec_15),
    .io_state_bits_flushPipe(exceptionGen_io_state_bits_flushPipe),
    .io_state_bits_replayInst(exceptionGen_io_state_bits_replayInst),
    .io_state_bits_singleStep(exceptionGen_io_state_bits_singleStep),
    .io_state_bits_crossPageIPFFix(exceptionGen_io_state_bits_crossPageIPFFix),
    .io_state_bits_trigger_frontendHit_0(exceptionGen_io_state_bits_trigger_frontendHit_0),
    .io_state_bits_trigger_frontendHit_1(exceptionGen_io_state_bits_trigger_frontendHit_1),
    .io_state_bits_trigger_frontendHit_2(exceptionGen_io_state_bits_trigger_frontendHit_2),
    .io_state_bits_trigger_frontendHit_3(exceptionGen_io_state_bits_trigger_frontendHit_3),
    .io_state_bits_trigger_backendHit_0(exceptionGen_io_state_bits_trigger_backendHit_0),
    .io_state_bits_trigger_backendHit_1(exceptionGen_io_state_bits_trigger_backendHit_1),
    .io_state_bits_trigger_backendHit_2(exceptionGen_io_state_bits_trigger_backendHit_2),
    .io_state_bits_trigger_backendHit_3(exceptionGen_io_state_bits_trigger_backendHit_3),
    .io_state_bits_trigger_backendHit_4(exceptionGen_io_state_bits_trigger_backendHit_4),
    .io_state_bits_trigger_backendHit_5(exceptionGen_io_state_bits_trigger_backendHit_5)
  );
  RobDeqPtrWrapper deqPtrGenModule ( // @[Rob.scala 774:31]
    .clock(deqPtrGenModule_clock),
    .reset(deqPtrGenModule_reset),
    .io_state(deqPtrGenModule_io_state),
    .io_deq_v_0(deqPtrGenModule_io_deq_v_0),
    .io_deq_v_1(deqPtrGenModule_io_deq_v_1),
    .io_deq_w0(deqPtrGenModule_io_deq_w0),
    .io_deq_w1(deqPtrGenModule_io_deq_w1),
    .io_exception_state_valid(deqPtrGenModule_io_exception_state_valid),
    .io_exception_state_bits_robIdx_flag(deqPtrGenModule_io_exception_state_bits_robIdx_flag),
    .io_exception_state_bits_robIdx_value(deqPtrGenModule_io_exception_state_bits_robIdx_value),
    .io_exception_state_bits_exceptionVec_0(deqPtrGenModule_io_exception_state_bits_exceptionVec_0),
    .io_exception_state_bits_exceptionVec_1(deqPtrGenModule_io_exception_state_bits_exceptionVec_1),
    .io_exception_state_bits_exceptionVec_2(deqPtrGenModule_io_exception_state_bits_exceptionVec_2),
    .io_exception_state_bits_exceptionVec_3(deqPtrGenModule_io_exception_state_bits_exceptionVec_3),
    .io_exception_state_bits_exceptionVec_4(deqPtrGenModule_io_exception_state_bits_exceptionVec_4),
    .io_exception_state_bits_exceptionVec_5(deqPtrGenModule_io_exception_state_bits_exceptionVec_5),
    .io_exception_state_bits_exceptionVec_6(deqPtrGenModule_io_exception_state_bits_exceptionVec_6),
    .io_exception_state_bits_exceptionVec_7(deqPtrGenModule_io_exception_state_bits_exceptionVec_7),
    .io_exception_state_bits_exceptionVec_8(deqPtrGenModule_io_exception_state_bits_exceptionVec_8),
    .io_exception_state_bits_exceptionVec_9(deqPtrGenModule_io_exception_state_bits_exceptionVec_9),
    .io_exception_state_bits_exceptionVec_10(deqPtrGenModule_io_exception_state_bits_exceptionVec_10),
    .io_exception_state_bits_exceptionVec_11(deqPtrGenModule_io_exception_state_bits_exceptionVec_11),
    .io_exception_state_bits_exceptionVec_12(deqPtrGenModule_io_exception_state_bits_exceptionVec_12),
    .io_exception_state_bits_exceptionVec_13(deqPtrGenModule_io_exception_state_bits_exceptionVec_13),
    .io_exception_state_bits_exceptionVec_14(deqPtrGenModule_io_exception_state_bits_exceptionVec_14),
    .io_exception_state_bits_exceptionVec_15(deqPtrGenModule_io_exception_state_bits_exceptionVec_15),
    .io_exception_state_bits_replayInst(deqPtrGenModule_io_exception_state_bits_replayInst),
    .io_exception_state_bits_singleStep(deqPtrGenModule_io_exception_state_bits_singleStep),
    .io_exception_state_bits_trigger_frontendHit_0(deqPtrGenModule_io_exception_state_bits_trigger_frontendHit_0),
    .io_exception_state_bits_trigger_frontendHit_1(deqPtrGenModule_io_exception_state_bits_trigger_frontendHit_1),
    .io_exception_state_bits_trigger_frontendHit_2(deqPtrGenModule_io_exception_state_bits_trigger_frontendHit_2),
    .io_exception_state_bits_trigger_frontendHit_3(deqPtrGenModule_io_exception_state_bits_trigger_frontendHit_3),
    .io_exception_state_bits_trigger_backendHit_0(deqPtrGenModule_io_exception_state_bits_trigger_backendHit_0),
    .io_exception_state_bits_trigger_backendHit_1(deqPtrGenModule_io_exception_state_bits_trigger_backendHit_1),
    .io_exception_state_bits_trigger_backendHit_2(deqPtrGenModule_io_exception_state_bits_trigger_backendHit_2),
    .io_exception_state_bits_trigger_backendHit_3(deqPtrGenModule_io_exception_state_bits_trigger_backendHit_3),
    .io_exception_state_bits_trigger_backendHit_4(deqPtrGenModule_io_exception_state_bits_trigger_backendHit_4),
    .io_exception_state_bits_trigger_backendHit_5(deqPtrGenModule_io_exception_state_bits_trigger_backendHit_5),
    .io_intrBitSetReg(deqPtrGenModule_io_intrBitSetReg),
    .io_hasNoSpecExec(deqPtrGenModule_io_hasNoSpecExec),
    .io_interrupt_safe(deqPtrGenModule_io_interrupt_safe),
    .io_blockCommit(deqPtrGenModule_io_blockCommit),
    .io_out_0_flag(deqPtrGenModule_io_out_0_flag),
    .io_out_0_value(deqPtrGenModule_io_out_0_value),
    .io_out_1_flag(deqPtrGenModule_io_out_1_flag),
    .io_out_1_value(deqPtrGenModule_io_out_1_value),
    .io_next_out_0_flag(deqPtrGenModule_io_next_out_0_flag),
    .io_next_out_0_value(deqPtrGenModule_io_next_out_0_value),
    .io_next_out_1_flag(deqPtrGenModule_io_next_out_1_flag),
    .io_next_out_1_value(deqPtrGenModule_io_next_out_1_value)
  );
  RobEnqPtrWrapper enqPtrGenModule ( // @[Rob.scala 786:31]
    .clock(enqPtrGenModule_clock),
    .reset(enqPtrGenModule_reset),
    .io_redirect_valid(enqPtrGenModule_io_redirect_valid),
    .io_redirect_bits_robIdx_flag(enqPtrGenModule_io_redirect_bits_robIdx_flag),
    .io_redirect_bits_robIdx_value(enqPtrGenModule_io_redirect_bits_robIdx_value),
    .io_redirect_bits_level(enqPtrGenModule_io_redirect_bits_level),
    .io_allowEnqueue(enqPtrGenModule_io_allowEnqueue),
    .io_hasBlockBackward(enqPtrGenModule_io_hasBlockBackward),
    .io_enq_0(enqPtrGenModule_io_enq_0),
    .io_enq_1(enqPtrGenModule_io_enq_1),
    .io_out_0_flag(enqPtrGenModule_io_out_0_flag),
    .io_out_0_value(enqPtrGenModule_io_out_0_value),
    .io_out_1_value(enqPtrGenModule_io_out_1_value)
  );
  SyncDataModuleTemplate__32entry_1 fflagsDataModule ( // @[Rob.scala 1007:32]
    .clock(fflagsDataModule_clock),
    .io_raddr_0(fflagsDataModule_io_raddr_0),
    .io_raddr_1(fflagsDataModule_io_raddr_1),
    .io_rdata_0(fflagsDataModule_io_rdata_0),
    .io_rdata_1(fflagsDataModule_io_rdata_1),
    .io_wen_0(fflagsDataModule_io_wen_0),
    .io_wen_1(fflagsDataModule_io_wen_1),
    .io_wen_2(fflagsDataModule_io_wen_2),
    .io_waddr_0(fflagsDataModule_io_waddr_0),
    .io_waddr_1(fflagsDataModule_io_waddr_1),
    .io_waddr_2(fflagsDataModule_io_waddr_2),
    .io_wdata_0(fflagsDataModule_io_wdata_0),
    .io_wdata_1(fflagsDataModule_io_wdata_1),
    .io_wdata_2(fflagsDataModule_io_wdata_2)
  );
`ifndef SYNTHESIS
  DifftestBasicInstrCommit difftest ( // @[Rob.scala 1235:28]
    .io_clock(difftest_io_clock),
    .io_coreid(difftest_io_coreid),
    .io_index(difftest_io_index),
    .io_valid(difftest_io_valid),
    .io_special(difftest_io_special),
    .io_skip(difftest_io_skip),
    .io_isRVC(difftest_io_isRVC),
    .io_rfwen(difftest_io_rfwen),
    .io_fpwen(difftest_io_fpwen),
    .io_wpdest(difftest_io_wpdest),
    .io_wdest(difftest_io_wdest)
  );
`endif
`ifndef SYNTHESIS
  DifftestBasicInstrCommit difftest_1 ( // @[Rob.scala 1235:28]
    .io_clock(difftest_1_io_clock),
    .io_coreid(difftest_1_io_coreid),
    .io_index(difftest_1_io_index),
    .io_valid(difftest_1_io_valid),
    .io_special(difftest_1_io_special),
    .io_skip(difftest_1_io_skip),
    .io_isRVC(difftest_1_io_isRVC),
    .io_rfwen(difftest_1_io_rfwen),
    .io_fpwen(difftest_1_io_fpwen),
    .io_wpdest(difftest_1_io_wpdest),
    .io_wdest(difftest_1_io_wdest)
  );
`endif
`ifndef SYNTHESIS
  DifftestBasicTrapEvent difftest_2 ( // @[Rob.scala 1298:26]
    .io_clock(difftest_2_io_clock),
    .io_coreid(difftest_2_io_coreid),
    .io_valid(difftest_2_io_valid),
    .io_cycleCnt(difftest_2_io_cycleCnt),
    .io_instrCnt(difftest_2_io_instrCnt),
    .io_hasWFI(difftest_2_io_hasWFI)
  );
`endif
  assign writebacked_exceptionEnable_MPORT_en = 1'h1;
  assign writebacked_exceptionEnable_MPORT_addr = deqPtrGenModule_io_out_0_value;
  assign writebacked_exceptionEnable_MPORT_data = writebacked[writebacked_exceptionEnable_MPORT_addr]; // @[Rob.scala 428:24]
  assign writebacked_isFlushPipe_MPORT_en = 1'h1;
  assign writebacked_isFlushPipe_MPORT_addr = deqPtrGenModule_io_out_0_value;
  assign writebacked_isFlushPipe_MPORT_data = writebacked[writebacked_isFlushPipe_MPORT_addr]; // @[Rob.scala 428:24]
  assign writebacked_commit_wMPORT_en = 1'h1;
  assign writebacked_commit_wMPORT_addr = deqPtrGenModule_io_out_0_value;
  assign writebacked_commit_wMPORT_data = writebacked[writebacked_commit_wMPORT_addr]; // @[Rob.scala 428:24]
  assign writebacked_commit_wMPORT_2_en = 1'h1;
  assign writebacked_commit_wMPORT_2_addr = deqPtrGenModule_io_out_1_value;
  assign writebacked_commit_wMPORT_2_data = writebacked[writebacked_commit_wMPORT_2_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_113_en = 1'h1;
  assign writebacked_MPORT_113_addr = 5'h0;
  assign writebacked_MPORT_113_data = writebacked[writebacked_MPORT_113_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_114_en = 1'h1;
  assign writebacked_MPORT_114_addr = 5'h0;
  assign writebacked_MPORT_114_data = writebacked[writebacked_MPORT_114_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_115_en = 1'h1;
  assign writebacked_MPORT_115_addr = 5'h1;
  assign writebacked_MPORT_115_data = writebacked[writebacked_MPORT_115_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_116_en = 1'h1;
  assign writebacked_MPORT_116_addr = 5'h1;
  assign writebacked_MPORT_116_data = writebacked[writebacked_MPORT_116_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_117_en = 1'h1;
  assign writebacked_MPORT_117_addr = 5'h2;
  assign writebacked_MPORT_117_data = writebacked[writebacked_MPORT_117_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_118_en = 1'h1;
  assign writebacked_MPORT_118_addr = 5'h2;
  assign writebacked_MPORT_118_data = writebacked[writebacked_MPORT_118_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_119_en = 1'h1;
  assign writebacked_MPORT_119_addr = 5'h3;
  assign writebacked_MPORT_119_data = writebacked[writebacked_MPORT_119_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_120_en = 1'h1;
  assign writebacked_MPORT_120_addr = 5'h3;
  assign writebacked_MPORT_120_data = writebacked[writebacked_MPORT_120_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_121_en = 1'h1;
  assign writebacked_MPORT_121_addr = 5'h4;
  assign writebacked_MPORT_121_data = writebacked[writebacked_MPORT_121_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_122_en = 1'h1;
  assign writebacked_MPORT_122_addr = 5'h4;
  assign writebacked_MPORT_122_data = writebacked[writebacked_MPORT_122_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_123_en = 1'h1;
  assign writebacked_MPORT_123_addr = 5'h5;
  assign writebacked_MPORT_123_data = writebacked[writebacked_MPORT_123_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_124_en = 1'h1;
  assign writebacked_MPORT_124_addr = 5'h5;
  assign writebacked_MPORT_124_data = writebacked[writebacked_MPORT_124_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_125_en = 1'h1;
  assign writebacked_MPORT_125_addr = 5'h6;
  assign writebacked_MPORT_125_data = writebacked[writebacked_MPORT_125_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_126_en = 1'h1;
  assign writebacked_MPORT_126_addr = 5'h6;
  assign writebacked_MPORT_126_data = writebacked[writebacked_MPORT_126_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_127_en = 1'h1;
  assign writebacked_MPORT_127_addr = 5'h7;
  assign writebacked_MPORT_127_data = writebacked[writebacked_MPORT_127_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_128_en = 1'h1;
  assign writebacked_MPORT_128_addr = 5'h7;
  assign writebacked_MPORT_128_data = writebacked[writebacked_MPORT_128_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_129_en = 1'h1;
  assign writebacked_MPORT_129_addr = 5'h8;
  assign writebacked_MPORT_129_data = writebacked[writebacked_MPORT_129_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_130_en = 1'h1;
  assign writebacked_MPORT_130_addr = 5'h8;
  assign writebacked_MPORT_130_data = writebacked[writebacked_MPORT_130_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_131_en = 1'h1;
  assign writebacked_MPORT_131_addr = 5'h9;
  assign writebacked_MPORT_131_data = writebacked[writebacked_MPORT_131_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_132_en = 1'h1;
  assign writebacked_MPORT_132_addr = 5'h9;
  assign writebacked_MPORT_132_data = writebacked[writebacked_MPORT_132_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_133_en = 1'h1;
  assign writebacked_MPORT_133_addr = 5'ha;
  assign writebacked_MPORT_133_data = writebacked[writebacked_MPORT_133_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_134_en = 1'h1;
  assign writebacked_MPORT_134_addr = 5'ha;
  assign writebacked_MPORT_134_data = writebacked[writebacked_MPORT_134_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_135_en = 1'h1;
  assign writebacked_MPORT_135_addr = 5'hb;
  assign writebacked_MPORT_135_data = writebacked[writebacked_MPORT_135_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_136_en = 1'h1;
  assign writebacked_MPORT_136_addr = 5'hb;
  assign writebacked_MPORT_136_data = writebacked[writebacked_MPORT_136_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_137_en = 1'h1;
  assign writebacked_MPORT_137_addr = 5'hc;
  assign writebacked_MPORT_137_data = writebacked[writebacked_MPORT_137_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_138_en = 1'h1;
  assign writebacked_MPORT_138_addr = 5'hc;
  assign writebacked_MPORT_138_data = writebacked[writebacked_MPORT_138_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_139_en = 1'h1;
  assign writebacked_MPORT_139_addr = 5'hd;
  assign writebacked_MPORT_139_data = writebacked[writebacked_MPORT_139_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_140_en = 1'h1;
  assign writebacked_MPORT_140_addr = 5'hd;
  assign writebacked_MPORT_140_data = writebacked[writebacked_MPORT_140_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_141_en = 1'h1;
  assign writebacked_MPORT_141_addr = 5'he;
  assign writebacked_MPORT_141_data = writebacked[writebacked_MPORT_141_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_142_en = 1'h1;
  assign writebacked_MPORT_142_addr = 5'he;
  assign writebacked_MPORT_142_data = writebacked[writebacked_MPORT_142_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_143_en = 1'h1;
  assign writebacked_MPORT_143_addr = 5'hf;
  assign writebacked_MPORT_143_data = writebacked[writebacked_MPORT_143_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_144_en = 1'h1;
  assign writebacked_MPORT_144_addr = 5'hf;
  assign writebacked_MPORT_144_data = writebacked[writebacked_MPORT_144_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_145_en = 1'h1;
  assign writebacked_MPORT_145_addr = 5'h10;
  assign writebacked_MPORT_145_data = writebacked[writebacked_MPORT_145_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_146_en = 1'h1;
  assign writebacked_MPORT_146_addr = 5'h10;
  assign writebacked_MPORT_146_data = writebacked[writebacked_MPORT_146_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_147_en = 1'h1;
  assign writebacked_MPORT_147_addr = 5'h11;
  assign writebacked_MPORT_147_data = writebacked[writebacked_MPORT_147_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_148_en = 1'h1;
  assign writebacked_MPORT_148_addr = 5'h11;
  assign writebacked_MPORT_148_data = writebacked[writebacked_MPORT_148_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_149_en = 1'h1;
  assign writebacked_MPORT_149_addr = 5'h12;
  assign writebacked_MPORT_149_data = writebacked[writebacked_MPORT_149_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_150_en = 1'h1;
  assign writebacked_MPORT_150_addr = 5'h12;
  assign writebacked_MPORT_150_data = writebacked[writebacked_MPORT_150_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_151_en = 1'h1;
  assign writebacked_MPORT_151_addr = 5'h13;
  assign writebacked_MPORT_151_data = writebacked[writebacked_MPORT_151_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_152_en = 1'h1;
  assign writebacked_MPORT_152_addr = 5'h13;
  assign writebacked_MPORT_152_data = writebacked[writebacked_MPORT_152_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_153_en = 1'h1;
  assign writebacked_MPORT_153_addr = 5'h14;
  assign writebacked_MPORT_153_data = writebacked[writebacked_MPORT_153_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_154_en = 1'h1;
  assign writebacked_MPORT_154_addr = 5'h14;
  assign writebacked_MPORT_154_data = writebacked[writebacked_MPORT_154_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_155_en = 1'h1;
  assign writebacked_MPORT_155_addr = 5'h15;
  assign writebacked_MPORT_155_data = writebacked[writebacked_MPORT_155_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_156_en = 1'h1;
  assign writebacked_MPORT_156_addr = 5'h15;
  assign writebacked_MPORT_156_data = writebacked[writebacked_MPORT_156_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_157_en = 1'h1;
  assign writebacked_MPORT_157_addr = 5'h16;
  assign writebacked_MPORT_157_data = writebacked[writebacked_MPORT_157_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_158_en = 1'h1;
  assign writebacked_MPORT_158_addr = 5'h16;
  assign writebacked_MPORT_158_data = writebacked[writebacked_MPORT_158_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_159_en = 1'h1;
  assign writebacked_MPORT_159_addr = 5'h17;
  assign writebacked_MPORT_159_data = writebacked[writebacked_MPORT_159_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_160_en = 1'h1;
  assign writebacked_MPORT_160_addr = 5'h17;
  assign writebacked_MPORT_160_data = writebacked[writebacked_MPORT_160_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_161_en = 1'h1;
  assign writebacked_MPORT_161_addr = 5'h18;
  assign writebacked_MPORT_161_data = writebacked[writebacked_MPORT_161_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_162_en = 1'h1;
  assign writebacked_MPORT_162_addr = 5'h18;
  assign writebacked_MPORT_162_data = writebacked[writebacked_MPORT_162_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_163_en = 1'h1;
  assign writebacked_MPORT_163_addr = 5'h19;
  assign writebacked_MPORT_163_data = writebacked[writebacked_MPORT_163_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_164_en = 1'h1;
  assign writebacked_MPORT_164_addr = 5'h19;
  assign writebacked_MPORT_164_data = writebacked[writebacked_MPORT_164_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_165_en = 1'h1;
  assign writebacked_MPORT_165_addr = 5'h1a;
  assign writebacked_MPORT_165_data = writebacked[writebacked_MPORT_165_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_166_en = 1'h1;
  assign writebacked_MPORT_166_addr = 5'h1a;
  assign writebacked_MPORT_166_data = writebacked[writebacked_MPORT_166_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_167_en = 1'h1;
  assign writebacked_MPORT_167_addr = 5'h1b;
  assign writebacked_MPORT_167_data = writebacked[writebacked_MPORT_167_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_168_en = 1'h1;
  assign writebacked_MPORT_168_addr = 5'h1b;
  assign writebacked_MPORT_168_data = writebacked[writebacked_MPORT_168_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_169_en = 1'h1;
  assign writebacked_MPORT_169_addr = 5'h1c;
  assign writebacked_MPORT_169_data = writebacked[writebacked_MPORT_169_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_170_en = 1'h1;
  assign writebacked_MPORT_170_addr = 5'h1c;
  assign writebacked_MPORT_170_data = writebacked[writebacked_MPORT_170_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_171_en = 1'h1;
  assign writebacked_MPORT_171_addr = 5'h1d;
  assign writebacked_MPORT_171_data = writebacked[writebacked_MPORT_171_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_172_en = 1'h1;
  assign writebacked_MPORT_172_addr = 5'h1d;
  assign writebacked_MPORT_172_data = writebacked[writebacked_MPORT_172_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_173_en = 1'h1;
  assign writebacked_MPORT_173_addr = 5'h1e;
  assign writebacked_MPORT_173_data = writebacked[writebacked_MPORT_173_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_174_en = 1'h1;
  assign writebacked_MPORT_174_addr = 5'h1e;
  assign writebacked_MPORT_174_data = writebacked[writebacked_MPORT_174_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_175_en = 1'h1;
  assign writebacked_MPORT_175_addr = 5'h1f;
  assign writebacked_MPORT_175_data = writebacked[writebacked_MPORT_175_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_176_en = 1'h1;
  assign writebacked_MPORT_176_addr = 5'h1f;
  assign writebacked_MPORT_176_data = writebacked[writebacked_MPORT_176_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_178_en = 1'h1;
  assign writebacked_MPORT_178_addr = 5'h0;
  assign writebacked_MPORT_178_data = writebacked[writebacked_MPORT_178_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_179_en = 1'h1;
  assign writebacked_MPORT_179_addr = 5'h0;
  assign writebacked_MPORT_179_data = writebacked[writebacked_MPORT_179_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_181_en = 1'h1;
  assign writebacked_MPORT_181_addr = 5'h1;
  assign writebacked_MPORT_181_data = writebacked[writebacked_MPORT_181_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_182_en = 1'h1;
  assign writebacked_MPORT_182_addr = 5'h1;
  assign writebacked_MPORT_182_data = writebacked[writebacked_MPORT_182_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_184_en = 1'h1;
  assign writebacked_MPORT_184_addr = 5'h2;
  assign writebacked_MPORT_184_data = writebacked[writebacked_MPORT_184_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_185_en = 1'h1;
  assign writebacked_MPORT_185_addr = 5'h2;
  assign writebacked_MPORT_185_data = writebacked[writebacked_MPORT_185_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_187_en = 1'h1;
  assign writebacked_MPORT_187_addr = 5'h3;
  assign writebacked_MPORT_187_data = writebacked[writebacked_MPORT_187_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_188_en = 1'h1;
  assign writebacked_MPORT_188_addr = 5'h3;
  assign writebacked_MPORT_188_data = writebacked[writebacked_MPORT_188_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_190_en = 1'h1;
  assign writebacked_MPORT_190_addr = 5'h4;
  assign writebacked_MPORT_190_data = writebacked[writebacked_MPORT_190_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_191_en = 1'h1;
  assign writebacked_MPORT_191_addr = 5'h4;
  assign writebacked_MPORT_191_data = writebacked[writebacked_MPORT_191_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_193_en = 1'h1;
  assign writebacked_MPORT_193_addr = 5'h5;
  assign writebacked_MPORT_193_data = writebacked[writebacked_MPORT_193_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_194_en = 1'h1;
  assign writebacked_MPORT_194_addr = 5'h5;
  assign writebacked_MPORT_194_data = writebacked[writebacked_MPORT_194_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_196_en = 1'h1;
  assign writebacked_MPORT_196_addr = 5'h6;
  assign writebacked_MPORT_196_data = writebacked[writebacked_MPORT_196_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_197_en = 1'h1;
  assign writebacked_MPORT_197_addr = 5'h6;
  assign writebacked_MPORT_197_data = writebacked[writebacked_MPORT_197_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_199_en = 1'h1;
  assign writebacked_MPORT_199_addr = 5'h7;
  assign writebacked_MPORT_199_data = writebacked[writebacked_MPORT_199_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_200_en = 1'h1;
  assign writebacked_MPORT_200_addr = 5'h7;
  assign writebacked_MPORT_200_data = writebacked[writebacked_MPORT_200_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_202_en = 1'h1;
  assign writebacked_MPORT_202_addr = 5'h8;
  assign writebacked_MPORT_202_data = writebacked[writebacked_MPORT_202_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_203_en = 1'h1;
  assign writebacked_MPORT_203_addr = 5'h8;
  assign writebacked_MPORT_203_data = writebacked[writebacked_MPORT_203_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_205_en = 1'h1;
  assign writebacked_MPORT_205_addr = 5'h9;
  assign writebacked_MPORT_205_data = writebacked[writebacked_MPORT_205_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_206_en = 1'h1;
  assign writebacked_MPORT_206_addr = 5'h9;
  assign writebacked_MPORT_206_data = writebacked[writebacked_MPORT_206_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_208_en = 1'h1;
  assign writebacked_MPORT_208_addr = 5'ha;
  assign writebacked_MPORT_208_data = writebacked[writebacked_MPORT_208_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_209_en = 1'h1;
  assign writebacked_MPORT_209_addr = 5'ha;
  assign writebacked_MPORT_209_data = writebacked[writebacked_MPORT_209_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_211_en = 1'h1;
  assign writebacked_MPORT_211_addr = 5'hb;
  assign writebacked_MPORT_211_data = writebacked[writebacked_MPORT_211_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_212_en = 1'h1;
  assign writebacked_MPORT_212_addr = 5'hb;
  assign writebacked_MPORT_212_data = writebacked[writebacked_MPORT_212_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_214_en = 1'h1;
  assign writebacked_MPORT_214_addr = 5'hc;
  assign writebacked_MPORT_214_data = writebacked[writebacked_MPORT_214_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_215_en = 1'h1;
  assign writebacked_MPORT_215_addr = 5'hc;
  assign writebacked_MPORT_215_data = writebacked[writebacked_MPORT_215_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_217_en = 1'h1;
  assign writebacked_MPORT_217_addr = 5'hd;
  assign writebacked_MPORT_217_data = writebacked[writebacked_MPORT_217_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_218_en = 1'h1;
  assign writebacked_MPORT_218_addr = 5'hd;
  assign writebacked_MPORT_218_data = writebacked[writebacked_MPORT_218_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_220_en = 1'h1;
  assign writebacked_MPORT_220_addr = 5'he;
  assign writebacked_MPORT_220_data = writebacked[writebacked_MPORT_220_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_221_en = 1'h1;
  assign writebacked_MPORT_221_addr = 5'he;
  assign writebacked_MPORT_221_data = writebacked[writebacked_MPORT_221_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_223_en = 1'h1;
  assign writebacked_MPORT_223_addr = 5'hf;
  assign writebacked_MPORT_223_data = writebacked[writebacked_MPORT_223_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_224_en = 1'h1;
  assign writebacked_MPORT_224_addr = 5'hf;
  assign writebacked_MPORT_224_data = writebacked[writebacked_MPORT_224_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_226_en = 1'h1;
  assign writebacked_MPORT_226_addr = 5'h10;
  assign writebacked_MPORT_226_data = writebacked[writebacked_MPORT_226_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_227_en = 1'h1;
  assign writebacked_MPORT_227_addr = 5'h10;
  assign writebacked_MPORT_227_data = writebacked[writebacked_MPORT_227_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_229_en = 1'h1;
  assign writebacked_MPORT_229_addr = 5'h11;
  assign writebacked_MPORT_229_data = writebacked[writebacked_MPORT_229_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_230_en = 1'h1;
  assign writebacked_MPORT_230_addr = 5'h11;
  assign writebacked_MPORT_230_data = writebacked[writebacked_MPORT_230_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_232_en = 1'h1;
  assign writebacked_MPORT_232_addr = 5'h12;
  assign writebacked_MPORT_232_data = writebacked[writebacked_MPORT_232_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_233_en = 1'h1;
  assign writebacked_MPORT_233_addr = 5'h12;
  assign writebacked_MPORT_233_data = writebacked[writebacked_MPORT_233_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_235_en = 1'h1;
  assign writebacked_MPORT_235_addr = 5'h13;
  assign writebacked_MPORT_235_data = writebacked[writebacked_MPORT_235_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_236_en = 1'h1;
  assign writebacked_MPORT_236_addr = 5'h13;
  assign writebacked_MPORT_236_data = writebacked[writebacked_MPORT_236_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_238_en = 1'h1;
  assign writebacked_MPORT_238_addr = 5'h14;
  assign writebacked_MPORT_238_data = writebacked[writebacked_MPORT_238_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_239_en = 1'h1;
  assign writebacked_MPORT_239_addr = 5'h14;
  assign writebacked_MPORT_239_data = writebacked[writebacked_MPORT_239_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_241_en = 1'h1;
  assign writebacked_MPORT_241_addr = 5'h15;
  assign writebacked_MPORT_241_data = writebacked[writebacked_MPORT_241_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_242_en = 1'h1;
  assign writebacked_MPORT_242_addr = 5'h15;
  assign writebacked_MPORT_242_data = writebacked[writebacked_MPORT_242_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_244_en = 1'h1;
  assign writebacked_MPORT_244_addr = 5'h16;
  assign writebacked_MPORT_244_data = writebacked[writebacked_MPORT_244_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_245_en = 1'h1;
  assign writebacked_MPORT_245_addr = 5'h16;
  assign writebacked_MPORT_245_data = writebacked[writebacked_MPORT_245_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_247_en = 1'h1;
  assign writebacked_MPORT_247_addr = 5'h17;
  assign writebacked_MPORT_247_data = writebacked[writebacked_MPORT_247_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_248_en = 1'h1;
  assign writebacked_MPORT_248_addr = 5'h17;
  assign writebacked_MPORT_248_data = writebacked[writebacked_MPORT_248_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_250_en = 1'h1;
  assign writebacked_MPORT_250_addr = 5'h18;
  assign writebacked_MPORT_250_data = writebacked[writebacked_MPORT_250_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_251_en = 1'h1;
  assign writebacked_MPORT_251_addr = 5'h18;
  assign writebacked_MPORT_251_data = writebacked[writebacked_MPORT_251_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_253_en = 1'h1;
  assign writebacked_MPORT_253_addr = 5'h19;
  assign writebacked_MPORT_253_data = writebacked[writebacked_MPORT_253_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_254_en = 1'h1;
  assign writebacked_MPORT_254_addr = 5'h19;
  assign writebacked_MPORT_254_data = writebacked[writebacked_MPORT_254_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_256_en = 1'h1;
  assign writebacked_MPORT_256_addr = 5'h1a;
  assign writebacked_MPORT_256_data = writebacked[writebacked_MPORT_256_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_257_en = 1'h1;
  assign writebacked_MPORT_257_addr = 5'h1a;
  assign writebacked_MPORT_257_data = writebacked[writebacked_MPORT_257_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_259_en = 1'h1;
  assign writebacked_MPORT_259_addr = 5'h1b;
  assign writebacked_MPORT_259_data = writebacked[writebacked_MPORT_259_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_260_en = 1'h1;
  assign writebacked_MPORT_260_addr = 5'h1b;
  assign writebacked_MPORT_260_data = writebacked[writebacked_MPORT_260_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_262_en = 1'h1;
  assign writebacked_MPORT_262_addr = 5'h1c;
  assign writebacked_MPORT_262_data = writebacked[writebacked_MPORT_262_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_263_en = 1'h1;
  assign writebacked_MPORT_263_addr = 5'h1c;
  assign writebacked_MPORT_263_data = writebacked[writebacked_MPORT_263_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_265_en = 1'h1;
  assign writebacked_MPORT_265_addr = 5'h1d;
  assign writebacked_MPORT_265_data = writebacked[writebacked_MPORT_265_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_266_en = 1'h1;
  assign writebacked_MPORT_266_addr = 5'h1d;
  assign writebacked_MPORT_266_data = writebacked[writebacked_MPORT_266_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_268_en = 1'h1;
  assign writebacked_MPORT_268_addr = 5'h1e;
  assign writebacked_MPORT_268_data = writebacked[writebacked_MPORT_268_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_269_en = 1'h1;
  assign writebacked_MPORT_269_addr = 5'h1e;
  assign writebacked_MPORT_269_data = writebacked[writebacked_MPORT_269_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_271_en = 1'h1;
  assign writebacked_MPORT_271_addr = 5'h1f;
  assign writebacked_MPORT_271_data = writebacked[writebacked_MPORT_271_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_272_en = 1'h1;
  assign writebacked_MPORT_272_addr = 5'h1f;
  assign writebacked_MPORT_272_data = writebacked[writebacked_MPORT_272_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_273_en = 1'h1;
  assign writebacked_MPORT_273_addr = 5'h0;
  assign writebacked_MPORT_273_data = writebacked[writebacked_MPORT_273_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_274_en = 1'h1;
  assign writebacked_MPORT_274_addr = 5'h1;
  assign writebacked_MPORT_274_data = writebacked[writebacked_MPORT_274_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_275_en = 1'h1;
  assign writebacked_MPORT_275_addr = 5'h2;
  assign writebacked_MPORT_275_data = writebacked[writebacked_MPORT_275_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_276_en = 1'h1;
  assign writebacked_MPORT_276_addr = 5'h3;
  assign writebacked_MPORT_276_data = writebacked[writebacked_MPORT_276_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_277_en = 1'h1;
  assign writebacked_MPORT_277_addr = 5'h4;
  assign writebacked_MPORT_277_data = writebacked[writebacked_MPORT_277_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_278_en = 1'h1;
  assign writebacked_MPORT_278_addr = 5'h5;
  assign writebacked_MPORT_278_data = writebacked[writebacked_MPORT_278_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_279_en = 1'h1;
  assign writebacked_MPORT_279_addr = 5'h6;
  assign writebacked_MPORT_279_data = writebacked[writebacked_MPORT_279_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_280_en = 1'h1;
  assign writebacked_MPORT_280_addr = 5'h7;
  assign writebacked_MPORT_280_data = writebacked[writebacked_MPORT_280_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_281_en = 1'h1;
  assign writebacked_MPORT_281_addr = 5'h8;
  assign writebacked_MPORT_281_data = writebacked[writebacked_MPORT_281_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_282_en = 1'h1;
  assign writebacked_MPORT_282_addr = 5'h9;
  assign writebacked_MPORT_282_data = writebacked[writebacked_MPORT_282_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_283_en = 1'h1;
  assign writebacked_MPORT_283_addr = 5'ha;
  assign writebacked_MPORT_283_data = writebacked[writebacked_MPORT_283_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_284_en = 1'h1;
  assign writebacked_MPORT_284_addr = 5'hb;
  assign writebacked_MPORT_284_data = writebacked[writebacked_MPORT_284_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_285_en = 1'h1;
  assign writebacked_MPORT_285_addr = 5'hc;
  assign writebacked_MPORT_285_data = writebacked[writebacked_MPORT_285_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_286_en = 1'h1;
  assign writebacked_MPORT_286_addr = 5'hd;
  assign writebacked_MPORT_286_data = writebacked[writebacked_MPORT_286_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_287_en = 1'h1;
  assign writebacked_MPORT_287_addr = 5'he;
  assign writebacked_MPORT_287_data = writebacked[writebacked_MPORT_287_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_288_en = 1'h1;
  assign writebacked_MPORT_288_addr = 5'hf;
  assign writebacked_MPORT_288_data = writebacked[writebacked_MPORT_288_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_289_en = 1'h1;
  assign writebacked_MPORT_289_addr = 5'h10;
  assign writebacked_MPORT_289_data = writebacked[writebacked_MPORT_289_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_290_en = 1'h1;
  assign writebacked_MPORT_290_addr = 5'h11;
  assign writebacked_MPORT_290_data = writebacked[writebacked_MPORT_290_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_291_en = 1'h1;
  assign writebacked_MPORT_291_addr = 5'h12;
  assign writebacked_MPORT_291_data = writebacked[writebacked_MPORT_291_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_292_en = 1'h1;
  assign writebacked_MPORT_292_addr = 5'h13;
  assign writebacked_MPORT_292_data = writebacked[writebacked_MPORT_292_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_293_en = 1'h1;
  assign writebacked_MPORT_293_addr = 5'h14;
  assign writebacked_MPORT_293_data = writebacked[writebacked_MPORT_293_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_294_en = 1'h1;
  assign writebacked_MPORT_294_addr = 5'h15;
  assign writebacked_MPORT_294_data = writebacked[writebacked_MPORT_294_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_295_en = 1'h1;
  assign writebacked_MPORT_295_addr = 5'h16;
  assign writebacked_MPORT_295_data = writebacked[writebacked_MPORT_295_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_296_en = 1'h1;
  assign writebacked_MPORT_296_addr = 5'h17;
  assign writebacked_MPORT_296_data = writebacked[writebacked_MPORT_296_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_297_en = 1'h1;
  assign writebacked_MPORT_297_addr = 5'h18;
  assign writebacked_MPORT_297_data = writebacked[writebacked_MPORT_297_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_298_en = 1'h1;
  assign writebacked_MPORT_298_addr = 5'h19;
  assign writebacked_MPORT_298_data = writebacked[writebacked_MPORT_298_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_299_en = 1'h1;
  assign writebacked_MPORT_299_addr = 5'h1a;
  assign writebacked_MPORT_299_data = writebacked[writebacked_MPORT_299_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_300_en = 1'h1;
  assign writebacked_MPORT_300_addr = 5'h1b;
  assign writebacked_MPORT_300_data = writebacked[writebacked_MPORT_300_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_301_en = 1'h1;
  assign writebacked_MPORT_301_addr = 5'h1c;
  assign writebacked_MPORT_301_data = writebacked[writebacked_MPORT_301_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_302_en = 1'h1;
  assign writebacked_MPORT_302_addr = 5'h1d;
  assign writebacked_MPORT_302_data = writebacked[writebacked_MPORT_302_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_303_en = 1'h1;
  assign writebacked_MPORT_303_addr = 5'h1e;
  assign writebacked_MPORT_303_data = writebacked[writebacked_MPORT_303_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_304_en = 1'h1;
  assign writebacked_MPORT_304_addr = 5'h1f;
  assign writebacked_MPORT_304_data = writebacked[writebacked_MPORT_304_addr]; // @[Rob.scala 428:24]
  assign writebacked_deqNotWritebacked_MPORT_en = 1'h1;
  assign writebacked_deqNotWritebacked_MPORT_addr = deqPtrGenModule_io_out_0_value;
  assign writebacked_deqNotWritebacked_MPORT_data = writebacked[writebacked_deqNotWritebacked_MPORT_addr]; // @[Rob.scala 428:24]
  assign writebacked_MPORT_92_data = _T_149 & _T_11;
  assign writebacked_MPORT_92_addr = enqPtrGenModule_io_out_0_value;
  assign writebacked_MPORT_92_mask = 1'h1;
  assign writebacked_MPORT_92_en = io_enq_req_0_valid & io_enq_canAccept;
  assign writebacked_MPORT_94_data = _T_154 & _T_50;
  assign writebacked_MPORT_94_addr = io_enq_needAlloc_0 ? enqPtrVec_1_value : enqPtrVec_0_value;
  assign writebacked_MPORT_94_mask = 1'h1;
  assign writebacked_MPORT_94_en = io_enq_req_1_valid & io_enq_canAccept;
  assign writebacked_MPORT_96_data = 1'h1;
  assign writebacked_MPORT_96_addr = exceptionGen_io_out_bits_robIdx_value;
  assign writebacked_MPORT_96_mask = 1'h1;
  assign writebacked_MPORT_96_en = exceptionGen_io_out_valid;
  assign writebacked_MPORT_98_data = 1'h1;
  assign writebacked_MPORT_98_addr = io_writeback_1_0_bits_uop_robIdx_value;
  assign writebacked_MPORT_98_mask = 1'h1;
  assign writebacked_MPORT_98_en = io_writeback_1_0_valid;
  assign writebacked_MPORT_99_data = 1'h1;
  assign writebacked_MPORT_99_addr = io_writeback_1_1_bits_uop_robIdx_value;
  assign writebacked_MPORT_99_mask = 1'h1;
  assign writebacked_MPORT_99_en = io_writeback_1_1_valid;
  assign writebacked_MPORT_100_data = ~block_wb_2;
  assign writebacked_MPORT_100_addr = io_writeback_1_2_bits_uop_robIdx_value;
  assign writebacked_MPORT_100_mask = 1'h1;
  assign writebacked_MPORT_100_en = io_writeback_1_2_valid;
  assign writebacked_MPORT_101_data = ~block_wb_3;
  assign writebacked_MPORT_101_addr = io_writeback_1_3_bits_uop_robIdx_value;
  assign writebacked_MPORT_101_mask = 1'h1;
  assign writebacked_MPORT_101_en = io_writeback_1_3_valid;
  assign writebacked_MPORT_102_data = ~block_wb_4;
  assign writebacked_MPORT_102_addr = io_writeback_1_4_bits_uop_robIdx_value;
  assign writebacked_MPORT_102_mask = 1'h1;
  assign writebacked_MPORT_102_en = io_writeback_1_4_valid;
  assign writebacked_MPORT_103_data = ~wbHasTriggerHit_5;
  assign writebacked_MPORT_103_addr = io_writeback_1_5_bits_uop_robIdx_value;
  assign writebacked_MPORT_103_mask = 1'h1;
  assign writebacked_MPORT_103_en = io_writeback_1_5_valid;
  assign writebacked_MPORT_104_data = ~block_wb_6;
  assign writebacked_MPORT_104_addr = io_writeback_1_6_bits_uop_robIdx_value;
  assign writebacked_MPORT_104_mask = 1'h1;
  assign writebacked_MPORT_104_en = io_writeback_1_6_valid;
  assign writebacked_MPORT_105_data = ~block_wb_7;
  assign writebacked_MPORT_105_addr = io_writeback_1_7_bits_uop_robIdx_value;
  assign writebacked_MPORT_105_mask = 1'h1;
  assign writebacked_MPORT_105_en = io_writeback_1_7_valid;
  assign writebacked_MPORT_106_data = ~block_wb_8;
  assign writebacked_MPORT_106_addr = io_writeback_1_8_bits_uop_robIdx_value;
  assign writebacked_MPORT_106_mask = 1'h1;
  assign writebacked_MPORT_106_en = io_writeback_1_8_valid;
  assign store_data_writebacked_commit_wMPORT_1_en = 1'h1;
  assign store_data_writebacked_commit_wMPORT_1_addr = deqPtrGenModule_io_out_0_value;
  assign store_data_writebacked_commit_wMPORT_1_data =
    store_data_writebacked[store_data_writebacked_commit_wMPORT_1_addr]; // @[Rob.scala 429:35]
  assign store_data_writebacked_commit_wMPORT_3_en = 1'h1;
  assign store_data_writebacked_commit_wMPORT_3_addr = deqPtrGenModule_io_out_1_value;
  assign store_data_writebacked_commit_wMPORT_3_data =
    store_data_writebacked[store_data_writebacked_commit_wMPORT_3_addr]; // @[Rob.scala 429:35]
  assign store_data_writebacked_MPORT_93_data = ~isStu;
  assign store_data_writebacked_MPORT_93_addr = enqPtrGenModule_io_out_0_value;
  assign store_data_writebacked_MPORT_93_mask = 1'h1;
  assign store_data_writebacked_MPORT_93_en = io_enq_req_0_valid & io_enq_canAccept;
  assign store_data_writebacked_MPORT_95_data = ~isStu_1;
  assign store_data_writebacked_MPORT_95_addr = io_enq_needAlloc_0 ? enqPtrVec_1_value : enqPtrVec_0_value;
  assign store_data_writebacked_MPORT_95_mask = 1'h1;
  assign store_data_writebacked_MPORT_95_en = io_enq_req_1_valid & io_enq_canAccept;
  assign store_data_writebacked_MPORT_97_data = 1'h1;
  assign store_data_writebacked_MPORT_97_addr = exceptionGen_io_out_bits_robIdx_value;
  assign store_data_writebacked_MPORT_97_mask = 1'h1;
  assign store_data_writebacked_MPORT_97_en = exceptionGen_io_out_valid;
  assign store_data_writebacked_MPORT_107_data = 1'h1;
  assign store_data_writebacked_MPORT_107_addr = REG_8;
  assign store_data_writebacked_MPORT_107_mask = 1'h1;
  assign store_data_writebacked_MPORT_107_en = REG_7;
  assign store_data_writebacked_MPORT_108_data = 1'h1;
  assign store_data_writebacked_MPORT_108_addr = REG_10;
  assign store_data_writebacked_MPORT_108_mask = 1'h1;
  assign store_data_writebacked_MPORT_108_en = REG_9;
  assign interrupt_safe_intrEnable_MPORT_en = 1'h1;
  assign interrupt_safe_intrEnable_MPORT_addr = deqPtrGenModule_io_out_0_value;
  assign interrupt_safe_intrEnable_MPORT_data = interrupt_safe[interrupt_safe_intrEnable_MPORT_addr]; // @[Rob.scala 436:27]
  assign interrupt_safe_deqPtrGenModule_io_interrupt_safe_MPORT_en = 1'h1;
  assign interrupt_safe_deqPtrGenModule_io_interrupt_safe_MPORT_addr = deqPtrGenModule_io_out_0_value;
  assign interrupt_safe_deqPtrGenModule_io_interrupt_safe_MPORT_data =
    interrupt_safe[interrupt_safe_deqPtrGenModule_io_interrupt_safe_MPORT_addr]; // @[Rob.scala 436:27]
  assign interrupt_safe_MPORT_111_data = REG_13;
  assign interrupt_safe_MPORT_111_addr = REG_12;
  assign interrupt_safe_MPORT_111_mask = 1'h1;
  assign interrupt_safe_MPORT_111_en = REG_11;
  assign interrupt_safe_MPORT_112_data = REG_16;
  assign interrupt_safe_MPORT_112_addr = REG_15;
  assign interrupt_safe_MPORT_112_mask = 1'h1;
  assign interrupt_safe_MPORT_112_en = REG_14;
  assign debug_microOp_cf_loadWaitBit_debug_deqUop_en = 1'h1;
  assign debug_microOp_cf_loadWaitBit_debug_deqUop_addr = deqPtrGenModule_io_out_0_value;
  assign debug_microOp_cf_loadWaitBit_debug_deqUop_data =
    debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_debug_deqUop_addr]; // @[Rob.scala 440:26]
  assign debug_microOp_cf_loadWaitBit_commitDebugUop_0_en = 1'h1;
  assign debug_microOp_cf_loadWaitBit_commitDebugUop_0_addr = deqPtrGenModule_io_out_0_value;
  assign debug_microOp_cf_loadWaitBit_commitDebugUop_0_data =
    debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_commitDebugUop_0_addr]; // @[Rob.scala 440:26]
  assign debug_microOp_cf_loadWaitBit_commitDebugUop_1_en = 1'h1;
  assign debug_microOp_cf_loadWaitBit_commitDebugUop_1_addr = deqPtrGenModule_io_out_1_value;
  assign debug_microOp_cf_loadWaitBit_commitDebugUop_1_data =
    debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_commitDebugUop_1_addr]; // @[Rob.scala 440:26]
  assign debug_microOp_cf_loadWaitBit_MPORT_data = io_enq_req_0_bits_cf_loadWaitBit;
  assign debug_microOp_cf_loadWaitBit_MPORT_addr = enqPtrGenModule_io_out_0_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_mask = 1'h1;
  assign debug_microOp_cf_loadWaitBit_MPORT_en = io_enq_req_0_valid & io_enq_canAccept;
  assign debug_microOp_cf_loadWaitBit_MPORT_1_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_1_addr = enqPtrGenModule_io_out_0_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_1_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_1_en = io_enq_req_0_valid & io_enq_canAccept;
  assign debug_microOp_cf_loadWaitBit_MPORT_2_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_2_addr = enqPtrGenModule_io_out_0_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_2_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_2_en = io_enq_req_0_valid & io_enq_canAccept;
  assign debug_microOp_cf_loadWaitBit_MPORT_3_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_3_addr = enqPtrGenModule_io_out_0_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_3_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_3_en = io_enq_req_0_valid & io_enq_canAccept;
  assign debug_microOp_cf_loadWaitBit_MPORT_4_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_4_addr = enqPtrGenModule_io_out_0_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_4_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_4_en = io_enq_req_0_valid & io_enq_canAccept;
  assign debug_microOp_cf_loadWaitBit_MPORT_5_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_5_addr = enqPtrGenModule_io_out_0_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_5_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_5_en = io_enq_req_0_valid & io_enq_canAccept;
  assign debug_microOp_cf_loadWaitBit_MPORT_6_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_6_addr = enqPtrGenModule_io_out_0_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_6_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_6_en = io_enq_req_0_valid & io_enq_canAccept;
  assign debug_microOp_cf_loadWaitBit_MPORT_7_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_7_addr = enqPtrGenModule_io_out_0_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_7_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_7_en = io_enq_req_0_valid & io_enq_canAccept;
  assign debug_microOp_cf_loadWaitBit_MPORT_8_data = io_enq_req_1_bits_cf_loadWaitBit;
  assign debug_microOp_cf_loadWaitBit_MPORT_8_addr = io_enq_needAlloc_0 ? enqPtrVec_1_value : enqPtrVec_0_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_8_mask = 1'h1;
  assign debug_microOp_cf_loadWaitBit_MPORT_8_en = io_enq_req_1_valid & io_enq_canAccept;
  assign debug_microOp_cf_loadWaitBit_MPORT_9_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_9_addr = io_enq_needAlloc_0 ? enqPtrVec_1_value : enqPtrVec_0_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_9_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_9_en = io_enq_req_1_valid & io_enq_canAccept;
  assign debug_microOp_cf_loadWaitBit_MPORT_10_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_10_addr = io_enq_needAlloc_0 ? enqPtrVec_1_value : enqPtrVec_0_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_10_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_10_en = io_enq_req_1_valid & io_enq_canAccept;
  assign debug_microOp_cf_loadWaitBit_MPORT_11_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_11_addr = io_enq_needAlloc_0 ? enqPtrVec_1_value : enqPtrVec_0_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_11_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_11_en = io_enq_req_1_valid & io_enq_canAccept;
  assign debug_microOp_cf_loadWaitBit_MPORT_12_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_12_addr = io_enq_needAlloc_0 ? enqPtrVec_1_value : enqPtrVec_0_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_12_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_12_en = io_enq_req_1_valid & io_enq_canAccept;
  assign debug_microOp_cf_loadWaitBit_MPORT_13_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_13_addr = io_enq_needAlloc_0 ? enqPtrVec_1_value : enqPtrVec_0_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_13_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_13_en = io_enq_req_1_valid & io_enq_canAccept;
  assign debug_microOp_cf_loadWaitBit_MPORT_14_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_14_addr = io_enq_needAlloc_0 ? enqPtrVec_1_value : enqPtrVec_0_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_14_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_14_en = io_enq_req_1_valid & io_enq_canAccept;
  assign debug_microOp_cf_loadWaitBit_MPORT_15_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_15_addr = io_enq_needAlloc_0 ? enqPtrVec_1_value : enqPtrVec_0_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_15_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_15_en = io_enq_req_1_valid & io_enq_canAccept;
  assign debug_microOp_cf_loadWaitBit_MPORT_16_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_16_addr = io_writeback_1_0_bits_uop_robIdx_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_16_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_16_en = io_writeback_1_0_valid;
  assign debug_microOp_cf_loadWaitBit_MPORT_17_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_17_addr = io_writeback_1_0_bits_uop_robIdx_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_17_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_17_en = io_writeback_1_0_valid;
  assign debug_microOp_cf_loadWaitBit_MPORT_18_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_18_addr = io_writeback_1_0_bits_uop_robIdx_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_18_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_18_en = io_writeback_1_0_valid;
  assign debug_microOp_cf_loadWaitBit_MPORT_19_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_19_addr = io_writeback_1_0_bits_uop_robIdx_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_19_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_19_en = io_writeback_1_0_valid;
  assign debug_microOp_cf_loadWaitBit_MPORT_20_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_20_addr = io_writeback_1_0_bits_uop_robIdx_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_20_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_20_en = io_writeback_1_0_valid;
  assign debug_microOp_cf_loadWaitBit_MPORT_21_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_21_addr = io_writeback_1_0_bits_uop_robIdx_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_21_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_21_en = io_writeback_1_0_valid;
  assign debug_microOp_cf_loadWaitBit_MPORT_22_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_22_addr = io_writeback_1_0_bits_uop_robIdx_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_22_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_22_en = io_writeback_1_0_valid;
  assign debug_microOp_cf_loadWaitBit_MPORT_23_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_23_addr = io_writeback_1_0_bits_uop_robIdx_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_23_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_23_en = io_writeback_1_0_valid;
  assign debug_microOp_cf_loadWaitBit_MPORT_24_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_24_addr = io_writeback_1_1_bits_uop_robIdx_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_24_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_24_en = io_writeback_1_1_valid;
  assign debug_microOp_cf_loadWaitBit_MPORT_25_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_25_addr = io_writeback_1_1_bits_uop_robIdx_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_25_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_25_en = io_writeback_1_1_valid;
  assign debug_microOp_cf_loadWaitBit_MPORT_26_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_26_addr = io_writeback_1_1_bits_uop_robIdx_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_26_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_26_en = io_writeback_1_1_valid;
  assign debug_microOp_cf_loadWaitBit_MPORT_27_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_27_addr = io_writeback_1_1_bits_uop_robIdx_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_27_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_27_en = io_writeback_1_1_valid;
  assign debug_microOp_cf_loadWaitBit_MPORT_28_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_28_addr = io_writeback_1_1_bits_uop_robIdx_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_28_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_28_en = io_writeback_1_1_valid;
  assign debug_microOp_cf_loadWaitBit_MPORT_29_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_29_addr = io_writeback_1_1_bits_uop_robIdx_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_29_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_29_en = io_writeback_1_1_valid;
  assign debug_microOp_cf_loadWaitBit_MPORT_30_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_30_addr = io_writeback_1_1_bits_uop_robIdx_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_30_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_30_en = io_writeback_1_1_valid;
  assign debug_microOp_cf_loadWaitBit_MPORT_31_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_31_addr = io_writeback_1_1_bits_uop_robIdx_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_31_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_31_en = io_writeback_1_1_valid;
  assign debug_microOp_cf_loadWaitBit_MPORT_32_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_32_addr = io_writeback_1_2_bits_uop_robIdx_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_32_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_32_en = io_writeback_1_2_valid;
  assign debug_microOp_cf_loadWaitBit_MPORT_33_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_33_addr = io_writeback_1_2_bits_uop_robIdx_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_33_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_33_en = io_writeback_1_2_valid;
  assign debug_microOp_cf_loadWaitBit_MPORT_34_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_34_addr = io_writeback_1_2_bits_uop_robIdx_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_34_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_34_en = io_writeback_1_2_valid;
  assign debug_microOp_cf_loadWaitBit_MPORT_35_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_35_addr = io_writeback_1_2_bits_uop_robIdx_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_35_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_35_en = io_writeback_1_2_valid;
  assign debug_microOp_cf_loadWaitBit_MPORT_36_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_36_addr = io_writeback_1_2_bits_uop_robIdx_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_36_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_36_en = io_writeback_1_2_valid;
  assign debug_microOp_cf_loadWaitBit_MPORT_37_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_37_addr = io_writeback_1_2_bits_uop_robIdx_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_37_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_37_en = io_writeback_1_2_valid;
  assign debug_microOp_cf_loadWaitBit_MPORT_38_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_38_addr = io_writeback_1_2_bits_uop_robIdx_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_38_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_38_en = io_writeback_1_2_valid;
  assign debug_microOp_cf_loadWaitBit_MPORT_39_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_39_addr = io_writeback_1_2_bits_uop_robIdx_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_39_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_39_en = io_writeback_1_2_valid;
  assign debug_microOp_cf_loadWaitBit_MPORT_40_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_40_addr = io_writeback_1_3_bits_uop_robIdx_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_40_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_40_en = io_writeback_1_3_valid;
  assign debug_microOp_cf_loadWaitBit_MPORT_41_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_41_addr = io_writeback_1_3_bits_uop_robIdx_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_41_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_41_en = io_writeback_1_3_valid;
  assign debug_microOp_cf_loadWaitBit_MPORT_42_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_42_addr = io_writeback_1_3_bits_uop_robIdx_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_42_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_42_en = io_writeback_1_3_valid;
  assign debug_microOp_cf_loadWaitBit_MPORT_43_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_43_addr = io_writeback_1_3_bits_uop_robIdx_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_43_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_43_en = io_writeback_1_3_valid;
  assign debug_microOp_cf_loadWaitBit_MPORT_44_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_44_addr = io_writeback_1_3_bits_uop_robIdx_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_44_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_44_en = io_writeback_1_3_valid;
  assign debug_microOp_cf_loadWaitBit_MPORT_45_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_45_addr = io_writeback_1_3_bits_uop_robIdx_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_45_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_45_en = io_writeback_1_3_valid;
  assign debug_microOp_cf_loadWaitBit_MPORT_46_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_46_addr = io_writeback_1_3_bits_uop_robIdx_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_46_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_46_en = io_writeback_1_3_valid;
  assign debug_microOp_cf_loadWaitBit_MPORT_47_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_47_addr = io_writeback_1_3_bits_uop_robIdx_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_47_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_47_en = io_writeback_1_3_valid;
  assign debug_microOp_cf_loadWaitBit_MPORT_48_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_48_addr = io_writeback_1_4_bits_uop_robIdx_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_48_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_48_en = io_writeback_1_4_valid;
  assign debug_microOp_cf_loadWaitBit_MPORT_49_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_49_addr = io_writeback_1_4_bits_uop_robIdx_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_49_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_49_en = io_writeback_1_4_valid;
  assign debug_microOp_cf_loadWaitBit_MPORT_50_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_50_addr = io_writeback_1_4_bits_uop_robIdx_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_50_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_50_en = io_writeback_1_4_valid;
  assign debug_microOp_cf_loadWaitBit_MPORT_51_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_51_addr = io_writeback_1_4_bits_uop_robIdx_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_51_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_51_en = io_writeback_1_4_valid;
  assign debug_microOp_cf_loadWaitBit_MPORT_52_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_52_addr = io_writeback_1_4_bits_uop_robIdx_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_52_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_52_en = io_writeback_1_4_valid;
  assign debug_microOp_cf_loadWaitBit_MPORT_53_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_53_addr = io_writeback_1_4_bits_uop_robIdx_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_53_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_53_en = io_writeback_1_4_valid;
  assign debug_microOp_cf_loadWaitBit_MPORT_54_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_54_addr = io_writeback_1_4_bits_uop_robIdx_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_54_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_54_en = io_writeback_1_4_valid;
  assign debug_microOp_cf_loadWaitBit_MPORT_55_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_55_addr = io_writeback_1_4_bits_uop_robIdx_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_55_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_55_en = io_writeback_1_4_valid;
  assign debug_microOp_cf_loadWaitBit_MPORT_56_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_56_addr = io_writeback_1_5_bits_uop_robIdx_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_56_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_56_en = io_writeback_1_5_valid;
  assign debug_microOp_cf_loadWaitBit_MPORT_57_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_57_addr = io_writeback_1_5_bits_uop_robIdx_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_57_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_57_en = io_writeback_1_5_valid;
  assign debug_microOp_cf_loadWaitBit_MPORT_58_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_58_addr = io_writeback_1_5_bits_uop_robIdx_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_58_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_58_en = io_writeback_1_5_valid;
  assign debug_microOp_cf_loadWaitBit_MPORT_59_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_59_addr = io_writeback_1_5_bits_uop_robIdx_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_59_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_59_en = io_writeback_1_5_valid;
  assign debug_microOp_cf_loadWaitBit_MPORT_60_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_60_addr = io_writeback_1_5_bits_uop_robIdx_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_60_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_60_en = io_writeback_1_5_valid;
  assign debug_microOp_cf_loadWaitBit_MPORT_61_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_61_addr = io_writeback_1_5_bits_uop_robIdx_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_61_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_61_en = io_writeback_1_5_valid;
  assign debug_microOp_cf_loadWaitBit_MPORT_62_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_62_addr = io_writeback_1_5_bits_uop_robIdx_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_62_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_62_en = io_writeback_1_5_valid;
  assign debug_microOp_cf_loadWaitBit_MPORT_63_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_63_addr = io_writeback_1_5_bits_uop_robIdx_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_63_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_63_en = io_writeback_1_5_valid;
  assign debug_microOp_cf_loadWaitBit_MPORT_64_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_64_addr = io_writeback_1_6_bits_uop_robIdx_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_64_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_64_en = io_writeback_1_6_valid;
  assign debug_microOp_cf_loadWaitBit_MPORT_65_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_65_addr = io_writeback_1_6_bits_uop_robIdx_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_65_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_65_en = io_writeback_1_6_valid;
  assign debug_microOp_cf_loadWaitBit_MPORT_66_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_66_addr = io_writeback_1_6_bits_uop_robIdx_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_66_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_66_en = io_writeback_1_6_valid;
  assign debug_microOp_cf_loadWaitBit_MPORT_67_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_67_addr = io_writeback_1_6_bits_uop_robIdx_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_67_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_67_en = io_writeback_1_6_valid;
  assign debug_microOp_cf_loadWaitBit_MPORT_68_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_68_addr = io_writeback_1_6_bits_uop_robIdx_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_68_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_68_en = io_writeback_1_6_valid;
  assign debug_microOp_cf_loadWaitBit_MPORT_69_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_69_addr = io_writeback_1_6_bits_uop_robIdx_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_69_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_69_en = io_writeback_1_6_valid;
  assign debug_microOp_cf_loadWaitBit_MPORT_70_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_70_addr = io_writeback_1_6_bits_uop_robIdx_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_70_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_70_en = io_writeback_1_6_valid;
  assign debug_microOp_cf_loadWaitBit_MPORT_71_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_71_addr = io_writeback_1_6_bits_uop_robIdx_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_71_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_71_en = io_writeback_1_6_valid;
  assign debug_microOp_cf_loadWaitBit_MPORT_72_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_72_addr = io_writeback_1_7_bits_uop_robIdx_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_72_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_72_en = io_writeback_1_7_valid;
  assign debug_microOp_cf_loadWaitBit_MPORT_73_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_73_addr = io_writeback_1_7_bits_uop_robIdx_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_73_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_73_en = io_writeback_1_7_valid;
  assign debug_microOp_cf_loadWaitBit_MPORT_74_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_74_addr = io_writeback_1_7_bits_uop_robIdx_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_74_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_74_en = io_writeback_1_7_valid;
  assign debug_microOp_cf_loadWaitBit_MPORT_75_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_75_addr = io_writeback_1_7_bits_uop_robIdx_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_75_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_75_en = io_writeback_1_7_valid;
  assign debug_microOp_cf_loadWaitBit_MPORT_76_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_76_addr = io_writeback_1_7_bits_uop_robIdx_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_76_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_76_en = io_writeback_1_7_valid;
  assign debug_microOp_cf_loadWaitBit_MPORT_77_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_77_addr = io_writeback_1_7_bits_uop_robIdx_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_77_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_77_en = io_writeback_1_7_valid;
  assign debug_microOp_cf_loadWaitBit_MPORT_78_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_78_addr = io_writeback_1_7_bits_uop_robIdx_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_78_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_78_en = io_writeback_1_7_valid;
  assign debug_microOp_cf_loadWaitBit_MPORT_79_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_79_addr = io_writeback_1_7_bits_uop_robIdx_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_79_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_79_en = io_writeback_1_7_valid;
  assign debug_microOp_cf_loadWaitBit_MPORT_80_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_80_addr = io_writeback_1_8_bits_uop_robIdx_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_80_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_80_en = io_writeback_1_8_valid;
  assign debug_microOp_cf_loadWaitBit_MPORT_81_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_81_addr = io_writeback_1_8_bits_uop_robIdx_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_81_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_81_en = io_writeback_1_8_valid;
  assign debug_microOp_cf_loadWaitBit_MPORT_82_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_82_addr = io_writeback_1_8_bits_uop_robIdx_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_82_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_82_en = io_writeback_1_8_valid;
  assign debug_microOp_cf_loadWaitBit_MPORT_83_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_83_addr = io_writeback_1_8_bits_uop_robIdx_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_83_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_83_en = io_writeback_1_8_valid;
  assign debug_microOp_cf_loadWaitBit_MPORT_84_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_84_addr = io_writeback_1_8_bits_uop_robIdx_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_84_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_84_en = io_writeback_1_8_valid;
  assign debug_microOp_cf_loadWaitBit_MPORT_85_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_85_addr = io_writeback_1_8_bits_uop_robIdx_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_85_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_85_en = io_writeback_1_8_valid;
  assign debug_microOp_cf_loadWaitBit_MPORT_86_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_86_addr = io_writeback_1_8_bits_uop_robIdx_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_86_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_86_en = io_writeback_1_8_valid;
  assign debug_microOp_cf_loadWaitBit_MPORT_87_data = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_87_addr = io_writeback_1_8_bits_uop_robIdx_value;
  assign debug_microOp_cf_loadWaitBit_MPORT_87_mask = 1'h0;
  assign debug_microOp_cf_loadWaitBit_MPORT_87_en = io_writeback_1_8_valid;
  assign debug_microOp_ctrl_isMove_debug_deqUop_en = 1'h1;
  assign debug_microOp_ctrl_isMove_debug_deqUop_addr = deqPtrGenModule_io_out_0_value;
  assign debug_microOp_ctrl_isMove_debug_deqUop_data =
    debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_debug_deqUop_addr]; // @[Rob.scala 440:26]
  assign debug_microOp_ctrl_isMove_commitDebugUop_0_en = 1'h1;
  assign debug_microOp_ctrl_isMove_commitDebugUop_0_addr = deqPtrGenModule_io_out_0_value;
  assign debug_microOp_ctrl_isMove_commitDebugUop_0_data =
    debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_commitDebugUop_0_addr]; // @[Rob.scala 440:26]
  assign debug_microOp_ctrl_isMove_commitDebugUop_1_en = 1'h1;
  assign debug_microOp_ctrl_isMove_commitDebugUop_1_addr = deqPtrGenModule_io_out_1_value;
  assign debug_microOp_ctrl_isMove_commitDebugUop_1_data =
    debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_commitDebugUop_1_addr]; // @[Rob.scala 440:26]
  assign debug_microOp_ctrl_isMove_MPORT_data = io_enq_req_0_bits_ctrl_isMove;
  assign debug_microOp_ctrl_isMove_MPORT_addr = enqPtrGenModule_io_out_0_value;
  assign debug_microOp_ctrl_isMove_MPORT_mask = 1'h1;
  assign debug_microOp_ctrl_isMove_MPORT_en = io_enq_req_0_valid & io_enq_canAccept;
  assign debug_microOp_ctrl_isMove_MPORT_1_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_1_addr = enqPtrGenModule_io_out_0_value;
  assign debug_microOp_ctrl_isMove_MPORT_1_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_1_en = io_enq_req_0_valid & io_enq_canAccept;
  assign debug_microOp_ctrl_isMove_MPORT_2_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_2_addr = enqPtrGenModule_io_out_0_value;
  assign debug_microOp_ctrl_isMove_MPORT_2_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_2_en = io_enq_req_0_valid & io_enq_canAccept;
  assign debug_microOp_ctrl_isMove_MPORT_3_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_3_addr = enqPtrGenModule_io_out_0_value;
  assign debug_microOp_ctrl_isMove_MPORT_3_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_3_en = io_enq_req_0_valid & io_enq_canAccept;
  assign debug_microOp_ctrl_isMove_MPORT_4_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_4_addr = enqPtrGenModule_io_out_0_value;
  assign debug_microOp_ctrl_isMove_MPORT_4_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_4_en = io_enq_req_0_valid & io_enq_canAccept;
  assign debug_microOp_ctrl_isMove_MPORT_5_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_5_addr = enqPtrGenModule_io_out_0_value;
  assign debug_microOp_ctrl_isMove_MPORT_5_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_5_en = io_enq_req_0_valid & io_enq_canAccept;
  assign debug_microOp_ctrl_isMove_MPORT_6_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_6_addr = enqPtrGenModule_io_out_0_value;
  assign debug_microOp_ctrl_isMove_MPORT_6_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_6_en = io_enq_req_0_valid & io_enq_canAccept;
  assign debug_microOp_ctrl_isMove_MPORT_7_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_7_addr = enqPtrGenModule_io_out_0_value;
  assign debug_microOp_ctrl_isMove_MPORT_7_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_7_en = io_enq_req_0_valid & io_enq_canAccept;
  assign debug_microOp_ctrl_isMove_MPORT_8_data = io_enq_req_1_bits_ctrl_isMove;
  assign debug_microOp_ctrl_isMove_MPORT_8_addr = io_enq_needAlloc_0 ? enqPtrVec_1_value : enqPtrVec_0_value;
  assign debug_microOp_ctrl_isMove_MPORT_8_mask = 1'h1;
  assign debug_microOp_ctrl_isMove_MPORT_8_en = io_enq_req_1_valid & io_enq_canAccept;
  assign debug_microOp_ctrl_isMove_MPORT_9_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_9_addr = io_enq_needAlloc_0 ? enqPtrVec_1_value : enqPtrVec_0_value;
  assign debug_microOp_ctrl_isMove_MPORT_9_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_9_en = io_enq_req_1_valid & io_enq_canAccept;
  assign debug_microOp_ctrl_isMove_MPORT_10_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_10_addr = io_enq_needAlloc_0 ? enqPtrVec_1_value : enqPtrVec_0_value;
  assign debug_microOp_ctrl_isMove_MPORT_10_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_10_en = io_enq_req_1_valid & io_enq_canAccept;
  assign debug_microOp_ctrl_isMove_MPORT_11_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_11_addr = io_enq_needAlloc_0 ? enqPtrVec_1_value : enqPtrVec_0_value;
  assign debug_microOp_ctrl_isMove_MPORT_11_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_11_en = io_enq_req_1_valid & io_enq_canAccept;
  assign debug_microOp_ctrl_isMove_MPORT_12_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_12_addr = io_enq_needAlloc_0 ? enqPtrVec_1_value : enqPtrVec_0_value;
  assign debug_microOp_ctrl_isMove_MPORT_12_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_12_en = io_enq_req_1_valid & io_enq_canAccept;
  assign debug_microOp_ctrl_isMove_MPORT_13_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_13_addr = io_enq_needAlloc_0 ? enqPtrVec_1_value : enqPtrVec_0_value;
  assign debug_microOp_ctrl_isMove_MPORT_13_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_13_en = io_enq_req_1_valid & io_enq_canAccept;
  assign debug_microOp_ctrl_isMove_MPORT_14_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_14_addr = io_enq_needAlloc_0 ? enqPtrVec_1_value : enqPtrVec_0_value;
  assign debug_microOp_ctrl_isMove_MPORT_14_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_14_en = io_enq_req_1_valid & io_enq_canAccept;
  assign debug_microOp_ctrl_isMove_MPORT_15_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_15_addr = io_enq_needAlloc_0 ? enqPtrVec_1_value : enqPtrVec_0_value;
  assign debug_microOp_ctrl_isMove_MPORT_15_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_15_en = io_enq_req_1_valid & io_enq_canAccept;
  assign debug_microOp_ctrl_isMove_MPORT_16_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_16_addr = io_writeback_1_0_bits_uop_robIdx_value;
  assign debug_microOp_ctrl_isMove_MPORT_16_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_16_en = io_writeback_1_0_valid;
  assign debug_microOp_ctrl_isMove_MPORT_17_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_17_addr = io_writeback_1_0_bits_uop_robIdx_value;
  assign debug_microOp_ctrl_isMove_MPORT_17_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_17_en = io_writeback_1_0_valid;
  assign debug_microOp_ctrl_isMove_MPORT_18_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_18_addr = io_writeback_1_0_bits_uop_robIdx_value;
  assign debug_microOp_ctrl_isMove_MPORT_18_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_18_en = io_writeback_1_0_valid;
  assign debug_microOp_ctrl_isMove_MPORT_19_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_19_addr = io_writeback_1_0_bits_uop_robIdx_value;
  assign debug_microOp_ctrl_isMove_MPORT_19_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_19_en = io_writeback_1_0_valid;
  assign debug_microOp_ctrl_isMove_MPORT_20_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_20_addr = io_writeback_1_0_bits_uop_robIdx_value;
  assign debug_microOp_ctrl_isMove_MPORT_20_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_20_en = io_writeback_1_0_valid;
  assign debug_microOp_ctrl_isMove_MPORT_21_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_21_addr = io_writeback_1_0_bits_uop_robIdx_value;
  assign debug_microOp_ctrl_isMove_MPORT_21_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_21_en = io_writeback_1_0_valid;
  assign debug_microOp_ctrl_isMove_MPORT_22_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_22_addr = io_writeback_1_0_bits_uop_robIdx_value;
  assign debug_microOp_ctrl_isMove_MPORT_22_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_22_en = io_writeback_1_0_valid;
  assign debug_microOp_ctrl_isMove_MPORT_23_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_23_addr = io_writeback_1_0_bits_uop_robIdx_value;
  assign debug_microOp_ctrl_isMove_MPORT_23_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_23_en = io_writeback_1_0_valid;
  assign debug_microOp_ctrl_isMove_MPORT_24_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_24_addr = io_writeback_1_1_bits_uop_robIdx_value;
  assign debug_microOp_ctrl_isMove_MPORT_24_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_24_en = io_writeback_1_1_valid;
  assign debug_microOp_ctrl_isMove_MPORT_25_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_25_addr = io_writeback_1_1_bits_uop_robIdx_value;
  assign debug_microOp_ctrl_isMove_MPORT_25_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_25_en = io_writeback_1_1_valid;
  assign debug_microOp_ctrl_isMove_MPORT_26_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_26_addr = io_writeback_1_1_bits_uop_robIdx_value;
  assign debug_microOp_ctrl_isMove_MPORT_26_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_26_en = io_writeback_1_1_valid;
  assign debug_microOp_ctrl_isMove_MPORT_27_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_27_addr = io_writeback_1_1_bits_uop_robIdx_value;
  assign debug_microOp_ctrl_isMove_MPORT_27_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_27_en = io_writeback_1_1_valid;
  assign debug_microOp_ctrl_isMove_MPORT_28_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_28_addr = io_writeback_1_1_bits_uop_robIdx_value;
  assign debug_microOp_ctrl_isMove_MPORT_28_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_28_en = io_writeback_1_1_valid;
  assign debug_microOp_ctrl_isMove_MPORT_29_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_29_addr = io_writeback_1_1_bits_uop_robIdx_value;
  assign debug_microOp_ctrl_isMove_MPORT_29_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_29_en = io_writeback_1_1_valid;
  assign debug_microOp_ctrl_isMove_MPORT_30_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_30_addr = io_writeback_1_1_bits_uop_robIdx_value;
  assign debug_microOp_ctrl_isMove_MPORT_30_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_30_en = io_writeback_1_1_valid;
  assign debug_microOp_ctrl_isMove_MPORT_31_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_31_addr = io_writeback_1_1_bits_uop_robIdx_value;
  assign debug_microOp_ctrl_isMove_MPORT_31_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_31_en = io_writeback_1_1_valid;
  assign debug_microOp_ctrl_isMove_MPORT_32_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_32_addr = io_writeback_1_2_bits_uop_robIdx_value;
  assign debug_microOp_ctrl_isMove_MPORT_32_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_32_en = io_writeback_1_2_valid;
  assign debug_microOp_ctrl_isMove_MPORT_33_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_33_addr = io_writeback_1_2_bits_uop_robIdx_value;
  assign debug_microOp_ctrl_isMove_MPORT_33_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_33_en = io_writeback_1_2_valid;
  assign debug_microOp_ctrl_isMove_MPORT_34_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_34_addr = io_writeback_1_2_bits_uop_robIdx_value;
  assign debug_microOp_ctrl_isMove_MPORT_34_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_34_en = io_writeback_1_2_valid;
  assign debug_microOp_ctrl_isMove_MPORT_35_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_35_addr = io_writeback_1_2_bits_uop_robIdx_value;
  assign debug_microOp_ctrl_isMove_MPORT_35_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_35_en = io_writeback_1_2_valid;
  assign debug_microOp_ctrl_isMove_MPORT_36_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_36_addr = io_writeback_1_2_bits_uop_robIdx_value;
  assign debug_microOp_ctrl_isMove_MPORT_36_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_36_en = io_writeback_1_2_valid;
  assign debug_microOp_ctrl_isMove_MPORT_37_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_37_addr = io_writeback_1_2_bits_uop_robIdx_value;
  assign debug_microOp_ctrl_isMove_MPORT_37_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_37_en = io_writeback_1_2_valid;
  assign debug_microOp_ctrl_isMove_MPORT_38_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_38_addr = io_writeback_1_2_bits_uop_robIdx_value;
  assign debug_microOp_ctrl_isMove_MPORT_38_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_38_en = io_writeback_1_2_valid;
  assign debug_microOp_ctrl_isMove_MPORT_39_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_39_addr = io_writeback_1_2_bits_uop_robIdx_value;
  assign debug_microOp_ctrl_isMove_MPORT_39_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_39_en = io_writeback_1_2_valid;
  assign debug_microOp_ctrl_isMove_MPORT_40_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_40_addr = io_writeback_1_3_bits_uop_robIdx_value;
  assign debug_microOp_ctrl_isMove_MPORT_40_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_40_en = io_writeback_1_3_valid;
  assign debug_microOp_ctrl_isMove_MPORT_41_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_41_addr = io_writeback_1_3_bits_uop_robIdx_value;
  assign debug_microOp_ctrl_isMove_MPORT_41_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_41_en = io_writeback_1_3_valid;
  assign debug_microOp_ctrl_isMove_MPORT_42_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_42_addr = io_writeback_1_3_bits_uop_robIdx_value;
  assign debug_microOp_ctrl_isMove_MPORT_42_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_42_en = io_writeback_1_3_valid;
  assign debug_microOp_ctrl_isMove_MPORT_43_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_43_addr = io_writeback_1_3_bits_uop_robIdx_value;
  assign debug_microOp_ctrl_isMove_MPORT_43_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_43_en = io_writeback_1_3_valid;
  assign debug_microOp_ctrl_isMove_MPORT_44_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_44_addr = io_writeback_1_3_bits_uop_robIdx_value;
  assign debug_microOp_ctrl_isMove_MPORT_44_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_44_en = io_writeback_1_3_valid;
  assign debug_microOp_ctrl_isMove_MPORT_45_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_45_addr = io_writeback_1_3_bits_uop_robIdx_value;
  assign debug_microOp_ctrl_isMove_MPORT_45_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_45_en = io_writeback_1_3_valid;
  assign debug_microOp_ctrl_isMove_MPORT_46_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_46_addr = io_writeback_1_3_bits_uop_robIdx_value;
  assign debug_microOp_ctrl_isMove_MPORT_46_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_46_en = io_writeback_1_3_valid;
  assign debug_microOp_ctrl_isMove_MPORT_47_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_47_addr = io_writeback_1_3_bits_uop_robIdx_value;
  assign debug_microOp_ctrl_isMove_MPORT_47_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_47_en = io_writeback_1_3_valid;
  assign debug_microOp_ctrl_isMove_MPORT_48_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_48_addr = io_writeback_1_4_bits_uop_robIdx_value;
  assign debug_microOp_ctrl_isMove_MPORT_48_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_48_en = io_writeback_1_4_valid;
  assign debug_microOp_ctrl_isMove_MPORT_49_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_49_addr = io_writeback_1_4_bits_uop_robIdx_value;
  assign debug_microOp_ctrl_isMove_MPORT_49_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_49_en = io_writeback_1_4_valid;
  assign debug_microOp_ctrl_isMove_MPORT_50_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_50_addr = io_writeback_1_4_bits_uop_robIdx_value;
  assign debug_microOp_ctrl_isMove_MPORT_50_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_50_en = io_writeback_1_4_valid;
  assign debug_microOp_ctrl_isMove_MPORT_51_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_51_addr = io_writeback_1_4_bits_uop_robIdx_value;
  assign debug_microOp_ctrl_isMove_MPORT_51_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_51_en = io_writeback_1_4_valid;
  assign debug_microOp_ctrl_isMove_MPORT_52_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_52_addr = io_writeback_1_4_bits_uop_robIdx_value;
  assign debug_microOp_ctrl_isMove_MPORT_52_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_52_en = io_writeback_1_4_valid;
  assign debug_microOp_ctrl_isMove_MPORT_53_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_53_addr = io_writeback_1_4_bits_uop_robIdx_value;
  assign debug_microOp_ctrl_isMove_MPORT_53_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_53_en = io_writeback_1_4_valid;
  assign debug_microOp_ctrl_isMove_MPORT_54_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_54_addr = io_writeback_1_4_bits_uop_robIdx_value;
  assign debug_microOp_ctrl_isMove_MPORT_54_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_54_en = io_writeback_1_4_valid;
  assign debug_microOp_ctrl_isMove_MPORT_55_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_55_addr = io_writeback_1_4_bits_uop_robIdx_value;
  assign debug_microOp_ctrl_isMove_MPORT_55_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_55_en = io_writeback_1_4_valid;
  assign debug_microOp_ctrl_isMove_MPORT_56_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_56_addr = io_writeback_1_5_bits_uop_robIdx_value;
  assign debug_microOp_ctrl_isMove_MPORT_56_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_56_en = io_writeback_1_5_valid;
  assign debug_microOp_ctrl_isMove_MPORT_57_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_57_addr = io_writeback_1_5_bits_uop_robIdx_value;
  assign debug_microOp_ctrl_isMove_MPORT_57_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_57_en = io_writeback_1_5_valid;
  assign debug_microOp_ctrl_isMove_MPORT_58_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_58_addr = io_writeback_1_5_bits_uop_robIdx_value;
  assign debug_microOp_ctrl_isMove_MPORT_58_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_58_en = io_writeback_1_5_valid;
  assign debug_microOp_ctrl_isMove_MPORT_59_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_59_addr = io_writeback_1_5_bits_uop_robIdx_value;
  assign debug_microOp_ctrl_isMove_MPORT_59_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_59_en = io_writeback_1_5_valid;
  assign debug_microOp_ctrl_isMove_MPORT_60_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_60_addr = io_writeback_1_5_bits_uop_robIdx_value;
  assign debug_microOp_ctrl_isMove_MPORT_60_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_60_en = io_writeback_1_5_valid;
  assign debug_microOp_ctrl_isMove_MPORT_61_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_61_addr = io_writeback_1_5_bits_uop_robIdx_value;
  assign debug_microOp_ctrl_isMove_MPORT_61_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_61_en = io_writeback_1_5_valid;
  assign debug_microOp_ctrl_isMove_MPORT_62_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_62_addr = io_writeback_1_5_bits_uop_robIdx_value;
  assign debug_microOp_ctrl_isMove_MPORT_62_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_62_en = io_writeback_1_5_valid;
  assign debug_microOp_ctrl_isMove_MPORT_63_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_63_addr = io_writeback_1_5_bits_uop_robIdx_value;
  assign debug_microOp_ctrl_isMove_MPORT_63_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_63_en = io_writeback_1_5_valid;
  assign debug_microOp_ctrl_isMove_MPORT_64_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_64_addr = io_writeback_1_6_bits_uop_robIdx_value;
  assign debug_microOp_ctrl_isMove_MPORT_64_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_64_en = io_writeback_1_6_valid;
  assign debug_microOp_ctrl_isMove_MPORT_65_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_65_addr = io_writeback_1_6_bits_uop_robIdx_value;
  assign debug_microOp_ctrl_isMove_MPORT_65_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_65_en = io_writeback_1_6_valid;
  assign debug_microOp_ctrl_isMove_MPORT_66_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_66_addr = io_writeback_1_6_bits_uop_robIdx_value;
  assign debug_microOp_ctrl_isMove_MPORT_66_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_66_en = io_writeback_1_6_valid;
  assign debug_microOp_ctrl_isMove_MPORT_67_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_67_addr = io_writeback_1_6_bits_uop_robIdx_value;
  assign debug_microOp_ctrl_isMove_MPORT_67_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_67_en = io_writeback_1_6_valid;
  assign debug_microOp_ctrl_isMove_MPORT_68_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_68_addr = io_writeback_1_6_bits_uop_robIdx_value;
  assign debug_microOp_ctrl_isMove_MPORT_68_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_68_en = io_writeback_1_6_valid;
  assign debug_microOp_ctrl_isMove_MPORT_69_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_69_addr = io_writeback_1_6_bits_uop_robIdx_value;
  assign debug_microOp_ctrl_isMove_MPORT_69_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_69_en = io_writeback_1_6_valid;
  assign debug_microOp_ctrl_isMove_MPORT_70_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_70_addr = io_writeback_1_6_bits_uop_robIdx_value;
  assign debug_microOp_ctrl_isMove_MPORT_70_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_70_en = io_writeback_1_6_valid;
  assign debug_microOp_ctrl_isMove_MPORT_71_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_71_addr = io_writeback_1_6_bits_uop_robIdx_value;
  assign debug_microOp_ctrl_isMove_MPORT_71_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_71_en = io_writeback_1_6_valid;
  assign debug_microOp_ctrl_isMove_MPORT_72_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_72_addr = io_writeback_1_7_bits_uop_robIdx_value;
  assign debug_microOp_ctrl_isMove_MPORT_72_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_72_en = io_writeback_1_7_valid;
  assign debug_microOp_ctrl_isMove_MPORT_73_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_73_addr = io_writeback_1_7_bits_uop_robIdx_value;
  assign debug_microOp_ctrl_isMove_MPORT_73_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_73_en = io_writeback_1_7_valid;
  assign debug_microOp_ctrl_isMove_MPORT_74_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_74_addr = io_writeback_1_7_bits_uop_robIdx_value;
  assign debug_microOp_ctrl_isMove_MPORT_74_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_74_en = io_writeback_1_7_valid;
  assign debug_microOp_ctrl_isMove_MPORT_75_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_75_addr = io_writeback_1_7_bits_uop_robIdx_value;
  assign debug_microOp_ctrl_isMove_MPORT_75_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_75_en = io_writeback_1_7_valid;
  assign debug_microOp_ctrl_isMove_MPORT_76_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_76_addr = io_writeback_1_7_bits_uop_robIdx_value;
  assign debug_microOp_ctrl_isMove_MPORT_76_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_76_en = io_writeback_1_7_valid;
  assign debug_microOp_ctrl_isMove_MPORT_77_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_77_addr = io_writeback_1_7_bits_uop_robIdx_value;
  assign debug_microOp_ctrl_isMove_MPORT_77_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_77_en = io_writeback_1_7_valid;
  assign debug_microOp_ctrl_isMove_MPORT_78_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_78_addr = io_writeback_1_7_bits_uop_robIdx_value;
  assign debug_microOp_ctrl_isMove_MPORT_78_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_78_en = io_writeback_1_7_valid;
  assign debug_microOp_ctrl_isMove_MPORT_79_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_79_addr = io_writeback_1_7_bits_uop_robIdx_value;
  assign debug_microOp_ctrl_isMove_MPORT_79_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_79_en = io_writeback_1_7_valid;
  assign debug_microOp_ctrl_isMove_MPORT_80_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_80_addr = io_writeback_1_8_bits_uop_robIdx_value;
  assign debug_microOp_ctrl_isMove_MPORT_80_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_80_en = io_writeback_1_8_valid;
  assign debug_microOp_ctrl_isMove_MPORT_81_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_81_addr = io_writeback_1_8_bits_uop_robIdx_value;
  assign debug_microOp_ctrl_isMove_MPORT_81_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_81_en = io_writeback_1_8_valid;
  assign debug_microOp_ctrl_isMove_MPORT_82_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_82_addr = io_writeback_1_8_bits_uop_robIdx_value;
  assign debug_microOp_ctrl_isMove_MPORT_82_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_82_en = io_writeback_1_8_valid;
  assign debug_microOp_ctrl_isMove_MPORT_83_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_83_addr = io_writeback_1_8_bits_uop_robIdx_value;
  assign debug_microOp_ctrl_isMove_MPORT_83_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_83_en = io_writeback_1_8_valid;
  assign debug_microOp_ctrl_isMove_MPORT_84_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_84_addr = io_writeback_1_8_bits_uop_robIdx_value;
  assign debug_microOp_ctrl_isMove_MPORT_84_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_84_en = io_writeback_1_8_valid;
  assign debug_microOp_ctrl_isMove_MPORT_85_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_85_addr = io_writeback_1_8_bits_uop_robIdx_value;
  assign debug_microOp_ctrl_isMove_MPORT_85_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_85_en = io_writeback_1_8_valid;
  assign debug_microOp_ctrl_isMove_MPORT_86_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_86_addr = io_writeback_1_8_bits_uop_robIdx_value;
  assign debug_microOp_ctrl_isMove_MPORT_86_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_86_en = io_writeback_1_8_valid;
  assign debug_microOp_ctrl_isMove_MPORT_87_data = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_87_addr = io_writeback_1_8_bits_uop_robIdx_value;
  assign debug_microOp_ctrl_isMove_MPORT_87_mask = 1'h0;
  assign debug_microOp_ctrl_isMove_MPORT_87_en = io_writeback_1_8_valid;
  assign dt_eliminatedMove_eliminatedMove_en = 1'h1;
  assign dt_eliminatedMove_eliminatedMove_addr = deqPtrGenModule_io_out_0_value;
  assign dt_eliminatedMove_eliminatedMove_data = dt_eliminatedMove[dt_eliminatedMove_eliminatedMove_addr]; // @[Rob.scala 1212:32]
  assign dt_eliminatedMove_eliminatedMove_1_en = 1'h1;
  assign dt_eliminatedMove_eliminatedMove_1_addr = deqPtrGenModule_io_out_1_value;
  assign dt_eliminatedMove_eliminatedMove_1_data = dt_eliminatedMove[dt_eliminatedMove_eliminatedMove_1_addr]; // @[Rob.scala 1212:32]
  assign dt_eliminatedMove_MPORT_305_data = io_enq_req_0_bits_eliminatedMove;
  assign dt_eliminatedMove_MPORT_305_addr = enqPtrGenModule_io_out_0_value;
  assign dt_eliminatedMove_MPORT_305_mask = 1'h1;
  assign dt_eliminatedMove_MPORT_305_en = io_enq_req_0_valid & io_enq_canAccept;
  assign dt_eliminatedMove_MPORT_307_data = io_enq_req_1_bits_eliminatedMove;
  assign dt_eliminatedMove_MPORT_307_addr = io_enq_needAlloc_0 ? enqPtrVec_1_value : enqPtrVec_0_value;
  assign dt_eliminatedMove_MPORT_307_mask = 1'h1;
  assign dt_eliminatedMove_MPORT_307_en = io_enq_req_1_valid & io_enq_canAccept;
  assign dt_isRVC_isRVC_en = 1'h1;
  assign dt_isRVC_isRVC_addr = deqPtrGenModule_io_out_0_value;
  assign dt_isRVC_isRVC_data = dt_isRVC[dt_isRVC_isRVC_addr]; // @[Rob.scala 1213:23]
  assign dt_isRVC_isRVC_1_en = 1'h1;
  assign dt_isRVC_isRVC_1_addr = deqPtrGenModule_io_out_1_value;
  assign dt_isRVC_isRVC_1_data = dt_isRVC[dt_isRVC_isRVC_1_addr]; // @[Rob.scala 1213:23]
  assign dt_isRVC_MPORT_306_data = io_enq_req_0_bits_cf_pd_isRVC;
  assign dt_isRVC_MPORT_306_addr = enqPtrGenModule_io_out_0_value;
  assign dt_isRVC_MPORT_306_mask = 1'h1;
  assign dt_isRVC_MPORT_306_en = io_enq_req_0_valid & io_enq_canAccept;
  assign dt_isRVC_MPORT_308_data = io_enq_req_1_bits_cf_pd_isRVC;
  assign dt_isRVC_MPORT_308_addr = io_enq_needAlloc_0 ? enqPtrVec_1_value : enqPtrVec_0_value;
  assign dt_isRVC_MPORT_308_mask = 1'h1;
  assign dt_isRVC_MPORT_308_en = io_enq_req_1_valid & io_enq_canAccept;
  assign dt_isXSTrap_trapVec_MPORT_en = 1'h1;
  assign dt_isXSTrap_trapVec_MPORT_addr = deqPtrGenModule_io_out_0_value;
  assign dt_isXSTrap_trapVec_MPORT_data = dt_isXSTrap[dt_isXSTrap_trapVec_MPORT_addr]; // @[Rob.scala 1290:26]
  assign dt_isXSTrap_trapVec_MPORT_1_en = 1'h1;
  assign dt_isXSTrap_trapVec_MPORT_1_addr = deqPtrGenModule_io_out_1_value;
  assign dt_isXSTrap_trapVec_MPORT_1_data = dt_isXSTrap[dt_isXSTrap_trapVec_MPORT_1_addr]; // @[Rob.scala 1290:26]
  assign dt_isXSTrap_MPORT_309_data = io_enq_req_0_bits_ctrl_isXSTrap;
  assign dt_isXSTrap_MPORT_309_addr = enqPtrGenModule_io_out_0_value;
  assign dt_isXSTrap_MPORT_309_mask = 1'h1;
  assign dt_isXSTrap_MPORT_309_en = io_enq_req_0_valid & io_enq_canAccept;
  assign dt_isXSTrap_MPORT_310_data = io_enq_req_1_bits_ctrl_isXSTrap;
  assign dt_isXSTrap_MPORT_310_addr = io_enq_needAlloc_0 ? enqPtrVec_1_value : enqPtrVec_0_value;
  assign dt_isXSTrap_MPORT_310_mask = 1'h1;
  assign dt_isXSTrap_MPORT_310_en = io_enq_req_1_valid & io_enq_canAccept;
  assign io_enq_canAccept = allowEnqueue & ~hasBlockBackward; // @[Rob.scala 517:36]
  assign io_enq_isEmpty = io_enq_isEmpty_REG; // @[Rob.scala 566:20]
  assign io_flushOut_valid = ~state & commit_v_0 & (intrEnable | exceptionEnable | isFlushPipe) & ~lastCycleFlush; // @[Rob.scala 636:116]
  assign io_flushOut_bits_robIdx_flag = deqPtrGenModule_io_out_0_flag; // @[Rob.scala 448:23 783:13]
  assign io_flushOut_bits_robIdx_value = deqPtrGenModule_io_out_0_value; // @[Rob.scala 448:23 783:13]
  assign io_flushOut_bits_ftqIdx_flag = dispatchData_io_rdata_0_ftqIdx_flag; // @[Rob.scala 639:27]
  assign io_flushOut_bits_ftqIdx_value = dispatchData_io_rdata_0_ftqIdx_value; // @[Rob.scala 639:27]
  assign io_flushOut_bits_ftqOffset = dispatchData_io_rdata_0_ftqOffset; // @[Rob.scala 640:30]
  assign io_flushOut_bits_level = deqHasReplayInst | intrEnable | exceptionEnable; // @[Rob.scala 641:64]
  assign io_exception_valid = io_exception_valid_REG; // @[Rob.scala 649:22]
  assign io_exception_bits_uop_cf_exceptionVec_0 = r_0; // @[Rob.scala 652:41]
  assign io_exception_bits_uop_cf_exceptionVec_1 = r_1; // @[Rob.scala 652:41]
  assign io_exception_bits_uop_cf_exceptionVec_2 = r_2; // @[Rob.scala 652:41]
  assign io_exception_bits_uop_cf_exceptionVec_3 = r_3; // @[Rob.scala 652:41]
  assign io_exception_bits_uop_cf_exceptionVec_4 = r_4; // @[Rob.scala 652:41]
  assign io_exception_bits_uop_cf_exceptionVec_5 = r_5; // @[Rob.scala 652:41]
  assign io_exception_bits_uop_cf_exceptionVec_6 = r_6; // @[Rob.scala 652:41]
  assign io_exception_bits_uop_cf_exceptionVec_7 = r_7; // @[Rob.scala 652:41]
  assign io_exception_bits_uop_cf_exceptionVec_8 = r_8; // @[Rob.scala 652:41]
  assign io_exception_bits_uop_cf_exceptionVec_9 = r_9; // @[Rob.scala 652:41]
  assign io_exception_bits_uop_cf_exceptionVec_11 = r_11; // @[Rob.scala 652:41]
  assign io_exception_bits_uop_cf_exceptionVec_12 = r_12; // @[Rob.scala 652:41]
  assign io_exception_bits_uop_cf_exceptionVec_13 = r_13; // @[Rob.scala 652:41]
  assign io_exception_bits_uop_cf_exceptionVec_15 = r_15; // @[Rob.scala 652:41]
  assign io_exception_bits_uop_cf_trigger_frontendHit_0 = io_exception_bits_uop_cf_trigger_rfrontendHit_0; // @[Rob.scala 656:36]
  assign io_exception_bits_uop_cf_trigger_frontendHit_1 = io_exception_bits_uop_cf_trigger_rfrontendHit_1; // @[Rob.scala 656:36]
  assign io_exception_bits_uop_cf_trigger_frontendHit_2 = io_exception_bits_uop_cf_trigger_rfrontendHit_2; // @[Rob.scala 656:36]
  assign io_exception_bits_uop_cf_trigger_frontendHit_3 = io_exception_bits_uop_cf_trigger_rfrontendHit_3; // @[Rob.scala 656:36]
  assign io_exception_bits_uop_cf_trigger_backendHit_0 = io_exception_bits_uop_cf_trigger_rbackendHit_0; // @[Rob.scala 656:36]
  assign io_exception_bits_uop_cf_trigger_backendHit_1 = io_exception_bits_uop_cf_trigger_rbackendHit_1; // @[Rob.scala 656:36]
  assign io_exception_bits_uop_cf_trigger_backendHit_2 = io_exception_bits_uop_cf_trigger_rbackendHit_2; // @[Rob.scala 656:36]
  assign io_exception_bits_uop_cf_trigger_backendHit_3 = io_exception_bits_uop_cf_trigger_rbackendHit_3; // @[Rob.scala 656:36]
  assign io_exception_bits_uop_cf_trigger_backendHit_4 = io_exception_bits_uop_cf_trigger_rbackendHit_4; // @[Rob.scala 656:36]
  assign io_exception_bits_uop_cf_trigger_backendHit_5 = io_exception_bits_uop_cf_trigger_rbackendHit_5; // @[Rob.scala 656:36]
  assign io_exception_bits_uop_cf_crossPageIPFFix = io_exception_bits_uop_cf_crossPageIPFFix_r; // @[Rob.scala 654:44]
  assign io_exception_bits_uop_ctrl_commitType = io_exception_bits_uop_ctrl_commitType_r; // @[Rob.scala 651:41]
  assign io_exception_bits_uop_ctrl_singleStep = io_exception_bits_uop_ctrl_singleStep_r; // @[Rob.scala 653:41]
  assign io_exception_bits_isInterrupt = io_exception_bits_isInterrupt_r; // @[Rob.scala 655:33]
  assign io_commits_isCommit = _io_flushOut_valid_T & ~blockCommit; // @[Rob.scala 701:43]
  assign io_commits_commitValid_0 = commit_v_0 & commit_w0 & ~isBlocked; // @[Rob.scala 714:61]
  assign io_commits_commitValid_1 = commit_v_1 & commit_w1 & ~isBlocked_1; // @[Rob.scala 714:61]
  assign io_commits_isWalk = state; // @[Rob.scala 700:30]
  assign io_commits_walkValid_0 = 6'h0 < walkCounter; // @[Rob.scala 669:61]
  assign io_commits_walkValid_1 = 6'h1 < walkCounter; // @[Rob.scala 669:61]
  assign io_commits_info_0_ldest = dispatchData_io_rdata_0_ldest; // @[Rob.scala 715:25]
  assign io_commits_info_0_rfWen = dispatchData_io_rdata_0_rfWen; // @[Rob.scala 715:25]
  assign io_commits_info_0_fpWen = dispatchData_io_rdata_0_fpWen; // @[Rob.scala 715:25]
  assign io_commits_info_0_wflags = dispatchData_io_rdata_0_wflags; // @[Rob.scala 715:25]
  assign io_commits_info_0_commitType = dispatchData_io_rdata_0_commitType; // @[Rob.scala 715:25]
  assign io_commits_info_0_pdest = dispatchData_io_rdata_0_pdest; // @[Rob.scala 715:25]
  assign io_commits_info_0_old_pdest = dispatchData_io_rdata_0_old_pdest; // @[Rob.scala 715:25]
  assign io_commits_info_0_ftqIdx_flag = dispatchData_io_rdata_0_ftqIdx_flag; // @[Rob.scala 715:25]
  assign io_commits_info_0_ftqIdx_value = dispatchData_io_rdata_0_ftqIdx_value; // @[Rob.scala 715:25]
  assign io_commits_info_0_ftqOffset = dispatchData_io_rdata_0_ftqOffset; // @[Rob.scala 715:25]
  assign io_commits_info_0_isMove = dispatchData_io_rdata_0_isMove; // @[Rob.scala 715:25]
  assign io_commits_info_1_ldest = dispatchData_io_rdata_1_ldest; // @[Rob.scala 715:25]
  assign io_commits_info_1_rfWen = dispatchData_io_rdata_1_rfWen; // @[Rob.scala 715:25]
  assign io_commits_info_1_fpWen = dispatchData_io_rdata_1_fpWen; // @[Rob.scala 715:25]
  assign io_commits_info_1_wflags = dispatchData_io_rdata_1_wflags; // @[Rob.scala 715:25]
  assign io_commits_info_1_commitType = dispatchData_io_rdata_1_commitType; // @[Rob.scala 715:25]
  assign io_commits_info_1_pdest = dispatchData_io_rdata_1_pdest; // @[Rob.scala 715:25]
  assign io_commits_info_1_old_pdest = dispatchData_io_rdata_1_old_pdest; // @[Rob.scala 715:25]
  assign io_commits_info_1_ftqIdx_flag = dispatchData_io_rdata_1_ftqIdx_flag; // @[Rob.scala 715:25]
  assign io_commits_info_1_ftqIdx_value = dispatchData_io_rdata_1_ftqIdx_value; // @[Rob.scala 715:25]
  assign io_commits_info_1_ftqOffset = dispatchData_io_rdata_1_ftqOffset; // @[Rob.scala 715:25]
  assign io_commits_info_1_isMove = dispatchData_io_rdata_1_isMove; // @[Rob.scala 715:25]
  assign io_lsq_scommit = io_lsq_scommit_REG; // @[Rob.scala 753:18]
  assign io_lsq_pendingld = io_lsq_pendingld_REG; // @[Rob.scala 755:20]
  assign io_lsq_pendingst = io_lsq_pendingst_REG; // @[Rob.scala 756:20]
  assign io_lsq_commit = io_lsq_commit_REG; // @[Rob.scala 757:17]
  assign io_csr_fflags_valid = io_csr_fflags_REG_valid; // @[Rob.scala 746:17]
  assign io_csr_fflags_bits = io_csr_fflags_REG_bits; // @[Rob.scala 746:17]
  assign io_csr_dirty_fs = io_csr_dirty_fs_REG; // @[Rob.scala 747:19]
  assign io_csr_perfinfo_retiredInstr = retireCounter_REG ? trueCommitCnt : 3'h0; // @[Rob.scala 1021:26]
  assign io_cpu_halt = hasWFI; // @[Rob.scala 503:15]
  assign io_perf_0_value = {{5'd0}, io_perf_0_value_REG_1}; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_1_value = {{5'd0}, io_perf_1_value_REG_1}; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_2_value = {{5'd0}, io_perf_2_value_REG_1}; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_3_value = {{5'd0}, io_perf_3_value_REG_1}; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_4_value = {{4'd0}, io_perf_4_value_REG_1}; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_5_value = {{3'd0}, io_perf_5_value_REG_1}; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_6_value = {{4'd0}, io_perf_6_value_REG_1}; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_7_value = {{4'd0}, io_perf_7_value_REG_1}; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_8_value = {{4'd0}, io_perf_8_value_REG_1}; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_9_value = {{4'd0}, io_perf_9_value_REG_1}; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_10_value = {{4'd0}, io_perf_10_value_REG_1}; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_11_value = {{4'd0}, io_perf_11_value_REG_1}; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_12_value = {{4'd0}, io_perf_12_value_REG_1}; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_13_value = {{5'd0}, io_perf_13_value_REG_1}; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_14_value = {{5'd0}, io_perf_14_value_REG_1}; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_15_value = {{5'd0}, io_perf_15_value_REG_1}; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_16_value = {{5'd0}, io_perf_16_value_REG_1}; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_17_value = {{5'd0}, io_perf_17_value_REG_1}; // @[PerfCounterUtils.scala 188:17]
  assign dispatchData_clock = clock;
  assign dispatchData_io_raddr_0 = _T_129 ? _commitReadAddr_next_WIRE__0 : walkPtrVec_next_0_value; // @[Rob.scala 950:32]
  assign dispatchData_io_raddr_1 = _T_129 ? _commitReadAddr_next_WIRE__1 : walkPtrVec_next_1_value; // @[Rob.scala 950:32]
  assign dispatchData_io_wen_0 = io_enq_req_0_valid & io_enq_canAccept; // @[Rob.scala 519:51]
  assign dispatchData_io_wen_1 = io_enq_req_1_valid & io_enq_canAccept; // @[Rob.scala 519:51]
  assign dispatchData_io_waddr_0 = enqPtrGenModule_io_out_0_value; // @[Rob.scala 447:23 791:13]
  assign dispatchData_io_waddr_1 = io_enq_needAlloc_0 ? enqPtrVec_1_value : enqPtrVec_0_value; // @[Rob.scala 516:{31,31}]
  assign dispatchData_io_wdata_0_ldest = io_enq_req_0_bits_ctrl_ldest; // @[Rob.scala 958:17]
  assign dispatchData_io_wdata_0_rfWen = io_enq_req_0_bits_ctrl_rfWen; // @[Rob.scala 959:17]
  assign dispatchData_io_wdata_0_fpWen = io_enq_req_0_bits_ctrl_fpWen; // @[Rob.scala 960:17]
  assign dispatchData_io_wdata_0_wflags = io_enq_req_0_bits_ctrl_fpu_wflags; // @[Rob.scala 961:18]
  assign dispatchData_io_wdata_0_commitType = io_enq_req_0_bits_ctrl_commitType; // @[Rob.scala 962:22]
  assign dispatchData_io_wdata_0_pdest = io_enq_req_0_bits_pdest; // @[Rob.scala 963:17]
  assign dispatchData_io_wdata_0_old_pdest = io_enq_req_0_bits_old_pdest; // @[Rob.scala 964:21]
  assign dispatchData_io_wdata_0_ftqIdx_flag = io_enq_req_0_bits_cf_ftqPtr_flag; // @[Rob.scala 965:18]
  assign dispatchData_io_wdata_0_ftqIdx_value = io_enq_req_0_bits_cf_ftqPtr_value; // @[Rob.scala 965:18]
  assign dispatchData_io_wdata_0_ftqOffset = io_enq_req_0_bits_cf_ftqOffset; // @[Rob.scala 966:21]
  assign dispatchData_io_wdata_0_isMove = io_enq_req_0_bits_eliminatedMove; // @[Rob.scala 967:18]
  assign dispatchData_io_wdata_1_ldest = io_enq_req_1_bits_ctrl_ldest; // @[Rob.scala 958:17]
  assign dispatchData_io_wdata_1_rfWen = io_enq_req_1_bits_ctrl_rfWen; // @[Rob.scala 959:17]
  assign dispatchData_io_wdata_1_fpWen = io_enq_req_1_bits_ctrl_fpWen; // @[Rob.scala 960:17]
  assign dispatchData_io_wdata_1_wflags = io_enq_req_1_bits_ctrl_fpu_wflags; // @[Rob.scala 961:18]
  assign dispatchData_io_wdata_1_commitType = io_enq_req_1_bits_ctrl_commitType; // @[Rob.scala 962:22]
  assign dispatchData_io_wdata_1_pdest = io_enq_req_1_bits_pdest; // @[Rob.scala 963:17]
  assign dispatchData_io_wdata_1_old_pdest = io_enq_req_1_bits_old_pdest; // @[Rob.scala 964:21]
  assign dispatchData_io_wdata_1_ftqIdx_flag = io_enq_req_1_bits_cf_ftqPtr_flag; // @[Rob.scala 965:18]
  assign dispatchData_io_wdata_1_ftqIdx_value = io_enq_req_1_bits_cf_ftqPtr_value; // @[Rob.scala 965:18]
  assign dispatchData_io_wdata_1_ftqOffset = io_enq_req_1_bits_cf_ftqOffset; // @[Rob.scala 966:21]
  assign dispatchData_io_wdata_1_isMove = io_enq_req_1_bits_eliminatedMove; // @[Rob.scala 967:18]
  assign exceptionGen_clock = clock;
  assign exceptionGen_reset = reset;
  assign exceptionGen_io_redirect_valid = io_redirect_valid; // @[Rob.scala 972:28]
  assign exceptionGen_io_redirect_bits_robIdx_flag = io_redirect_bits_robIdx_flag; // @[Rob.scala 972:28]
  assign exceptionGen_io_redirect_bits_robIdx_value = io_redirect_bits_robIdx_value; // @[Rob.scala 972:28]
  assign exceptionGen_io_redirect_bits_level = io_redirect_bits_level; // @[Rob.scala 972:28]
  assign exceptionGen_io_flush = io_flushOut_valid; // @[Rob.scala 973:25]
  assign exceptionGen_io_enq_0_valid = io_enq_req_0_valid & io_enq_canAccept; // @[Rob.scala 519:51]
  assign exceptionGen_io_enq_0_bits_robIdx_flag = io_enq_req_0_bits_robIdx_flag; // @[Rob.scala 976:40]
  assign exceptionGen_io_enq_0_bits_robIdx_value = io_enq_req_0_bits_robIdx_value; // @[Rob.scala 976:40]
  assign exceptionGen_io_enq_0_bits_exceptionVec_1 = io_enq_req_0_bits_cf_exceptionVec_1; // @[package.scala 549:25 551:38]
  assign exceptionGen_io_enq_0_bits_exceptionVec_2 = io_enq_req_0_bits_cf_exceptionVec_2; // @[package.scala 549:25 551:38]
  assign exceptionGen_io_enq_0_bits_exceptionVec_12 = io_enq_req_0_bits_cf_exceptionVec_12; // @[package.scala 549:25 551:38]
  assign exceptionGen_io_enq_0_bits_flushPipe = io_enq_req_0_bits_ctrl_flushPipe; // @[Rob.scala 978:43]
  assign exceptionGen_io_enq_0_bits_singleStep = io_enq_req_0_bits_ctrl_singleStep; // @[Rob.scala 981:44]
  assign exceptionGen_io_enq_0_bits_crossPageIPFFix = io_enq_req_0_bits_cf_crossPageIPFFix; // @[Rob.scala 982:49]
  assign exceptionGen_io_enq_0_bits_trigger_frontendHit_0 = io_enq_req_0_bits_cf_trigger_frontendHit_0; // @[Rob.scala 984:53]
  assign exceptionGen_io_enq_0_bits_trigger_frontendHit_1 = io_enq_req_0_bits_cf_trigger_frontendHit_1; // @[Rob.scala 984:53]
  assign exceptionGen_io_enq_0_bits_trigger_frontendHit_2 = io_enq_req_0_bits_cf_trigger_frontendHit_2; // @[Rob.scala 984:53]
  assign exceptionGen_io_enq_0_bits_trigger_frontendHit_3 = io_enq_req_0_bits_cf_trigger_frontendHit_3; // @[Rob.scala 984:53]
  assign exceptionGen_io_enq_1_valid = io_enq_req_1_valid & io_enq_canAccept; // @[Rob.scala 519:51]
  assign exceptionGen_io_enq_1_bits_robIdx_flag = io_enq_req_1_bits_robIdx_flag; // @[Rob.scala 976:40]
  assign exceptionGen_io_enq_1_bits_robIdx_value = io_enq_req_1_bits_robIdx_value; // @[Rob.scala 976:40]
  assign exceptionGen_io_enq_1_bits_exceptionVec_1 = io_enq_req_1_bits_cf_exceptionVec_1; // @[package.scala 549:25 551:38]
  assign exceptionGen_io_enq_1_bits_exceptionVec_2 = io_enq_req_1_bits_cf_exceptionVec_2; // @[package.scala 549:25 551:38]
  assign exceptionGen_io_enq_1_bits_exceptionVec_12 = io_enq_req_1_bits_cf_exceptionVec_12; // @[package.scala 549:25 551:38]
  assign exceptionGen_io_enq_1_bits_flushPipe = io_enq_req_1_bits_ctrl_flushPipe; // @[Rob.scala 978:43]
  assign exceptionGen_io_enq_1_bits_singleStep = io_enq_req_1_bits_ctrl_singleStep; // @[Rob.scala 981:44]
  assign exceptionGen_io_enq_1_bits_crossPageIPFFix = io_enq_req_1_bits_cf_crossPageIPFFix; // @[Rob.scala 982:49]
  assign exceptionGen_io_enq_1_bits_trigger_frontendHit_0 = io_enq_req_1_bits_cf_trigger_frontendHit_0; // @[Rob.scala 984:53]
  assign exceptionGen_io_enq_1_bits_trigger_frontendHit_1 = io_enq_req_1_bits_cf_trigger_frontendHit_1; // @[Rob.scala 984:53]
  assign exceptionGen_io_enq_1_bits_trigger_frontendHit_2 = io_enq_req_1_bits_cf_trigger_frontendHit_2; // @[Rob.scala 984:53]
  assign exceptionGen_io_enq_1_bits_trigger_frontendHit_3 = io_enq_req_1_bits_cf_trigger_frontendHit_3; // @[Rob.scala 984:53]
  assign exceptionGen_io_wb_0_valid = io_writeback_0_3_valid; // @[Rob.scala 991:33]
  assign exceptionGen_io_wb_0_bits_robIdx_flag = io_writeback_0_3_bits_uop_robIdx_flag; // @[Rob.scala 992:33]
  assign exceptionGen_io_wb_0_bits_robIdx_value = io_writeback_0_3_bits_uop_robIdx_value; // @[Rob.scala 992:33]
  assign exceptionGen_io_wb_0_bits_exceptionVec_2 = io_writeback_0_3_bits_uop_cf_exceptionVec_2; // @[package.scala 549:25 551:38]
  assign exceptionGen_io_wb_0_bits_exceptionVec_3 = io_writeback_0_3_bits_uop_cf_exceptionVec_3; // @[package.scala 549:25 551:38]
  assign exceptionGen_io_wb_0_bits_exceptionVec_8 = io_writeback_0_3_bits_uop_cf_exceptionVec_8; // @[package.scala 549:25 551:38]
  assign exceptionGen_io_wb_0_bits_exceptionVec_9 = io_writeback_0_3_bits_uop_cf_exceptionVec_9; // @[package.scala 549:25 551:38]
  assign exceptionGen_io_wb_0_bits_exceptionVec_11 = io_writeback_0_3_bits_uop_cf_exceptionVec_11; // @[package.scala 549:25 551:38]
  assign exceptionGen_io_wb_0_bits_flushPipe = io_writeback_0_3_bits_uop_ctrl_flushPipe; // @[Rob.scala 994:66]
  assign exceptionGen_io_wb_1_valid = io_writeback_0_6_valid; // @[Rob.scala 991:33]
  assign exceptionGen_io_wb_1_bits_robIdx_flag = io_writeback_0_6_bits_uop_robIdx_flag; // @[Rob.scala 992:33]
  assign exceptionGen_io_wb_1_bits_robIdx_value = io_writeback_0_6_bits_uop_robIdx_value; // @[Rob.scala 992:33]
  assign exceptionGen_io_wb_1_bits_exceptionVec_4 = io_writeback_0_6_bits_uop_cf_exceptionVec_4; // @[package.scala 549:25 551:38]
  assign exceptionGen_io_wb_1_bits_exceptionVec_5 = io_writeback_0_6_bits_uop_cf_exceptionVec_5; // @[package.scala 549:25 551:38]
  assign exceptionGen_io_wb_1_bits_exceptionVec_13 = io_writeback_0_6_bits_uop_cf_exceptionVec_13; // @[package.scala 549:25 551:38]
  assign exceptionGen_io_wb_1_bits_flushPipe = io_writeback_0_6_bits_uop_ctrl_flushPipe; // @[Rob.scala 994:66]
  assign exceptionGen_io_wb_1_bits_replayInst = io_writeback_0_6_bits_uop_ctrl_replayInst; // @[Rob.scala 995:67]
  assign exceptionGen_io_wb_1_bits_trigger_backendHit_0 = io_writeback_0_6_bits_uop_cf_trigger_backendHit_0; // @[Rob.scala 1000:36]
  assign exceptionGen_io_wb_1_bits_trigger_backendHit_1 = io_writeback_0_6_bits_uop_cf_trigger_backendHit_1; // @[Rob.scala 1000:36]
  assign exceptionGen_io_wb_1_bits_trigger_backendHit_2 = io_writeback_0_6_bits_uop_cf_trigger_backendHit_2; // @[Rob.scala 1000:36]
  assign exceptionGen_io_wb_1_bits_trigger_backendHit_3 = io_writeback_0_6_bits_uop_cf_trigger_backendHit_3; // @[Rob.scala 1000:36]
  assign exceptionGen_io_wb_1_bits_trigger_backendHit_4 = io_writeback_0_6_bits_uop_cf_trigger_backendHit_4; // @[Rob.scala 1000:36]
  assign exceptionGen_io_wb_1_bits_trigger_backendHit_5 = io_writeback_0_6_bits_uop_cf_trigger_backendHit_5; // @[Rob.scala 1000:36]
  assign exceptionGen_io_wb_2_valid = io_writeback_0_7_valid; // @[Rob.scala 991:33]
  assign exceptionGen_io_wb_2_bits_robIdx_flag = io_writeback_0_7_bits_uop_robIdx_flag; // @[Rob.scala 992:33]
  assign exceptionGen_io_wb_2_bits_robIdx_value = io_writeback_0_7_bits_uop_robIdx_value; // @[Rob.scala 992:33]
  assign exceptionGen_io_wb_2_bits_exceptionVec_4 = io_writeback_0_7_bits_uop_cf_exceptionVec_4; // @[package.scala 549:25 551:38]
  assign exceptionGen_io_wb_2_bits_exceptionVec_5 = io_writeback_0_7_bits_uop_cf_exceptionVec_5; // @[package.scala 549:25 551:38]
  assign exceptionGen_io_wb_2_bits_exceptionVec_13 = io_writeback_0_7_bits_uop_cf_exceptionVec_13; // @[package.scala 549:25 551:38]
  assign exceptionGen_io_wb_2_bits_flushPipe = io_writeback_0_7_bits_uop_ctrl_flushPipe; // @[Rob.scala 994:66]
  assign exceptionGen_io_wb_2_bits_replayInst = io_writeback_0_7_bits_uop_ctrl_replayInst; // @[Rob.scala 995:67]
  assign exceptionGen_io_wb_2_bits_trigger_backendHit_0 = io_writeback_0_7_bits_uop_cf_trigger_backendHit_0; // @[Rob.scala 1000:36]
  assign exceptionGen_io_wb_2_bits_trigger_backendHit_1 = io_writeback_0_7_bits_uop_cf_trigger_backendHit_1; // @[Rob.scala 1000:36]
  assign exceptionGen_io_wb_2_bits_trigger_backendHit_2 = io_writeback_0_7_bits_uop_cf_trigger_backendHit_2; // @[Rob.scala 1000:36]
  assign exceptionGen_io_wb_2_bits_trigger_backendHit_3 = io_writeback_0_7_bits_uop_cf_trigger_backendHit_3; // @[Rob.scala 1000:36]
  assign exceptionGen_io_wb_2_bits_trigger_backendHit_4 = io_writeback_0_7_bits_uop_cf_trigger_backendHit_4; // @[Rob.scala 1000:36]
  assign exceptionGen_io_wb_2_bits_trigger_backendHit_5 = io_writeback_0_7_bits_uop_cf_trigger_backendHit_5; // @[Rob.scala 1000:36]
  assign exceptionGen_io_wb_3_valid = io_writeback_0_8_valid; // @[Rob.scala 991:33]
  assign exceptionGen_io_wb_3_bits_robIdx_flag = io_writeback_0_8_bits_uop_robIdx_flag; // @[Rob.scala 992:33]
  assign exceptionGen_io_wb_3_bits_robIdx_value = io_writeback_0_8_bits_uop_robIdx_value; // @[Rob.scala 992:33]
  assign exceptionGen_io_wb_3_bits_exceptionVec_4 = io_writeback_0_8_bits_uop_cf_exceptionVec_4; // @[package.scala 549:25 551:38]
  assign exceptionGen_io_wb_3_bits_exceptionVec_5 = io_writeback_0_8_bits_uop_cf_exceptionVec_5; // @[package.scala 549:25 551:38]
  assign exceptionGen_io_wb_3_bits_exceptionVec_6 = io_writeback_0_8_bits_uop_cf_exceptionVec_6; // @[package.scala 549:25 551:38]
  assign exceptionGen_io_wb_3_bits_exceptionVec_7 = io_writeback_0_8_bits_uop_cf_exceptionVec_7; // @[package.scala 549:25 551:38]
  assign exceptionGen_io_wb_3_bits_exceptionVec_13 = io_writeback_0_8_bits_uop_cf_exceptionVec_13; // @[package.scala 549:25 551:38]
  assign exceptionGen_io_wb_3_bits_exceptionVec_15 = io_writeback_0_8_bits_uop_cf_exceptionVec_15; // @[package.scala 549:25 551:38]
  assign exceptionGen_io_wb_3_bits_trigger_backendHit_0 = io_writeback_0_8_bits_uop_cf_trigger_backendHit_0; // @[Rob.scala 1000:36]
  assign exceptionGen_io_wb_3_bits_trigger_backendHit_1 = io_writeback_0_8_bits_uop_cf_trigger_backendHit_1; // @[Rob.scala 1000:36]
  assign exceptionGen_io_wb_3_bits_trigger_backendHit_2 = io_writeback_0_8_bits_uop_cf_trigger_backendHit_2; // @[Rob.scala 1000:36]
  assign exceptionGen_io_wb_3_bits_trigger_backendHit_3 = io_writeback_0_8_bits_uop_cf_trigger_backendHit_3; // @[Rob.scala 1000:36]
  assign exceptionGen_io_wb_3_bits_trigger_backendHit_4 = io_writeback_0_8_bits_uop_cf_trigger_backendHit_4; // @[Rob.scala 1000:36]
  assign exceptionGen_io_wb_3_bits_trigger_backendHit_5 = io_writeback_0_8_bits_uop_cf_trigger_backendHit_5; // @[Rob.scala 1000:36]
  assign exceptionGen_io_wb_4_valid = io_writeback_0_9_valid; // @[Rob.scala 991:33]
  assign exceptionGen_io_wb_4_bits_robIdx_flag = io_writeback_0_9_bits_uop_robIdx_flag; // @[Rob.scala 992:33]
  assign exceptionGen_io_wb_4_bits_robIdx_value = io_writeback_0_9_bits_uop_robIdx_value; // @[Rob.scala 992:33]
  assign exceptionGen_io_wb_4_bits_exceptionVec_6 = io_writeback_0_9_bits_uop_cf_exceptionVec_6; // @[package.scala 549:25 551:38]
  assign exceptionGen_io_wb_4_bits_exceptionVec_7 = io_writeback_0_9_bits_uop_cf_exceptionVec_7; // @[package.scala 549:25 551:38]
  assign exceptionGen_io_wb_4_bits_exceptionVec_15 = io_writeback_0_9_bits_uop_cf_exceptionVec_15; // @[package.scala 549:25 551:38]
  assign exceptionGen_io_wb_4_bits_trigger_backendHit_0 = io_writeback_0_9_bits_uop_cf_trigger_backendHit_0; // @[Rob.scala 1000:36]
  assign exceptionGen_io_wb_4_bits_trigger_backendHit_1 = io_writeback_0_9_bits_uop_cf_trigger_backendHit_1; // @[Rob.scala 1000:36]
  assign exceptionGen_io_wb_4_bits_trigger_backendHit_4 = io_writeback_0_9_bits_uop_cf_trigger_backendHit_4; // @[Rob.scala 1000:36]
  assign deqPtrGenModule_clock = clock;
  assign deqPtrGenModule_reset = reset;
  assign deqPtrGenModule_io_state = {{1'd0}, state}; // @[Rob.scala 775:28]
  assign deqPtrGenModule_io_deq_v_0 = 5'h1f == deqPtrVec_0_value ? valid_31 : _GEN_4837; // @[Rob.scala 636:{43,43}]
  assign deqPtrGenModule_io_deq_v_1 = 5'h1f == deqPtrVec_1_value ? valid_31 : _GEN_5073; // @[Rob.scala 703:{25,25}]
  assign deqPtrGenModule_io_deq_w0 = writebacked_commit_wMPORT_data & store_data_writebacked_commit_wMPORT_1_data; // @[Rob.scala 705:70]
  assign deqPtrGenModule_io_deq_w1 = writebacked_commit_wMPORT_2_data & store_data_writebacked_commit_wMPORT_3_data; // @[Rob.scala 705:70]
  assign deqPtrGenModule_io_exception_state_valid = exceptionGen_io_state_valid; // @[Rob.scala 778:38]
  assign deqPtrGenModule_io_exception_state_bits_robIdx_flag = exceptionGen_io_state_bits_robIdx_flag; // @[Rob.scala 778:38]
  assign deqPtrGenModule_io_exception_state_bits_robIdx_value = exceptionGen_io_state_bits_robIdx_value; // @[Rob.scala 778:38]
  assign deqPtrGenModule_io_exception_state_bits_exceptionVec_0 = exceptionGen_io_state_bits_exceptionVec_0; // @[Rob.scala 778:38]
  assign deqPtrGenModule_io_exception_state_bits_exceptionVec_1 = exceptionGen_io_state_bits_exceptionVec_1; // @[Rob.scala 778:38]
  assign deqPtrGenModule_io_exception_state_bits_exceptionVec_2 = exceptionGen_io_state_bits_exceptionVec_2; // @[Rob.scala 778:38]
  assign deqPtrGenModule_io_exception_state_bits_exceptionVec_3 = exceptionGen_io_state_bits_exceptionVec_3; // @[Rob.scala 778:38]
  assign deqPtrGenModule_io_exception_state_bits_exceptionVec_4 = exceptionGen_io_state_bits_exceptionVec_4; // @[Rob.scala 778:38]
  assign deqPtrGenModule_io_exception_state_bits_exceptionVec_5 = exceptionGen_io_state_bits_exceptionVec_5; // @[Rob.scala 778:38]
  assign deqPtrGenModule_io_exception_state_bits_exceptionVec_6 = exceptionGen_io_state_bits_exceptionVec_6; // @[Rob.scala 778:38]
  assign deqPtrGenModule_io_exception_state_bits_exceptionVec_7 = exceptionGen_io_state_bits_exceptionVec_7; // @[Rob.scala 778:38]
  assign deqPtrGenModule_io_exception_state_bits_exceptionVec_8 = exceptionGen_io_state_bits_exceptionVec_8; // @[Rob.scala 778:38]
  assign deqPtrGenModule_io_exception_state_bits_exceptionVec_9 = exceptionGen_io_state_bits_exceptionVec_9; // @[Rob.scala 778:38]
  assign deqPtrGenModule_io_exception_state_bits_exceptionVec_10 = exceptionGen_io_state_bits_exceptionVec_10; // @[Rob.scala 778:38]
  assign deqPtrGenModule_io_exception_state_bits_exceptionVec_11 = exceptionGen_io_state_bits_exceptionVec_11; // @[Rob.scala 778:38]
  assign deqPtrGenModule_io_exception_state_bits_exceptionVec_12 = exceptionGen_io_state_bits_exceptionVec_12; // @[Rob.scala 778:38]
  assign deqPtrGenModule_io_exception_state_bits_exceptionVec_13 = exceptionGen_io_state_bits_exceptionVec_13; // @[Rob.scala 778:38]
  assign deqPtrGenModule_io_exception_state_bits_exceptionVec_14 = exceptionGen_io_state_bits_exceptionVec_14; // @[Rob.scala 778:38]
  assign deqPtrGenModule_io_exception_state_bits_exceptionVec_15 = exceptionGen_io_state_bits_exceptionVec_15; // @[Rob.scala 778:38]
  assign deqPtrGenModule_io_exception_state_bits_replayInst = exceptionGen_io_state_bits_replayInst; // @[Rob.scala 778:38]
  assign deqPtrGenModule_io_exception_state_bits_singleStep = exceptionGen_io_state_bits_singleStep; // @[Rob.scala 778:38]
  assign deqPtrGenModule_io_exception_state_bits_trigger_frontendHit_0 =
    exceptionGen_io_state_bits_trigger_frontendHit_0; // @[Rob.scala 778:38]
  assign deqPtrGenModule_io_exception_state_bits_trigger_frontendHit_1 =
    exceptionGen_io_state_bits_trigger_frontendHit_1; // @[Rob.scala 778:38]
  assign deqPtrGenModule_io_exception_state_bits_trigger_frontendHit_2 =
    exceptionGen_io_state_bits_trigger_frontendHit_2; // @[Rob.scala 778:38]
  assign deqPtrGenModule_io_exception_state_bits_trigger_frontendHit_3 =
    exceptionGen_io_state_bits_trigger_frontendHit_3; // @[Rob.scala 778:38]
  assign deqPtrGenModule_io_exception_state_bits_trigger_backendHit_0 = exceptionGen_io_state_bits_trigger_backendHit_0; // @[Rob.scala 778:38]
  assign deqPtrGenModule_io_exception_state_bits_trigger_backendHit_1 = exceptionGen_io_state_bits_trigger_backendHit_1; // @[Rob.scala 778:38]
  assign deqPtrGenModule_io_exception_state_bits_trigger_backendHit_2 = exceptionGen_io_state_bits_trigger_backendHit_2; // @[Rob.scala 778:38]
  assign deqPtrGenModule_io_exception_state_bits_trigger_backendHit_3 = exceptionGen_io_state_bits_trigger_backendHit_3; // @[Rob.scala 778:38]
  assign deqPtrGenModule_io_exception_state_bits_trigger_backendHit_4 = exceptionGen_io_state_bits_trigger_backendHit_4; // @[Rob.scala 778:38]
  assign deqPtrGenModule_io_exception_state_bits_trigger_backendHit_5 = exceptionGen_io_state_bits_trigger_backendHit_5; // @[Rob.scala 778:38]
  assign deqPtrGenModule_io_intrBitSetReg = intrBitSetReg; // @[Rob.scala 779:36]
  assign deqPtrGenModule_io_hasNoSpecExec = hasNoSpecExec; // @[Rob.scala 780:36]
  assign deqPtrGenModule_io_interrupt_safe = interrupt_safe_deqPtrGenModule_io_interrupt_safe_MPORT_data; // @[Rob.scala 781:37]
  assign deqPtrGenModule_io_blockCommit = misPredBlock | isReplaying | lastCycleFlush | hasWFI; // @[Rob.scala 698:67]
  assign enqPtrGenModule_clock = clock;
  assign enqPtrGenModule_reset = reset;
  assign enqPtrGenModule_io_redirect_valid = io_redirect_valid; // @[Rob.scala 787:31]
  assign enqPtrGenModule_io_redirect_bits_robIdx_flag = io_redirect_bits_robIdx_flag; // @[Rob.scala 787:31]
  assign enqPtrGenModule_io_redirect_bits_robIdx_value = io_redirect_bits_robIdx_value; // @[Rob.scala 787:31]
  assign enqPtrGenModule_io_redirect_bits_level = io_redirect_bits_level; // @[Rob.scala 787:31]
  assign enqPtrGenModule_io_allowEnqueue = allowEnqueue; // @[Rob.scala 788:35]
  assign enqPtrGenModule_io_hasBlockBackward = hasBlockBackward; // @[Rob.scala 789:39]
  assign enqPtrGenModule_io_enq_0 = io_enq_req_0_valid; // @[Rob.scala 790:{36,36}]
  assign enqPtrGenModule_io_enq_1 = io_enq_req_1_valid; // @[Rob.scala 790:{36,36}]
  assign fflagsDataModule_clock = clock;
  assign fflagsDataModule_io_raddr_0 = deqPtrGenModule_io_next_out_0_value; // @[Rob.scala 1015:{39,39}]
  assign fflagsDataModule_io_raddr_1 = deqPtrGenModule_io_next_out_1_value; // @[Rob.scala 1015:{39,39}]
  assign fflagsDataModule_io_wen_0 = io_writeback_0_3_valid; // @[Rob.scala 1011:34]
  assign fflagsDataModule_io_wen_1 = io_writeback_0_4_valid; // @[Rob.scala 1011:34]
  assign fflagsDataModule_io_wen_2 = io_writeback_0_5_valid; // @[Rob.scala 1011:34]
  assign fflagsDataModule_io_waddr_0 = io_writeback_0_3_bits_uop_robIdx_value; // @[Rob.scala 1012:34]
  assign fflagsDataModule_io_waddr_1 = io_writeback_0_4_bits_uop_robIdx_value; // @[Rob.scala 1012:34]
  assign fflagsDataModule_io_waddr_2 = io_writeback_0_5_bits_uop_robIdx_value; // @[Rob.scala 1012:34]
  assign fflagsDataModule_io_wdata_0 = io_writeback_0_3_bits_fflags; // @[Rob.scala 1013:34]
  assign fflagsDataModule_io_wdata_1 = io_writeback_0_4_bits_fflags; // @[Rob.scala 1013:34]
  assign fflagsDataModule_io_wdata_2 = io_writeback_0_5_bits_fflags; // @[Rob.scala 1013:34]
  assign difftest_io_clock = clock; // @[Rob.scala 1236:27]
  assign difftest_io_coreid = io_hartId; // @[Rob.scala 1237:27]
  assign difftest_io_index = 8'h0; // @[Rob.scala 1238:27]
  assign difftest_io_valid = difftest_io_valid_REG_2; // @[Rob.scala 1239:27]
  assign difftest_io_special = {{7'd0}, difftest_io_special_REG_2}; // @[Rob.scala 1240:27]
  assign difftest_io_skip = difftest_io_skip_REG_2; // @[Rob.scala 1241:27]
  assign difftest_io_isRVC = difftest_io_isRVC_REG_2; // @[Rob.scala 1242:27]
  assign difftest_io_rfwen = difftest_io_rfwen_REG_2; // @[Rob.scala 1243:27]
  assign difftest_io_fpwen = difftest_io_fpwen_REG_2; // @[Rob.scala 1244:27]
  assign difftest_io_wpdest = {{26'd0}, difftest_io_wpdest_REG_2}; // @[Rob.scala 1245:27]
  assign difftest_io_wdest = {{3'd0}, difftest_io_wdest_REG_2}; // @[Rob.scala 1246:27]
  assign difftest_1_io_clock = clock; // @[Rob.scala 1236:27]
  assign difftest_1_io_coreid = io_hartId; // @[Rob.scala 1237:27]
  assign difftest_1_io_index = 8'h1; // @[Rob.scala 1238:27]
  assign difftest_1_io_valid = difftest_io_valid_REG_5; // @[Rob.scala 1239:27]
  assign difftest_1_io_special = {{7'd0}, difftest_io_special_REG_5}; // @[Rob.scala 1240:27]
  assign difftest_1_io_skip = difftest_io_skip_REG_5; // @[Rob.scala 1241:27]
  assign difftest_1_io_isRVC = difftest_io_isRVC_REG_5; // @[Rob.scala 1242:27]
  assign difftest_1_io_rfwen = difftest_io_rfwen_REG_5; // @[Rob.scala 1243:27]
  assign difftest_1_io_fpwen = difftest_io_fpwen_REG_5; // @[Rob.scala 1244:27]
  assign difftest_1_io_wpdest = {{26'd0}, difftest_io_wpdest_REG_5}; // @[Rob.scala 1245:27]
  assign difftest_1_io_wdest = {{3'd0}, difftest_io_wdest_REG_5}; // @[Rob.scala 1246:27]
  assign difftest_2_io_clock = clock; // @[Rob.scala 1299:26]
  assign difftest_2_io_coreid = io_hartId; // @[Rob.scala 1300:26]
  assign difftest_2_io_valid = trapVec_0 | trapVec_1; // @[Rob.scala 1297:35]
  assign difftest_2_io_cycleCnt = timer; // @[Rob.scala 1302:26]
  assign difftest_2_io_instrCnt = instrCntReg + _GEN_11347; // @[Rob.scala 1022:30]
  assign difftest_2_io_hasWFI = 1'h0;
  always @(posedge clock) begin
    if (writebacked_MPORT_92_en & writebacked_MPORT_92_mask) begin
      writebacked[writebacked_MPORT_92_addr] <= writebacked_MPORT_92_data; // @[Rob.scala 428:24]
    end
    if (writebacked_MPORT_94_en & writebacked_MPORT_94_mask) begin
      writebacked[writebacked_MPORT_94_addr] <= writebacked_MPORT_94_data; // @[Rob.scala 428:24]
    end
    if (writebacked_MPORT_96_en & writebacked_MPORT_96_mask) begin
      writebacked[writebacked_MPORT_96_addr] <= writebacked_MPORT_96_data; // @[Rob.scala 428:24]
    end
    if (writebacked_MPORT_98_en & writebacked_MPORT_98_mask) begin
      writebacked[writebacked_MPORT_98_addr] <= writebacked_MPORT_98_data; // @[Rob.scala 428:24]
    end
    if (writebacked_MPORT_99_en & writebacked_MPORT_99_mask) begin
      writebacked[writebacked_MPORT_99_addr] <= writebacked_MPORT_99_data; // @[Rob.scala 428:24]
    end
    if (writebacked_MPORT_100_en & writebacked_MPORT_100_mask) begin
      writebacked[writebacked_MPORT_100_addr] <= writebacked_MPORT_100_data; // @[Rob.scala 428:24]
    end
    if (writebacked_MPORT_101_en & writebacked_MPORT_101_mask) begin
      writebacked[writebacked_MPORT_101_addr] <= writebacked_MPORT_101_data; // @[Rob.scala 428:24]
    end
    if (writebacked_MPORT_102_en & writebacked_MPORT_102_mask) begin
      writebacked[writebacked_MPORT_102_addr] <= writebacked_MPORT_102_data; // @[Rob.scala 428:24]
    end
    if (writebacked_MPORT_103_en & writebacked_MPORT_103_mask) begin
      writebacked[writebacked_MPORT_103_addr] <= writebacked_MPORT_103_data; // @[Rob.scala 428:24]
    end
    if (writebacked_MPORT_104_en & writebacked_MPORT_104_mask) begin
      writebacked[writebacked_MPORT_104_addr] <= writebacked_MPORT_104_data; // @[Rob.scala 428:24]
    end
    if (writebacked_MPORT_105_en & writebacked_MPORT_105_mask) begin
      writebacked[writebacked_MPORT_105_addr] <= writebacked_MPORT_105_data; // @[Rob.scala 428:24]
    end
    if (writebacked_MPORT_106_en & writebacked_MPORT_106_mask) begin
      writebacked[writebacked_MPORT_106_addr] <= writebacked_MPORT_106_data; // @[Rob.scala 428:24]
    end
    if (store_data_writebacked_MPORT_93_en & store_data_writebacked_MPORT_93_mask) begin
      store_data_writebacked[store_data_writebacked_MPORT_93_addr] <= store_data_writebacked_MPORT_93_data; // @[Rob.scala 429:35]
    end
    if (store_data_writebacked_MPORT_95_en & store_data_writebacked_MPORT_95_mask) begin
      store_data_writebacked[store_data_writebacked_MPORT_95_addr] <= store_data_writebacked_MPORT_95_data; // @[Rob.scala 429:35]
    end
    if (store_data_writebacked_MPORT_97_en & store_data_writebacked_MPORT_97_mask) begin
      store_data_writebacked[store_data_writebacked_MPORT_97_addr] <= store_data_writebacked_MPORT_97_data; // @[Rob.scala 429:35]
    end
    if (store_data_writebacked_MPORT_107_en & store_data_writebacked_MPORT_107_mask) begin
      store_data_writebacked[store_data_writebacked_MPORT_107_addr] <= store_data_writebacked_MPORT_107_data; // @[Rob.scala 429:35]
    end
    if (store_data_writebacked_MPORT_108_en & store_data_writebacked_MPORT_108_mask) begin
      store_data_writebacked[store_data_writebacked_MPORT_108_addr] <= store_data_writebacked_MPORT_108_data; // @[Rob.scala 429:35]
    end
    if (interrupt_safe_MPORT_111_en & interrupt_safe_MPORT_111_mask) begin
      interrupt_safe[interrupt_safe_MPORT_111_addr] <= interrupt_safe_MPORT_111_data; // @[Rob.scala 436:27]
    end
    if (interrupt_safe_MPORT_112_en & interrupt_safe_MPORT_112_mask) begin
      interrupt_safe[interrupt_safe_MPORT_112_addr] <= interrupt_safe_MPORT_112_data; // @[Rob.scala 436:27]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_en & debug_microOp_cf_loadWaitBit_MPORT_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_addr] <= debug_microOp_cf_loadWaitBit_MPORT_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_1_en & debug_microOp_cf_loadWaitBit_MPORT_1_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_1_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_1_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_2_en & debug_microOp_cf_loadWaitBit_MPORT_2_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_2_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_2_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_3_en & debug_microOp_cf_loadWaitBit_MPORT_3_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_3_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_3_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_4_en & debug_microOp_cf_loadWaitBit_MPORT_4_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_4_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_4_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_5_en & debug_microOp_cf_loadWaitBit_MPORT_5_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_5_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_5_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_6_en & debug_microOp_cf_loadWaitBit_MPORT_6_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_6_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_6_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_7_en & debug_microOp_cf_loadWaitBit_MPORT_7_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_7_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_7_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_8_en & debug_microOp_cf_loadWaitBit_MPORT_8_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_8_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_8_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_9_en & debug_microOp_cf_loadWaitBit_MPORT_9_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_9_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_9_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_10_en & debug_microOp_cf_loadWaitBit_MPORT_10_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_10_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_10_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_11_en & debug_microOp_cf_loadWaitBit_MPORT_11_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_11_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_11_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_12_en & debug_microOp_cf_loadWaitBit_MPORT_12_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_12_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_12_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_13_en & debug_microOp_cf_loadWaitBit_MPORT_13_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_13_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_13_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_14_en & debug_microOp_cf_loadWaitBit_MPORT_14_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_14_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_14_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_15_en & debug_microOp_cf_loadWaitBit_MPORT_15_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_15_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_15_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_16_en & debug_microOp_cf_loadWaitBit_MPORT_16_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_16_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_16_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_17_en & debug_microOp_cf_loadWaitBit_MPORT_17_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_17_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_17_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_18_en & debug_microOp_cf_loadWaitBit_MPORT_18_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_18_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_18_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_19_en & debug_microOp_cf_loadWaitBit_MPORT_19_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_19_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_19_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_20_en & debug_microOp_cf_loadWaitBit_MPORT_20_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_20_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_20_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_21_en & debug_microOp_cf_loadWaitBit_MPORT_21_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_21_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_21_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_22_en & debug_microOp_cf_loadWaitBit_MPORT_22_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_22_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_22_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_23_en & debug_microOp_cf_loadWaitBit_MPORT_23_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_23_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_23_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_24_en & debug_microOp_cf_loadWaitBit_MPORT_24_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_24_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_24_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_25_en & debug_microOp_cf_loadWaitBit_MPORT_25_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_25_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_25_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_26_en & debug_microOp_cf_loadWaitBit_MPORT_26_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_26_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_26_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_27_en & debug_microOp_cf_loadWaitBit_MPORT_27_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_27_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_27_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_28_en & debug_microOp_cf_loadWaitBit_MPORT_28_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_28_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_28_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_29_en & debug_microOp_cf_loadWaitBit_MPORT_29_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_29_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_29_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_30_en & debug_microOp_cf_loadWaitBit_MPORT_30_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_30_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_30_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_31_en & debug_microOp_cf_loadWaitBit_MPORT_31_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_31_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_31_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_32_en & debug_microOp_cf_loadWaitBit_MPORT_32_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_32_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_32_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_33_en & debug_microOp_cf_loadWaitBit_MPORT_33_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_33_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_33_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_34_en & debug_microOp_cf_loadWaitBit_MPORT_34_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_34_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_34_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_35_en & debug_microOp_cf_loadWaitBit_MPORT_35_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_35_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_35_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_36_en & debug_microOp_cf_loadWaitBit_MPORT_36_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_36_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_36_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_37_en & debug_microOp_cf_loadWaitBit_MPORT_37_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_37_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_37_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_38_en & debug_microOp_cf_loadWaitBit_MPORT_38_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_38_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_38_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_39_en & debug_microOp_cf_loadWaitBit_MPORT_39_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_39_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_39_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_40_en & debug_microOp_cf_loadWaitBit_MPORT_40_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_40_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_40_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_41_en & debug_microOp_cf_loadWaitBit_MPORT_41_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_41_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_41_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_42_en & debug_microOp_cf_loadWaitBit_MPORT_42_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_42_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_42_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_43_en & debug_microOp_cf_loadWaitBit_MPORT_43_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_43_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_43_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_44_en & debug_microOp_cf_loadWaitBit_MPORT_44_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_44_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_44_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_45_en & debug_microOp_cf_loadWaitBit_MPORT_45_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_45_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_45_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_46_en & debug_microOp_cf_loadWaitBit_MPORT_46_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_46_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_46_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_47_en & debug_microOp_cf_loadWaitBit_MPORT_47_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_47_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_47_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_48_en & debug_microOp_cf_loadWaitBit_MPORT_48_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_48_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_48_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_49_en & debug_microOp_cf_loadWaitBit_MPORT_49_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_49_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_49_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_50_en & debug_microOp_cf_loadWaitBit_MPORT_50_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_50_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_50_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_51_en & debug_microOp_cf_loadWaitBit_MPORT_51_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_51_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_51_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_52_en & debug_microOp_cf_loadWaitBit_MPORT_52_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_52_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_52_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_53_en & debug_microOp_cf_loadWaitBit_MPORT_53_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_53_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_53_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_54_en & debug_microOp_cf_loadWaitBit_MPORT_54_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_54_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_54_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_55_en & debug_microOp_cf_loadWaitBit_MPORT_55_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_55_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_55_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_56_en & debug_microOp_cf_loadWaitBit_MPORT_56_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_56_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_56_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_57_en & debug_microOp_cf_loadWaitBit_MPORT_57_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_57_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_57_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_58_en & debug_microOp_cf_loadWaitBit_MPORT_58_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_58_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_58_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_59_en & debug_microOp_cf_loadWaitBit_MPORT_59_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_59_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_59_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_60_en & debug_microOp_cf_loadWaitBit_MPORT_60_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_60_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_60_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_61_en & debug_microOp_cf_loadWaitBit_MPORT_61_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_61_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_61_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_62_en & debug_microOp_cf_loadWaitBit_MPORT_62_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_62_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_62_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_63_en & debug_microOp_cf_loadWaitBit_MPORT_63_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_63_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_63_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_64_en & debug_microOp_cf_loadWaitBit_MPORT_64_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_64_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_64_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_65_en & debug_microOp_cf_loadWaitBit_MPORT_65_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_65_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_65_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_66_en & debug_microOp_cf_loadWaitBit_MPORT_66_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_66_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_66_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_67_en & debug_microOp_cf_loadWaitBit_MPORT_67_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_67_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_67_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_68_en & debug_microOp_cf_loadWaitBit_MPORT_68_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_68_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_68_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_69_en & debug_microOp_cf_loadWaitBit_MPORT_69_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_69_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_69_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_70_en & debug_microOp_cf_loadWaitBit_MPORT_70_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_70_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_70_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_71_en & debug_microOp_cf_loadWaitBit_MPORT_71_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_71_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_71_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_72_en & debug_microOp_cf_loadWaitBit_MPORT_72_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_72_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_72_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_73_en & debug_microOp_cf_loadWaitBit_MPORT_73_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_73_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_73_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_74_en & debug_microOp_cf_loadWaitBit_MPORT_74_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_74_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_74_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_75_en & debug_microOp_cf_loadWaitBit_MPORT_75_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_75_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_75_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_76_en & debug_microOp_cf_loadWaitBit_MPORT_76_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_76_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_76_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_77_en & debug_microOp_cf_loadWaitBit_MPORT_77_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_77_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_77_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_78_en & debug_microOp_cf_loadWaitBit_MPORT_78_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_78_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_78_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_79_en & debug_microOp_cf_loadWaitBit_MPORT_79_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_79_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_79_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_80_en & debug_microOp_cf_loadWaitBit_MPORT_80_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_80_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_80_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_81_en & debug_microOp_cf_loadWaitBit_MPORT_81_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_81_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_81_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_82_en & debug_microOp_cf_loadWaitBit_MPORT_82_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_82_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_82_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_83_en & debug_microOp_cf_loadWaitBit_MPORT_83_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_83_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_83_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_84_en & debug_microOp_cf_loadWaitBit_MPORT_84_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_84_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_84_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_85_en & debug_microOp_cf_loadWaitBit_MPORT_85_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_85_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_85_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_86_en & debug_microOp_cf_loadWaitBit_MPORT_86_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_86_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_86_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_cf_loadWaitBit_MPORT_87_en & debug_microOp_cf_loadWaitBit_MPORT_87_mask) begin
      debug_microOp_cf_loadWaitBit[debug_microOp_cf_loadWaitBit_MPORT_87_addr] <=
        debug_microOp_cf_loadWaitBit_MPORT_87_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_en & debug_microOp_ctrl_isMove_MPORT_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_addr] <= debug_microOp_ctrl_isMove_MPORT_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_1_en & debug_microOp_ctrl_isMove_MPORT_1_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_1_addr] <= debug_microOp_ctrl_isMove_MPORT_1_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_2_en & debug_microOp_ctrl_isMove_MPORT_2_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_2_addr] <= debug_microOp_ctrl_isMove_MPORT_2_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_3_en & debug_microOp_ctrl_isMove_MPORT_3_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_3_addr] <= debug_microOp_ctrl_isMove_MPORT_3_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_4_en & debug_microOp_ctrl_isMove_MPORT_4_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_4_addr] <= debug_microOp_ctrl_isMove_MPORT_4_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_5_en & debug_microOp_ctrl_isMove_MPORT_5_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_5_addr] <= debug_microOp_ctrl_isMove_MPORT_5_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_6_en & debug_microOp_ctrl_isMove_MPORT_6_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_6_addr] <= debug_microOp_ctrl_isMove_MPORT_6_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_7_en & debug_microOp_ctrl_isMove_MPORT_7_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_7_addr] <= debug_microOp_ctrl_isMove_MPORT_7_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_8_en & debug_microOp_ctrl_isMove_MPORT_8_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_8_addr] <= debug_microOp_ctrl_isMove_MPORT_8_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_9_en & debug_microOp_ctrl_isMove_MPORT_9_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_9_addr] <= debug_microOp_ctrl_isMove_MPORT_9_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_10_en & debug_microOp_ctrl_isMove_MPORT_10_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_10_addr] <= debug_microOp_ctrl_isMove_MPORT_10_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_11_en & debug_microOp_ctrl_isMove_MPORT_11_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_11_addr] <= debug_microOp_ctrl_isMove_MPORT_11_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_12_en & debug_microOp_ctrl_isMove_MPORT_12_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_12_addr] <= debug_microOp_ctrl_isMove_MPORT_12_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_13_en & debug_microOp_ctrl_isMove_MPORT_13_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_13_addr] <= debug_microOp_ctrl_isMove_MPORT_13_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_14_en & debug_microOp_ctrl_isMove_MPORT_14_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_14_addr] <= debug_microOp_ctrl_isMove_MPORT_14_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_15_en & debug_microOp_ctrl_isMove_MPORT_15_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_15_addr] <= debug_microOp_ctrl_isMove_MPORT_15_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_16_en & debug_microOp_ctrl_isMove_MPORT_16_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_16_addr] <= debug_microOp_ctrl_isMove_MPORT_16_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_17_en & debug_microOp_ctrl_isMove_MPORT_17_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_17_addr] <= debug_microOp_ctrl_isMove_MPORT_17_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_18_en & debug_microOp_ctrl_isMove_MPORT_18_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_18_addr] <= debug_microOp_ctrl_isMove_MPORT_18_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_19_en & debug_microOp_ctrl_isMove_MPORT_19_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_19_addr] <= debug_microOp_ctrl_isMove_MPORT_19_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_20_en & debug_microOp_ctrl_isMove_MPORT_20_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_20_addr] <= debug_microOp_ctrl_isMove_MPORT_20_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_21_en & debug_microOp_ctrl_isMove_MPORT_21_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_21_addr] <= debug_microOp_ctrl_isMove_MPORT_21_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_22_en & debug_microOp_ctrl_isMove_MPORT_22_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_22_addr] <= debug_microOp_ctrl_isMove_MPORT_22_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_23_en & debug_microOp_ctrl_isMove_MPORT_23_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_23_addr] <= debug_microOp_ctrl_isMove_MPORT_23_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_24_en & debug_microOp_ctrl_isMove_MPORT_24_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_24_addr] <= debug_microOp_ctrl_isMove_MPORT_24_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_25_en & debug_microOp_ctrl_isMove_MPORT_25_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_25_addr] <= debug_microOp_ctrl_isMove_MPORT_25_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_26_en & debug_microOp_ctrl_isMove_MPORT_26_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_26_addr] <= debug_microOp_ctrl_isMove_MPORT_26_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_27_en & debug_microOp_ctrl_isMove_MPORT_27_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_27_addr] <= debug_microOp_ctrl_isMove_MPORT_27_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_28_en & debug_microOp_ctrl_isMove_MPORT_28_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_28_addr] <= debug_microOp_ctrl_isMove_MPORT_28_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_29_en & debug_microOp_ctrl_isMove_MPORT_29_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_29_addr] <= debug_microOp_ctrl_isMove_MPORT_29_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_30_en & debug_microOp_ctrl_isMove_MPORT_30_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_30_addr] <= debug_microOp_ctrl_isMove_MPORT_30_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_31_en & debug_microOp_ctrl_isMove_MPORT_31_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_31_addr] <= debug_microOp_ctrl_isMove_MPORT_31_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_32_en & debug_microOp_ctrl_isMove_MPORT_32_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_32_addr] <= debug_microOp_ctrl_isMove_MPORT_32_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_33_en & debug_microOp_ctrl_isMove_MPORT_33_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_33_addr] <= debug_microOp_ctrl_isMove_MPORT_33_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_34_en & debug_microOp_ctrl_isMove_MPORT_34_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_34_addr] <= debug_microOp_ctrl_isMove_MPORT_34_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_35_en & debug_microOp_ctrl_isMove_MPORT_35_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_35_addr] <= debug_microOp_ctrl_isMove_MPORT_35_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_36_en & debug_microOp_ctrl_isMove_MPORT_36_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_36_addr] <= debug_microOp_ctrl_isMove_MPORT_36_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_37_en & debug_microOp_ctrl_isMove_MPORT_37_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_37_addr] <= debug_microOp_ctrl_isMove_MPORT_37_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_38_en & debug_microOp_ctrl_isMove_MPORT_38_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_38_addr] <= debug_microOp_ctrl_isMove_MPORT_38_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_39_en & debug_microOp_ctrl_isMove_MPORT_39_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_39_addr] <= debug_microOp_ctrl_isMove_MPORT_39_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_40_en & debug_microOp_ctrl_isMove_MPORT_40_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_40_addr] <= debug_microOp_ctrl_isMove_MPORT_40_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_41_en & debug_microOp_ctrl_isMove_MPORT_41_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_41_addr] <= debug_microOp_ctrl_isMove_MPORT_41_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_42_en & debug_microOp_ctrl_isMove_MPORT_42_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_42_addr] <= debug_microOp_ctrl_isMove_MPORT_42_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_43_en & debug_microOp_ctrl_isMove_MPORT_43_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_43_addr] <= debug_microOp_ctrl_isMove_MPORT_43_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_44_en & debug_microOp_ctrl_isMove_MPORT_44_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_44_addr] <= debug_microOp_ctrl_isMove_MPORT_44_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_45_en & debug_microOp_ctrl_isMove_MPORT_45_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_45_addr] <= debug_microOp_ctrl_isMove_MPORT_45_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_46_en & debug_microOp_ctrl_isMove_MPORT_46_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_46_addr] <= debug_microOp_ctrl_isMove_MPORT_46_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_47_en & debug_microOp_ctrl_isMove_MPORT_47_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_47_addr] <= debug_microOp_ctrl_isMove_MPORT_47_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_48_en & debug_microOp_ctrl_isMove_MPORT_48_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_48_addr] <= debug_microOp_ctrl_isMove_MPORT_48_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_49_en & debug_microOp_ctrl_isMove_MPORT_49_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_49_addr] <= debug_microOp_ctrl_isMove_MPORT_49_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_50_en & debug_microOp_ctrl_isMove_MPORT_50_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_50_addr] <= debug_microOp_ctrl_isMove_MPORT_50_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_51_en & debug_microOp_ctrl_isMove_MPORT_51_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_51_addr] <= debug_microOp_ctrl_isMove_MPORT_51_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_52_en & debug_microOp_ctrl_isMove_MPORT_52_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_52_addr] <= debug_microOp_ctrl_isMove_MPORT_52_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_53_en & debug_microOp_ctrl_isMove_MPORT_53_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_53_addr] <= debug_microOp_ctrl_isMove_MPORT_53_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_54_en & debug_microOp_ctrl_isMove_MPORT_54_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_54_addr] <= debug_microOp_ctrl_isMove_MPORT_54_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_55_en & debug_microOp_ctrl_isMove_MPORT_55_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_55_addr] <= debug_microOp_ctrl_isMove_MPORT_55_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_56_en & debug_microOp_ctrl_isMove_MPORT_56_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_56_addr] <= debug_microOp_ctrl_isMove_MPORT_56_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_57_en & debug_microOp_ctrl_isMove_MPORT_57_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_57_addr] <= debug_microOp_ctrl_isMove_MPORT_57_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_58_en & debug_microOp_ctrl_isMove_MPORT_58_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_58_addr] <= debug_microOp_ctrl_isMove_MPORT_58_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_59_en & debug_microOp_ctrl_isMove_MPORT_59_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_59_addr] <= debug_microOp_ctrl_isMove_MPORT_59_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_60_en & debug_microOp_ctrl_isMove_MPORT_60_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_60_addr] <= debug_microOp_ctrl_isMove_MPORT_60_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_61_en & debug_microOp_ctrl_isMove_MPORT_61_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_61_addr] <= debug_microOp_ctrl_isMove_MPORT_61_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_62_en & debug_microOp_ctrl_isMove_MPORT_62_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_62_addr] <= debug_microOp_ctrl_isMove_MPORT_62_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_63_en & debug_microOp_ctrl_isMove_MPORT_63_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_63_addr] <= debug_microOp_ctrl_isMove_MPORT_63_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_64_en & debug_microOp_ctrl_isMove_MPORT_64_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_64_addr] <= debug_microOp_ctrl_isMove_MPORT_64_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_65_en & debug_microOp_ctrl_isMove_MPORT_65_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_65_addr] <= debug_microOp_ctrl_isMove_MPORT_65_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_66_en & debug_microOp_ctrl_isMove_MPORT_66_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_66_addr] <= debug_microOp_ctrl_isMove_MPORT_66_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_67_en & debug_microOp_ctrl_isMove_MPORT_67_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_67_addr] <= debug_microOp_ctrl_isMove_MPORT_67_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_68_en & debug_microOp_ctrl_isMove_MPORT_68_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_68_addr] <= debug_microOp_ctrl_isMove_MPORT_68_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_69_en & debug_microOp_ctrl_isMove_MPORT_69_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_69_addr] <= debug_microOp_ctrl_isMove_MPORT_69_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_70_en & debug_microOp_ctrl_isMove_MPORT_70_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_70_addr] <= debug_microOp_ctrl_isMove_MPORT_70_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_71_en & debug_microOp_ctrl_isMove_MPORT_71_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_71_addr] <= debug_microOp_ctrl_isMove_MPORT_71_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_72_en & debug_microOp_ctrl_isMove_MPORT_72_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_72_addr] <= debug_microOp_ctrl_isMove_MPORT_72_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_73_en & debug_microOp_ctrl_isMove_MPORT_73_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_73_addr] <= debug_microOp_ctrl_isMove_MPORT_73_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_74_en & debug_microOp_ctrl_isMove_MPORT_74_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_74_addr] <= debug_microOp_ctrl_isMove_MPORT_74_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_75_en & debug_microOp_ctrl_isMove_MPORT_75_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_75_addr] <= debug_microOp_ctrl_isMove_MPORT_75_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_76_en & debug_microOp_ctrl_isMove_MPORT_76_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_76_addr] <= debug_microOp_ctrl_isMove_MPORT_76_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_77_en & debug_microOp_ctrl_isMove_MPORT_77_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_77_addr] <= debug_microOp_ctrl_isMove_MPORT_77_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_78_en & debug_microOp_ctrl_isMove_MPORT_78_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_78_addr] <= debug_microOp_ctrl_isMove_MPORT_78_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_79_en & debug_microOp_ctrl_isMove_MPORT_79_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_79_addr] <= debug_microOp_ctrl_isMove_MPORT_79_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_80_en & debug_microOp_ctrl_isMove_MPORT_80_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_80_addr] <= debug_microOp_ctrl_isMove_MPORT_80_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_81_en & debug_microOp_ctrl_isMove_MPORT_81_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_81_addr] <= debug_microOp_ctrl_isMove_MPORT_81_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_82_en & debug_microOp_ctrl_isMove_MPORT_82_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_82_addr] <= debug_microOp_ctrl_isMove_MPORT_82_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_83_en & debug_microOp_ctrl_isMove_MPORT_83_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_83_addr] <= debug_microOp_ctrl_isMove_MPORT_83_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_84_en & debug_microOp_ctrl_isMove_MPORT_84_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_84_addr] <= debug_microOp_ctrl_isMove_MPORT_84_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_85_en & debug_microOp_ctrl_isMove_MPORT_85_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_85_addr] <= debug_microOp_ctrl_isMove_MPORT_85_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_86_en & debug_microOp_ctrl_isMove_MPORT_86_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_86_addr] <= debug_microOp_ctrl_isMove_MPORT_86_data; // @[Rob.scala 440:26]
    end
    if (debug_microOp_ctrl_isMove_MPORT_87_en & debug_microOp_ctrl_isMove_MPORT_87_mask) begin
      debug_microOp_ctrl_isMove[debug_microOp_ctrl_isMove_MPORT_87_addr] <= debug_microOp_ctrl_isMove_MPORT_87_data; // @[Rob.scala 440:26]
    end
    if (dt_eliminatedMove_MPORT_305_en & dt_eliminatedMove_MPORT_305_mask) begin
      dt_eliminatedMove[dt_eliminatedMove_MPORT_305_addr] <= dt_eliminatedMove_MPORT_305_data; // @[Rob.scala 1212:32]
    end
    if (dt_eliminatedMove_MPORT_307_en & dt_eliminatedMove_MPORT_307_mask) begin
      dt_eliminatedMove[dt_eliminatedMove_MPORT_307_addr] <= dt_eliminatedMove_MPORT_307_data; // @[Rob.scala 1212:32]
    end
    if (dt_isRVC_MPORT_306_en & dt_isRVC_MPORT_306_mask) begin
      dt_isRVC[dt_isRVC_MPORT_306_addr] <= dt_isRVC_MPORT_306_data; // @[Rob.scala 1213:23]
    end
    if (dt_isRVC_MPORT_308_en & dt_isRVC_MPORT_308_mask) begin
      dt_isRVC[dt_isRVC_MPORT_308_addr] <= dt_isRVC_MPORT_308_data; // @[Rob.scala 1213:23]
    end
    if (dt_isXSTrap_MPORT_309_en & dt_isXSTrap_MPORT_309_mask) begin
      dt_isXSTrap[dt_isXSTrap_MPORT_309_addr] <= dt_isXSTrap_MPORT_309_data; // @[Rob.scala 1290:26]
    end
    if (dt_isXSTrap_MPORT_310_en & dt_isXSTrap_MPORT_310_mask) begin
      dt_isXSTrap[dt_isXSTrap_MPORT_310_addr] <= dt_isXSTrap_MPORT_310_data; // @[Rob.scala 1290:26]
    end
    if (io_redirect_valid) begin // @[Rob.scala 797:28]
      walkPtrVec_0_flag <= deqPtrGenModule_io_next_out_0_flag;
    end else if (state) begin // @[Rob.scala 799:8]
      walkPtrVec_0_flag <= walkPtrVec_next_new_ptr_flag;
    end
    if (io_redirect_valid) begin // @[Rob.scala 797:28]
      walkPtrVec_0_value <= deqPtrGenModule_io_next_out_0_value;
    end else if (state) begin // @[Rob.scala 799:8]
      walkPtrVec_0_value <= walkPtrVec_next_new_ptr_value;
    end
    if (io_redirect_valid) begin // @[Rob.scala 797:28]
      walkPtrVec_1_flag <= deqPtrGenModule_io_next_out_1_flag;
    end else if (state) begin // @[Rob.scala 799:8]
      walkPtrVec_1_flag <= walkPtrVec_next_new_ptr_1_flag;
    end
    if (io_redirect_valid) begin // @[Rob.scala 797:28]
      walkPtrVec_1_value <= deqPtrGenModule_io_next_out_1_value;
    end else if (state) begin // @[Rob.scala 799:8]
      walkPtrVec_1_value <= walkPtrVec_next_new_ptr_1_value;
    end
    REG <= hasWFI; // @[Rob.scala 508:33]
    REG_1 <= io_csr_wfiEvent; // @[Rob.scala 512:24]
    REG_2 <= REG_1; // @[Rob.scala 512:16]
    io_enq_isEmpty_REG <= isEmpty & ~(|_io_enq_isEmpty_T); // @[Rob.scala 566:39]
    REG_3 <= io_lsq_isMMIO_0; // @[Rob.scala 606:18]
    REG_4 <= io_lsq_uop_0_robIdx_value; // @[Rob.scala 607:19]
    REG_5 <= io_lsq_isMMIO_1; // @[Rob.scala 606:18]
    REG_6 <= io_lsq_uop_1_robIdx_value; // @[Rob.scala 607:19]
    intrBitSetReg <= io_csr_intrBitSet; // @[Rob.scala 617:30]
    lastCycleFlush <= io_flushOut_valid; // @[Rob.scala 634:31]
    io_exception_valid_REG <= _io_flushOut_valid_T_1 & _io_flushOut_valid_T_2 & _io_flushOut_valid_T_5; // @[Rob.scala 648:102]
    if (exceptionHappen) begin // @[Reg.scala 17:18]
      io_exception_bits_uop_ctrl_commitType_r <= dispatchData_io_rdata_0_commitType; // @[Reg.scala 17:22]
    end
    if (exceptionHappen) begin // @[Reg.scala 17:18]
      r_0 <= exceptionGen_io_state_bits_exceptionVec_0; // @[Reg.scala 17:22]
    end
    if (exceptionHappen) begin // @[Reg.scala 17:18]
      r_1 <= exceptionGen_io_state_bits_exceptionVec_1; // @[Reg.scala 17:22]
    end
    if (exceptionHappen) begin // @[Reg.scala 17:18]
      r_2 <= exceptionGen_io_state_bits_exceptionVec_2; // @[Reg.scala 17:22]
    end
    if (exceptionHappen) begin // @[Reg.scala 17:18]
      r_3 <= exceptionGen_io_state_bits_exceptionVec_3; // @[Reg.scala 17:22]
    end
    if (exceptionHappen) begin // @[Reg.scala 17:18]
      r_4 <= exceptionGen_io_state_bits_exceptionVec_4; // @[Reg.scala 17:22]
    end
    if (exceptionHappen) begin // @[Reg.scala 17:18]
      r_5 <= exceptionGen_io_state_bits_exceptionVec_5; // @[Reg.scala 17:22]
    end
    if (exceptionHappen) begin // @[Reg.scala 17:18]
      r_6 <= exceptionGen_io_state_bits_exceptionVec_6; // @[Reg.scala 17:22]
    end
    if (exceptionHappen) begin // @[Reg.scala 17:18]
      r_7 <= exceptionGen_io_state_bits_exceptionVec_7; // @[Reg.scala 17:22]
    end
    if (exceptionHappen) begin // @[Reg.scala 17:18]
      r_8 <= exceptionGen_io_state_bits_exceptionVec_8; // @[Reg.scala 17:22]
    end
    if (exceptionHappen) begin // @[Reg.scala 17:18]
      r_9 <= exceptionGen_io_state_bits_exceptionVec_9; // @[Reg.scala 17:22]
    end
    if (exceptionHappen) begin // @[Reg.scala 17:18]
      r_11 <= exceptionGen_io_state_bits_exceptionVec_11; // @[Reg.scala 17:22]
    end
    if (exceptionHappen) begin // @[Reg.scala 17:18]
      r_12 <= exceptionGen_io_state_bits_exceptionVec_12; // @[Reg.scala 17:22]
    end
    if (exceptionHappen) begin // @[Reg.scala 17:18]
      r_13 <= exceptionGen_io_state_bits_exceptionVec_13; // @[Reg.scala 17:22]
    end
    if (exceptionHappen) begin // @[Reg.scala 17:18]
      r_15 <= exceptionGen_io_state_bits_exceptionVec_15; // @[Reg.scala 17:22]
    end
    if (exceptionHappen) begin // @[Reg.scala 17:18]
      io_exception_bits_uop_ctrl_singleStep_r <= exceptionGen_io_state_bits_singleStep; // @[Reg.scala 17:22]
    end
    if (exceptionHappen) begin // @[Reg.scala 17:18]
      io_exception_bits_uop_cf_crossPageIPFFix_r <= exceptionGen_io_state_bits_crossPageIPFFix; // @[Reg.scala 17:22]
    end
    if (exceptionHappen) begin // @[Reg.scala 17:18]
      io_exception_bits_isInterrupt_r <= intrEnable; // @[Reg.scala 17:22]
    end
    if (exceptionHappen) begin // @[Reg.scala 17:18]
      io_exception_bits_uop_cf_trigger_rfrontendHit_0 <= exceptionGen_io_state_bits_trigger_frontendHit_0; // @[Reg.scala 17:22]
    end
    if (exceptionHappen) begin // @[Reg.scala 17:18]
      io_exception_bits_uop_cf_trigger_rfrontendHit_1 <= exceptionGen_io_state_bits_trigger_frontendHit_1; // @[Reg.scala 17:22]
    end
    if (exceptionHappen) begin // @[Reg.scala 17:18]
      io_exception_bits_uop_cf_trigger_rfrontendHit_2 <= exceptionGen_io_state_bits_trigger_frontendHit_2; // @[Reg.scala 17:22]
    end
    if (exceptionHappen) begin // @[Reg.scala 17:18]
      io_exception_bits_uop_cf_trigger_rfrontendHit_3 <= exceptionGen_io_state_bits_trigger_frontendHit_3; // @[Reg.scala 17:22]
    end
    if (exceptionHappen) begin // @[Reg.scala 17:18]
      io_exception_bits_uop_cf_trigger_rbackendHit_0 <= exceptionGen_io_state_bits_trigger_backendHit_0; // @[Reg.scala 17:22]
    end
    if (exceptionHappen) begin // @[Reg.scala 17:18]
      io_exception_bits_uop_cf_trigger_rbackendHit_1 <= exceptionGen_io_state_bits_trigger_backendHit_1; // @[Reg.scala 17:22]
    end
    if (exceptionHappen) begin // @[Reg.scala 17:18]
      io_exception_bits_uop_cf_trigger_rbackendHit_2 <= exceptionGen_io_state_bits_trigger_backendHit_2; // @[Reg.scala 17:22]
    end
    if (exceptionHappen) begin // @[Reg.scala 17:18]
      io_exception_bits_uop_cf_trigger_rbackendHit_3 <= exceptionGen_io_state_bits_trigger_backendHit_3; // @[Reg.scala 17:22]
    end
    if (exceptionHappen) begin // @[Reg.scala 17:18]
      io_exception_bits_uop_cf_trigger_rbackendHit_4 <= exceptionGen_io_state_bits_trigger_backendHit_4; // @[Reg.scala 17:22]
    end
    if (exceptionHappen) begin // @[Reg.scala 17:18]
      io_exception_bits_uop_cf_trigger_rbackendHit_5 <= exceptionGen_io_state_bits_trigger_backendHit_5; // @[Reg.scala 17:22]
    end
    walkCounter <= _GEN_5110[5:0];
    if (misPredWb) begin // @[Rob.scala 693:29]
      misPredBlockCounter <= 3'h7;
    end else begin
      misPredBlockCounter <= _misPredBlockCounter_T;
    end
    io_csr_fflags_REG_valid <= io_commits_isCommit & |_fflags_valid_T; // @[Rob.scala 681:39]
    io_csr_fflags_REG_bits <= _fflags_bits_T | _fflags_bits_T_1; // @[Rob.scala 684:14]
    io_csr_dirty_fs_REG <= io_commits_isCommit & |_dirty_fs_T; // @[Rob.scala 685:38]
    if (io_commits_isCommit) begin // @[Rob.scala 753:32]
      io_lsq_scommit_REG <= _io_lsq_scommit_T;
    end else begin
      io_lsq_scommit_REG <= 2'h0;
    end
    io_lsq_pendingld_REG <= io_commits_isCommit & _ldCommitVec_T & commit_v_0 & _GEN_5108; // @[Rob.scala 755:127]
    io_lsq_pendingst_REG <= io_commits_isCommit & _stCommitVec_T & commit_v_0; // @[Rob.scala 756:105]
    io_lsq_commit_REG <= io_commits_isCommit & io_commits_commitValid_0; // @[Rob.scala 757:48]
    if (io_redirect_valid) begin // @[Rob.scala 858:27]
      if (io_redirect_bits_level) begin // @[Rob.scala 864:26]
        redirectHeadVec_0_flag <= redirectHeadVec_0_new_ptr_1_flag;
      end else begin
        redirectHeadVec_0_flag <= redirectHeadVec_0_new_ptr_2_flag;
      end
    end else if (redirectState) begin // @[Rob.scala 847:40]
      redirectHeadVec_0_flag <= redirectHeadVec_0_new_ptr_flag; // @[Rob.scala 848:58]
    end
    if (io_redirect_valid) begin // @[Rob.scala 858:27]
      if (io_redirect_bits_level) begin // @[Rob.scala 864:26]
        redirectHeadVec_0_value <= redirectHeadVec_0_new_ptr_1_value;
      end else begin
        redirectHeadVec_0_value <= redirectHeadVec_0_new_ptr_2_value;
      end
    end else if (redirectState) begin // @[Rob.scala 847:40]
      redirectHeadVec_0_value <= redirectHeadVec_0_new_ptr_value; // @[Rob.scala 848:58]
    end
    if (io_redirect_valid) begin // @[Rob.scala 858:27]
      if (io_redirect_bits_level) begin // @[Rob.scala 864:26]
        redirectHeadVec_1_flag <= redirectHeadVec_0_new_ptr_2_flag;
      end else begin
        redirectHeadVec_1_flag <= redirectHeadVec_1_new_ptr_2_flag;
      end
    end else if (redirectState) begin // @[Rob.scala 847:40]
      redirectHeadVec_1_flag <= redirectHeadVec_1_new_ptr_flag; // @[Rob.scala 848:58]
    end
    if (io_redirect_valid) begin // @[Rob.scala 858:27]
      if (io_redirect_bits_level) begin // @[Rob.scala 864:26]
        redirectHeadVec_1_value <= redirectHeadVec_0_new_ptr_2_value;
      end else begin
        redirectHeadVec_1_value <= redirectHeadVec_1_new_ptr_2_value;
      end
    end else if (redirectState) begin // @[Rob.scala 847:40]
      redirectHeadVec_1_value <= redirectHeadVec_1_new_ptr_value; // @[Rob.scala 848:58]
    end
    if (io_redirect_valid) begin // @[Rob.scala 858:27]
      if (~redirectState) begin // @[Rob.scala 860:42]
        redirectTail_flag <= enqPtrVec_0_flag; // @[Rob.scala 861:20]
      end
    end
    if (io_redirect_valid) begin // @[Rob.scala 858:27]
      if (~redirectState) begin // @[Rob.scala 860:42]
        redirectTail_value <= enqPtrVec_0_value; // @[Rob.scala 861:20]
      end
    end
    REG_7 <= io_writeback_1_9_valid; // @[Rob.scala 918:17]
    REG_8 <= io_writeback_1_9_bits_uop_robIdx_value; // @[Rob.scala 919:37]
    REG_9 <= io_writeback_1_10_valid; // @[Rob.scala 918:17]
    REG_10 <= io_writeback_1_10_bits_uop_robIdx_value; // @[Rob.scala 919:37]
    REG_11 <= io_enq_req_0_valid & io_enq_canAccept; // @[Rob.scala 519:51]
    REG_12 <= enqPtrGenModule_io_out_0_value; // @[Rob.scala 447:23 791:13]
    REG_13 <= ~_allow_interrupts_T_3; // @[Rob.scala 942:30]
    REG_14 <= io_enq_req_1_valid & io_enq_canAccept; // @[Rob.scala 519:51]
    if (io_enq_needAlloc_0) begin // @[Rob.scala 516:31]
      REG_15 <= enqPtrVec_1_value; // @[Rob.scala 516:31]
    end else begin
      REG_15 <= enqPtrVec_0_value;
    end
    REG_16 <= ~_allow_interrupts_T_7; // @[Rob.scala 942:30]
    fuseCommitCnt_REG <= io_commits_commitValid_0 & io_commits_info_0_commitType[2]; // @[Rob.scala 1019:106]
    fuseCommitCnt_REG_1 <= io_commits_commitValid_1 & io_commits_info_1_commitType[2]; // @[Rob.scala 1019:106]
    trueCommitCnt_REG <= io_commits_commitValid_0 + io_commits_commitValid_1; // @[Bitwise.scala 48:55]
    retireCounter_REG <= io_commits_isCommit; // @[Rob.scala 1021:34]
    if (io_writeback_1_8_valid) begin // @[Rob.scala 1222:23]
      if (5'h0 == io_writeback_1_8_bits_uop_robIdx_value) begin // @[Rob.scala 1224:28]
        dt_exuDebug_0_isMMIO <= io_writeback_1_8_bits_debug_isMMIO; // @[Rob.scala 1224:28]
      end else begin
        dt_exuDebug_0_isMMIO <= _GEN_10635;
      end
    end else begin
      dt_exuDebug_0_isMMIO <= _GEN_10635;
    end
    if (io_writeback_1_8_valid) begin // @[Rob.scala 1222:23]
      if (5'h0 == io_writeback_1_8_bits_uop_robIdx_value) begin // @[Rob.scala 1224:28]
        dt_exuDebug_0_isPerfCnt <= io_writeback_1_8_bits_debug_isPerfCnt; // @[Rob.scala 1224:28]
      end else begin
        dt_exuDebug_0_isPerfCnt <= _GEN_10667;
      end
    end else begin
      dt_exuDebug_0_isPerfCnt <= _GEN_10667;
    end
    if (io_writeback_1_8_valid) begin // @[Rob.scala 1222:23]
      if (5'h1 == io_writeback_1_8_bits_uop_robIdx_value) begin // @[Rob.scala 1224:28]
        dt_exuDebug_1_isMMIO <= io_writeback_1_8_bits_debug_isMMIO; // @[Rob.scala 1224:28]
      end else begin
        dt_exuDebug_1_isMMIO <= _GEN_10636;
      end
    end else begin
      dt_exuDebug_1_isMMIO <= _GEN_10636;
    end
    if (io_writeback_1_8_valid) begin // @[Rob.scala 1222:23]
      if (5'h1 == io_writeback_1_8_bits_uop_robIdx_value) begin // @[Rob.scala 1224:28]
        dt_exuDebug_1_isPerfCnt <= io_writeback_1_8_bits_debug_isPerfCnt; // @[Rob.scala 1224:28]
      end else begin
        dt_exuDebug_1_isPerfCnt <= _GEN_10668;
      end
    end else begin
      dt_exuDebug_1_isPerfCnt <= _GEN_10668;
    end
    if (io_writeback_1_8_valid) begin // @[Rob.scala 1222:23]
      if (5'h2 == io_writeback_1_8_bits_uop_robIdx_value) begin // @[Rob.scala 1224:28]
        dt_exuDebug_2_isMMIO <= io_writeback_1_8_bits_debug_isMMIO; // @[Rob.scala 1224:28]
      end else begin
        dt_exuDebug_2_isMMIO <= _GEN_10637;
      end
    end else begin
      dt_exuDebug_2_isMMIO <= _GEN_10637;
    end
    if (io_writeback_1_8_valid) begin // @[Rob.scala 1222:23]
      if (5'h2 == io_writeback_1_8_bits_uop_robIdx_value) begin // @[Rob.scala 1224:28]
        dt_exuDebug_2_isPerfCnt <= io_writeback_1_8_bits_debug_isPerfCnt; // @[Rob.scala 1224:28]
      end else begin
        dt_exuDebug_2_isPerfCnt <= _GEN_10669;
      end
    end else begin
      dt_exuDebug_2_isPerfCnt <= _GEN_10669;
    end
    if (io_writeback_1_8_valid) begin // @[Rob.scala 1222:23]
      if (5'h3 == io_writeback_1_8_bits_uop_robIdx_value) begin // @[Rob.scala 1224:28]
        dt_exuDebug_3_isMMIO <= io_writeback_1_8_bits_debug_isMMIO; // @[Rob.scala 1224:28]
      end else begin
        dt_exuDebug_3_isMMIO <= _GEN_10638;
      end
    end else begin
      dt_exuDebug_3_isMMIO <= _GEN_10638;
    end
    if (io_writeback_1_8_valid) begin // @[Rob.scala 1222:23]
      if (5'h3 == io_writeback_1_8_bits_uop_robIdx_value) begin // @[Rob.scala 1224:28]
        dt_exuDebug_3_isPerfCnt <= io_writeback_1_8_bits_debug_isPerfCnt; // @[Rob.scala 1224:28]
      end else begin
        dt_exuDebug_3_isPerfCnt <= _GEN_10670;
      end
    end else begin
      dt_exuDebug_3_isPerfCnt <= _GEN_10670;
    end
    if (io_writeback_1_8_valid) begin // @[Rob.scala 1222:23]
      if (5'h4 == io_writeback_1_8_bits_uop_robIdx_value) begin // @[Rob.scala 1224:28]
        dt_exuDebug_4_isMMIO <= io_writeback_1_8_bits_debug_isMMIO; // @[Rob.scala 1224:28]
      end else begin
        dt_exuDebug_4_isMMIO <= _GEN_10639;
      end
    end else begin
      dt_exuDebug_4_isMMIO <= _GEN_10639;
    end
    if (io_writeback_1_8_valid) begin // @[Rob.scala 1222:23]
      if (5'h4 == io_writeback_1_8_bits_uop_robIdx_value) begin // @[Rob.scala 1224:28]
        dt_exuDebug_4_isPerfCnt <= io_writeback_1_8_bits_debug_isPerfCnt; // @[Rob.scala 1224:28]
      end else begin
        dt_exuDebug_4_isPerfCnt <= _GEN_10671;
      end
    end else begin
      dt_exuDebug_4_isPerfCnt <= _GEN_10671;
    end
    if (io_writeback_1_8_valid) begin // @[Rob.scala 1222:23]
      if (5'h5 == io_writeback_1_8_bits_uop_robIdx_value) begin // @[Rob.scala 1224:28]
        dt_exuDebug_5_isMMIO <= io_writeback_1_8_bits_debug_isMMIO; // @[Rob.scala 1224:28]
      end else begin
        dt_exuDebug_5_isMMIO <= _GEN_10640;
      end
    end else begin
      dt_exuDebug_5_isMMIO <= _GEN_10640;
    end
    if (io_writeback_1_8_valid) begin // @[Rob.scala 1222:23]
      if (5'h5 == io_writeback_1_8_bits_uop_robIdx_value) begin // @[Rob.scala 1224:28]
        dt_exuDebug_5_isPerfCnt <= io_writeback_1_8_bits_debug_isPerfCnt; // @[Rob.scala 1224:28]
      end else begin
        dt_exuDebug_5_isPerfCnt <= _GEN_10672;
      end
    end else begin
      dt_exuDebug_5_isPerfCnt <= _GEN_10672;
    end
    if (io_writeback_1_8_valid) begin // @[Rob.scala 1222:23]
      if (5'h6 == io_writeback_1_8_bits_uop_robIdx_value) begin // @[Rob.scala 1224:28]
        dt_exuDebug_6_isMMIO <= io_writeback_1_8_bits_debug_isMMIO; // @[Rob.scala 1224:28]
      end else begin
        dt_exuDebug_6_isMMIO <= _GEN_10641;
      end
    end else begin
      dt_exuDebug_6_isMMIO <= _GEN_10641;
    end
    if (io_writeback_1_8_valid) begin // @[Rob.scala 1222:23]
      if (5'h6 == io_writeback_1_8_bits_uop_robIdx_value) begin // @[Rob.scala 1224:28]
        dt_exuDebug_6_isPerfCnt <= io_writeback_1_8_bits_debug_isPerfCnt; // @[Rob.scala 1224:28]
      end else begin
        dt_exuDebug_6_isPerfCnt <= _GEN_10673;
      end
    end else begin
      dt_exuDebug_6_isPerfCnt <= _GEN_10673;
    end
    if (io_writeback_1_8_valid) begin // @[Rob.scala 1222:23]
      if (5'h7 == io_writeback_1_8_bits_uop_robIdx_value) begin // @[Rob.scala 1224:28]
        dt_exuDebug_7_isMMIO <= io_writeback_1_8_bits_debug_isMMIO; // @[Rob.scala 1224:28]
      end else begin
        dt_exuDebug_7_isMMIO <= _GEN_10642;
      end
    end else begin
      dt_exuDebug_7_isMMIO <= _GEN_10642;
    end
    if (io_writeback_1_8_valid) begin // @[Rob.scala 1222:23]
      if (5'h7 == io_writeback_1_8_bits_uop_robIdx_value) begin // @[Rob.scala 1224:28]
        dt_exuDebug_7_isPerfCnt <= io_writeback_1_8_bits_debug_isPerfCnt; // @[Rob.scala 1224:28]
      end else begin
        dt_exuDebug_7_isPerfCnt <= _GEN_10674;
      end
    end else begin
      dt_exuDebug_7_isPerfCnt <= _GEN_10674;
    end
    if (io_writeback_1_8_valid) begin // @[Rob.scala 1222:23]
      if (5'h8 == io_writeback_1_8_bits_uop_robIdx_value) begin // @[Rob.scala 1224:28]
        dt_exuDebug_8_isMMIO <= io_writeback_1_8_bits_debug_isMMIO; // @[Rob.scala 1224:28]
      end else begin
        dt_exuDebug_8_isMMIO <= _GEN_10643;
      end
    end else begin
      dt_exuDebug_8_isMMIO <= _GEN_10643;
    end
    if (io_writeback_1_8_valid) begin // @[Rob.scala 1222:23]
      if (5'h8 == io_writeback_1_8_bits_uop_robIdx_value) begin // @[Rob.scala 1224:28]
        dt_exuDebug_8_isPerfCnt <= io_writeback_1_8_bits_debug_isPerfCnt; // @[Rob.scala 1224:28]
      end else begin
        dt_exuDebug_8_isPerfCnt <= _GEN_10675;
      end
    end else begin
      dt_exuDebug_8_isPerfCnt <= _GEN_10675;
    end
    if (io_writeback_1_8_valid) begin // @[Rob.scala 1222:23]
      if (5'h9 == io_writeback_1_8_bits_uop_robIdx_value) begin // @[Rob.scala 1224:28]
        dt_exuDebug_9_isMMIO <= io_writeback_1_8_bits_debug_isMMIO; // @[Rob.scala 1224:28]
      end else begin
        dt_exuDebug_9_isMMIO <= _GEN_10644;
      end
    end else begin
      dt_exuDebug_9_isMMIO <= _GEN_10644;
    end
    if (io_writeback_1_8_valid) begin // @[Rob.scala 1222:23]
      if (5'h9 == io_writeback_1_8_bits_uop_robIdx_value) begin // @[Rob.scala 1224:28]
        dt_exuDebug_9_isPerfCnt <= io_writeback_1_8_bits_debug_isPerfCnt; // @[Rob.scala 1224:28]
      end else begin
        dt_exuDebug_9_isPerfCnt <= _GEN_10676;
      end
    end else begin
      dt_exuDebug_9_isPerfCnt <= _GEN_10676;
    end
    if (io_writeback_1_8_valid) begin // @[Rob.scala 1222:23]
      if (5'ha == io_writeback_1_8_bits_uop_robIdx_value) begin // @[Rob.scala 1224:28]
        dt_exuDebug_10_isMMIO <= io_writeback_1_8_bits_debug_isMMIO; // @[Rob.scala 1224:28]
      end else begin
        dt_exuDebug_10_isMMIO <= _GEN_10645;
      end
    end else begin
      dt_exuDebug_10_isMMIO <= _GEN_10645;
    end
    if (io_writeback_1_8_valid) begin // @[Rob.scala 1222:23]
      if (5'ha == io_writeback_1_8_bits_uop_robIdx_value) begin // @[Rob.scala 1224:28]
        dt_exuDebug_10_isPerfCnt <= io_writeback_1_8_bits_debug_isPerfCnt; // @[Rob.scala 1224:28]
      end else begin
        dt_exuDebug_10_isPerfCnt <= _GEN_10677;
      end
    end else begin
      dt_exuDebug_10_isPerfCnt <= _GEN_10677;
    end
    if (io_writeback_1_8_valid) begin // @[Rob.scala 1222:23]
      if (5'hb == io_writeback_1_8_bits_uop_robIdx_value) begin // @[Rob.scala 1224:28]
        dt_exuDebug_11_isMMIO <= io_writeback_1_8_bits_debug_isMMIO; // @[Rob.scala 1224:28]
      end else begin
        dt_exuDebug_11_isMMIO <= _GEN_10646;
      end
    end else begin
      dt_exuDebug_11_isMMIO <= _GEN_10646;
    end
    if (io_writeback_1_8_valid) begin // @[Rob.scala 1222:23]
      if (5'hb == io_writeback_1_8_bits_uop_robIdx_value) begin // @[Rob.scala 1224:28]
        dt_exuDebug_11_isPerfCnt <= io_writeback_1_8_bits_debug_isPerfCnt; // @[Rob.scala 1224:28]
      end else begin
        dt_exuDebug_11_isPerfCnt <= _GEN_10678;
      end
    end else begin
      dt_exuDebug_11_isPerfCnt <= _GEN_10678;
    end
    if (io_writeback_1_8_valid) begin // @[Rob.scala 1222:23]
      if (5'hc == io_writeback_1_8_bits_uop_robIdx_value) begin // @[Rob.scala 1224:28]
        dt_exuDebug_12_isMMIO <= io_writeback_1_8_bits_debug_isMMIO; // @[Rob.scala 1224:28]
      end else begin
        dt_exuDebug_12_isMMIO <= _GEN_10647;
      end
    end else begin
      dt_exuDebug_12_isMMIO <= _GEN_10647;
    end
    if (io_writeback_1_8_valid) begin // @[Rob.scala 1222:23]
      if (5'hc == io_writeback_1_8_bits_uop_robIdx_value) begin // @[Rob.scala 1224:28]
        dt_exuDebug_12_isPerfCnt <= io_writeback_1_8_bits_debug_isPerfCnt; // @[Rob.scala 1224:28]
      end else begin
        dt_exuDebug_12_isPerfCnt <= _GEN_10679;
      end
    end else begin
      dt_exuDebug_12_isPerfCnt <= _GEN_10679;
    end
    if (io_writeback_1_8_valid) begin // @[Rob.scala 1222:23]
      if (5'hd == io_writeback_1_8_bits_uop_robIdx_value) begin // @[Rob.scala 1224:28]
        dt_exuDebug_13_isMMIO <= io_writeback_1_8_bits_debug_isMMIO; // @[Rob.scala 1224:28]
      end else begin
        dt_exuDebug_13_isMMIO <= _GEN_10648;
      end
    end else begin
      dt_exuDebug_13_isMMIO <= _GEN_10648;
    end
    if (io_writeback_1_8_valid) begin // @[Rob.scala 1222:23]
      if (5'hd == io_writeback_1_8_bits_uop_robIdx_value) begin // @[Rob.scala 1224:28]
        dt_exuDebug_13_isPerfCnt <= io_writeback_1_8_bits_debug_isPerfCnt; // @[Rob.scala 1224:28]
      end else begin
        dt_exuDebug_13_isPerfCnt <= _GEN_10680;
      end
    end else begin
      dt_exuDebug_13_isPerfCnt <= _GEN_10680;
    end
    if (io_writeback_1_8_valid) begin // @[Rob.scala 1222:23]
      if (5'he == io_writeback_1_8_bits_uop_robIdx_value) begin // @[Rob.scala 1224:28]
        dt_exuDebug_14_isMMIO <= io_writeback_1_8_bits_debug_isMMIO; // @[Rob.scala 1224:28]
      end else begin
        dt_exuDebug_14_isMMIO <= _GEN_10649;
      end
    end else begin
      dt_exuDebug_14_isMMIO <= _GEN_10649;
    end
    if (io_writeback_1_8_valid) begin // @[Rob.scala 1222:23]
      if (5'he == io_writeback_1_8_bits_uop_robIdx_value) begin // @[Rob.scala 1224:28]
        dt_exuDebug_14_isPerfCnt <= io_writeback_1_8_bits_debug_isPerfCnt; // @[Rob.scala 1224:28]
      end else begin
        dt_exuDebug_14_isPerfCnt <= _GEN_10681;
      end
    end else begin
      dt_exuDebug_14_isPerfCnt <= _GEN_10681;
    end
    if (io_writeback_1_8_valid) begin // @[Rob.scala 1222:23]
      if (5'hf == io_writeback_1_8_bits_uop_robIdx_value) begin // @[Rob.scala 1224:28]
        dt_exuDebug_15_isMMIO <= io_writeback_1_8_bits_debug_isMMIO; // @[Rob.scala 1224:28]
      end else begin
        dt_exuDebug_15_isMMIO <= _GEN_10650;
      end
    end else begin
      dt_exuDebug_15_isMMIO <= _GEN_10650;
    end
    if (io_writeback_1_8_valid) begin // @[Rob.scala 1222:23]
      if (5'hf == io_writeback_1_8_bits_uop_robIdx_value) begin // @[Rob.scala 1224:28]
        dt_exuDebug_15_isPerfCnt <= io_writeback_1_8_bits_debug_isPerfCnt; // @[Rob.scala 1224:28]
      end else begin
        dt_exuDebug_15_isPerfCnt <= _GEN_10682;
      end
    end else begin
      dt_exuDebug_15_isPerfCnt <= _GEN_10682;
    end
    if (io_writeback_1_8_valid) begin // @[Rob.scala 1222:23]
      if (5'h10 == io_writeback_1_8_bits_uop_robIdx_value) begin // @[Rob.scala 1224:28]
        dt_exuDebug_16_isMMIO <= io_writeback_1_8_bits_debug_isMMIO; // @[Rob.scala 1224:28]
      end else begin
        dt_exuDebug_16_isMMIO <= _GEN_10651;
      end
    end else begin
      dt_exuDebug_16_isMMIO <= _GEN_10651;
    end
    if (io_writeback_1_8_valid) begin // @[Rob.scala 1222:23]
      if (5'h10 == io_writeback_1_8_bits_uop_robIdx_value) begin // @[Rob.scala 1224:28]
        dt_exuDebug_16_isPerfCnt <= io_writeback_1_8_bits_debug_isPerfCnt; // @[Rob.scala 1224:28]
      end else begin
        dt_exuDebug_16_isPerfCnt <= _GEN_10683;
      end
    end else begin
      dt_exuDebug_16_isPerfCnt <= _GEN_10683;
    end
    if (io_writeback_1_8_valid) begin // @[Rob.scala 1222:23]
      if (5'h11 == io_writeback_1_8_bits_uop_robIdx_value) begin // @[Rob.scala 1224:28]
        dt_exuDebug_17_isMMIO <= io_writeback_1_8_bits_debug_isMMIO; // @[Rob.scala 1224:28]
      end else begin
        dt_exuDebug_17_isMMIO <= _GEN_10652;
      end
    end else begin
      dt_exuDebug_17_isMMIO <= _GEN_10652;
    end
    if (io_writeback_1_8_valid) begin // @[Rob.scala 1222:23]
      if (5'h11 == io_writeback_1_8_bits_uop_robIdx_value) begin // @[Rob.scala 1224:28]
        dt_exuDebug_17_isPerfCnt <= io_writeback_1_8_bits_debug_isPerfCnt; // @[Rob.scala 1224:28]
      end else begin
        dt_exuDebug_17_isPerfCnt <= _GEN_10684;
      end
    end else begin
      dt_exuDebug_17_isPerfCnt <= _GEN_10684;
    end
    if (io_writeback_1_8_valid) begin // @[Rob.scala 1222:23]
      if (5'h12 == io_writeback_1_8_bits_uop_robIdx_value) begin // @[Rob.scala 1224:28]
        dt_exuDebug_18_isMMIO <= io_writeback_1_8_bits_debug_isMMIO; // @[Rob.scala 1224:28]
      end else begin
        dt_exuDebug_18_isMMIO <= _GEN_10653;
      end
    end else begin
      dt_exuDebug_18_isMMIO <= _GEN_10653;
    end
    if (io_writeback_1_8_valid) begin // @[Rob.scala 1222:23]
      if (5'h12 == io_writeback_1_8_bits_uop_robIdx_value) begin // @[Rob.scala 1224:28]
        dt_exuDebug_18_isPerfCnt <= io_writeback_1_8_bits_debug_isPerfCnt; // @[Rob.scala 1224:28]
      end else begin
        dt_exuDebug_18_isPerfCnt <= _GEN_10685;
      end
    end else begin
      dt_exuDebug_18_isPerfCnt <= _GEN_10685;
    end
    if (io_writeback_1_8_valid) begin // @[Rob.scala 1222:23]
      if (5'h13 == io_writeback_1_8_bits_uop_robIdx_value) begin // @[Rob.scala 1224:28]
        dt_exuDebug_19_isMMIO <= io_writeback_1_8_bits_debug_isMMIO; // @[Rob.scala 1224:28]
      end else begin
        dt_exuDebug_19_isMMIO <= _GEN_10654;
      end
    end else begin
      dt_exuDebug_19_isMMIO <= _GEN_10654;
    end
    if (io_writeback_1_8_valid) begin // @[Rob.scala 1222:23]
      if (5'h13 == io_writeback_1_8_bits_uop_robIdx_value) begin // @[Rob.scala 1224:28]
        dt_exuDebug_19_isPerfCnt <= io_writeback_1_8_bits_debug_isPerfCnt; // @[Rob.scala 1224:28]
      end else begin
        dt_exuDebug_19_isPerfCnt <= _GEN_10686;
      end
    end else begin
      dt_exuDebug_19_isPerfCnt <= _GEN_10686;
    end
    if (io_writeback_1_8_valid) begin // @[Rob.scala 1222:23]
      if (5'h14 == io_writeback_1_8_bits_uop_robIdx_value) begin // @[Rob.scala 1224:28]
        dt_exuDebug_20_isMMIO <= io_writeback_1_8_bits_debug_isMMIO; // @[Rob.scala 1224:28]
      end else begin
        dt_exuDebug_20_isMMIO <= _GEN_10655;
      end
    end else begin
      dt_exuDebug_20_isMMIO <= _GEN_10655;
    end
    if (io_writeback_1_8_valid) begin // @[Rob.scala 1222:23]
      if (5'h14 == io_writeback_1_8_bits_uop_robIdx_value) begin // @[Rob.scala 1224:28]
        dt_exuDebug_20_isPerfCnt <= io_writeback_1_8_bits_debug_isPerfCnt; // @[Rob.scala 1224:28]
      end else begin
        dt_exuDebug_20_isPerfCnt <= _GEN_10687;
      end
    end else begin
      dt_exuDebug_20_isPerfCnt <= _GEN_10687;
    end
    if (io_writeback_1_8_valid) begin // @[Rob.scala 1222:23]
      if (5'h15 == io_writeback_1_8_bits_uop_robIdx_value) begin // @[Rob.scala 1224:28]
        dt_exuDebug_21_isMMIO <= io_writeback_1_8_bits_debug_isMMIO; // @[Rob.scala 1224:28]
      end else begin
        dt_exuDebug_21_isMMIO <= _GEN_10656;
      end
    end else begin
      dt_exuDebug_21_isMMIO <= _GEN_10656;
    end
    if (io_writeback_1_8_valid) begin // @[Rob.scala 1222:23]
      if (5'h15 == io_writeback_1_8_bits_uop_robIdx_value) begin // @[Rob.scala 1224:28]
        dt_exuDebug_21_isPerfCnt <= io_writeback_1_8_bits_debug_isPerfCnt; // @[Rob.scala 1224:28]
      end else begin
        dt_exuDebug_21_isPerfCnt <= _GEN_10688;
      end
    end else begin
      dt_exuDebug_21_isPerfCnt <= _GEN_10688;
    end
    if (io_writeback_1_8_valid) begin // @[Rob.scala 1222:23]
      if (5'h16 == io_writeback_1_8_bits_uop_robIdx_value) begin // @[Rob.scala 1224:28]
        dt_exuDebug_22_isMMIO <= io_writeback_1_8_bits_debug_isMMIO; // @[Rob.scala 1224:28]
      end else begin
        dt_exuDebug_22_isMMIO <= _GEN_10657;
      end
    end else begin
      dt_exuDebug_22_isMMIO <= _GEN_10657;
    end
    if (io_writeback_1_8_valid) begin // @[Rob.scala 1222:23]
      if (5'h16 == io_writeback_1_8_bits_uop_robIdx_value) begin // @[Rob.scala 1224:28]
        dt_exuDebug_22_isPerfCnt <= io_writeback_1_8_bits_debug_isPerfCnt; // @[Rob.scala 1224:28]
      end else begin
        dt_exuDebug_22_isPerfCnt <= _GEN_10689;
      end
    end else begin
      dt_exuDebug_22_isPerfCnt <= _GEN_10689;
    end
    if (io_writeback_1_8_valid) begin // @[Rob.scala 1222:23]
      if (5'h17 == io_writeback_1_8_bits_uop_robIdx_value) begin // @[Rob.scala 1224:28]
        dt_exuDebug_23_isMMIO <= io_writeback_1_8_bits_debug_isMMIO; // @[Rob.scala 1224:28]
      end else begin
        dt_exuDebug_23_isMMIO <= _GEN_10658;
      end
    end else begin
      dt_exuDebug_23_isMMIO <= _GEN_10658;
    end
    if (io_writeback_1_8_valid) begin // @[Rob.scala 1222:23]
      if (5'h17 == io_writeback_1_8_bits_uop_robIdx_value) begin // @[Rob.scala 1224:28]
        dt_exuDebug_23_isPerfCnt <= io_writeback_1_8_bits_debug_isPerfCnt; // @[Rob.scala 1224:28]
      end else begin
        dt_exuDebug_23_isPerfCnt <= _GEN_10690;
      end
    end else begin
      dt_exuDebug_23_isPerfCnt <= _GEN_10690;
    end
    if (io_writeback_1_8_valid) begin // @[Rob.scala 1222:23]
      if (5'h18 == io_writeback_1_8_bits_uop_robIdx_value) begin // @[Rob.scala 1224:28]
        dt_exuDebug_24_isMMIO <= io_writeback_1_8_bits_debug_isMMIO; // @[Rob.scala 1224:28]
      end else begin
        dt_exuDebug_24_isMMIO <= _GEN_10659;
      end
    end else begin
      dt_exuDebug_24_isMMIO <= _GEN_10659;
    end
    if (io_writeback_1_8_valid) begin // @[Rob.scala 1222:23]
      if (5'h18 == io_writeback_1_8_bits_uop_robIdx_value) begin // @[Rob.scala 1224:28]
        dt_exuDebug_24_isPerfCnt <= io_writeback_1_8_bits_debug_isPerfCnt; // @[Rob.scala 1224:28]
      end else begin
        dt_exuDebug_24_isPerfCnt <= _GEN_10691;
      end
    end else begin
      dt_exuDebug_24_isPerfCnt <= _GEN_10691;
    end
    if (io_writeback_1_8_valid) begin // @[Rob.scala 1222:23]
      if (5'h19 == io_writeback_1_8_bits_uop_robIdx_value) begin // @[Rob.scala 1224:28]
        dt_exuDebug_25_isMMIO <= io_writeback_1_8_bits_debug_isMMIO; // @[Rob.scala 1224:28]
      end else begin
        dt_exuDebug_25_isMMIO <= _GEN_10660;
      end
    end else begin
      dt_exuDebug_25_isMMIO <= _GEN_10660;
    end
    if (io_writeback_1_8_valid) begin // @[Rob.scala 1222:23]
      if (5'h19 == io_writeback_1_8_bits_uop_robIdx_value) begin // @[Rob.scala 1224:28]
        dt_exuDebug_25_isPerfCnt <= io_writeback_1_8_bits_debug_isPerfCnt; // @[Rob.scala 1224:28]
      end else begin
        dt_exuDebug_25_isPerfCnt <= _GEN_10692;
      end
    end else begin
      dt_exuDebug_25_isPerfCnt <= _GEN_10692;
    end
    if (io_writeback_1_8_valid) begin // @[Rob.scala 1222:23]
      if (5'h1a == io_writeback_1_8_bits_uop_robIdx_value) begin // @[Rob.scala 1224:28]
        dt_exuDebug_26_isMMIO <= io_writeback_1_8_bits_debug_isMMIO; // @[Rob.scala 1224:28]
      end else begin
        dt_exuDebug_26_isMMIO <= _GEN_10661;
      end
    end else begin
      dt_exuDebug_26_isMMIO <= _GEN_10661;
    end
    if (io_writeback_1_8_valid) begin // @[Rob.scala 1222:23]
      if (5'h1a == io_writeback_1_8_bits_uop_robIdx_value) begin // @[Rob.scala 1224:28]
        dt_exuDebug_26_isPerfCnt <= io_writeback_1_8_bits_debug_isPerfCnt; // @[Rob.scala 1224:28]
      end else begin
        dt_exuDebug_26_isPerfCnt <= _GEN_10693;
      end
    end else begin
      dt_exuDebug_26_isPerfCnt <= _GEN_10693;
    end
    if (io_writeback_1_8_valid) begin // @[Rob.scala 1222:23]
      if (5'h1b == io_writeback_1_8_bits_uop_robIdx_value) begin // @[Rob.scala 1224:28]
        dt_exuDebug_27_isMMIO <= io_writeback_1_8_bits_debug_isMMIO; // @[Rob.scala 1224:28]
      end else begin
        dt_exuDebug_27_isMMIO <= _GEN_10662;
      end
    end else begin
      dt_exuDebug_27_isMMIO <= _GEN_10662;
    end
    if (io_writeback_1_8_valid) begin // @[Rob.scala 1222:23]
      if (5'h1b == io_writeback_1_8_bits_uop_robIdx_value) begin // @[Rob.scala 1224:28]
        dt_exuDebug_27_isPerfCnt <= io_writeback_1_8_bits_debug_isPerfCnt; // @[Rob.scala 1224:28]
      end else begin
        dt_exuDebug_27_isPerfCnt <= _GEN_10694;
      end
    end else begin
      dt_exuDebug_27_isPerfCnt <= _GEN_10694;
    end
    if (io_writeback_1_8_valid) begin // @[Rob.scala 1222:23]
      if (5'h1c == io_writeback_1_8_bits_uop_robIdx_value) begin // @[Rob.scala 1224:28]
        dt_exuDebug_28_isMMIO <= io_writeback_1_8_bits_debug_isMMIO; // @[Rob.scala 1224:28]
      end else begin
        dt_exuDebug_28_isMMIO <= _GEN_10663;
      end
    end else begin
      dt_exuDebug_28_isMMIO <= _GEN_10663;
    end
    if (io_writeback_1_8_valid) begin // @[Rob.scala 1222:23]
      if (5'h1c == io_writeback_1_8_bits_uop_robIdx_value) begin // @[Rob.scala 1224:28]
        dt_exuDebug_28_isPerfCnt <= io_writeback_1_8_bits_debug_isPerfCnt; // @[Rob.scala 1224:28]
      end else begin
        dt_exuDebug_28_isPerfCnt <= _GEN_10695;
      end
    end else begin
      dt_exuDebug_28_isPerfCnt <= _GEN_10695;
    end
    if (io_writeback_1_8_valid) begin // @[Rob.scala 1222:23]
      if (5'h1d == io_writeback_1_8_bits_uop_robIdx_value) begin // @[Rob.scala 1224:28]
        dt_exuDebug_29_isMMIO <= io_writeback_1_8_bits_debug_isMMIO; // @[Rob.scala 1224:28]
      end else begin
        dt_exuDebug_29_isMMIO <= _GEN_10664;
      end
    end else begin
      dt_exuDebug_29_isMMIO <= _GEN_10664;
    end
    if (io_writeback_1_8_valid) begin // @[Rob.scala 1222:23]
      if (5'h1d == io_writeback_1_8_bits_uop_robIdx_value) begin // @[Rob.scala 1224:28]
        dt_exuDebug_29_isPerfCnt <= io_writeback_1_8_bits_debug_isPerfCnt; // @[Rob.scala 1224:28]
      end else begin
        dt_exuDebug_29_isPerfCnt <= _GEN_10696;
      end
    end else begin
      dt_exuDebug_29_isPerfCnt <= _GEN_10696;
    end
    if (io_writeback_1_8_valid) begin // @[Rob.scala 1222:23]
      if (5'h1e == io_writeback_1_8_bits_uop_robIdx_value) begin // @[Rob.scala 1224:28]
        dt_exuDebug_30_isMMIO <= io_writeback_1_8_bits_debug_isMMIO; // @[Rob.scala 1224:28]
      end else begin
        dt_exuDebug_30_isMMIO <= _GEN_10665;
      end
    end else begin
      dt_exuDebug_30_isMMIO <= _GEN_10665;
    end
    if (io_writeback_1_8_valid) begin // @[Rob.scala 1222:23]
      if (5'h1e == io_writeback_1_8_bits_uop_robIdx_value) begin // @[Rob.scala 1224:28]
        dt_exuDebug_30_isPerfCnt <= io_writeback_1_8_bits_debug_isPerfCnt; // @[Rob.scala 1224:28]
      end else begin
        dt_exuDebug_30_isPerfCnt <= _GEN_10697;
      end
    end else begin
      dt_exuDebug_30_isPerfCnt <= _GEN_10697;
    end
    if (io_writeback_1_8_valid) begin // @[Rob.scala 1222:23]
      if (5'h1f == io_writeback_1_8_bits_uop_robIdx_value) begin // @[Rob.scala 1224:28]
        dt_exuDebug_31_isMMIO <= io_writeback_1_8_bits_debug_isMMIO; // @[Rob.scala 1224:28]
      end else begin
        dt_exuDebug_31_isMMIO <= _GEN_10666;
      end
    end else begin
      dt_exuDebug_31_isMMIO <= _GEN_10666;
    end
    if (io_writeback_1_8_valid) begin // @[Rob.scala 1222:23]
      if (5'h1f == io_writeback_1_8_bits_uop_robIdx_value) begin // @[Rob.scala 1224:28]
        dt_exuDebug_31_isPerfCnt <= io_writeback_1_8_bits_debug_isPerfCnt; // @[Rob.scala 1224:28]
      end else begin
        dt_exuDebug_31_isPerfCnt <= _GEN_10698;
      end
    end else begin
      dt_exuDebug_31_isPerfCnt <= _GEN_10698;
    end
    difftest_io_valid_REG <= io_commits_commitValid_0 & io_commits_isCommit; // @[Rob.scala 1239:80]
    difftest_io_valid_REG_1 <= difftest_io_valid_REG; // @[Rob.scala 1239:45]
    difftest_io_valid_REG_2 <= difftest_io_valid_REG_1; // @[Rob.scala 1239:37]
    difftest_io_special_REG <= io_commits_info_0_commitType[2]; // @[package.scala 134:53]
    difftest_io_special_REG_1 <= difftest_io_special_REG; // @[Rob.scala 1240:45]
    difftest_io_special_REG_2 <= difftest_io_special_REG_1; // @[Rob.scala 1240:37]
    if (dt_eliminatedMove_eliminatedMove_data) begin // @[Rob.scala 1241:57]
      difftest_io_skip_REG <= 1'h0;
    end else begin
      difftest_io_skip_REG <= _GEN_11050 | _GEN_11082;
    end
    difftest_io_skip_REG_1 <= difftest_io_skip_REG; // @[Rob.scala 1241:45]
    difftest_io_skip_REG_2 <= difftest_io_skip_REG_1; // @[Rob.scala 1241:37]
    difftest_io_isRVC_REG <= dt_isRVC_isRVC_data; // @[Rob.scala 1242:53]
    difftest_io_isRVC_REG_1 <= difftest_io_isRVC_REG; // @[Rob.scala 1242:45]
    difftest_io_isRVC_REG_2 <= difftest_io_isRVC_REG_1; // @[Rob.scala 1242:37]
    difftest_io_rfwen_REG <= io_commits_commitValid_0 & io_commits_info_0_rfWen & io_commits_info_0_ldest != 5'h0; // @[Rob.scala 1243:100]
    difftest_io_rfwen_REG_1 <= difftest_io_rfwen_REG; // @[Rob.scala 1243:45]
    difftest_io_rfwen_REG_2 <= difftest_io_rfwen_REG_1; // @[Rob.scala 1243:37]
    difftest_io_fpwen_REG <= io_commits_commitValid_0 & io_commits_info_0_fpWen; // @[Rob.scala 1244:80]
    difftest_io_fpwen_REG_1 <= difftest_io_fpwen_REG; // @[Rob.scala 1244:45]
    difftest_io_fpwen_REG_2 <= difftest_io_fpwen_REG_1; // @[Rob.scala 1244:37]
    difftest_io_wpdest_REG <= io_commits_info_0_pdest; // @[Rob.scala 1245:53]
    difftest_io_wpdest_REG_1 <= difftest_io_wpdest_REG; // @[Rob.scala 1245:45]
    difftest_io_wpdest_REG_2 <= difftest_io_wpdest_REG_1; // @[Rob.scala 1245:37]
    difftest_io_wdest_REG <= io_commits_info_0_ldest; // @[Rob.scala 1246:53]
    difftest_io_wdest_REG_1 <= difftest_io_wdest_REG; // @[Rob.scala 1246:45]
    difftest_io_wdest_REG_2 <= difftest_io_wdest_REG_1; // @[Rob.scala 1246:37]
    difftest_io_valid_REG_3 <= io_commits_commitValid_1 & io_commits_isCommit; // @[Rob.scala 1239:80]
    difftest_io_valid_REG_4 <= difftest_io_valid_REG_3; // @[Rob.scala 1239:45]
    difftest_io_valid_REG_5 <= difftest_io_valid_REG_4; // @[Rob.scala 1239:37]
    difftest_io_special_REG_3 <= io_commits_info_1_commitType[2]; // @[package.scala 134:53]
    difftest_io_special_REG_4 <= difftest_io_special_REG_3; // @[Rob.scala 1240:45]
    difftest_io_special_REG_5 <= difftest_io_special_REG_4; // @[Rob.scala 1240:37]
    if (dt_eliminatedMove_eliminatedMove_1_data) begin // @[Rob.scala 1241:57]
      difftest_io_skip_REG_3 <= 1'h0;
    end else begin
      difftest_io_skip_REG_3 <= _GEN_11114 | _GEN_11146;
    end
    difftest_io_skip_REG_4 <= difftest_io_skip_REG_3; // @[Rob.scala 1241:45]
    difftest_io_skip_REG_5 <= difftest_io_skip_REG_4; // @[Rob.scala 1241:37]
    difftest_io_isRVC_REG_3 <= dt_isRVC_isRVC_1_data; // @[Rob.scala 1242:53]
    difftest_io_isRVC_REG_4 <= difftest_io_isRVC_REG_3; // @[Rob.scala 1242:45]
    difftest_io_isRVC_REG_5 <= difftest_io_isRVC_REG_4; // @[Rob.scala 1242:37]
    difftest_io_rfwen_REG_3 <= io_commits_commitValid_1 & io_commits_info_1_rfWen & io_commits_info_1_ldest != 5'h0; // @[Rob.scala 1243:100]
    difftest_io_rfwen_REG_4 <= difftest_io_rfwen_REG_3; // @[Rob.scala 1243:45]
    difftest_io_rfwen_REG_5 <= difftest_io_rfwen_REG_4; // @[Rob.scala 1243:37]
    difftest_io_fpwen_REG_3 <= io_commits_commitValid_1 & io_commits_info_1_fpWen; // @[Rob.scala 1244:80]
    difftest_io_fpwen_REG_4 <= difftest_io_fpwen_REG_3; // @[Rob.scala 1244:45]
    difftest_io_fpwen_REG_5 <= difftest_io_fpwen_REG_4; // @[Rob.scala 1244:37]
    difftest_io_wpdest_REG_3 <= io_commits_info_1_pdest; // @[Rob.scala 1245:53]
    difftest_io_wpdest_REG_4 <= difftest_io_wpdest_REG_3; // @[Rob.scala 1245:45]
    difftest_io_wpdest_REG_5 <= difftest_io_wpdest_REG_4; // @[Rob.scala 1245:37]
    difftest_io_wdest_REG_3 <= io_commits_info_1_ldest; // @[Rob.scala 1246:53]
    difftest_io_wdest_REG_4 <= difftest_io_wdest_REG_3; // @[Rob.scala 1246:45]
    difftest_io_wdest_REG_5 <= difftest_io_wdest_REG_4; // @[Rob.scala 1246:37]
    validEntriesBanks_0 <= _T_461 + _T_491; // @[Bitwise.scala 48:55]
    validEntries <= validEntriesBanks_0; // @[Rob.scala 1307:29]
    REG_19 <= io_commits_isCommit; // @[Rob.scala 1049:53]
    REG_20_0 <= io_commits_commitValid_0 & debug_microOp_ctrl_isMove_commitDebugUop_0_data; // @[Rob.scala 1308:94]
    REG_20_1 <= io_commits_commitValid_1 & debug_microOp_ctrl_isMove_commitDebugUop_1_data; // @[Rob.scala 1308:94]
    REG_21 <= io_commits_isCommit; // @[Rob.scala 1049:53]
    REG_22 <= io_commits_isCommit; // @[Rob.scala 1049:53]
    REG_23_0 <= io_commits_commitValid_0 & _ldCommitVec_T; // @[Rob.scala 1064:88]
    REG_23_1 <= io_commits_commitValid_1 & _ldCommitVec_T_2; // @[Rob.scala 1064:88]
    REG_24 <= io_commits_isCommit; // @[Rob.scala 1049:53]
    REG_25_0 <= io_commits_commitValid_0 & commitIsBranch_0; // @[Rob.scala 1067:92]
    REG_25_1 <= io_commits_commitValid_1 & commitIsBranch_1; // @[Rob.scala 1067:92]
    REG_26 <= io_commits_isCommit; // @[Rob.scala 1049:53]
    REG_27_0 <= ldCommitVec_0 & debug_microOp_cf_loadWaitBit_commitDebugUop_0_data; // @[Rob.scala 1311:96]
    REG_27_1 <= ldCommitVec_1 & debug_microOp_cf_loadWaitBit_commitDebugUop_1_data; // @[Rob.scala 1311:96]
    REG_28 <= io_commits_isCommit; // @[Rob.scala 1049:53]
    REG_29_0 <= io_commits_commitValid_0 & _stCommitVec_T; // @[Rob.scala 1312:96]
    REG_29_1 <= io_commits_commitValid_1 & _stCommitVec_T_2; // @[Rob.scala 1312:96]
    REG_30 <= io_commits_isCommit; // @[Rob.scala 1049:53]
    io_perf_0_value_REG <= io_flushOut_valid & intrEnable; // @[Rob.scala 1314:51]
    io_perf_0_value_REG_1 <= io_perf_0_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_1_value_REG <= io_flushOut_valid & exceptionEnable; // @[Rob.scala 1315:51]
    io_perf_1_value_REG_1 <= io_perf_1_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_2_value_REG <= io_flushOut_valid & isFlushPipe; // @[Rob.scala 1316:51]
    io_perf_2_value_REG_1 <= io_perf_2_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_3_value_REG <= _T_108 & deqHasReplayInst; // @[Rob.scala 1317:66]
    io_perf_3_value_REG_1 <= io_perf_3_value_REG; // @[PerfCounterUtils.scala 188:27]
    if (io_commits_isCommit) begin // @[Rob.scala 1048:42]
      io_perf_4_value_REG <= commitCnt;
    end else begin
      io_perf_4_value_REG <= 2'h0;
    end
    io_perf_4_value_REG_1 <= io_perf_4_value_REG; // @[PerfCounterUtils.scala 188:27]
    if (REG_19) begin // @[Rob.scala 1049:45]
      io_perf_5_value_REG <= trueCommitCnt;
    end else begin
      io_perf_5_value_REG <= 3'h0;
    end
    io_perf_5_value_REG_1 <= io_perf_5_value_REG; // @[PerfCounterUtils.scala 188:27]
    if (REG_21) begin // @[Rob.scala 1049:45]
      io_perf_6_value_REG <= _T_1083;
    end else begin
      io_perf_6_value_REG <= 2'h0;
    end
    io_perf_6_value_REG_1 <= io_perf_6_value_REG; // @[PerfCounterUtils.scala 188:27]
    if (REG_22) begin // @[Rob.scala 1049:45]
      io_perf_7_value_REG <= fuseCommitCnt;
    end else begin
      io_perf_7_value_REG <= 2'h0;
    end
    io_perf_7_value_REG_1 <= io_perf_7_value_REG; // @[PerfCounterUtils.scala 188:27]
    if (REG_24) begin // @[Rob.scala 1049:45]
      io_perf_8_value_REG <= _T_1087;
    end else begin
      io_perf_8_value_REG <= 2'h0;
    end
    io_perf_8_value_REG_1 <= io_perf_8_value_REG; // @[PerfCounterUtils.scala 188:27]
    if (REG_26) begin // @[Rob.scala 1049:45]
      io_perf_9_value_REG <= _T_1090;
    end else begin
      io_perf_9_value_REG <= 2'h0;
    end
    io_perf_9_value_REG_1 <= io_perf_9_value_REG; // @[PerfCounterUtils.scala 188:27]
    if (REG_28) begin // @[Rob.scala 1049:45]
      io_perf_10_value_REG <= _T_1093;
    end else begin
      io_perf_10_value_REG <= 2'h0;
    end
    io_perf_10_value_REG_1 <= io_perf_10_value_REG; // @[PerfCounterUtils.scala 188:27]
    if (REG_30) begin // @[Rob.scala 1049:45]
      io_perf_11_value_REG <= _T_1096;
    end else begin
      io_perf_11_value_REG <= 2'h0;
    end
    io_perf_11_value_REG_1 <= io_perf_11_value_REG; // @[PerfCounterUtils.scala 188:27]
    if (io_commits_isWalk) begin // @[Rob.scala 1326:36]
      io_perf_12_value_REG <= _T_619;
    end else begin
      io_perf_12_value_REG <= 2'h0;
    end
    io_perf_12_value_REG_1 <= io_perf_12_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_13_value_REG <= state; // @[Rob.scala 1327:40]
    io_perf_13_value_REG_1 <= io_perf_13_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_14_value_REG <= validEntries <= 6'h8; // @[Rob.scala 1328:46]
    io_perf_14_value_REG_1 <= io_perf_14_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_15_value_REG <= validEntries > 6'h8 & validEntries <= 6'h10; // @[Rob.scala 1329:65]
    io_perf_15_value_REG_1 <= io_perf_15_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_16_value_REG <= validEntries > 6'h10 & validEntries <= 6'h18; // @[Rob.scala 1330:65]
    io_perf_16_value_REG_1 <= io_perf_16_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_17_value_REG <= validEntries > 6'h18; // @[Rob.scala 1331:46]
    io_perf_17_value_REG_1 <= io_perf_17_value_REG; // @[PerfCounterUtils.scala 188:27]
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Rob.scala 876:24]
      valid_0 <= 1'h0; // @[Rob.scala 877:{32,32}]
    end else if (_T_125) begin
      if (5'h0 == commitReadAddr_1) begin
        valid_0 <= 1'h0;
      end else begin
        valid_0 <= _GEN_5446;
      end
    end else begin
      valid_0 <= _GEN_5446;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Rob.scala 876:24]
      valid_1 <= 1'h0; // @[Rob.scala 877:{32,32}]
    end else if (_T_125) begin
      if (5'h1 == commitReadAddr_1) begin
        valid_1 <= 1'h0;
      end else begin
        valid_1 <= _GEN_5447;
      end
    end else begin
      valid_1 <= _GEN_5447;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Rob.scala 876:24]
      valid_2 <= 1'h0; // @[Rob.scala 877:{32,32}]
    end else if (_T_125) begin
      if (5'h2 == commitReadAddr_1) begin
        valid_2 <= 1'h0;
      end else begin
        valid_2 <= _GEN_5448;
      end
    end else begin
      valid_2 <= _GEN_5448;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Rob.scala 876:24]
      valid_3 <= 1'h0; // @[Rob.scala 877:{32,32}]
    end else if (_T_125) begin
      if (5'h3 == commitReadAddr_1) begin
        valid_3 <= 1'h0;
      end else begin
        valid_3 <= _GEN_5449;
      end
    end else begin
      valid_3 <= _GEN_5449;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Rob.scala 876:24]
      valid_4 <= 1'h0; // @[Rob.scala 877:{32,32}]
    end else if (_T_125) begin
      if (5'h4 == commitReadAddr_1) begin
        valid_4 <= 1'h0;
      end else begin
        valid_4 <= _GEN_5450;
      end
    end else begin
      valid_4 <= _GEN_5450;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Rob.scala 876:24]
      valid_5 <= 1'h0; // @[Rob.scala 877:{32,32}]
    end else if (_T_125) begin
      if (5'h5 == commitReadAddr_1) begin
        valid_5 <= 1'h0;
      end else begin
        valid_5 <= _GEN_5451;
      end
    end else begin
      valid_5 <= _GEN_5451;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Rob.scala 876:24]
      valid_6 <= 1'h0; // @[Rob.scala 877:{32,32}]
    end else if (_T_125) begin
      if (5'h6 == commitReadAddr_1) begin
        valid_6 <= 1'h0;
      end else begin
        valid_6 <= _GEN_5452;
      end
    end else begin
      valid_6 <= _GEN_5452;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Rob.scala 876:24]
      valid_7 <= 1'h0; // @[Rob.scala 877:{32,32}]
    end else if (_T_125) begin
      if (5'h7 == commitReadAddr_1) begin
        valid_7 <= 1'h0;
      end else begin
        valid_7 <= _GEN_5453;
      end
    end else begin
      valid_7 <= _GEN_5453;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Rob.scala 876:24]
      valid_8 <= 1'h0; // @[Rob.scala 877:{32,32}]
    end else if (_T_125) begin
      if (5'h8 == commitReadAddr_1) begin
        valid_8 <= 1'h0;
      end else begin
        valid_8 <= _GEN_5454;
      end
    end else begin
      valid_8 <= _GEN_5454;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Rob.scala 876:24]
      valid_9 <= 1'h0; // @[Rob.scala 877:{32,32}]
    end else if (_T_125) begin
      if (5'h9 == commitReadAddr_1) begin
        valid_9 <= 1'h0;
      end else begin
        valid_9 <= _GEN_5455;
      end
    end else begin
      valid_9 <= _GEN_5455;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Rob.scala 876:24]
      valid_10 <= 1'h0; // @[Rob.scala 877:{32,32}]
    end else if (_T_125) begin
      if (5'ha == commitReadAddr_1) begin
        valid_10 <= 1'h0;
      end else begin
        valid_10 <= _GEN_5456;
      end
    end else begin
      valid_10 <= _GEN_5456;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Rob.scala 876:24]
      valid_11 <= 1'h0; // @[Rob.scala 877:{32,32}]
    end else if (_T_125) begin
      if (5'hb == commitReadAddr_1) begin
        valid_11 <= 1'h0;
      end else begin
        valid_11 <= _GEN_5457;
      end
    end else begin
      valid_11 <= _GEN_5457;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Rob.scala 876:24]
      valid_12 <= 1'h0; // @[Rob.scala 877:{32,32}]
    end else if (_T_125) begin
      if (5'hc == commitReadAddr_1) begin
        valid_12 <= 1'h0;
      end else begin
        valid_12 <= _GEN_5458;
      end
    end else begin
      valid_12 <= _GEN_5458;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Rob.scala 876:24]
      valid_13 <= 1'h0; // @[Rob.scala 877:{32,32}]
    end else if (_T_125) begin
      if (5'hd == commitReadAddr_1) begin
        valid_13 <= 1'h0;
      end else begin
        valid_13 <= _GEN_5459;
      end
    end else begin
      valid_13 <= _GEN_5459;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Rob.scala 876:24]
      valid_14 <= 1'h0; // @[Rob.scala 877:{32,32}]
    end else if (_T_125) begin
      if (5'he == commitReadAddr_1) begin
        valid_14 <= 1'h0;
      end else begin
        valid_14 <= _GEN_5460;
      end
    end else begin
      valid_14 <= _GEN_5460;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Rob.scala 876:24]
      valid_15 <= 1'h0; // @[Rob.scala 877:{32,32}]
    end else if (_T_125) begin
      if (5'hf == commitReadAddr_1) begin
        valid_15 <= 1'h0;
      end else begin
        valid_15 <= _GEN_5461;
      end
    end else begin
      valid_15 <= _GEN_5461;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Rob.scala 876:24]
      valid_16 <= 1'h0; // @[Rob.scala 877:{32,32}]
    end else if (_T_125) begin
      if (5'h10 == commitReadAddr_1) begin
        valid_16 <= 1'h0;
      end else begin
        valid_16 <= _GEN_5462;
      end
    end else begin
      valid_16 <= _GEN_5462;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Rob.scala 876:24]
      valid_17 <= 1'h0; // @[Rob.scala 877:{32,32}]
    end else if (_T_125) begin
      if (5'h11 == commitReadAddr_1) begin
        valid_17 <= 1'h0;
      end else begin
        valid_17 <= _GEN_5463;
      end
    end else begin
      valid_17 <= _GEN_5463;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Rob.scala 876:24]
      valid_18 <= 1'h0; // @[Rob.scala 877:{32,32}]
    end else if (_T_125) begin
      if (5'h12 == commitReadAddr_1) begin
        valid_18 <= 1'h0;
      end else begin
        valid_18 <= _GEN_5464;
      end
    end else begin
      valid_18 <= _GEN_5464;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Rob.scala 876:24]
      valid_19 <= 1'h0; // @[Rob.scala 877:{32,32}]
    end else if (_T_125) begin
      if (5'h13 == commitReadAddr_1) begin
        valid_19 <= 1'h0;
      end else begin
        valid_19 <= _GEN_5465;
      end
    end else begin
      valid_19 <= _GEN_5465;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Rob.scala 876:24]
      valid_20 <= 1'h0; // @[Rob.scala 877:{32,32}]
    end else if (_T_125) begin
      if (5'h14 == commitReadAddr_1) begin
        valid_20 <= 1'h0;
      end else begin
        valid_20 <= _GEN_5466;
      end
    end else begin
      valid_20 <= _GEN_5466;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Rob.scala 876:24]
      valid_21 <= 1'h0; // @[Rob.scala 877:{32,32}]
    end else if (_T_125) begin
      if (5'h15 == commitReadAddr_1) begin
        valid_21 <= 1'h0;
      end else begin
        valid_21 <= _GEN_5467;
      end
    end else begin
      valid_21 <= _GEN_5467;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Rob.scala 876:24]
      valid_22 <= 1'h0; // @[Rob.scala 877:{32,32}]
    end else if (_T_125) begin
      if (5'h16 == commitReadAddr_1) begin
        valid_22 <= 1'h0;
      end else begin
        valid_22 <= _GEN_5468;
      end
    end else begin
      valid_22 <= _GEN_5468;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Rob.scala 876:24]
      valid_23 <= 1'h0; // @[Rob.scala 877:{32,32}]
    end else if (_T_125) begin
      if (5'h17 == commitReadAddr_1) begin
        valid_23 <= 1'h0;
      end else begin
        valid_23 <= _GEN_5469;
      end
    end else begin
      valid_23 <= _GEN_5469;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Rob.scala 876:24]
      valid_24 <= 1'h0; // @[Rob.scala 877:{32,32}]
    end else if (_T_125) begin
      if (5'h18 == commitReadAddr_1) begin
        valid_24 <= 1'h0;
      end else begin
        valid_24 <= _GEN_5470;
      end
    end else begin
      valid_24 <= _GEN_5470;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Rob.scala 876:24]
      valid_25 <= 1'h0; // @[Rob.scala 877:{32,32}]
    end else if (_T_125) begin
      if (5'h19 == commitReadAddr_1) begin
        valid_25 <= 1'h0;
      end else begin
        valid_25 <= _GEN_5471;
      end
    end else begin
      valid_25 <= _GEN_5471;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Rob.scala 876:24]
      valid_26 <= 1'h0; // @[Rob.scala 877:{32,32}]
    end else if (_T_125) begin
      if (5'h1a == commitReadAddr_1) begin
        valid_26 <= 1'h0;
      end else begin
        valid_26 <= _GEN_5472;
      end
    end else begin
      valid_26 <= _GEN_5472;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Rob.scala 876:24]
      valid_27 <= 1'h0; // @[Rob.scala 877:{32,32}]
    end else if (_T_125) begin
      if (5'h1b == commitReadAddr_1) begin
        valid_27 <= 1'h0;
      end else begin
        valid_27 <= _GEN_5473;
      end
    end else begin
      valid_27 <= _GEN_5473;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Rob.scala 876:24]
      valid_28 <= 1'h0; // @[Rob.scala 877:{32,32}]
    end else if (_T_125) begin
      if (5'h1c == commitReadAddr_1) begin
        valid_28 <= 1'h0;
      end else begin
        valid_28 <= _GEN_5474;
      end
    end else begin
      valid_28 <= _GEN_5474;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Rob.scala 876:24]
      valid_29 <= 1'h0; // @[Rob.scala 877:{32,32}]
    end else if (_T_125) begin
      if (5'h1d == commitReadAddr_1) begin
        valid_29 <= 1'h0;
      end else begin
        valid_29 <= _GEN_5475;
      end
    end else begin
      valid_29 <= _GEN_5475;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Rob.scala 876:24]
      valid_30 <= 1'h0; // @[Rob.scala 877:{32,32}]
    end else if (_T_125) begin
      if (5'h1e == commitReadAddr_1) begin
        valid_30 <= 1'h0;
      end else begin
        valid_30 <= _GEN_5476;
      end
    end else begin
      valid_30 <= _GEN_5476;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Rob.scala 876:24]
      valid_31 <= 1'h0; // @[Rob.scala 877:{32,32}]
    end else if (_T_125) begin
      if (5'h1f == commitReadAddr_1) begin
        valid_31 <= 1'h0;
      end else begin
        valid_31 <= _GEN_5477;
      end
    end else begin
      valid_31 <= _GEN_5477;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Rob.scala 606:38]
      mmio_0 <= 1'h0;
    end else if (REG_5) begin // @[Rob.scala 606:38]
      mmio_0 <= _GEN_4743;
    end else if (REG_3) begin // @[Rob.scala 523:26]
      mmio_0 <= _GEN_4679; // @[Rob.scala 562:{22,22}]
    end else if (canEnqueue_1) begin
      if (5'h0 == allocatePtrVec_1_value) begin
        mmio_0 <= 1'h0;
      end else begin
        mmio_0 <= _GEN_804;
      end
    end else begin
      mmio_0 <= _GEN_804;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Rob.scala 606:38]
      mmio_1 <= 1'h0;
    end else if (REG_5) begin // @[Rob.scala 606:38]
      mmio_1 <= _GEN_4744;
    end else if (REG_3) begin // @[Rob.scala 523:26]
      mmio_1 <= _GEN_4680; // @[Rob.scala 562:{22,22}]
    end else if (canEnqueue_1) begin
      if (5'h1 == allocatePtrVec_1_value) begin
        mmio_1 <= 1'h0;
      end else begin
        mmio_1 <= _GEN_805;
      end
    end else begin
      mmio_1 <= _GEN_805;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Rob.scala 606:38]
      mmio_2 <= 1'h0;
    end else if (REG_5) begin // @[Rob.scala 606:38]
      mmio_2 <= _GEN_4745;
    end else if (REG_3) begin // @[Rob.scala 523:26]
      mmio_2 <= _GEN_4681; // @[Rob.scala 562:{22,22}]
    end else if (canEnqueue_1) begin
      if (5'h2 == allocatePtrVec_1_value) begin
        mmio_2 <= 1'h0;
      end else begin
        mmio_2 <= _GEN_806;
      end
    end else begin
      mmio_2 <= _GEN_806;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Rob.scala 606:38]
      mmio_3 <= 1'h0;
    end else if (REG_5) begin // @[Rob.scala 606:38]
      mmio_3 <= _GEN_4746;
    end else if (REG_3) begin // @[Rob.scala 523:26]
      mmio_3 <= _GEN_4682; // @[Rob.scala 562:{22,22}]
    end else if (canEnqueue_1) begin
      if (5'h3 == allocatePtrVec_1_value) begin
        mmio_3 <= 1'h0;
      end else begin
        mmio_3 <= _GEN_807;
      end
    end else begin
      mmio_3 <= _GEN_807;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Rob.scala 606:38]
      mmio_4 <= 1'h0;
    end else if (REG_5) begin // @[Rob.scala 606:38]
      mmio_4 <= _GEN_4747;
    end else if (REG_3) begin // @[Rob.scala 523:26]
      mmio_4 <= _GEN_4683; // @[Rob.scala 562:{22,22}]
    end else if (canEnqueue_1) begin
      if (5'h4 == allocatePtrVec_1_value) begin
        mmio_4 <= 1'h0;
      end else begin
        mmio_4 <= _GEN_808;
      end
    end else begin
      mmio_4 <= _GEN_808;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Rob.scala 606:38]
      mmio_5 <= 1'h0;
    end else if (REG_5) begin // @[Rob.scala 606:38]
      mmio_5 <= _GEN_4748;
    end else if (REG_3) begin // @[Rob.scala 523:26]
      mmio_5 <= _GEN_4684; // @[Rob.scala 562:{22,22}]
    end else if (canEnqueue_1) begin
      if (5'h5 == allocatePtrVec_1_value) begin
        mmio_5 <= 1'h0;
      end else begin
        mmio_5 <= _GEN_809;
      end
    end else begin
      mmio_5 <= _GEN_809;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Rob.scala 606:38]
      mmio_6 <= 1'h0;
    end else if (REG_5) begin // @[Rob.scala 606:38]
      mmio_6 <= _GEN_4749;
    end else if (REG_3) begin // @[Rob.scala 523:26]
      mmio_6 <= _GEN_4685; // @[Rob.scala 562:{22,22}]
    end else if (canEnqueue_1) begin
      if (5'h6 == allocatePtrVec_1_value) begin
        mmio_6 <= 1'h0;
      end else begin
        mmio_6 <= _GEN_810;
      end
    end else begin
      mmio_6 <= _GEN_810;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Rob.scala 606:38]
      mmio_7 <= 1'h0;
    end else if (REG_5) begin // @[Rob.scala 606:38]
      mmio_7 <= _GEN_4750;
    end else if (REG_3) begin // @[Rob.scala 523:26]
      mmio_7 <= _GEN_4686; // @[Rob.scala 562:{22,22}]
    end else if (canEnqueue_1) begin
      if (5'h7 == allocatePtrVec_1_value) begin
        mmio_7 <= 1'h0;
      end else begin
        mmio_7 <= _GEN_811;
      end
    end else begin
      mmio_7 <= _GEN_811;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Rob.scala 606:38]
      mmio_8 <= 1'h0;
    end else if (REG_5) begin // @[Rob.scala 606:38]
      mmio_8 <= _GEN_4751;
    end else if (REG_3) begin // @[Rob.scala 523:26]
      mmio_8 <= _GEN_4687; // @[Rob.scala 562:{22,22}]
    end else if (canEnqueue_1) begin
      if (5'h8 == allocatePtrVec_1_value) begin
        mmio_8 <= 1'h0;
      end else begin
        mmio_8 <= _GEN_812;
      end
    end else begin
      mmio_8 <= _GEN_812;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Rob.scala 606:38]
      mmio_9 <= 1'h0;
    end else if (REG_5) begin // @[Rob.scala 606:38]
      mmio_9 <= _GEN_4752;
    end else if (REG_3) begin // @[Rob.scala 523:26]
      mmio_9 <= _GEN_4688; // @[Rob.scala 562:{22,22}]
    end else if (canEnqueue_1) begin
      if (5'h9 == allocatePtrVec_1_value) begin
        mmio_9 <= 1'h0;
      end else begin
        mmio_9 <= _GEN_813;
      end
    end else begin
      mmio_9 <= _GEN_813;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Rob.scala 606:38]
      mmio_10 <= 1'h0;
    end else if (REG_5) begin // @[Rob.scala 606:38]
      mmio_10 <= _GEN_4753;
    end else if (REG_3) begin // @[Rob.scala 523:26]
      mmio_10 <= _GEN_4689; // @[Rob.scala 562:{22,22}]
    end else if (canEnqueue_1) begin
      if (5'ha == allocatePtrVec_1_value) begin
        mmio_10 <= 1'h0;
      end else begin
        mmio_10 <= _GEN_814;
      end
    end else begin
      mmio_10 <= _GEN_814;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Rob.scala 606:38]
      mmio_11 <= 1'h0;
    end else if (REG_5) begin // @[Rob.scala 606:38]
      mmio_11 <= _GEN_4754;
    end else if (REG_3) begin // @[Rob.scala 523:26]
      mmio_11 <= _GEN_4690; // @[Rob.scala 562:{22,22}]
    end else if (canEnqueue_1) begin
      if (5'hb == allocatePtrVec_1_value) begin
        mmio_11 <= 1'h0;
      end else begin
        mmio_11 <= _GEN_815;
      end
    end else begin
      mmio_11 <= _GEN_815;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Rob.scala 606:38]
      mmio_12 <= 1'h0;
    end else if (REG_5) begin // @[Rob.scala 606:38]
      mmio_12 <= _GEN_4755;
    end else if (REG_3) begin // @[Rob.scala 523:26]
      mmio_12 <= _GEN_4691; // @[Rob.scala 562:{22,22}]
    end else if (canEnqueue_1) begin
      if (5'hc == allocatePtrVec_1_value) begin
        mmio_12 <= 1'h0;
      end else begin
        mmio_12 <= _GEN_816;
      end
    end else begin
      mmio_12 <= _GEN_816;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Rob.scala 606:38]
      mmio_13 <= 1'h0;
    end else if (REG_5) begin // @[Rob.scala 606:38]
      mmio_13 <= _GEN_4756;
    end else if (REG_3) begin // @[Rob.scala 523:26]
      mmio_13 <= _GEN_4692; // @[Rob.scala 562:{22,22}]
    end else if (canEnqueue_1) begin
      if (5'hd == allocatePtrVec_1_value) begin
        mmio_13 <= 1'h0;
      end else begin
        mmio_13 <= _GEN_817;
      end
    end else begin
      mmio_13 <= _GEN_817;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Rob.scala 606:38]
      mmio_14 <= 1'h0;
    end else if (REG_5) begin // @[Rob.scala 606:38]
      mmio_14 <= _GEN_4757;
    end else if (REG_3) begin // @[Rob.scala 523:26]
      mmio_14 <= _GEN_4693; // @[Rob.scala 562:{22,22}]
    end else if (canEnqueue_1) begin
      if (5'he == allocatePtrVec_1_value) begin
        mmio_14 <= 1'h0;
      end else begin
        mmio_14 <= _GEN_818;
      end
    end else begin
      mmio_14 <= _GEN_818;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Rob.scala 606:38]
      mmio_15 <= 1'h0;
    end else if (REG_5) begin // @[Rob.scala 606:38]
      mmio_15 <= _GEN_4758;
    end else if (REG_3) begin // @[Rob.scala 523:26]
      mmio_15 <= _GEN_4694; // @[Rob.scala 562:{22,22}]
    end else if (canEnqueue_1) begin
      if (5'hf == allocatePtrVec_1_value) begin
        mmio_15 <= 1'h0;
      end else begin
        mmio_15 <= _GEN_819;
      end
    end else begin
      mmio_15 <= _GEN_819;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Rob.scala 606:38]
      mmio_16 <= 1'h0;
    end else if (REG_5) begin // @[Rob.scala 606:38]
      mmio_16 <= _GEN_4759;
    end else if (REG_3) begin // @[Rob.scala 523:26]
      mmio_16 <= _GEN_4695; // @[Rob.scala 562:{22,22}]
    end else if (canEnqueue_1) begin
      if (5'h10 == allocatePtrVec_1_value) begin
        mmio_16 <= 1'h0;
      end else begin
        mmio_16 <= _GEN_820;
      end
    end else begin
      mmio_16 <= _GEN_820;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Rob.scala 606:38]
      mmio_17 <= 1'h0;
    end else if (REG_5) begin // @[Rob.scala 606:38]
      mmio_17 <= _GEN_4760;
    end else if (REG_3) begin // @[Rob.scala 523:26]
      mmio_17 <= _GEN_4696; // @[Rob.scala 562:{22,22}]
    end else if (canEnqueue_1) begin
      if (5'h11 == allocatePtrVec_1_value) begin
        mmio_17 <= 1'h0;
      end else begin
        mmio_17 <= _GEN_821;
      end
    end else begin
      mmio_17 <= _GEN_821;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Rob.scala 606:38]
      mmio_18 <= 1'h0;
    end else if (REG_5) begin // @[Rob.scala 606:38]
      mmio_18 <= _GEN_4761;
    end else if (REG_3) begin // @[Rob.scala 523:26]
      mmio_18 <= _GEN_4697; // @[Rob.scala 562:{22,22}]
    end else if (canEnqueue_1) begin
      if (5'h12 == allocatePtrVec_1_value) begin
        mmio_18 <= 1'h0;
      end else begin
        mmio_18 <= _GEN_822;
      end
    end else begin
      mmio_18 <= _GEN_822;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Rob.scala 606:38]
      mmio_19 <= 1'h0;
    end else if (REG_5) begin // @[Rob.scala 606:38]
      mmio_19 <= _GEN_4762;
    end else if (REG_3) begin // @[Rob.scala 523:26]
      mmio_19 <= _GEN_4698; // @[Rob.scala 562:{22,22}]
    end else if (canEnqueue_1) begin
      if (5'h13 == allocatePtrVec_1_value) begin
        mmio_19 <= 1'h0;
      end else begin
        mmio_19 <= _GEN_823;
      end
    end else begin
      mmio_19 <= _GEN_823;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Rob.scala 606:38]
      mmio_20 <= 1'h0;
    end else if (REG_5) begin // @[Rob.scala 606:38]
      mmio_20 <= _GEN_4763;
    end else if (REG_3) begin // @[Rob.scala 523:26]
      mmio_20 <= _GEN_4699; // @[Rob.scala 562:{22,22}]
    end else if (canEnqueue_1) begin
      if (5'h14 == allocatePtrVec_1_value) begin
        mmio_20 <= 1'h0;
      end else begin
        mmio_20 <= _GEN_824;
      end
    end else begin
      mmio_20 <= _GEN_824;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Rob.scala 606:38]
      mmio_21 <= 1'h0;
    end else if (REG_5) begin // @[Rob.scala 606:38]
      mmio_21 <= _GEN_4764;
    end else if (REG_3) begin // @[Rob.scala 523:26]
      mmio_21 <= _GEN_4700; // @[Rob.scala 562:{22,22}]
    end else if (canEnqueue_1) begin
      if (5'h15 == allocatePtrVec_1_value) begin
        mmio_21 <= 1'h0;
      end else begin
        mmio_21 <= _GEN_825;
      end
    end else begin
      mmio_21 <= _GEN_825;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Rob.scala 606:38]
      mmio_22 <= 1'h0;
    end else if (REG_5) begin // @[Rob.scala 606:38]
      mmio_22 <= _GEN_4765;
    end else if (REG_3) begin // @[Rob.scala 523:26]
      mmio_22 <= _GEN_4701; // @[Rob.scala 562:{22,22}]
    end else if (canEnqueue_1) begin
      if (5'h16 == allocatePtrVec_1_value) begin
        mmio_22 <= 1'h0;
      end else begin
        mmio_22 <= _GEN_826;
      end
    end else begin
      mmio_22 <= _GEN_826;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Rob.scala 606:38]
      mmio_23 <= 1'h0;
    end else if (REG_5) begin // @[Rob.scala 606:38]
      mmio_23 <= _GEN_4766;
    end else if (REG_3) begin // @[Rob.scala 523:26]
      mmio_23 <= _GEN_4702; // @[Rob.scala 562:{22,22}]
    end else if (canEnqueue_1) begin
      if (5'h17 == allocatePtrVec_1_value) begin
        mmio_23 <= 1'h0;
      end else begin
        mmio_23 <= _GEN_827;
      end
    end else begin
      mmio_23 <= _GEN_827;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Rob.scala 606:38]
      mmio_24 <= 1'h0;
    end else if (REG_5) begin // @[Rob.scala 606:38]
      mmio_24 <= _GEN_4767;
    end else if (REG_3) begin // @[Rob.scala 523:26]
      mmio_24 <= _GEN_4703; // @[Rob.scala 562:{22,22}]
    end else if (canEnqueue_1) begin
      if (5'h18 == allocatePtrVec_1_value) begin
        mmio_24 <= 1'h0;
      end else begin
        mmio_24 <= _GEN_828;
      end
    end else begin
      mmio_24 <= _GEN_828;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Rob.scala 606:38]
      mmio_25 <= 1'h0;
    end else if (REG_5) begin // @[Rob.scala 606:38]
      mmio_25 <= _GEN_4768;
    end else if (REG_3) begin // @[Rob.scala 523:26]
      mmio_25 <= _GEN_4704; // @[Rob.scala 562:{22,22}]
    end else if (canEnqueue_1) begin
      if (5'h19 == allocatePtrVec_1_value) begin
        mmio_25 <= 1'h0;
      end else begin
        mmio_25 <= _GEN_829;
      end
    end else begin
      mmio_25 <= _GEN_829;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Rob.scala 606:38]
      mmio_26 <= 1'h0;
    end else if (REG_5) begin // @[Rob.scala 606:38]
      mmio_26 <= _GEN_4769;
    end else if (REG_3) begin // @[Rob.scala 523:26]
      mmio_26 <= _GEN_4705; // @[Rob.scala 562:{22,22}]
    end else if (canEnqueue_1) begin
      if (5'h1a == allocatePtrVec_1_value) begin
        mmio_26 <= 1'h0;
      end else begin
        mmio_26 <= _GEN_830;
      end
    end else begin
      mmio_26 <= _GEN_830;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Rob.scala 606:38]
      mmio_27 <= 1'h0;
    end else if (REG_5) begin // @[Rob.scala 606:38]
      mmio_27 <= _GEN_4770;
    end else if (REG_3) begin // @[Rob.scala 523:26]
      mmio_27 <= _GEN_4706; // @[Rob.scala 562:{22,22}]
    end else if (canEnqueue_1) begin
      if (5'h1b == allocatePtrVec_1_value) begin
        mmio_27 <= 1'h0;
      end else begin
        mmio_27 <= _GEN_831;
      end
    end else begin
      mmio_27 <= _GEN_831;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Rob.scala 606:38]
      mmio_28 <= 1'h0;
    end else if (REG_5) begin // @[Rob.scala 606:38]
      mmio_28 <= _GEN_4771;
    end else if (REG_3) begin // @[Rob.scala 523:26]
      mmio_28 <= _GEN_4707; // @[Rob.scala 562:{22,22}]
    end else if (canEnqueue_1) begin
      if (5'h1c == allocatePtrVec_1_value) begin
        mmio_28 <= 1'h0;
      end else begin
        mmio_28 <= _GEN_832;
      end
    end else begin
      mmio_28 <= _GEN_832;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Rob.scala 606:38]
      mmio_29 <= 1'h0;
    end else if (REG_5) begin // @[Rob.scala 606:38]
      mmio_29 <= _GEN_4772;
    end else if (REG_3) begin // @[Rob.scala 523:26]
      mmio_29 <= _GEN_4708; // @[Rob.scala 562:{22,22}]
    end else if (canEnqueue_1) begin
      if (5'h1d == allocatePtrVec_1_value) begin
        mmio_29 <= 1'h0;
      end else begin
        mmio_29 <= _GEN_833;
      end
    end else begin
      mmio_29 <= _GEN_833;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Rob.scala 606:38]
      mmio_30 <= 1'h0;
    end else if (REG_5) begin // @[Rob.scala 606:38]
      mmio_30 <= _GEN_4773;
    end else if (REG_3) begin // @[Rob.scala 523:26]
      mmio_30 <= _GEN_4709; // @[Rob.scala 562:{22,22}]
    end else if (canEnqueue_1) begin
      if (5'h1e == allocatePtrVec_1_value) begin
        mmio_30 <= 1'h0;
      end else begin
        mmio_30 <= _GEN_834;
      end
    end else begin
      mmio_30 <= _GEN_834;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Rob.scala 606:38]
      mmio_31 <= 1'h0;
    end else if (REG_5) begin // @[Rob.scala 606:38]
      mmio_31 <= _GEN_4774;
    end else if (REG_3) begin // @[Rob.scala 523:26]
      mmio_31 <= _GEN_4710; // @[Rob.scala 562:{22,22}]
    end else if (canEnqueue_1) begin
      if (5'h1f == allocatePtrVec_1_value) begin
        mmio_31 <= 1'h0;
      end else begin
        mmio_31 <= _GEN_835;
      end
    end else begin
      mmio_31 <= _GEN_835;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Rob.scala 806:49]
      allowEnqueue <= 1'h1;
    end else begin
      allowEnqueue <= _allowEnqueue_T_1 <= 6'h1e;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Rob.scala 764:23]
      state <= 1'h0;
    end else begin
      state <= io_redirect_valid | _state_next_T_2;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Rob.scala 523:26]
      hasBlockBackward <= 1'h0;
    end else if (canEnqueue_1) begin // @[Rob.scala 523:26]
      hasBlockBackward <= _GEN_1156;
    end else if (canEnqueue_0) begin // @[Rob.scala 495:18]
      hasBlockBackward <= _GEN_329; // @[Rob.scala 495:36]
    end else if (isEmpty) begin // @[Rob.scala 490:33]
      hasBlockBackward <= 1'h0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Rob.scala 523:26]
      hasNoSpecExec <= 1'h0;
    end else if (canEnqueue_1) begin // @[Rob.scala 523:26]
      hasNoSpecExec <= _GEN_1157;
    end else if (canEnqueue_0) begin // @[Rob.scala 497:63]
      hasNoSpecExec <= _GEN_330; // @[Rob.scala 497:78]
    end else if (_T_2 | _T_5) begin // @[Rob.scala 491:30]
      hasNoSpecExec <= 1'h0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Rob.scala 568:25]
      hasWFI <= 1'h0; // @[Rob.scala 569:12]
    end else if (~io_wfi_enable) begin // @[Rob.scala 523:26]
      hasWFI <= 1'h0;
    end else if (canEnqueue_1) begin // @[Rob.scala 523:26]
      hasWFI <= _GEN_1160;
    end else if (canEnqueue_0) begin // @[Rob.scala 512:80]
      hasWFI <= _GEN_333; // @[Rob.scala 513:12]
    end else if (REG_2 | io_flushOut_valid | wfi_timeout) begin // @[Rob.scala 502:23]
      hasWFI <= 1'h0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Rob.scala 506:17]
      wfi_cycles <= 20'h0; // @[Rob.scala 507:16]
    end else if (hasWFI) begin // @[Rob.scala 508:43]
      wfi_cycles <= _wfi_cycles_T_1; // @[Rob.scala 509:16]
    end else if (~hasWFI & REG) begin // @[Rob.scala 505:27]
      wfi_cycles <= 20'h0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[GTimer.scala 24:12]
      timer <= 64'h0;
    end else begin
      timer <= timer + 64'h1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Rob.scala 858:27]
      redirectState <= 1'h0; // @[Rob.scala 859:19]
    end else begin
      redirectState <= io_redirect_valid | _GEN_5276;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Rob.scala 1022:30]
      instrCntReg <= 64'h0;
    end else begin
      instrCntReg <= instrCntReg + _GEN_11347;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    writebacked[initvar] = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    store_data_writebacked[initvar] = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    interrupt_safe[initvar] = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    debug_microOp_cf_loadWaitBit[initvar] = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    debug_microOp_ctrl_isMove[initvar] = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    dt_eliminatedMove[initvar] = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    dt_isRVC[initvar] = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    dt_isXSTrap[initvar] = _RAND_7[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  valid_0 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  valid_1 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  valid_2 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  valid_3 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  valid_4 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  valid_5 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  valid_6 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  valid_7 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  valid_8 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  valid_9 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  valid_10 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  valid_11 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  valid_12 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  valid_13 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  valid_14 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  valid_15 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  valid_16 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  valid_17 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  valid_18 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  valid_19 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  valid_20 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  valid_21 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  valid_22 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  valid_23 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  valid_24 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  valid_25 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  valid_26 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  valid_27 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  valid_28 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  valid_29 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  valid_30 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  valid_31 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  mmio_0 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  mmio_1 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  mmio_2 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  mmio_3 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  mmio_4 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  mmio_5 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  mmio_6 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  mmio_7 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  mmio_8 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  mmio_9 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  mmio_10 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  mmio_11 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  mmio_12 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  mmio_13 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  mmio_14 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  mmio_15 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  mmio_16 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  mmio_17 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  mmio_18 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  mmio_19 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  mmio_20 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  mmio_21 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  mmio_22 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  mmio_23 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  mmio_24 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  mmio_25 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  mmio_26 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  mmio_27 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  mmio_28 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  mmio_29 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  mmio_30 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  mmio_31 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  walkPtrVec_0_flag = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  walkPtrVec_0_value = _RAND_73[4:0];
  _RAND_74 = {1{`RANDOM}};
  walkPtrVec_1_flag = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  walkPtrVec_1_value = _RAND_75[4:0];
  _RAND_76 = {1{`RANDOM}};
  allowEnqueue = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  state = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  hasBlockBackward = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  hasNoSpecExec = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  hasWFI = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  wfi_cycles = _RAND_81[19:0];
  _RAND_82 = {1{`RANDOM}};
  REG = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  REG_1 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  REG_2 = _RAND_84[0:0];
  _RAND_85 = {2{`RANDOM}};
  timer = _RAND_85[63:0];
  _RAND_86 = {1{`RANDOM}};
  io_enq_isEmpty_REG = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  REG_3 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  REG_4 = _RAND_88[4:0];
  _RAND_89 = {1{`RANDOM}};
  REG_5 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  REG_6 = _RAND_90[4:0];
  _RAND_91 = {1{`RANDOM}};
  intrBitSetReg = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  lastCycleFlush = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  io_exception_valid_REG = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  io_exception_bits_uop_ctrl_commitType_r = _RAND_94[2:0];
  _RAND_95 = {1{`RANDOM}};
  r_0 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  r_1 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  r_2 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  r_3 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  r_4 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  r_5 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  r_6 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  r_7 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  r_8 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  r_9 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  r_11 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  r_12 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  r_13 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  r_15 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  io_exception_bits_uop_ctrl_singleStep_r = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  io_exception_bits_uop_cf_crossPageIPFFix_r = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  io_exception_bits_isInterrupt_r = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  io_exception_bits_uop_cf_trigger_rfrontendHit_0 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  io_exception_bits_uop_cf_trigger_rfrontendHit_1 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  io_exception_bits_uop_cf_trigger_rfrontendHit_2 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  io_exception_bits_uop_cf_trigger_rfrontendHit_3 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  io_exception_bits_uop_cf_trigger_rbackendHit_0 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  io_exception_bits_uop_cf_trigger_rbackendHit_1 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  io_exception_bits_uop_cf_trigger_rbackendHit_2 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  io_exception_bits_uop_cf_trigger_rbackendHit_3 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  io_exception_bits_uop_cf_trigger_rbackendHit_4 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  io_exception_bits_uop_cf_trigger_rbackendHit_5 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  walkCounter = _RAND_122[5:0];
  _RAND_123 = {1{`RANDOM}};
  misPredBlockCounter = _RAND_123[2:0];
  _RAND_124 = {1{`RANDOM}};
  io_csr_fflags_REG_valid = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  io_csr_fflags_REG_bits = _RAND_125[4:0];
  _RAND_126 = {1{`RANDOM}};
  io_csr_dirty_fs_REG = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  io_lsq_scommit_REG = _RAND_127[1:0];
  _RAND_128 = {1{`RANDOM}};
  io_lsq_pendingld_REG = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  io_lsq_pendingst_REG = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  io_lsq_commit_REG = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  redirectHeadVec_0_flag = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  redirectHeadVec_0_value = _RAND_132[4:0];
  _RAND_133 = {1{`RANDOM}};
  redirectHeadVec_1_flag = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  redirectHeadVec_1_value = _RAND_134[4:0];
  _RAND_135 = {1{`RANDOM}};
  redirectTail_flag = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  redirectTail_value = _RAND_136[4:0];
  _RAND_137 = {1{`RANDOM}};
  redirectState = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  REG_7 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  REG_8 = _RAND_139[4:0];
  _RAND_140 = {1{`RANDOM}};
  REG_9 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  REG_10 = _RAND_141[4:0];
  _RAND_142 = {1{`RANDOM}};
  REG_11 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  REG_12 = _RAND_143[4:0];
  _RAND_144 = {1{`RANDOM}};
  REG_13 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  REG_14 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  REG_15 = _RAND_146[4:0];
  _RAND_147 = {1{`RANDOM}};
  REG_16 = _RAND_147[0:0];
  _RAND_148 = {2{`RANDOM}};
  instrCntReg = _RAND_148[63:0];
  _RAND_149 = {1{`RANDOM}};
  fuseCommitCnt_REG = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  fuseCommitCnt_REG_1 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  trueCommitCnt_REG = _RAND_151[1:0];
  _RAND_152 = {1{`RANDOM}};
  retireCounter_REG = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  dt_exuDebug_0_isMMIO = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  dt_exuDebug_0_isPerfCnt = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  dt_exuDebug_1_isMMIO = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  dt_exuDebug_1_isPerfCnt = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  dt_exuDebug_2_isMMIO = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  dt_exuDebug_2_isPerfCnt = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  dt_exuDebug_3_isMMIO = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  dt_exuDebug_3_isPerfCnt = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  dt_exuDebug_4_isMMIO = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  dt_exuDebug_4_isPerfCnt = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  dt_exuDebug_5_isMMIO = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  dt_exuDebug_5_isPerfCnt = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  dt_exuDebug_6_isMMIO = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  dt_exuDebug_6_isPerfCnt = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  dt_exuDebug_7_isMMIO = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  dt_exuDebug_7_isPerfCnt = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  dt_exuDebug_8_isMMIO = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  dt_exuDebug_8_isPerfCnt = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  dt_exuDebug_9_isMMIO = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  dt_exuDebug_9_isPerfCnt = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  dt_exuDebug_10_isMMIO = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  dt_exuDebug_10_isPerfCnt = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  dt_exuDebug_11_isMMIO = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  dt_exuDebug_11_isPerfCnt = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  dt_exuDebug_12_isMMIO = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  dt_exuDebug_12_isPerfCnt = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  dt_exuDebug_13_isMMIO = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  dt_exuDebug_13_isPerfCnt = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  dt_exuDebug_14_isMMIO = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  dt_exuDebug_14_isPerfCnt = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  dt_exuDebug_15_isMMIO = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  dt_exuDebug_15_isPerfCnt = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  dt_exuDebug_16_isMMIO = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  dt_exuDebug_16_isPerfCnt = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  dt_exuDebug_17_isMMIO = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  dt_exuDebug_17_isPerfCnt = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  dt_exuDebug_18_isMMIO = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  dt_exuDebug_18_isPerfCnt = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  dt_exuDebug_19_isMMIO = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  dt_exuDebug_19_isPerfCnt = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  dt_exuDebug_20_isMMIO = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  dt_exuDebug_20_isPerfCnt = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  dt_exuDebug_21_isMMIO = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  dt_exuDebug_21_isPerfCnt = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  dt_exuDebug_22_isMMIO = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  dt_exuDebug_22_isPerfCnt = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  dt_exuDebug_23_isMMIO = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  dt_exuDebug_23_isPerfCnt = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  dt_exuDebug_24_isMMIO = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  dt_exuDebug_24_isPerfCnt = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  dt_exuDebug_25_isMMIO = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  dt_exuDebug_25_isPerfCnt = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  dt_exuDebug_26_isMMIO = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  dt_exuDebug_26_isPerfCnt = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  dt_exuDebug_27_isMMIO = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  dt_exuDebug_27_isPerfCnt = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  dt_exuDebug_28_isMMIO = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  dt_exuDebug_28_isPerfCnt = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  dt_exuDebug_29_isMMIO = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  dt_exuDebug_29_isPerfCnt = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  dt_exuDebug_30_isMMIO = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  dt_exuDebug_30_isPerfCnt = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  dt_exuDebug_31_isMMIO = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  dt_exuDebug_31_isPerfCnt = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  difftest_io_valid_REG = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  difftest_io_valid_REG_1 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  difftest_io_valid_REG_2 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  difftest_io_special_REG = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  difftest_io_special_REG_1 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  difftest_io_special_REG_2 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  difftest_io_skip_REG = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  difftest_io_skip_REG_1 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  difftest_io_skip_REG_2 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  difftest_io_isRVC_REG = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  difftest_io_isRVC_REG_1 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  difftest_io_isRVC_REG_2 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  difftest_io_rfwen_REG = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  difftest_io_rfwen_REG_1 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  difftest_io_rfwen_REG_2 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  difftest_io_fpwen_REG = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  difftest_io_fpwen_REG_1 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  difftest_io_fpwen_REG_2 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  difftest_io_wpdest_REG = _RAND_235[5:0];
  _RAND_236 = {1{`RANDOM}};
  difftest_io_wpdest_REG_1 = _RAND_236[5:0];
  _RAND_237 = {1{`RANDOM}};
  difftest_io_wpdest_REG_2 = _RAND_237[5:0];
  _RAND_238 = {1{`RANDOM}};
  difftest_io_wdest_REG = _RAND_238[4:0];
  _RAND_239 = {1{`RANDOM}};
  difftest_io_wdest_REG_1 = _RAND_239[4:0];
  _RAND_240 = {1{`RANDOM}};
  difftest_io_wdest_REG_2 = _RAND_240[4:0];
  _RAND_241 = {1{`RANDOM}};
  difftest_io_valid_REG_3 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  difftest_io_valid_REG_4 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  difftest_io_valid_REG_5 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  difftest_io_special_REG_3 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  difftest_io_special_REG_4 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  difftest_io_special_REG_5 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  difftest_io_skip_REG_3 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  difftest_io_skip_REG_4 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  difftest_io_skip_REG_5 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  difftest_io_isRVC_REG_3 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  difftest_io_isRVC_REG_4 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  difftest_io_isRVC_REG_5 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  difftest_io_rfwen_REG_3 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  difftest_io_rfwen_REG_4 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  difftest_io_rfwen_REG_5 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  difftest_io_fpwen_REG_3 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  difftest_io_fpwen_REG_4 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  difftest_io_fpwen_REG_5 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  difftest_io_wpdest_REG_3 = _RAND_259[5:0];
  _RAND_260 = {1{`RANDOM}};
  difftest_io_wpdest_REG_4 = _RAND_260[5:0];
  _RAND_261 = {1{`RANDOM}};
  difftest_io_wpdest_REG_5 = _RAND_261[5:0];
  _RAND_262 = {1{`RANDOM}};
  difftest_io_wdest_REG_3 = _RAND_262[4:0];
  _RAND_263 = {1{`RANDOM}};
  difftest_io_wdest_REG_4 = _RAND_263[4:0];
  _RAND_264 = {1{`RANDOM}};
  difftest_io_wdest_REG_5 = _RAND_264[4:0];
  _RAND_265 = {1{`RANDOM}};
  validEntriesBanks_0 = _RAND_265[5:0];
  _RAND_266 = {1{`RANDOM}};
  validEntries = _RAND_266[5:0];
  _RAND_267 = {1{`RANDOM}};
  REG_19 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  REG_20_0 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  REG_20_1 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  REG_21 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  REG_22 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  REG_23_0 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  REG_23_1 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  REG_24 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  REG_25_0 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  REG_25_1 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  REG_26 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  REG_27_0 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  REG_27_1 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  REG_28 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  REG_29_0 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  REG_29_1 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  REG_30 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  io_perf_0_value_REG = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  io_perf_0_value_REG_1 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  io_perf_1_value_REG = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  io_perf_1_value_REG_1 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  io_perf_2_value_REG = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  io_perf_2_value_REG_1 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  io_perf_3_value_REG = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  io_perf_3_value_REG_1 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  io_perf_4_value_REG = _RAND_292[1:0];
  _RAND_293 = {1{`RANDOM}};
  io_perf_4_value_REG_1 = _RAND_293[1:0];
  _RAND_294 = {1{`RANDOM}};
  io_perf_5_value_REG = _RAND_294[2:0];
  _RAND_295 = {1{`RANDOM}};
  io_perf_5_value_REG_1 = _RAND_295[2:0];
  _RAND_296 = {1{`RANDOM}};
  io_perf_6_value_REG = _RAND_296[1:0];
  _RAND_297 = {1{`RANDOM}};
  io_perf_6_value_REG_1 = _RAND_297[1:0];
  _RAND_298 = {1{`RANDOM}};
  io_perf_7_value_REG = _RAND_298[1:0];
  _RAND_299 = {1{`RANDOM}};
  io_perf_7_value_REG_1 = _RAND_299[1:0];
  _RAND_300 = {1{`RANDOM}};
  io_perf_8_value_REG = _RAND_300[1:0];
  _RAND_301 = {1{`RANDOM}};
  io_perf_8_value_REG_1 = _RAND_301[1:0];
  _RAND_302 = {1{`RANDOM}};
  io_perf_9_value_REG = _RAND_302[1:0];
  _RAND_303 = {1{`RANDOM}};
  io_perf_9_value_REG_1 = _RAND_303[1:0];
  _RAND_304 = {1{`RANDOM}};
  io_perf_10_value_REG = _RAND_304[1:0];
  _RAND_305 = {1{`RANDOM}};
  io_perf_10_value_REG_1 = _RAND_305[1:0];
  _RAND_306 = {1{`RANDOM}};
  io_perf_11_value_REG = _RAND_306[1:0];
  _RAND_307 = {1{`RANDOM}};
  io_perf_11_value_REG_1 = _RAND_307[1:0];
  _RAND_308 = {1{`RANDOM}};
  io_perf_12_value_REG = _RAND_308[1:0];
  _RAND_309 = {1{`RANDOM}};
  io_perf_12_value_REG_1 = _RAND_309[1:0];
  _RAND_310 = {1{`RANDOM}};
  io_perf_13_value_REG = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  io_perf_13_value_REG_1 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  io_perf_14_value_REG = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  io_perf_14_value_REG_1 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  io_perf_15_value_REG = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  io_perf_15_value_REG_1 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  io_perf_16_value_REG = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  io_perf_16_value_REG_1 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  io_perf_17_value_REG = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  io_perf_17_value_REG_1 = _RAND_319[0:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    valid_0 = 1'h0;
  end
  if (reset) begin
    valid_1 = 1'h0;
  end
  if (reset) begin
    valid_2 = 1'h0;
  end
  if (reset) begin
    valid_3 = 1'h0;
  end
  if (reset) begin
    valid_4 = 1'h0;
  end
  if (reset) begin
    valid_5 = 1'h0;
  end
  if (reset) begin
    valid_6 = 1'h0;
  end
  if (reset) begin
    valid_7 = 1'h0;
  end
  if (reset) begin
    valid_8 = 1'h0;
  end
  if (reset) begin
    valid_9 = 1'h0;
  end
  if (reset) begin
    valid_10 = 1'h0;
  end
  if (reset) begin
    valid_11 = 1'h0;
  end
  if (reset) begin
    valid_12 = 1'h0;
  end
  if (reset) begin
    valid_13 = 1'h0;
  end
  if (reset) begin
    valid_14 = 1'h0;
  end
  if (reset) begin
    valid_15 = 1'h0;
  end
  if (reset) begin
    valid_16 = 1'h0;
  end
  if (reset) begin
    valid_17 = 1'h0;
  end
  if (reset) begin
    valid_18 = 1'h0;
  end
  if (reset) begin
    valid_19 = 1'h0;
  end
  if (reset) begin
    valid_20 = 1'h0;
  end
  if (reset) begin
    valid_21 = 1'h0;
  end
  if (reset) begin
    valid_22 = 1'h0;
  end
  if (reset) begin
    valid_23 = 1'h0;
  end
  if (reset) begin
    valid_24 = 1'h0;
  end
  if (reset) begin
    valid_25 = 1'h0;
  end
  if (reset) begin
    valid_26 = 1'h0;
  end
  if (reset) begin
    valid_27 = 1'h0;
  end
  if (reset) begin
    valid_28 = 1'h0;
  end
  if (reset) begin
    valid_29 = 1'h0;
  end
  if (reset) begin
    valid_30 = 1'h0;
  end
  if (reset) begin
    valid_31 = 1'h0;
  end
  if (reset) begin
    mmio_0 = 1'h0;
  end
  if (reset) begin
    mmio_1 = 1'h0;
  end
  if (reset) begin
    mmio_2 = 1'h0;
  end
  if (reset) begin
    mmio_3 = 1'h0;
  end
  if (reset) begin
    mmio_4 = 1'h0;
  end
  if (reset) begin
    mmio_5 = 1'h0;
  end
  if (reset) begin
    mmio_6 = 1'h0;
  end
  if (reset) begin
    mmio_7 = 1'h0;
  end
  if (reset) begin
    mmio_8 = 1'h0;
  end
  if (reset) begin
    mmio_9 = 1'h0;
  end
  if (reset) begin
    mmio_10 = 1'h0;
  end
  if (reset) begin
    mmio_11 = 1'h0;
  end
  if (reset) begin
    mmio_12 = 1'h0;
  end
  if (reset) begin
    mmio_13 = 1'h0;
  end
  if (reset) begin
    mmio_14 = 1'h0;
  end
  if (reset) begin
    mmio_15 = 1'h0;
  end
  if (reset) begin
    mmio_16 = 1'h0;
  end
  if (reset) begin
    mmio_17 = 1'h0;
  end
  if (reset) begin
    mmio_18 = 1'h0;
  end
  if (reset) begin
    mmio_19 = 1'h0;
  end
  if (reset) begin
    mmio_20 = 1'h0;
  end
  if (reset) begin
    mmio_21 = 1'h0;
  end
  if (reset) begin
    mmio_22 = 1'h0;
  end
  if (reset) begin
    mmio_23 = 1'h0;
  end
  if (reset) begin
    mmio_24 = 1'h0;
  end
  if (reset) begin
    mmio_25 = 1'h0;
  end
  if (reset) begin
    mmio_26 = 1'h0;
  end
  if (reset) begin
    mmio_27 = 1'h0;
  end
  if (reset) begin
    mmio_28 = 1'h0;
  end
  if (reset) begin
    mmio_29 = 1'h0;
  end
  if (reset) begin
    mmio_30 = 1'h0;
  end
  if (reset) begin
    mmio_31 = 1'h0;
  end
  if (reset) begin
    allowEnqueue = 1'h1;
  end
  if (reset) begin
    state = 1'h0;
  end
  if (reset) begin
    hasBlockBackward = 1'h0;
  end
  if (reset) begin
    hasNoSpecExec = 1'h0;
  end
  if (reset) begin
    hasWFI = 1'h0;
  end
  if (reset) begin
    wfi_cycles = 20'h0;
  end
  if (reset) begin
    timer = 64'h0;
  end
  if (reset) begin
    redirectState = 1'h0;
  end
  if (reset) begin
    instrCntReg = 64'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule

