module DelayN_114(
  input  [3:0] io_in,
  output [3:0] io_out
);
  assign io_out = io_in; // @[Hold.scala 92:10]
endmodule

